VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO map9v3
  CLASS BLOCK ;
  FOREIGN map9v3 ;
  ORIGIN 1.900 4.000 ;
  SIZE 231.000 BY 208.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 200.400 226.800 201.600 ;
        RECT 1.200 191.800 2.000 200.400 ;
        RECT 5.400 195.800 6.200 200.400 ;
        RECT 10.800 191.800 11.600 200.400 ;
        RECT 12.400 195.800 13.200 200.400 ;
        RECT 15.600 195.800 16.400 200.400 ;
        RECT 17.200 195.800 18.000 200.400 ;
        RECT 23.600 193.000 24.400 200.400 ;
        RECT 28.400 196.200 29.200 200.400 ;
        RECT 31.600 195.800 32.400 200.400 ;
        RECT 33.200 195.800 34.000 200.400 ;
        RECT 36.400 195.800 37.200 200.400 ;
        RECT 42.800 191.800 43.600 200.400 ;
        RECT 45.000 195.800 45.800 200.400 ;
        RECT 49.200 191.800 50.000 200.400 ;
        RECT 50.800 191.800 51.600 200.400 ;
        RECT 55.600 193.000 56.400 200.400 ;
        RECT 60.400 195.800 61.200 200.400 ;
        RECT 63.600 195.800 64.400 200.400 ;
        RECT 65.200 191.800 66.000 200.400 ;
        RECT 70.000 191.800 70.800 200.400 ;
        RECT 74.200 195.800 75.000 200.400 ;
        RECT 78.000 193.000 78.800 200.400 ;
        RECT 81.200 195.800 82.000 200.400 ;
        RECT 84.400 195.800 85.200 200.400 ;
        RECT 88.200 195.800 89.000 200.400 ;
        RECT 92.400 191.800 93.200 200.400 ;
        RECT 95.600 195.800 96.400 200.400 ;
        RECT 97.200 191.800 98.000 200.400 ;
        RECT 102.000 195.800 102.800 200.400 ;
        RECT 105.200 195.800 106.000 200.400 ;
        RECT 108.400 195.800 109.200 200.400 ;
        RECT 111.600 193.000 112.400 200.400 ;
        RECT 114.800 195.800 115.600 200.400 ;
        RECT 118.000 195.800 118.800 200.400 ;
        RECT 121.200 195.800 122.000 200.400 ;
        RECT 124.400 195.800 125.200 200.400 ;
        RECT 132.400 195.800 133.200 200.400 ;
        RECT 135.600 195.800 136.400 200.400 ;
        RECT 142.000 195.800 142.800 200.400 ;
        RECT 145.200 195.800 146.000 200.400 ;
        RECT 148.400 195.800 149.200 200.400 ;
        RECT 153.200 193.000 154.000 200.400 ;
        RECT 158.000 193.000 158.800 200.400 ;
        RECT 161.200 195.800 162.000 200.400 ;
        RECT 164.400 195.800 165.200 200.400 ;
        RECT 167.600 195.800 168.400 200.400 ;
        RECT 174.000 195.800 174.800 200.400 ;
        RECT 177.200 195.800 178.000 200.400 ;
        RECT 185.200 195.800 186.000 200.400 ;
        RECT 188.400 195.800 189.200 200.400 ;
        RECT 191.600 195.800 192.400 200.400 ;
        RECT 194.800 195.800 195.600 200.400 ;
        RECT 199.600 193.000 200.400 200.400 ;
        RECT 206.000 193.000 206.800 200.400 ;
        RECT 141.800 191.800 142.600 192.000 ;
        RECT 145.200 191.800 146.000 192.400 ;
        RECT 119.000 191.200 146.000 191.800 ;
        RECT 164.400 191.800 165.200 192.400 ;
        RECT 167.600 191.800 168.600 192.000 ;
        RECT 212.400 191.800 213.200 200.400 ;
        RECT 215.600 195.800 216.400 200.400 ;
        RECT 218.800 193.000 219.600 200.400 ;
        RECT 164.400 191.200 191.400 191.800 ;
        RECT 119.000 191.000 119.800 191.200 ;
        RECT 190.600 191.000 191.400 191.200 ;
        RECT 18.200 170.800 19.000 171.000 ;
        RECT 157.000 170.800 157.800 171.000 ;
        RECT 221.000 170.800 221.800 171.000 ;
        RECT 18.200 170.200 45.200 170.800 ;
        RECT 130.800 170.200 157.800 170.800 ;
        RECT 194.800 170.200 221.800 170.800 ;
        RECT 1.200 161.600 2.000 170.200 ;
        RECT 5.400 161.600 6.200 166.200 ;
        RECT 7.600 161.600 8.400 170.200 ;
        RECT 41.000 170.000 41.800 170.200 ;
        RECT 44.400 169.600 45.200 170.200 ;
        RECT 11.800 161.600 12.600 166.200 ;
        RECT 14.000 161.600 14.800 166.200 ;
        RECT 17.200 161.600 18.000 166.200 ;
        RECT 20.400 161.600 21.200 166.200 ;
        RECT 23.600 161.600 24.400 166.200 ;
        RECT 31.600 161.600 32.400 166.200 ;
        RECT 34.800 161.600 35.600 166.200 ;
        RECT 41.200 161.600 42.000 166.200 ;
        RECT 44.400 161.600 45.200 166.200 ;
        RECT 47.600 161.600 48.400 166.200 ;
        RECT 52.400 161.600 53.200 165.800 ;
        RECT 55.600 161.600 56.400 166.200 ;
        RECT 57.200 161.600 58.000 170.200 ;
        RECT 61.400 161.600 62.200 166.200 ;
        RECT 64.200 161.600 65.000 166.200 ;
        RECT 68.400 161.600 69.200 170.200 ;
        RECT 70.600 161.600 71.400 166.200 ;
        RECT 74.800 161.600 75.600 170.200 ;
        RECT 78.000 161.600 79.000 168.800 ;
        RECT 84.200 162.200 85.200 168.800 ;
        RECT 84.200 161.600 85.000 162.200 ;
        RECT 89.200 161.600 90.000 166.200 ;
        RECT 92.400 161.600 93.200 170.200 ;
        RECT 96.600 161.600 97.400 166.200 ;
        RECT 99.400 161.600 100.200 166.200 ;
        RECT 103.600 161.600 104.400 170.200 ;
        RECT 108.400 161.600 109.200 170.200 ;
        RECT 111.600 161.600 112.400 169.800 ;
        RECT 114.800 161.600 115.600 166.200 ;
        RECT 119.600 161.600 120.400 170.200 ;
        RECT 130.800 169.600 131.600 170.200 ;
        RECT 134.200 170.000 135.000 170.200 ;
        RECT 122.800 161.600 123.600 169.000 ;
        RECT 127.600 161.600 128.400 166.200 ;
        RECT 130.800 161.600 131.600 166.200 ;
        RECT 134.000 161.600 134.800 166.200 ;
        RECT 140.400 161.600 141.200 166.200 ;
        RECT 143.600 161.600 144.400 166.200 ;
        RECT 151.600 161.600 152.400 166.200 ;
        RECT 154.800 161.600 155.600 166.200 ;
        RECT 158.000 161.600 158.800 166.200 ;
        RECT 161.200 161.600 162.000 166.200 ;
        RECT 166.000 161.600 166.800 169.000 ;
        RECT 169.200 161.600 170.000 166.200 ;
        RECT 174.000 161.600 174.800 169.800 ;
        RECT 179.200 161.600 180.000 170.200 ;
        RECT 194.800 169.600 195.600 170.200 ;
        RECT 198.200 170.000 199.000 170.200 ;
        RECT 183.600 161.600 184.400 169.000 ;
        RECT 188.400 161.600 189.200 166.200 ;
        RECT 191.600 161.600 192.400 166.200 ;
        RECT 194.800 161.600 195.600 166.200 ;
        RECT 198.000 161.600 198.800 166.200 ;
        RECT 204.400 161.600 205.200 166.200 ;
        RECT 207.600 161.600 208.400 166.200 ;
        RECT 215.600 161.600 216.400 166.200 ;
        RECT 218.800 161.600 219.600 166.200 ;
        RECT 222.000 161.600 222.800 166.200 ;
        RECT 225.200 161.600 226.000 166.200 ;
        RECT 0.400 160.400 226.800 161.600 ;
        RECT 2.800 153.000 3.600 160.400 ;
        RECT 9.200 151.800 10.000 160.400 ;
        RECT 10.800 151.800 11.600 160.400 ;
        RECT 15.000 155.800 15.800 160.400 ;
        RECT 17.200 155.800 18.000 160.400 ;
        RECT 20.400 155.800 21.200 160.400 ;
        RECT 23.600 155.800 24.400 160.400 ;
        RECT 30.000 155.800 30.800 160.400 ;
        RECT 33.200 155.800 34.000 160.400 ;
        RECT 41.200 155.800 42.000 160.400 ;
        RECT 44.400 155.800 45.200 160.400 ;
        RECT 47.600 155.800 48.400 160.400 ;
        RECT 50.800 155.800 51.600 160.400 ;
        RECT 54.600 155.800 55.400 160.400 ;
        RECT 20.400 151.800 21.200 152.400 ;
        RECT 23.800 151.800 24.600 152.000 ;
        RECT 58.800 151.800 59.600 160.400 ;
        RECT 62.000 152.200 62.800 160.400 ;
        RECT 65.200 155.800 66.000 160.400 ;
        RECT 66.800 151.800 67.600 160.400 ;
        RECT 73.200 155.800 74.000 160.400 ;
        RECT 76.400 155.800 77.200 160.400 ;
        RECT 79.600 155.800 80.400 160.400 ;
        RECT 86.000 155.800 86.800 160.400 ;
        RECT 89.200 155.800 90.000 160.400 ;
        RECT 97.200 155.800 98.000 160.400 ;
        RECT 100.400 155.800 101.200 160.400 ;
        RECT 103.600 155.800 104.400 160.400 ;
        RECT 106.800 155.800 107.600 160.400 ;
        RECT 76.400 151.800 77.200 152.400 ;
        RECT 79.600 151.800 80.600 152.000 ;
        RECT 108.400 151.800 109.200 160.400 ;
        RECT 111.600 151.800 112.400 160.400 ;
        RECT 114.800 151.800 115.600 160.400 ;
        RECT 118.000 151.800 118.800 160.400 ;
        RECT 121.200 151.800 122.000 160.400 ;
        RECT 124.400 155.800 125.200 160.400 ;
        RECT 127.600 155.800 128.400 160.400 ;
        RECT 130.800 155.800 131.600 160.400 ;
        RECT 137.200 155.800 138.000 160.400 ;
        RECT 140.400 155.800 141.200 160.400 ;
        RECT 148.400 155.800 149.200 160.400 ;
        RECT 151.600 155.800 152.400 160.400 ;
        RECT 154.800 155.800 155.600 160.400 ;
        RECT 158.000 155.800 158.800 160.400 ;
        RECT 161.400 159.800 162.200 160.400 ;
        RECT 161.200 153.200 162.200 159.800 ;
        RECT 167.400 153.200 168.400 160.400 ;
        RECT 127.600 151.800 128.400 152.400 ;
        RECT 172.400 152.200 173.200 160.400 ;
        RECT 131.000 151.800 131.800 152.000 ;
        RECT 177.600 151.800 178.400 160.400 ;
        RECT 182.000 155.800 182.800 160.400 ;
        RECT 185.200 155.800 186.000 160.400 ;
        RECT 188.400 155.800 189.200 160.400 ;
        RECT 191.600 155.800 192.400 160.400 ;
        RECT 198.000 155.800 198.800 160.400 ;
        RECT 201.200 155.800 202.000 160.400 ;
        RECT 209.200 155.800 210.000 160.400 ;
        RECT 212.400 155.800 213.200 160.400 ;
        RECT 215.600 155.800 216.400 160.400 ;
        RECT 218.800 155.800 219.600 160.400 ;
        RECT 222.000 153.000 222.800 160.400 ;
        RECT 188.400 151.800 189.200 152.400 ;
        RECT 191.600 151.800 192.600 152.000 ;
        RECT 20.400 151.200 47.400 151.800 ;
        RECT 76.400 151.200 103.400 151.800 ;
        RECT 127.600 151.200 154.600 151.800 ;
        RECT 188.400 151.200 215.400 151.800 ;
        RECT 46.600 151.000 47.400 151.200 ;
        RECT 102.600 151.000 103.400 151.200 ;
        RECT 153.800 151.000 154.600 151.200 ;
        RECT 214.600 151.000 215.400 151.200 ;
        RECT 72.600 130.800 73.400 131.000 ;
        RECT 186.200 130.800 187.000 131.000 ;
        RECT 72.600 130.200 99.600 130.800 ;
        RECT 186.200 130.200 213.200 130.800 ;
        RECT 1.800 121.600 2.600 126.200 ;
        RECT 6.000 121.600 6.800 130.200 ;
        RECT 7.600 121.600 8.400 126.200 ;
        RECT 12.400 121.600 13.200 129.000 ;
        RECT 22.000 121.600 22.800 129.000 ;
        RECT 26.800 121.600 27.600 128.200 ;
        RECT 39.600 121.600 40.400 126.200 ;
        RECT 42.800 121.600 43.600 130.200 ;
        RECT 95.400 130.000 96.200 130.200 ;
        RECT 98.800 129.600 99.600 130.200 ;
        RECT 47.600 121.600 48.400 126.200 ;
        RECT 50.800 121.600 51.600 125.800 ;
        RECT 54.000 121.600 54.800 126.200 ;
        RECT 57.200 121.600 58.000 125.800 ;
        RECT 62.000 121.600 62.800 126.200 ;
        RECT 65.200 121.600 66.000 129.000 ;
        RECT 68.400 121.600 69.200 126.200 ;
        RECT 71.600 121.600 72.400 126.200 ;
        RECT 74.800 121.600 75.600 126.200 ;
        RECT 78.000 121.600 78.800 126.200 ;
        RECT 86.000 121.600 86.800 126.200 ;
        RECT 89.200 121.600 90.000 126.200 ;
        RECT 95.600 121.600 96.400 126.200 ;
        RECT 98.800 121.600 99.600 126.200 ;
        RECT 102.000 121.600 102.800 126.200 ;
        RECT 105.200 121.600 106.000 130.200 ;
        RECT 108.400 121.600 109.200 130.200 ;
        RECT 111.600 121.600 112.400 130.200 ;
        RECT 114.800 121.600 115.600 130.200 ;
        RECT 118.000 121.600 118.800 130.200 ;
        RECT 119.600 121.600 120.400 130.200 ;
        RECT 122.800 121.600 123.600 130.200 ;
        RECT 126.000 121.600 126.800 130.200 ;
        RECT 129.200 121.600 130.000 130.200 ;
        RECT 132.400 121.600 133.200 130.200 ;
        RECT 135.600 121.600 136.400 129.000 ;
        RECT 138.800 121.600 139.600 130.200 ;
        RECT 143.600 121.600 144.400 129.000 ;
        RECT 150.000 121.600 150.800 126.200 ;
        RECT 152.200 121.600 153.000 126.200 ;
        RECT 156.400 121.600 157.200 130.200 ;
        RECT 158.000 121.600 158.800 130.200 ;
        RECT 162.200 121.600 163.000 126.200 ;
        RECT 165.000 121.600 165.800 126.200 ;
        RECT 169.200 121.600 170.000 130.200 ;
        RECT 209.000 130.000 209.800 130.200 ;
        RECT 212.400 129.600 213.200 130.200 ;
        RECT 174.000 121.600 174.800 129.000 ;
        RECT 178.800 121.600 179.600 126.200 ;
        RECT 182.000 121.600 182.800 126.200 ;
        RECT 185.200 121.600 186.000 126.200 ;
        RECT 188.400 121.600 189.200 126.200 ;
        RECT 191.600 121.600 192.400 126.200 ;
        RECT 199.600 121.600 200.400 126.200 ;
        RECT 202.800 121.600 203.600 126.200 ;
        RECT 209.200 121.600 210.000 126.200 ;
        RECT 212.400 121.600 213.200 126.200 ;
        RECT 215.600 121.600 216.400 126.200 ;
        RECT 218.800 121.600 219.600 129.000 ;
        RECT 0.400 120.400 226.800 121.600 ;
        RECT 2.800 113.000 3.600 120.400 ;
        RECT 6.000 115.800 6.800 120.400 ;
        RECT 9.200 115.800 10.000 120.400 ;
        RECT 12.400 115.800 13.200 120.400 ;
        RECT 15.600 115.800 16.400 120.400 ;
        RECT 23.600 115.800 24.400 120.400 ;
        RECT 26.800 115.800 27.600 120.400 ;
        RECT 33.200 115.800 34.000 120.400 ;
        RECT 36.400 115.800 37.200 120.400 ;
        RECT 39.600 115.800 40.400 120.400 ;
        RECT 42.800 115.800 43.600 120.400 ;
        RECT 50.800 113.000 51.600 120.400 ;
        RECT 33.000 111.800 33.800 112.000 ;
        RECT 36.400 111.800 37.200 112.400 ;
        RECT 54.000 111.800 54.800 120.400 ;
        RECT 58.800 115.800 59.600 120.400 ;
        RECT 62.000 115.800 62.800 120.400 ;
        RECT 65.200 116.200 66.000 120.400 ;
        RECT 68.400 115.800 69.200 120.400 ;
        RECT 70.000 115.800 70.800 120.400 ;
        RECT 73.200 116.200 74.000 120.400 ;
        RECT 76.400 111.800 77.200 120.400 ;
        RECT 79.600 111.800 80.400 120.400 ;
        RECT 81.200 111.800 82.000 120.400 ;
        RECT 84.400 113.000 85.200 120.400 ;
        RECT 89.200 111.800 90.000 120.400 ;
        RECT 92.400 111.800 93.200 120.400 ;
        RECT 95.600 111.800 96.400 120.400 ;
        RECT 97.200 111.800 98.000 120.400 ;
        RECT 100.400 113.000 101.200 120.400 ;
        RECT 103.600 115.800 104.400 120.400 ;
        RECT 108.400 113.000 109.200 120.400 ;
        RECT 111.600 111.800 112.400 120.400 ;
        RECT 114.400 111.800 115.200 120.400 ;
        RECT 119.600 112.200 120.400 120.400 ;
        RECT 124.400 113.000 125.200 120.400 ;
        RECT 127.600 111.800 128.400 120.400 ;
        RECT 130.800 113.000 131.600 120.400 ;
        RECT 134.000 111.800 134.800 120.400 ;
        RECT 137.200 115.800 138.000 120.400 ;
        RECT 140.400 115.800 141.200 120.400 ;
        RECT 143.600 115.800 144.400 120.400 ;
        RECT 150.000 115.800 150.800 120.400 ;
        RECT 153.200 115.800 154.000 120.400 ;
        RECT 161.200 115.800 162.000 120.400 ;
        RECT 164.400 115.800 165.200 120.400 ;
        RECT 167.600 115.800 168.400 120.400 ;
        RECT 170.800 115.800 171.600 120.400 ;
        RECT 175.600 113.000 176.400 120.400 ;
        RECT 180.400 115.800 181.200 120.400 ;
        RECT 183.600 115.800 184.400 120.400 ;
        RECT 186.800 115.800 187.600 120.400 ;
        RECT 193.200 115.800 194.000 120.400 ;
        RECT 196.400 115.800 197.200 120.400 ;
        RECT 204.400 115.800 205.200 120.400 ;
        RECT 207.600 115.800 208.400 120.400 ;
        RECT 210.800 115.800 211.600 120.400 ;
        RECT 214.000 115.800 214.800 120.400 ;
        RECT 217.200 115.800 218.000 120.400 ;
        RECT 220.400 113.000 221.200 120.400 ;
        RECT 140.400 111.800 141.200 112.400 ;
        RECT 143.600 111.800 144.600 112.000 ;
        RECT 183.600 111.800 184.400 112.400 ;
        RECT 187.000 111.800 187.800 112.000 ;
        RECT 10.200 111.200 37.200 111.800 ;
        RECT 140.400 111.200 167.400 111.800 ;
        RECT 183.600 111.200 210.600 111.800 ;
        RECT 10.200 111.000 11.000 111.200 ;
        RECT 166.600 111.000 167.400 111.200 ;
        RECT 209.800 111.000 210.600 111.200 ;
        RECT 64.600 90.800 65.400 91.000 ;
        RECT 106.200 90.800 107.000 91.000 ;
        RECT 211.400 90.800 212.200 91.000 ;
        RECT 64.600 90.200 91.600 90.800 ;
        RECT 106.200 90.200 133.200 90.800 ;
        RECT 185.200 90.200 212.200 90.800 ;
        RECT 1.200 81.600 2.000 86.200 ;
        RECT 5.000 81.600 5.800 86.200 ;
        RECT 9.200 81.600 10.000 90.200 ;
        RECT 10.800 81.600 11.600 86.200 ;
        RECT 14.000 81.600 14.800 85.800 ;
        RECT 18.800 81.600 19.600 85.800 ;
        RECT 22.000 81.600 22.800 86.200 ;
        RECT 25.200 81.600 26.000 86.200 ;
        RECT 28.400 81.600 29.200 86.200 ;
        RECT 30.000 81.600 30.800 90.200 ;
        RECT 34.200 81.600 35.000 86.200 ;
        RECT 38.000 81.600 38.800 86.200 ;
        RECT 41.200 81.600 42.000 90.200 ;
        RECT 45.400 81.600 46.200 86.200 ;
        RECT 48.200 81.600 49.000 86.200 ;
        RECT 52.400 81.600 53.200 90.200 ;
        RECT 87.400 90.000 88.200 90.200 ;
        RECT 54.000 81.600 54.800 86.200 ;
        RECT 57.200 81.600 58.000 89.800 ;
        RECT 90.800 89.600 91.600 90.200 ;
        RECT 129.000 90.000 130.000 90.200 ;
        RECT 132.400 89.600 133.200 90.200 ;
        RECT 60.400 81.600 61.200 86.200 ;
        RECT 63.600 81.600 64.400 86.200 ;
        RECT 66.800 81.600 67.600 86.200 ;
        RECT 70.000 81.600 70.800 86.200 ;
        RECT 78.000 81.600 78.800 86.200 ;
        RECT 81.200 81.600 82.000 86.200 ;
        RECT 87.600 81.600 88.400 86.200 ;
        RECT 90.800 81.600 91.600 86.200 ;
        RECT 94.000 81.600 94.800 86.200 ;
        RECT 98.800 81.600 99.600 89.000 ;
        RECT 102.000 81.600 102.800 86.200 ;
        RECT 105.200 81.600 106.000 86.200 ;
        RECT 108.400 81.600 109.200 86.200 ;
        RECT 111.600 81.600 112.400 86.200 ;
        RECT 119.600 81.600 120.400 86.200 ;
        RECT 122.800 81.600 123.600 86.200 ;
        RECT 129.200 81.600 130.000 86.200 ;
        RECT 132.400 81.600 133.200 86.200 ;
        RECT 135.600 81.600 136.400 86.200 ;
        RECT 139.400 81.600 140.200 86.200 ;
        RECT 143.600 81.600 144.400 90.200 ;
        RECT 148.400 81.600 149.200 89.000 ;
        RECT 154.800 81.600 155.600 90.200 ;
        RECT 158.000 81.600 159.000 88.800 ;
        RECT 164.200 82.200 165.200 88.800 ;
        RECT 164.200 81.600 165.000 82.200 ;
        RECT 167.600 81.600 168.400 90.200 ;
        RECT 171.800 81.600 172.600 86.200 ;
        RECT 174.000 81.600 174.800 90.200 ;
        RECT 185.200 89.600 186.000 90.200 ;
        RECT 188.400 90.000 189.400 90.200 ;
        RECT 178.200 81.600 179.000 86.200 ;
        RECT 182.000 81.600 182.800 86.200 ;
        RECT 185.200 81.600 186.000 86.200 ;
        RECT 188.400 81.600 189.200 86.200 ;
        RECT 194.800 81.600 195.600 86.200 ;
        RECT 198.000 81.600 198.800 86.200 ;
        RECT 206.000 81.600 206.800 86.200 ;
        RECT 209.200 81.600 210.000 86.200 ;
        RECT 212.400 81.600 213.200 86.200 ;
        RECT 215.600 81.600 216.400 86.200 ;
        RECT 218.800 81.600 219.600 89.800 ;
        RECT 224.000 81.600 224.800 90.200 ;
        RECT 0.400 80.400 226.800 81.600 ;
        RECT 2.800 73.000 3.600 80.400 ;
        RECT 7.600 73.000 8.400 80.400 ;
        RECT 10.800 75.800 11.600 80.400 ;
        RECT 14.000 75.800 14.800 80.400 ;
        RECT 17.200 75.800 18.000 80.400 ;
        RECT 20.400 75.800 21.200 80.400 ;
        RECT 28.400 75.800 29.200 80.400 ;
        RECT 31.600 75.800 32.400 80.400 ;
        RECT 38.000 75.800 38.800 80.400 ;
        RECT 41.200 75.800 42.000 80.400 ;
        RECT 44.400 75.800 45.200 80.400 ;
        RECT 47.600 75.800 48.400 80.400 ;
        RECT 52.400 76.200 53.200 80.400 ;
        RECT 55.600 75.800 56.400 80.400 ;
        RECT 57.200 75.800 58.000 80.400 ;
        RECT 60.400 76.200 61.200 80.400 ;
        RECT 64.200 75.800 65.000 80.400 ;
        RECT 37.800 71.800 38.600 72.000 ;
        RECT 41.200 71.800 42.000 72.400 ;
        RECT 68.400 71.800 69.200 80.400 ;
        RECT 70.000 71.800 70.800 80.400 ;
        RECT 74.200 75.800 75.000 80.400 ;
        RECT 76.400 75.800 77.200 80.400 ;
        RECT 79.600 75.800 80.400 80.400 ;
        RECT 81.200 71.800 82.000 80.400 ;
        RECT 84.400 73.000 85.200 80.400 ;
        RECT 89.200 75.800 90.000 80.400 ;
        RECT 92.400 75.800 93.200 80.400 ;
        RECT 95.600 75.800 96.400 80.400 ;
        RECT 102.000 75.800 102.800 80.400 ;
        RECT 105.200 75.800 106.000 80.400 ;
        RECT 113.200 75.800 114.000 80.400 ;
        RECT 116.400 75.800 117.200 80.400 ;
        RECT 119.600 75.800 120.400 80.400 ;
        RECT 122.800 75.800 123.600 80.400 ;
        RECT 126.000 75.800 126.800 80.400 ;
        RECT 129.200 75.800 130.000 80.400 ;
        RECT 132.400 75.800 133.200 80.400 ;
        RECT 138.800 75.800 139.600 80.400 ;
        RECT 142.000 75.800 142.800 80.400 ;
        RECT 150.000 75.800 150.800 80.400 ;
        RECT 153.200 75.800 154.000 80.400 ;
        RECT 156.400 75.800 157.200 80.400 ;
        RECT 159.600 75.800 160.400 80.400 ;
        RECT 161.200 75.800 162.000 80.400 ;
        RECT 164.400 75.800 165.200 80.400 ;
        RECT 167.600 75.800 168.400 80.400 ;
        RECT 174.000 75.800 174.800 80.400 ;
        RECT 177.200 75.800 178.000 80.400 ;
        RECT 185.200 75.800 186.000 80.400 ;
        RECT 188.400 75.800 189.200 80.400 ;
        RECT 191.600 75.800 192.400 80.400 ;
        RECT 194.800 75.800 195.600 80.400 ;
        RECT 198.000 75.800 198.800 80.400 ;
        RECT 202.800 73.000 203.600 80.400 ;
        RECT 92.400 71.800 93.200 72.400 ;
        RECT 95.600 71.800 96.600 72.000 ;
        RECT 129.200 71.800 130.000 72.400 ;
        RECT 132.600 71.800 133.400 72.000 ;
        RECT 164.400 71.800 165.200 72.400 ;
        RECT 167.600 71.800 168.600 72.000 ;
        RECT 207.600 71.800 208.400 80.400 ;
        RECT 214.000 73.000 214.800 80.400 ;
        RECT 218.800 73.000 219.600 80.400 ;
        RECT 15.000 71.200 42.000 71.800 ;
        RECT 92.400 71.200 119.400 71.800 ;
        RECT 129.200 71.200 156.200 71.800 ;
        RECT 164.400 71.200 191.400 71.800 ;
        RECT 15.000 71.000 15.800 71.200 ;
        RECT 118.600 71.000 119.400 71.200 ;
        RECT 155.400 71.000 156.200 71.200 ;
        RECT 190.600 71.000 191.400 71.200 ;
        RECT 10.200 50.800 11.000 51.000 ;
        RECT 69.400 50.800 70.200 51.000 ;
        RECT 131.800 50.800 132.600 51.000 ;
        RECT 216.200 50.800 217.000 51.000 ;
        RECT 10.200 50.200 37.200 50.800 ;
        RECT 69.400 50.200 96.400 50.800 ;
        RECT 131.800 50.200 158.800 50.800 ;
        RECT 190.000 50.200 217.000 50.800 ;
        RECT 33.000 50.000 34.000 50.200 ;
        RECT 36.400 49.600 37.200 50.200 ;
        RECT 92.200 50.000 93.200 50.200 ;
        RECT 95.600 49.600 96.400 50.200 ;
        RECT 2.800 41.600 3.600 49.000 ;
        RECT 6.000 41.600 6.800 46.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 12.400 41.600 13.200 46.200 ;
        RECT 15.600 41.600 16.400 46.200 ;
        RECT 23.600 41.600 24.400 46.200 ;
        RECT 26.800 41.600 27.600 46.200 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 42.800 41.600 43.600 46.200 ;
        RECT 49.200 41.600 50.000 49.000 ;
        RECT 54.000 41.600 54.800 46.200 ;
        RECT 55.600 41.600 56.400 46.200 ;
        RECT 58.800 41.600 59.600 45.800 ;
        RECT 63.600 41.600 64.400 46.200 ;
        RECT 65.200 41.600 66.000 46.200 ;
        RECT 68.400 41.600 69.200 46.200 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 74.800 41.600 75.600 46.200 ;
        RECT 82.800 41.600 83.600 46.200 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 92.400 41.600 93.200 46.200 ;
        RECT 95.600 41.600 96.400 46.200 ;
        RECT 98.800 41.600 99.600 46.200 ;
        RECT 102.000 41.600 102.800 46.200 ;
        RECT 105.200 41.600 106.000 50.200 ;
        RECT 108.400 41.600 109.200 50.200 ;
        RECT 111.600 41.600 112.400 50.200 ;
        RECT 114.800 41.600 115.600 50.200 ;
        RECT 118.000 41.600 118.800 50.200 ;
        RECT 154.600 50.000 155.600 50.200 ;
        RECT 158.000 49.600 158.800 50.200 ;
        RECT 121.200 41.600 122.000 45.800 ;
        RECT 124.400 41.600 125.200 46.200 ;
        RECT 127.600 41.600 128.400 46.200 ;
        RECT 130.800 41.600 131.600 46.200 ;
        RECT 134.000 41.600 134.800 46.200 ;
        RECT 137.200 41.600 138.000 46.200 ;
        RECT 145.200 41.600 146.000 46.200 ;
        RECT 148.400 41.600 149.200 46.200 ;
        RECT 154.800 41.600 155.600 46.200 ;
        RECT 158.000 41.600 158.800 46.200 ;
        RECT 161.200 41.600 162.000 46.200 ;
        RECT 162.800 41.600 163.600 46.200 ;
        RECT 167.600 41.600 168.400 49.000 ;
        RECT 173.000 41.600 173.800 46.200 ;
        RECT 177.200 41.600 178.000 50.200 ;
        RECT 178.800 41.600 179.600 50.200 ;
        RECT 190.000 49.600 190.800 50.200 ;
        RECT 193.400 50.000 194.200 50.200 ;
        RECT 183.000 41.600 183.800 46.200 ;
        RECT 186.800 41.600 187.600 46.200 ;
        RECT 190.000 41.600 190.800 46.200 ;
        RECT 193.200 41.600 194.000 46.200 ;
        RECT 199.600 41.600 200.400 46.200 ;
        RECT 202.800 41.600 203.600 46.200 ;
        RECT 210.800 41.600 211.600 46.200 ;
        RECT 214.000 41.600 214.800 46.200 ;
        RECT 217.200 41.600 218.000 46.200 ;
        RECT 220.400 41.600 221.200 46.200 ;
        RECT 222.000 41.600 222.800 46.200 ;
        RECT 0.400 40.400 226.800 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 4.400 35.800 5.200 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 10.800 35.800 11.600 40.400 ;
        RECT 18.800 35.800 19.600 40.400 ;
        RECT 22.000 35.600 22.800 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 39.600 32.200 40.400 40.400 ;
        RECT 42.800 35.800 43.600 40.400 ;
        RECT 44.400 35.800 45.200 40.400 ;
        RECT 47.600 31.800 48.400 40.400 ;
        RECT 51.800 35.800 52.600 40.400 ;
        RECT 54.000 35.800 54.800 40.400 ;
        RECT 57.200 35.800 58.000 40.400 ;
        RECT 60.400 35.800 61.200 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 71.600 35.800 72.400 40.400 ;
        RECT 74.800 35.800 75.600 40.400 ;
        RECT 81.200 35.800 82.000 40.400 ;
        RECT 84.400 35.800 85.200 40.400 ;
        RECT 87.600 35.800 88.400 40.400 ;
        RECT 81.000 31.800 82.000 32.000 ;
        RECT 84.400 31.800 85.200 32.400 ;
        RECT 90.800 31.800 91.600 40.400 ;
        RECT 94.000 33.000 94.800 40.400 ;
        RECT 98.800 33.000 99.600 40.400 ;
        RECT 102.000 31.800 102.800 40.400 ;
        RECT 103.600 31.800 104.400 40.400 ;
        RECT 106.800 31.800 107.600 40.400 ;
        RECT 110.000 31.800 110.800 40.400 ;
        RECT 111.600 35.800 112.400 40.400 ;
        RECT 114.800 35.800 115.600 40.400 ;
        RECT 118.000 35.800 118.800 40.400 ;
        RECT 124.400 35.800 125.200 40.400 ;
        RECT 127.600 35.800 128.400 40.400 ;
        RECT 135.600 35.800 136.400 40.400 ;
        RECT 138.800 35.800 139.600 40.400 ;
        RECT 142.000 35.800 142.800 40.400 ;
        RECT 145.200 35.800 146.000 40.400 ;
        RECT 148.400 35.800 149.200 40.400 ;
        RECT 114.800 31.800 115.600 32.400 ;
        RECT 118.200 31.800 119.000 32.000 ;
        RECT 152.800 31.800 153.600 40.400 ;
        RECT 158.000 32.200 158.800 40.400 ;
        RECT 161.200 35.800 162.000 40.400 ;
        RECT 164.400 35.800 165.200 40.400 ;
        RECT 167.600 35.800 168.400 40.400 ;
        RECT 170.800 35.800 171.600 40.400 ;
        RECT 178.800 35.800 179.600 40.400 ;
        RECT 182.000 35.800 182.800 40.400 ;
        RECT 188.400 35.800 189.200 40.400 ;
        RECT 191.600 35.800 192.400 40.400 ;
        RECT 194.800 35.800 195.600 40.400 ;
        RECT 201.200 33.000 202.000 40.400 ;
        RECT 206.000 35.800 206.800 40.400 ;
        RECT 188.200 31.800 189.000 32.000 ;
        RECT 191.600 31.800 192.400 32.400 ;
        RECT 209.200 32.200 210.000 40.400 ;
        RECT 214.400 31.800 215.200 40.400 ;
        RECT 218.800 35.800 219.600 40.400 ;
        RECT 222.000 33.000 222.800 40.400 ;
        RECT 58.200 31.200 85.200 31.800 ;
        RECT 114.800 31.200 141.800 31.800 ;
        RECT 58.200 31.000 59.000 31.200 ;
        RECT 141.000 31.000 141.800 31.200 ;
        RECT 165.400 31.200 192.400 31.800 ;
        RECT 165.400 31.000 166.200 31.200 ;
        RECT 10.800 30.000 34.200 30.600 ;
        RECT 10.800 29.400 11.600 30.000 ;
        RECT 22.000 29.600 22.800 30.000 ;
        RECT 28.400 29.600 29.200 30.000 ;
        RECT 33.400 29.800 34.200 30.000 ;
        RECT 5.400 10.800 6.200 11.000 ;
        RECT 50.200 10.800 51.000 11.000 ;
        RECT 126.600 10.800 127.400 11.000 ;
        RECT 213.000 10.800 213.800 11.000 ;
        RECT 5.400 10.200 32.400 10.800 ;
        RECT 50.200 10.200 77.200 10.800 ;
        RECT 100.400 10.200 127.400 10.800 ;
        RECT 186.800 10.200 213.800 10.800 ;
        RECT 28.200 10.000 29.200 10.200 ;
        RECT 31.600 9.600 32.400 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 10.800 1.600 11.600 6.200 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 22.000 1.600 22.800 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 38.000 1.600 38.800 10.200 ;
        RECT 73.000 10.000 74.000 10.200 ;
        RECT 76.400 9.600 77.200 10.200 ;
        RECT 44.400 1.600 45.200 6.200 ;
        RECT 46.000 1.600 46.800 6.200 ;
        RECT 49.200 1.600 50.000 6.200 ;
        RECT 52.400 1.600 53.200 6.200 ;
        RECT 55.600 1.600 56.400 6.200 ;
        RECT 63.600 1.600 64.400 6.200 ;
        RECT 66.800 1.600 67.600 6.200 ;
        RECT 73.200 1.600 74.000 6.200 ;
        RECT 76.400 1.600 77.200 6.200 ;
        RECT 79.600 1.600 80.400 6.200 ;
        RECT 82.800 1.600 83.600 10.200 ;
        RECT 86.000 1.600 86.800 10.200 ;
        RECT 89.200 1.600 90.000 10.200 ;
        RECT 92.400 1.600 93.200 10.200 ;
        RECT 95.600 1.600 96.400 10.200 ;
        RECT 100.400 9.600 101.200 10.200 ;
        RECT 103.600 10.000 104.600 10.200 ;
        RECT 97.200 1.600 98.000 6.200 ;
        RECT 100.400 1.600 101.200 6.200 ;
        RECT 103.600 1.600 104.400 6.200 ;
        RECT 110.000 1.600 110.800 6.200 ;
        RECT 113.200 1.600 114.000 6.200 ;
        RECT 121.200 1.600 122.000 6.200 ;
        RECT 124.400 1.600 125.200 6.200 ;
        RECT 127.600 1.600 128.400 6.200 ;
        RECT 130.800 1.600 131.600 6.200 ;
        RECT 134.000 1.600 134.800 9.000 ;
        RECT 138.800 1.600 139.600 6.200 ;
        RECT 143.200 1.600 144.000 10.200 ;
        RECT 148.400 1.600 149.200 9.800 ;
        RECT 153.200 1.600 154.000 9.000 ;
        RECT 158.000 1.600 158.800 6.200 ;
        RECT 161.200 1.600 162.000 9.000 ;
        RECT 166.000 1.600 166.800 9.000 ;
        RECT 172.400 1.600 173.200 9.000 ;
        RECT 176.200 1.600 177.000 6.200 ;
        RECT 180.400 1.600 181.200 10.200 ;
        RECT 186.800 9.600 187.600 10.200 ;
        RECT 190.200 10.000 191.000 10.200 ;
        RECT 183.600 1.600 184.400 6.200 ;
        RECT 186.800 1.600 187.600 6.200 ;
        RECT 190.000 1.600 190.800 6.200 ;
        RECT 196.400 1.600 197.200 6.200 ;
        RECT 199.600 1.600 200.400 6.200 ;
        RECT 207.600 1.600 208.400 6.200 ;
        RECT 210.800 1.600 211.600 6.200 ;
        RECT 214.000 1.600 214.800 6.200 ;
        RECT 217.200 1.600 218.000 6.200 ;
        RECT 220.400 1.600 221.200 9.000 ;
        RECT 0.400 0.400 226.800 1.600 ;
      LAYER via1 ;
        RECT 41.200 200.600 42.000 201.400 ;
        RECT 134.000 200.600 134.800 201.400 ;
        RECT 145.200 197.600 146.000 198.400 ;
        RECT 145.200 191.600 146.000 192.400 ;
        RECT 167.600 191.200 168.400 192.000 ;
        RECT 44.400 163.600 45.200 164.400 ;
        RECT 130.800 163.600 131.600 164.400 ;
        RECT 194.800 163.600 195.600 164.400 ;
        RECT 41.200 160.600 42.000 161.400 ;
        RECT 134.000 160.600 134.800 161.400 ;
        RECT 20.400 157.600 21.200 158.400 ;
        RECT 20.400 151.600 21.200 152.400 ;
        RECT 79.600 151.200 80.400 152.000 ;
        RECT 127.600 157.600 128.400 158.400 ;
        RECT 127.600 151.600 128.400 152.400 ;
        RECT 191.600 151.200 192.400 152.000 ;
        RECT 98.800 123.600 99.600 124.400 ;
        RECT 212.400 123.600 213.200 124.400 ;
        RECT 41.200 120.600 42.000 121.400 ;
        RECT 134.000 120.600 134.800 121.400 ;
        RECT 36.400 117.600 37.200 118.400 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 183.600 117.600 184.400 118.400 ;
        RECT 143.600 111.200 144.400 112.000 ;
        RECT 183.600 111.600 184.400 112.400 ;
        RECT 129.200 90.000 130.000 90.800 ;
        RECT 90.800 83.600 91.600 84.400 ;
        RECT 129.200 85.400 130.000 86.200 ;
        RECT 188.400 85.400 189.200 86.200 ;
        RECT 41.200 80.600 42.000 81.400 ;
        RECT 134.000 80.600 134.800 81.400 ;
        RECT 41.200 77.600 42.000 78.400 ;
        RECT 41.200 71.600 42.000 72.400 ;
        RECT 129.200 77.600 130.000 78.400 ;
        RECT 95.600 71.200 96.400 72.000 ;
        RECT 129.200 71.600 130.000 72.400 ;
        RECT 167.600 71.200 168.400 72.000 ;
        RECT 33.200 50.000 34.000 50.800 ;
        RECT 92.400 50.000 93.200 50.800 ;
        RECT 33.200 43.600 34.000 44.400 ;
        RECT 92.400 43.600 93.200 44.400 ;
        RECT 154.800 50.000 155.600 50.800 ;
        RECT 154.800 45.400 155.600 46.200 ;
        RECT 190.000 43.600 190.800 44.400 ;
        RECT 41.200 40.600 42.000 41.400 ;
        RECT 134.000 40.600 134.800 41.400 ;
        RECT 81.200 31.200 82.000 32.000 ;
        RECT 114.800 37.600 115.600 38.400 ;
        RECT 114.800 31.600 115.600 32.400 ;
        RECT 191.600 37.600 192.400 38.400 ;
        RECT 191.600 31.600 192.400 32.400 ;
        RECT 28.400 10.000 29.200 10.800 ;
        RECT 28.400 3.600 29.200 4.400 ;
        RECT 73.200 10.000 74.000 10.800 ;
        RECT 73.200 5.400 74.000 6.200 ;
        RECT 103.600 5.400 104.400 6.200 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 41.200 0.600 42.000 1.400 ;
        RECT 134.000 0.600 134.800 1.400 ;
      LAYER metal2 ;
        RECT 40.800 200.600 42.400 201.400 ;
        RECT 133.600 200.600 135.200 201.400 ;
        RECT 145.200 197.600 146.000 198.400 ;
        RECT 145.300 192.400 145.900 197.600 ;
        RECT 167.600 195.800 168.400 196.600 ;
        RECT 145.200 191.600 146.000 192.400 ;
        RECT 167.700 192.000 168.300 195.800 ;
        RECT 167.600 191.200 168.400 192.000 ;
        RECT 44.400 169.600 45.200 170.400 ;
        RECT 130.800 169.600 131.600 170.400 ;
        RECT 194.800 169.600 195.600 170.400 ;
        RECT 44.500 164.400 45.100 169.600 ;
        RECT 130.900 164.400 131.500 169.600 ;
        RECT 194.900 164.400 195.500 169.600 ;
        RECT 44.400 163.600 45.200 164.400 ;
        RECT 130.800 163.600 131.600 164.400 ;
        RECT 194.800 163.600 195.600 164.400 ;
        RECT 40.800 160.600 42.400 161.400 ;
        RECT 133.600 160.600 135.200 161.400 ;
        RECT 20.400 157.600 21.200 158.400 ;
        RECT 127.600 157.600 128.400 158.400 ;
        RECT 20.500 152.400 21.100 157.600 ;
        RECT 79.600 155.800 80.400 156.600 ;
        RECT 20.400 151.600 21.200 152.400 ;
        RECT 79.700 152.000 80.300 155.800 ;
        RECT 127.700 152.400 128.300 157.600 ;
        RECT 191.600 155.800 192.400 156.600 ;
        RECT 79.600 151.200 80.400 152.000 ;
        RECT 127.600 151.600 128.400 152.400 ;
        RECT 191.700 152.000 192.300 155.800 ;
        RECT 191.600 151.200 192.400 152.000 ;
        RECT 98.800 129.600 99.600 130.400 ;
        RECT 212.400 129.600 213.200 130.400 ;
        RECT 98.900 124.400 99.500 129.600 ;
        RECT 212.500 124.400 213.100 129.600 ;
        RECT 98.800 123.600 99.600 124.400 ;
        RECT 212.400 123.600 213.200 124.400 ;
        RECT 40.800 120.600 42.400 121.400 ;
        RECT 133.600 120.600 135.200 121.400 ;
        RECT 36.400 117.600 37.200 118.400 ;
        RECT 183.600 117.600 184.400 118.400 ;
        RECT 36.500 112.400 37.100 117.600 ;
        RECT 143.600 115.800 144.400 116.600 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 143.700 112.000 144.300 115.800 ;
        RECT 183.700 112.400 184.300 117.600 ;
        RECT 143.600 111.200 144.400 112.000 ;
        RECT 183.600 111.600 184.400 112.400 ;
        RECT 90.800 89.600 91.600 90.400 ;
        RECT 129.200 90.000 130.000 90.800 ;
        RECT 188.400 90.000 189.200 90.800 ;
        RECT 90.900 84.400 91.500 89.600 ;
        RECT 129.300 86.200 129.900 90.000 ;
        RECT 188.500 86.200 189.100 90.000 ;
        RECT 129.200 85.400 130.000 86.200 ;
        RECT 188.400 85.400 189.200 86.200 ;
        RECT 90.800 83.600 91.600 84.400 ;
        RECT 40.800 80.600 42.400 81.400 ;
        RECT 133.600 80.600 135.200 81.400 ;
        RECT 41.200 77.600 42.000 78.400 ;
        RECT 129.200 77.600 130.000 78.400 ;
        RECT 41.300 72.400 41.900 77.600 ;
        RECT 95.600 75.800 96.400 76.600 ;
        RECT 41.200 71.600 42.000 72.400 ;
        RECT 95.700 72.000 96.300 75.800 ;
        RECT 129.300 72.400 129.900 77.600 ;
        RECT 167.600 75.800 168.400 76.600 ;
        RECT 95.600 71.200 96.400 72.000 ;
        RECT 129.200 71.600 130.000 72.400 ;
        RECT 167.700 72.000 168.300 75.800 ;
        RECT 167.600 71.200 168.400 72.000 ;
        RECT 33.200 50.000 34.000 50.800 ;
        RECT 92.400 50.000 93.200 50.800 ;
        RECT 154.800 50.000 155.600 50.800 ;
        RECT 33.300 44.400 33.900 50.000 ;
        RECT 92.500 44.400 93.100 50.000 ;
        RECT 154.900 46.200 155.500 50.000 ;
        RECT 190.000 49.600 190.800 50.400 ;
        RECT 154.800 45.400 155.600 46.200 ;
        RECT 190.100 44.400 190.700 49.600 ;
        RECT 33.200 43.600 34.000 44.400 ;
        RECT 92.400 43.600 93.200 44.400 ;
        RECT 190.000 43.600 190.800 44.400 ;
        RECT 40.800 40.600 42.400 41.400 ;
        RECT 133.600 40.600 135.200 41.400 ;
        RECT 114.800 37.600 115.600 38.400 ;
        RECT 191.600 37.600 192.400 38.400 ;
        RECT 22.000 35.600 22.800 36.400 ;
        RECT 81.200 35.800 82.000 36.600 ;
        RECT 22.100 30.400 22.700 35.600 ;
        RECT 81.300 32.000 81.900 35.800 ;
        RECT 114.900 32.400 115.500 37.600 ;
        RECT 191.700 32.400 192.300 37.600 ;
        RECT 81.200 31.200 82.000 32.000 ;
        RECT 114.800 31.600 115.600 32.400 ;
        RECT 191.600 31.600 192.400 32.400 ;
        RECT 22.000 29.600 22.800 30.400 ;
        RECT 28.400 10.000 29.200 10.800 ;
        RECT 73.200 10.000 74.000 10.800 ;
        RECT 103.600 10.000 104.400 10.800 ;
        RECT 28.500 4.400 29.100 10.000 ;
        RECT 73.300 6.200 73.900 10.000 ;
        RECT 103.700 6.200 104.300 10.000 ;
        RECT 186.800 9.600 187.600 10.400 ;
        RECT 73.200 5.400 74.000 6.200 ;
        RECT 103.600 5.400 104.400 6.200 ;
        RECT 186.900 4.400 187.500 9.600 ;
        RECT 28.400 3.600 29.200 4.400 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 40.800 0.600 42.400 1.400 ;
        RECT 133.600 0.600 135.200 1.400 ;
      LAYER via2 ;
        RECT 41.200 200.600 42.000 201.400 ;
        RECT 134.000 200.600 134.800 201.400 ;
        RECT 41.200 160.600 42.000 161.400 ;
        RECT 134.000 160.600 134.800 161.400 ;
        RECT 41.200 120.600 42.000 121.400 ;
        RECT 134.000 120.600 134.800 121.400 ;
        RECT 41.200 80.600 42.000 81.400 ;
        RECT 134.000 80.600 134.800 81.400 ;
        RECT 41.200 40.600 42.000 41.400 ;
        RECT 134.000 40.600 134.800 41.400 ;
        RECT 41.200 0.600 42.000 1.400 ;
        RECT 134.000 0.600 134.800 1.400 ;
      LAYER metal3 ;
        RECT 40.800 200.400 42.400 201.600 ;
        RECT 133.600 200.400 135.200 201.600 ;
        RECT 40.800 160.400 42.400 161.600 ;
        RECT 133.600 160.400 135.200 161.600 ;
        RECT 40.800 120.400 42.400 121.600 ;
        RECT 133.600 120.400 135.200 121.600 ;
        RECT 40.800 80.400 42.400 81.600 ;
        RECT 133.600 80.400 135.200 81.600 ;
        RECT 40.800 40.400 42.400 41.600 ;
        RECT 133.600 40.400 135.200 41.600 ;
        RECT 40.800 0.400 42.400 1.600 ;
        RECT 133.600 0.400 135.200 1.600 ;
      LAYER via3 ;
        RECT 41.200 200.600 42.000 201.400 ;
        RECT 134.000 200.600 134.800 201.400 ;
        RECT 41.200 160.600 42.000 161.400 ;
        RECT 134.000 160.600 134.800 161.400 ;
        RECT 41.200 120.600 42.000 121.400 ;
        RECT 134.000 120.600 134.800 121.400 ;
        RECT 41.200 80.600 42.000 81.400 ;
        RECT 134.000 80.600 134.800 81.400 ;
        RECT 41.200 40.600 42.000 41.400 ;
        RECT 134.000 40.600 134.800 41.400 ;
        RECT 41.200 0.600 42.000 1.400 ;
        RECT 134.000 0.600 134.800 1.400 ;
      LAYER metal4 ;
        RECT 40.800 -4.000 42.400 204.000 ;
        RECT 133.600 -4.000 135.200 204.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.800 181.600 3.600 185.400 ;
        RECT 7.600 181.600 8.400 184.200 ;
        RECT 10.800 181.600 11.600 184.200 ;
        RECT 15.600 181.600 16.400 186.200 ;
        RECT 17.200 181.600 18.000 184.200 ;
        RECT 20.400 181.600 21.200 184.200 ;
        RECT 24.600 181.600 25.400 186.200 ;
        RECT 31.600 181.600 32.400 188.200 ;
        RECT 33.200 181.600 34.000 186.200 ;
        RECT 39.600 181.600 40.400 184.200 ;
        RECT 42.800 181.600 43.600 184.200 ;
        RECT 47.600 181.600 48.400 185.400 ;
        RECT 50.800 181.600 51.600 186.200 ;
        RECT 54.600 181.600 55.400 186.200 ;
        RECT 58.800 181.600 59.600 184.200 ;
        RECT 63.600 181.600 64.400 186.200 ;
        RECT 65.200 181.600 66.000 184.200 ;
        RECT 68.400 181.600 69.200 184.200 ;
        RECT 71.600 181.600 72.400 185.400 ;
        RECT 78.000 181.600 78.800 186.200 ;
        RECT 81.200 181.600 82.000 186.200 ;
        RECT 90.800 181.600 91.600 185.400 ;
        RECT 95.600 181.600 96.400 184.200 ;
        RECT 97.200 181.600 98.000 184.200 ;
        RECT 100.400 181.600 101.200 184.200 ;
        RECT 105.200 181.600 106.000 186.200 ;
        RECT 108.400 181.600 109.200 184.200 ;
        RECT 111.600 181.600 112.400 186.200 ;
        RECT 114.800 181.600 115.600 184.200 ;
        RECT 121.200 181.600 122.000 186.200 ;
        RECT 132.400 181.600 133.200 184.200 ;
        RECT 135.600 181.600 136.400 184.200 ;
        RECT 145.200 181.600 146.000 186.200 ;
        RECT 153.200 181.600 154.000 186.200 ;
        RECT 158.000 181.600 158.800 186.200 ;
        RECT 164.400 181.600 165.200 186.200 ;
        RECT 174.000 181.600 174.800 184.200 ;
        RECT 177.200 181.600 178.000 184.200 ;
        RECT 188.400 181.600 189.200 186.200 ;
        RECT 194.800 181.600 195.600 184.200 ;
        RECT 199.600 181.600 200.400 186.200 ;
        RECT 202.800 181.600 203.600 184.200 ;
        RECT 207.000 181.600 207.800 186.200 ;
        RECT 209.200 181.600 210.000 184.200 ;
        RECT 212.400 181.600 213.200 184.200 ;
        RECT 215.600 181.600 216.400 184.200 ;
        RECT 218.800 181.600 219.600 186.200 ;
        RECT 0.400 180.400 226.800 181.600 ;
        RECT 2.800 176.600 3.600 180.400 ;
        RECT 9.200 176.600 10.000 180.400 ;
        RECT 14.000 177.800 14.800 180.400 ;
        RECT 20.400 175.800 21.200 180.400 ;
        RECT 31.600 177.800 32.400 180.400 ;
        RECT 34.800 177.800 35.600 180.400 ;
        RECT 44.400 175.800 45.200 180.400 ;
        RECT 55.600 173.800 56.400 180.400 ;
        RECT 58.800 176.600 59.600 180.400 ;
        RECT 66.800 176.600 67.600 180.400 ;
        RECT 73.200 176.600 74.000 180.400 ;
        RECT 78.000 176.400 79.000 180.400 ;
        RECT 84.200 179.800 85.000 180.400 ;
        RECT 84.200 176.400 85.200 179.800 ;
        RECT 89.200 177.800 90.000 180.400 ;
        RECT 94.000 176.600 94.800 180.400 ;
        RECT 102.000 176.600 102.800 180.400 ;
        RECT 105.200 177.800 106.000 180.400 ;
        RECT 108.400 177.800 109.200 180.400 ;
        RECT 112.200 176.000 113.000 180.400 ;
        RECT 116.400 177.800 117.200 180.400 ;
        RECT 119.600 177.800 120.400 180.400 ;
        RECT 122.800 175.800 123.600 180.400 ;
        RECT 130.800 175.800 131.600 180.400 ;
        RECT 140.400 177.800 141.200 180.400 ;
        RECT 143.600 177.800 144.400 180.400 ;
        RECT 154.800 175.800 155.600 180.400 ;
        RECT 161.200 177.800 162.000 180.400 ;
        RECT 162.800 177.800 163.600 180.400 ;
        RECT 167.000 175.800 167.800 180.400 ;
        RECT 169.200 177.800 170.000 180.400 ;
        RECT 174.000 175.400 174.800 180.400 ;
        RECT 179.200 175.000 180.000 180.400 ;
        RECT 183.600 175.800 184.400 180.400 ;
        RECT 188.400 177.800 189.200 180.400 ;
        RECT 194.800 175.800 195.600 180.400 ;
        RECT 204.400 177.800 205.200 180.400 ;
        RECT 207.600 177.800 208.400 180.400 ;
        RECT 218.800 175.800 219.600 180.400 ;
        RECT 225.200 177.800 226.000 180.400 ;
        RECT 2.800 141.600 3.600 146.200 ;
        RECT 6.000 141.600 6.800 144.200 ;
        RECT 9.200 141.600 10.000 144.200 ;
        RECT 12.400 141.600 13.200 145.400 ;
        RECT 20.400 141.600 21.200 146.200 ;
        RECT 30.000 141.600 30.800 144.200 ;
        RECT 33.200 141.600 34.000 144.200 ;
        RECT 44.400 141.600 45.200 146.200 ;
        RECT 50.800 141.600 51.600 144.200 ;
        RECT 57.200 141.600 58.000 145.400 ;
        RECT 62.600 141.600 63.400 146.000 ;
        RECT 66.800 141.600 67.600 144.200 ;
        RECT 70.000 141.600 70.800 144.200 ;
        RECT 76.400 141.600 77.200 146.200 ;
        RECT 86.000 141.600 86.800 144.200 ;
        RECT 89.200 141.600 90.000 144.200 ;
        RECT 100.400 141.600 101.200 146.200 ;
        RECT 106.800 141.600 107.600 144.200 ;
        RECT 108.400 141.600 109.200 146.200 ;
        RECT 111.600 141.600 112.400 146.200 ;
        RECT 114.800 141.600 115.600 146.200 ;
        RECT 118.000 141.600 118.800 146.200 ;
        RECT 121.200 141.600 122.000 146.200 ;
        RECT 127.600 141.600 128.400 146.200 ;
        RECT 137.200 141.600 138.000 144.200 ;
        RECT 140.400 141.600 141.200 144.200 ;
        RECT 151.600 141.600 152.400 146.200 ;
        RECT 158.000 141.600 158.800 144.200 ;
        RECT 161.200 142.200 162.200 145.600 ;
        RECT 161.400 141.600 162.200 142.200 ;
        RECT 167.400 141.600 168.400 145.600 ;
        RECT 172.400 141.600 173.200 146.600 ;
        RECT 177.600 141.600 178.400 147.000 ;
        RECT 182.000 141.600 182.800 144.200 ;
        RECT 188.400 141.600 189.200 146.200 ;
        RECT 198.000 141.600 198.800 144.200 ;
        RECT 201.200 141.600 202.000 144.200 ;
        RECT 212.400 141.600 213.200 146.200 ;
        RECT 218.800 141.600 219.600 144.200 ;
        RECT 222.000 141.600 222.800 146.200 ;
        RECT 0.400 140.400 226.800 141.600 ;
        RECT 4.400 136.600 5.200 140.400 ;
        RECT 7.600 137.800 8.400 140.400 ;
        RECT 11.400 135.800 12.200 140.400 ;
        RECT 15.600 137.800 16.400 140.400 ;
        RECT 17.200 135.800 18.000 140.400 ;
        RECT 23.200 135.800 24.000 140.400 ;
        RECT 26.800 137.800 27.600 140.400 ;
        RECT 30.000 138.200 30.800 140.400 ;
        RECT 39.600 137.800 40.400 140.400 ;
        RECT 42.800 137.800 43.600 140.400 ;
        RECT 46.000 137.800 46.800 140.400 ;
        RECT 47.600 133.800 48.400 140.400 ;
        RECT 54.000 133.800 54.800 140.400 ;
        RECT 62.000 137.800 62.800 140.400 ;
        RECT 65.200 135.800 66.000 140.400 ;
        RECT 68.400 137.800 69.200 140.400 ;
        RECT 74.800 135.800 75.600 140.400 ;
        RECT 86.000 137.800 86.800 140.400 ;
        RECT 89.200 137.800 90.000 140.400 ;
        RECT 98.800 135.800 99.600 140.400 ;
        RECT 105.200 135.800 106.000 140.400 ;
        RECT 108.400 135.800 109.200 140.400 ;
        RECT 111.600 135.800 112.400 140.400 ;
        RECT 114.800 135.800 115.600 140.400 ;
        RECT 118.000 135.800 118.800 140.400 ;
        RECT 119.600 135.800 120.400 140.400 ;
        RECT 122.800 135.800 123.600 140.400 ;
        RECT 126.000 135.800 126.800 140.400 ;
        RECT 129.200 135.800 130.000 140.400 ;
        RECT 132.400 135.800 133.200 140.400 ;
        RECT 135.600 135.800 136.400 140.400 ;
        RECT 138.800 135.800 139.600 140.400 ;
        RECT 142.600 135.800 143.400 140.400 ;
        RECT 146.800 137.800 147.600 140.400 ;
        RECT 150.000 137.800 150.800 140.400 ;
        RECT 154.800 136.600 155.600 140.400 ;
        RECT 159.600 136.600 160.400 140.400 ;
        RECT 167.600 136.600 168.400 140.400 ;
        RECT 170.800 137.800 171.600 140.400 ;
        RECT 175.000 135.800 175.800 140.400 ;
        RECT 178.800 137.800 179.600 140.400 ;
        RECT 182.000 137.800 182.800 140.400 ;
        RECT 188.400 135.800 189.200 140.400 ;
        RECT 199.600 137.800 200.400 140.400 ;
        RECT 202.800 137.800 203.600 140.400 ;
        RECT 212.400 135.800 213.200 140.400 ;
        RECT 218.800 135.800 219.600 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 6.000 101.600 6.800 104.200 ;
        RECT 12.400 101.600 13.200 106.200 ;
        RECT 23.600 101.600 24.400 104.200 ;
        RECT 26.800 101.600 27.600 104.200 ;
        RECT 36.400 101.600 37.200 106.200 ;
        RECT 42.800 101.600 43.600 104.200 ;
        RECT 46.000 101.600 46.800 106.200 ;
        RECT 52.000 101.600 52.800 106.200 ;
        RECT 54.000 101.600 54.800 104.200 ;
        RECT 57.200 101.600 58.000 104.200 ;
        RECT 62.000 101.600 62.800 106.200 ;
        RECT 68.400 101.600 69.200 108.200 ;
        RECT 70.000 101.600 70.800 108.200 ;
        RECT 76.400 101.600 77.200 106.200 ;
        RECT 79.600 101.600 80.400 106.200 ;
        RECT 81.200 101.600 82.000 106.200 ;
        RECT 84.400 101.600 85.200 106.200 ;
        RECT 89.200 101.600 90.000 106.200 ;
        RECT 92.400 101.600 93.200 106.200 ;
        RECT 95.600 101.600 96.400 106.200 ;
        RECT 97.200 101.600 98.000 106.200 ;
        RECT 100.400 101.600 101.200 106.200 ;
        RECT 103.600 101.600 104.400 104.200 ;
        RECT 108.400 101.600 109.200 106.200 ;
        RECT 111.600 101.600 112.400 106.200 ;
        RECT 114.400 101.600 115.200 107.000 ;
        RECT 119.600 101.600 120.400 106.600 ;
        RECT 124.400 101.600 125.200 106.200 ;
        RECT 127.600 101.600 128.400 106.200 ;
        RECT 130.800 101.600 131.600 106.200 ;
        RECT 134.000 101.600 134.800 106.200 ;
        RECT 140.400 101.600 141.200 106.200 ;
        RECT 150.000 101.600 150.800 104.200 ;
        RECT 153.200 101.600 154.000 104.200 ;
        RECT 164.400 101.600 165.200 106.200 ;
        RECT 170.800 101.600 171.600 104.200 ;
        RECT 172.400 101.600 173.200 104.200 ;
        RECT 176.600 101.600 177.400 106.200 ;
        RECT 183.600 101.600 184.400 106.200 ;
        RECT 193.200 101.600 194.000 104.200 ;
        RECT 196.400 101.600 197.200 104.200 ;
        RECT 207.600 101.600 208.400 106.200 ;
        RECT 214.000 101.600 214.800 104.200 ;
        RECT 217.200 101.600 218.000 104.200 ;
        RECT 220.400 101.600 221.200 106.200 ;
        RECT 0.400 100.400 226.800 101.600 ;
        RECT 1.200 97.800 2.000 100.400 ;
        RECT 7.600 96.600 8.400 100.400 ;
        RECT 10.800 93.800 11.600 100.400 ;
        RECT 22.000 93.800 22.800 100.400 ;
        RECT 25.200 97.800 26.000 100.400 ;
        RECT 28.400 97.800 29.200 100.400 ;
        RECT 31.600 96.600 32.400 100.400 ;
        RECT 38.000 97.800 38.800 100.400 ;
        RECT 42.800 96.600 43.600 100.400 ;
        RECT 50.800 96.600 51.600 100.400 ;
        RECT 56.600 96.000 57.400 100.400 ;
        RECT 60.400 97.800 61.200 100.400 ;
        RECT 66.800 95.800 67.600 100.400 ;
        RECT 78.000 97.800 78.800 100.400 ;
        RECT 81.200 97.800 82.000 100.400 ;
        RECT 90.800 95.800 91.600 100.400 ;
        RECT 98.800 95.800 99.600 100.400 ;
        RECT 102.000 97.800 102.800 100.400 ;
        RECT 108.400 95.800 109.200 100.400 ;
        RECT 119.600 97.800 120.400 100.400 ;
        RECT 122.800 97.800 123.600 100.400 ;
        RECT 132.400 95.800 133.200 100.400 ;
        RECT 142.000 96.600 142.800 100.400 ;
        RECT 145.200 97.800 146.000 100.400 ;
        RECT 149.400 95.800 150.200 100.400 ;
        RECT 151.600 97.800 152.400 100.400 ;
        RECT 154.800 97.800 155.600 100.400 ;
        RECT 158.000 96.400 159.000 100.400 ;
        RECT 164.200 99.800 165.000 100.400 ;
        RECT 164.200 96.400 165.200 99.800 ;
        RECT 169.200 96.600 170.000 100.400 ;
        RECT 175.600 96.600 176.400 100.400 ;
        RECT 185.200 95.800 186.000 100.400 ;
        RECT 194.800 97.800 195.600 100.400 ;
        RECT 198.000 97.800 198.800 100.400 ;
        RECT 209.200 95.800 210.000 100.400 ;
        RECT 215.600 97.800 216.400 100.400 ;
        RECT 218.800 95.400 219.600 100.400 ;
        RECT 224.000 95.000 224.800 100.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 7.600 61.600 8.400 66.200 ;
        RECT 10.800 61.600 11.600 64.200 ;
        RECT 17.200 61.600 18.000 66.200 ;
        RECT 28.400 61.600 29.200 64.200 ;
        RECT 31.600 61.600 32.400 64.200 ;
        RECT 41.200 61.600 42.000 66.200 ;
        RECT 47.600 61.600 48.400 64.200 ;
        RECT 55.600 61.600 56.400 68.200 ;
        RECT 57.200 61.600 58.000 68.200 ;
        RECT 66.800 61.600 67.600 65.400 ;
        RECT 71.600 61.600 72.400 65.400 ;
        RECT 79.600 61.600 80.400 66.200 ;
        RECT 81.200 61.600 82.000 66.200 ;
        RECT 84.400 61.600 85.200 66.200 ;
        RECT 92.400 61.600 93.200 66.200 ;
        RECT 102.000 61.600 102.800 64.200 ;
        RECT 105.200 61.600 106.000 64.200 ;
        RECT 116.400 61.600 117.200 66.200 ;
        RECT 122.800 61.600 123.600 64.200 ;
        RECT 129.200 61.600 130.000 66.200 ;
        RECT 138.800 61.600 139.600 64.200 ;
        RECT 142.000 61.600 142.800 64.200 ;
        RECT 153.200 61.600 154.000 66.200 ;
        RECT 159.600 61.600 160.400 64.200 ;
        RECT 164.400 61.600 165.200 66.200 ;
        RECT 174.000 61.600 174.800 64.200 ;
        RECT 177.200 61.600 178.000 64.200 ;
        RECT 188.400 61.600 189.200 66.200 ;
        RECT 194.800 61.600 195.600 64.200 ;
        RECT 198.000 61.600 198.800 64.200 ;
        RECT 201.800 61.600 202.600 66.200 ;
        RECT 206.000 61.600 206.800 64.200 ;
        RECT 207.600 61.600 208.400 64.200 ;
        RECT 210.800 61.600 211.600 64.200 ;
        RECT 214.000 61.600 214.800 66.200 ;
        RECT 218.800 61.600 219.600 66.200 ;
        RECT 0.400 60.400 226.800 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 6.000 57.800 6.800 60.400 ;
        RECT 12.400 55.800 13.200 60.400 ;
        RECT 23.600 57.800 24.400 60.400 ;
        RECT 26.800 57.800 27.600 60.400 ;
        RECT 36.400 55.800 37.200 60.400 ;
        RECT 42.800 57.800 43.600 60.400 ;
        RECT 46.000 57.800 46.800 60.400 ;
        RECT 50.200 55.800 51.000 60.400 ;
        RECT 54.000 57.800 54.800 60.400 ;
        RECT 55.600 53.800 56.400 60.400 ;
        RECT 63.600 57.800 64.400 60.400 ;
        RECT 65.200 57.800 66.000 60.400 ;
        RECT 71.600 55.800 72.400 60.400 ;
        RECT 82.800 57.800 83.600 60.400 ;
        RECT 86.000 57.800 86.800 60.400 ;
        RECT 95.600 55.800 96.400 60.400 ;
        RECT 102.000 57.800 102.800 60.400 ;
        RECT 105.200 55.800 106.000 60.400 ;
        RECT 108.400 55.800 109.200 60.400 ;
        RECT 111.600 55.800 112.400 60.400 ;
        RECT 114.800 55.800 115.600 60.400 ;
        RECT 118.000 55.800 118.800 60.400 ;
        RECT 124.400 53.800 125.200 60.400 ;
        RECT 127.600 57.800 128.400 60.400 ;
        RECT 134.000 55.800 134.800 60.400 ;
        RECT 145.200 57.800 146.000 60.400 ;
        RECT 148.400 57.800 149.200 60.400 ;
        RECT 158.000 55.800 158.800 60.400 ;
        RECT 162.800 57.800 163.600 60.400 ;
        RECT 166.600 55.800 167.400 60.400 ;
        RECT 170.800 57.800 171.600 60.400 ;
        RECT 175.600 56.600 176.400 60.400 ;
        RECT 180.400 56.600 181.200 60.400 ;
        RECT 190.000 55.800 190.800 60.400 ;
        RECT 199.600 57.800 200.400 60.400 ;
        RECT 202.800 57.800 203.600 60.400 ;
        RECT 214.000 55.800 214.800 60.400 ;
        RECT 220.400 57.800 221.200 60.400 ;
        RECT 222.000 57.800 222.800 60.400 ;
        RECT 1.200 21.600 2.000 24.200 ;
        RECT 7.600 21.600 8.400 26.200 ;
        RECT 18.800 21.600 19.600 24.200 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 31.600 21.600 32.400 26.200 ;
        RECT 40.200 21.600 41.000 26.000 ;
        RECT 44.400 21.600 45.200 24.200 ;
        RECT 49.200 21.600 50.000 25.400 ;
        RECT 54.000 21.600 54.800 24.200 ;
        RECT 60.400 21.600 61.200 26.200 ;
        RECT 71.600 21.600 72.400 24.200 ;
        RECT 74.800 21.600 75.600 24.200 ;
        RECT 84.400 21.600 85.200 26.200 ;
        RECT 90.800 21.600 91.600 26.200 ;
        RECT 94.000 21.600 94.800 26.200 ;
        RECT 98.800 21.600 99.600 26.200 ;
        RECT 102.000 21.600 102.800 26.200 ;
        RECT 103.600 21.600 104.400 26.200 ;
        RECT 106.800 21.600 107.600 26.200 ;
        RECT 110.000 21.600 110.800 26.200 ;
        RECT 114.800 21.600 115.600 26.200 ;
        RECT 124.400 21.600 125.200 24.200 ;
        RECT 127.600 21.600 128.400 24.200 ;
        RECT 138.800 21.600 139.600 26.200 ;
        RECT 145.200 21.600 146.000 24.200 ;
        RECT 148.400 21.600 149.200 24.200 ;
        RECT 152.800 21.600 153.600 27.000 ;
        RECT 158.000 21.600 158.800 26.600 ;
        RECT 161.200 21.600 162.000 24.200 ;
        RECT 167.600 21.600 168.400 26.200 ;
        RECT 178.800 21.600 179.600 24.200 ;
        RECT 182.000 21.600 182.800 24.200 ;
        RECT 191.600 21.600 192.400 26.200 ;
        RECT 198.000 21.600 198.800 24.200 ;
        RECT 202.200 21.600 203.000 26.200 ;
        RECT 206.000 21.600 206.800 24.200 ;
        RECT 209.200 21.600 210.000 26.600 ;
        RECT 214.400 21.600 215.200 27.000 ;
        RECT 218.800 21.600 219.600 24.200 ;
        RECT 222.000 21.600 222.800 26.200 ;
        RECT 0.400 20.400 226.800 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 22.000 17.800 22.800 20.400 ;
        RECT 31.600 15.800 32.400 20.400 ;
        RECT 38.000 17.800 38.800 20.400 ;
        RECT 41.200 17.800 42.000 20.400 ;
        RECT 44.400 17.800 45.200 20.400 ;
        RECT 46.000 17.800 46.800 20.400 ;
        RECT 52.400 15.800 53.200 20.400 ;
        RECT 63.600 17.800 64.400 20.400 ;
        RECT 66.800 17.800 67.600 20.400 ;
        RECT 76.400 15.800 77.200 20.400 ;
        RECT 82.800 15.800 83.600 20.400 ;
        RECT 86.000 15.800 86.800 20.400 ;
        RECT 89.200 15.800 90.000 20.400 ;
        RECT 92.400 15.800 93.200 20.400 ;
        RECT 95.600 15.800 96.400 20.400 ;
        RECT 100.400 15.800 101.200 20.400 ;
        RECT 110.000 17.800 110.800 20.400 ;
        RECT 113.200 17.800 114.000 20.400 ;
        RECT 124.400 15.800 125.200 20.400 ;
        RECT 130.800 17.800 131.600 20.400 ;
        RECT 134.000 15.800 134.800 20.400 ;
        RECT 138.800 17.800 139.600 20.400 ;
        RECT 143.200 15.000 144.000 20.400 ;
        RECT 148.400 15.400 149.200 20.400 ;
        RECT 153.200 15.800 154.000 20.400 ;
        RECT 158.000 17.800 158.800 20.400 ;
        RECT 161.200 15.800 162.000 20.400 ;
        RECT 165.000 15.800 165.800 20.400 ;
        RECT 169.200 17.800 170.000 20.400 ;
        RECT 172.400 15.800 173.200 20.400 ;
        RECT 178.800 16.600 179.600 20.400 ;
        RECT 186.800 15.800 187.600 20.400 ;
        RECT 196.400 17.800 197.200 20.400 ;
        RECT 199.600 17.800 200.400 20.400 ;
        RECT 210.800 15.800 211.600 20.400 ;
        RECT 217.200 17.800 218.000 20.400 ;
        RECT 220.400 15.800 221.200 20.400 ;
      LAYER via1 ;
        RECT 87.600 180.600 88.400 181.400 ;
        RECT 186.800 180.600 187.600 181.400 ;
        RECT 87.600 140.600 88.400 141.400 ;
        RECT 186.800 140.600 187.600 141.400 ;
        RECT 87.600 100.600 88.400 101.400 ;
        RECT 186.800 100.600 187.600 101.400 ;
        RECT 87.600 60.600 88.400 61.400 ;
        RECT 186.800 60.600 187.600 61.400 ;
        RECT 87.600 20.600 88.400 21.400 ;
        RECT 186.800 20.600 187.600 21.400 ;
      LAYER metal2 ;
        RECT 87.200 180.600 88.800 181.400 ;
        RECT 186.400 180.600 188.000 181.400 ;
        RECT 87.200 140.600 88.800 141.400 ;
        RECT 186.400 140.600 188.000 141.400 ;
        RECT 87.200 100.600 88.800 101.400 ;
        RECT 186.400 100.600 188.000 101.400 ;
        RECT 87.200 60.600 88.800 61.400 ;
        RECT 186.400 60.600 188.000 61.400 ;
        RECT 87.200 20.600 88.800 21.400 ;
        RECT 186.400 20.600 188.000 21.400 ;
      LAYER via2 ;
        RECT 87.600 180.600 88.400 181.400 ;
        RECT 186.800 180.600 187.600 181.400 ;
        RECT 87.600 140.600 88.400 141.400 ;
        RECT 186.800 140.600 187.600 141.400 ;
        RECT 87.600 100.600 88.400 101.400 ;
        RECT 186.800 100.600 187.600 101.400 ;
        RECT 87.600 60.600 88.400 61.400 ;
        RECT 186.800 60.600 187.600 61.400 ;
        RECT 87.600 20.600 88.400 21.400 ;
        RECT 186.800 20.600 187.600 21.400 ;
      LAYER metal3 ;
        RECT 87.200 180.400 88.800 181.600 ;
        RECT 186.400 180.400 188.000 181.600 ;
        RECT 87.200 140.400 88.800 141.600 ;
        RECT 186.400 140.400 188.000 141.600 ;
        RECT 87.200 100.400 88.800 101.600 ;
        RECT 186.400 100.400 188.000 101.600 ;
        RECT 87.200 60.400 88.800 61.600 ;
        RECT 186.400 60.400 188.000 61.600 ;
        RECT 87.200 20.400 88.800 21.600 ;
        RECT 186.400 20.400 188.000 21.600 ;
      LAYER via3 ;
        RECT 87.600 180.600 88.400 181.400 ;
        RECT 186.800 180.600 187.600 181.400 ;
        RECT 87.600 140.600 88.400 141.400 ;
        RECT 186.800 140.600 187.600 141.400 ;
        RECT 87.600 100.600 88.400 101.400 ;
        RECT 186.800 100.600 187.600 101.400 ;
        RECT 87.600 60.600 88.400 61.400 ;
        RECT 186.800 60.600 187.600 61.400 ;
        RECT 87.600 20.600 88.400 21.400 ;
        RECT 186.800 20.600 187.600 21.400 ;
      LAYER metal4 ;
        RECT 87.200 -4.000 88.800 204.000 ;
        RECT 186.400 -4.000 188.000 204.000 ;
    END
  END gnd
  PIN clock
    PORT
      LAYER metal1 ;
        RECT 108.400 148.200 110.200 149.000 ;
        RECT 108.400 147.600 109.200 148.200 ;
        RECT 118.000 134.300 118.800 134.400 ;
        RECT 119.600 134.300 120.400 134.400 ;
        RECT 118.000 133.800 120.400 134.300 ;
        RECT 117.000 133.700 121.400 133.800 ;
        RECT 117.000 133.000 118.800 133.700 ;
        RECT 119.600 133.000 121.400 133.700 ;
        RECT 105.200 53.800 106.000 54.400 ;
        RECT 105.200 53.000 107.000 53.800 ;
        RECT 95.600 13.800 96.400 14.400 ;
        RECT 94.600 13.000 96.400 13.800 ;
      LAYER via1 ;
        RECT 118.000 133.600 118.800 134.400 ;
        RECT 105.200 53.600 106.000 54.400 ;
        RECT 95.600 13.600 96.400 14.400 ;
      LAYER metal2 ;
        RECT 108.400 147.600 109.200 148.400 ;
        RECT 108.500 144.400 109.100 147.600 ;
        RECT 108.400 143.600 109.200 144.400 ;
        RECT 118.000 143.600 118.800 144.400 ;
        RECT 118.100 134.400 118.700 143.600 ;
        RECT 118.000 133.600 118.800 134.400 ;
        RECT 118.100 106.400 118.700 133.600 ;
        RECT 118.000 105.600 118.800 106.400 ;
        RECT 105.200 61.600 106.000 62.400 ;
        RECT 105.300 54.400 105.900 61.600 ;
        RECT 105.200 54.300 106.000 54.400 ;
        RECT 103.700 53.700 106.000 54.300 ;
        RECT 103.700 16.400 104.300 53.700 ;
        RECT 105.200 53.600 106.000 53.700 ;
        RECT 95.600 15.600 96.400 16.400 ;
        RECT 103.600 15.600 104.400 16.400 ;
        RECT 95.700 14.400 96.300 15.600 ;
        RECT 95.600 13.600 96.400 14.400 ;
        RECT 95.700 -1.700 96.300 13.600 ;
        RECT 94.100 -2.300 96.300 -1.700 ;
      LAYER metal3 ;
        RECT 108.400 144.300 109.200 144.400 ;
        RECT 118.000 144.300 118.800 144.400 ;
        RECT 108.400 143.700 118.800 144.300 ;
        RECT 108.400 143.600 109.200 143.700 ;
        RECT 118.000 143.600 118.800 143.700 ;
        RECT 113.200 106.300 114.000 106.400 ;
        RECT 118.000 106.300 118.800 106.400 ;
        RECT 113.200 105.700 118.800 106.300 ;
        RECT 113.200 105.600 114.000 105.700 ;
        RECT 118.000 105.600 118.800 105.700 ;
        RECT 105.200 62.300 106.000 62.400 ;
        RECT 113.200 62.300 114.000 62.400 ;
        RECT 105.200 61.700 114.000 62.300 ;
        RECT 105.200 61.600 106.000 61.700 ;
        RECT 113.200 61.600 114.000 61.700 ;
        RECT 95.600 16.300 96.400 16.400 ;
        RECT 103.600 16.300 104.400 16.400 ;
        RECT 95.600 15.700 104.400 16.300 ;
        RECT 95.600 15.600 96.400 15.700 ;
        RECT 103.600 15.600 104.400 15.700 ;
      LAYER metal4 ;
        RECT 113.000 61.400 114.200 106.600 ;
    END
  END clock
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 102.000 28.300 102.800 28.400 ;
        RECT 103.600 28.300 104.400 28.400 ;
        RECT 102.000 27.700 104.400 28.300 ;
        RECT 102.000 27.600 102.800 27.700 ;
        RECT 103.600 26.800 104.400 27.700 ;
      LAYER metal2 ;
        RECT 102.000 27.600 102.800 28.400 ;
        RECT 102.100 2.400 102.700 27.600 ;
        RECT 102.000 1.600 102.800 2.400 ;
        RECT 106.800 1.600 107.600 2.400 ;
        RECT 106.900 -2.300 107.500 1.600 ;
      LAYER metal3 ;
        RECT 102.000 2.300 102.800 2.400 ;
        RECT 106.800 2.300 107.600 2.400 ;
        RECT 102.000 1.700 107.600 2.300 ;
        RECT 102.000 1.600 102.800 1.700 ;
        RECT 106.800 1.600 107.600 1.700 ;
    END
  END reset
  PIN start
    PORT
      LAYER metal1 ;
        RECT 66.800 13.600 67.600 15.200 ;
      LAYER metal2 ;
        RECT 66.800 13.600 67.600 14.400 ;
        RECT 66.900 2.400 67.500 13.600 ;
        RECT 62.000 1.600 62.800 2.400 ;
        RECT 66.800 1.600 67.600 2.400 ;
        RECT 62.100 -2.300 62.700 1.600 ;
      LAYER metal3 ;
        RECT 62.000 2.300 62.800 2.400 ;
        RECT 66.800 2.300 67.600 2.400 ;
        RECT 62.000 1.700 67.600 2.300 ;
        RECT 62.000 1.600 62.800 1.700 ;
        RECT 66.800 1.600 67.600 1.700 ;
    END
  END start
  PIN N[0]
    PORT
      LAYER metal1 ;
        RECT 212.400 184.800 213.200 186.400 ;
      LAYER via1 ;
        RECT 212.400 185.600 213.200 186.400 ;
      LAYER metal2 ;
        RECT 210.900 188.300 211.500 204.300 ;
        RECT 210.900 187.700 213.100 188.300 ;
        RECT 212.500 186.400 213.100 187.700 ;
        RECT 212.400 185.600 213.200 186.400 ;
    END
  END N[0]
  PIN N[1]
    PORT
      LAYER metal1 ;
        RECT 63.600 188.300 64.400 188.400 ;
        RECT 63.600 187.700 65.900 188.300 ;
        RECT 63.600 186.800 64.400 187.700 ;
        RECT 65.300 186.400 65.900 187.700 ;
        RECT 65.200 184.800 66.000 186.400 ;
        RECT 87.600 176.300 88.400 176.400 ;
        RECT 89.200 176.300 90.000 177.200 ;
        RECT 87.600 175.700 90.000 176.300 ;
        RECT 87.600 175.600 88.400 175.700 ;
        RECT 89.200 175.600 90.000 175.700 ;
      LAYER via1 ;
        RECT 65.200 185.600 66.000 186.400 ;
      LAYER metal2 ;
        RECT 65.300 186.400 65.900 204.300 ;
        RECT 65.200 185.600 66.000 186.400 ;
        RECT 65.300 176.400 65.900 185.600 ;
        RECT 65.200 175.600 66.000 176.400 ;
        RECT 87.600 175.600 88.400 176.400 ;
      LAYER metal3 ;
        RECT 65.200 176.300 66.000 176.400 ;
        RECT 87.600 176.300 88.400 176.400 ;
        RECT 65.200 175.700 88.400 176.300 ;
        RECT 65.200 175.600 66.000 175.700 ;
        RECT 87.600 175.600 88.400 175.700 ;
    END
  END N[1]
  PIN N[2]
    PORT
      LAYER metal1 ;
        RECT 60.400 191.600 61.200 193.200 ;
        RECT 68.400 189.600 69.200 191.200 ;
      LAYER metal2 ;
        RECT 60.400 191.600 61.200 192.400 ;
        RECT 60.500 190.300 61.100 191.600 ;
        RECT 62.100 190.400 62.700 204.300 ;
        RECT 62.000 190.300 62.800 190.400 ;
        RECT 60.500 189.700 62.800 190.300 ;
        RECT 62.000 189.600 62.800 189.700 ;
        RECT 68.400 189.600 69.200 190.400 ;
      LAYER metal3 ;
        RECT 62.000 190.300 62.800 190.400 ;
        RECT 68.400 190.300 69.200 190.400 ;
        RECT 62.000 189.700 69.200 190.300 ;
        RECT 62.000 189.600 62.800 189.700 ;
        RECT 68.400 189.600 69.200 189.700 ;
    END
  END N[2]
  PIN N[3]
    PORT
      LAYER metal1 ;
        RECT 49.200 188.200 50.000 188.400 ;
        RECT 48.400 187.600 50.000 188.200 ;
        RECT 55.600 187.600 56.400 189.200 ;
        RECT 48.400 187.200 49.200 187.600 ;
        RECT 42.800 184.800 43.600 186.400 ;
        RECT 58.000 174.400 58.800 174.800 ;
        RECT 57.200 173.800 58.800 174.400 ;
        RECT 57.200 173.600 58.000 173.800 ;
      LAYER via1 ;
        RECT 49.200 187.600 50.000 188.400 ;
        RECT 42.800 185.600 43.600 186.400 ;
      LAYER metal2 ;
        RECT 55.700 188.400 56.300 204.300 ;
        RECT 42.800 187.600 43.600 188.400 ;
        RECT 49.200 187.600 50.000 188.400 ;
        RECT 55.600 187.600 56.400 188.400 ;
        RECT 42.900 186.400 43.500 187.600 ;
        RECT 42.800 185.600 43.600 186.400 ;
        RECT 55.700 176.300 56.300 187.600 ;
        RECT 55.700 175.700 57.900 176.300 ;
        RECT 57.300 174.400 57.900 175.700 ;
        RECT 57.200 173.600 58.000 174.400 ;
      LAYER metal3 ;
        RECT 42.800 188.300 43.600 188.400 ;
        RECT 49.200 188.300 50.000 188.400 ;
        RECT 55.600 188.300 56.400 188.400 ;
        RECT 42.800 187.700 56.400 188.300 ;
        RECT 42.800 187.600 43.600 187.700 ;
        RECT 49.200 187.600 50.000 187.700 ;
        RECT 55.600 187.600 56.400 187.700 ;
    END
  END N[3]
  PIN N[4]
    PORT
      LAYER metal1 ;
        RECT 44.400 193.600 46.000 194.400 ;
        RECT 45.200 192.400 45.800 193.600 ;
        RECT 44.400 191.800 45.800 192.400 ;
        RECT 44.400 191.600 45.200 191.800 ;
        RECT 39.600 189.600 40.400 191.200 ;
      LAYER metal2 ;
        RECT 44.500 194.400 45.100 204.300 ;
        RECT 44.400 193.600 45.200 194.400 ;
        RECT 44.500 190.400 45.100 193.600 ;
        RECT 39.600 189.600 40.400 190.400 ;
        RECT 44.400 189.600 45.200 190.400 ;
      LAYER metal3 ;
        RECT 39.600 190.300 40.400 190.400 ;
        RECT 44.400 190.300 45.200 190.400 ;
        RECT 39.600 189.700 45.200 190.300 ;
        RECT 39.600 189.600 40.400 189.700 ;
        RECT 44.400 189.600 45.200 189.700 ;
    END
  END N[4]
  PIN N[5]
    PORT
      LAYER metal1 ;
        RECT 1.200 188.200 2.000 188.400 ;
        RECT 1.200 187.600 2.800 188.200 ;
        RECT 2.000 187.200 2.800 187.600 ;
        RECT 10.800 184.800 11.600 186.400 ;
        RECT 17.200 184.800 18.000 186.400 ;
        RECT 2.000 174.400 2.800 174.800 ;
        RECT 1.200 173.800 2.800 174.400 ;
        RECT 1.200 173.600 2.000 173.800 ;
      LAYER via1 ;
        RECT 10.800 185.600 11.600 186.400 ;
        RECT 17.200 185.600 18.000 186.400 ;
      LAYER metal2 ;
        RECT 1.200 187.600 2.000 188.400 ;
        RECT 1.300 174.400 1.900 187.600 ;
        RECT 10.800 185.600 11.600 186.400 ;
        RECT 17.200 185.600 18.000 186.400 ;
        RECT 1.200 173.600 2.000 174.400 ;
      LAYER metal3 ;
        RECT 1.200 188.300 2.000 188.400 ;
        RECT -1.900 187.700 11.500 188.300 ;
        RECT 1.200 187.600 2.000 187.700 ;
        RECT 10.900 186.400 11.500 187.700 ;
        RECT 10.800 186.300 11.600 186.400 ;
        RECT 17.200 186.300 18.000 186.400 ;
        RECT 10.800 185.700 18.000 186.300 ;
        RECT 10.800 185.600 11.600 185.700 ;
        RECT 17.200 185.600 18.000 185.700 ;
    END
  END N[5]
  PIN N[6]
    PORT
      LAYER metal1 ;
        RECT 5.200 193.600 6.000 194.400 ;
        RECT 5.400 192.400 6.000 193.600 ;
        RECT 5.400 191.800 6.800 192.400 ;
        RECT 6.000 191.600 6.800 191.800 ;
        RECT 6.100 190.300 6.700 191.600 ;
        RECT 7.600 190.300 8.400 191.200 ;
        RECT 6.100 189.700 8.400 190.300 ;
        RECT 7.600 189.600 8.400 189.700 ;
      LAYER metal2 ;
        RECT 6.000 191.600 6.800 192.400 ;
      LAYER metal3 ;
        RECT 6.000 192.300 6.800 192.400 ;
        RECT -1.900 191.700 6.800 192.300 ;
        RECT 6.000 191.600 6.800 191.700 ;
    END
  END N[6]
  PIN N[7]
    PORT
      LAYER metal1 ;
        RECT 28.400 95.600 29.200 97.200 ;
        RECT 8.400 94.400 9.200 94.800 ;
        RECT 28.500 94.400 29.100 95.600 ;
        RECT 30.800 94.400 31.600 94.800 ;
        RECT 8.400 93.800 10.000 94.400 ;
        RECT 9.200 93.600 10.000 93.800 ;
        RECT 28.400 94.300 29.200 94.400 ;
        RECT 30.000 94.300 31.600 94.400 ;
        RECT 28.400 93.800 31.600 94.300 ;
        RECT 28.400 93.700 30.800 93.800 ;
        RECT 28.400 93.600 29.200 93.700 ;
        RECT 30.000 93.600 30.800 93.700 ;
      LAYER metal2 ;
        RECT 9.200 93.600 10.000 94.400 ;
        RECT 28.400 93.600 29.200 94.400 ;
        RECT 9.300 90.400 9.900 93.600 ;
        RECT 28.500 90.400 29.100 93.600 ;
        RECT 9.200 89.600 10.000 90.400 ;
        RECT 28.400 89.600 29.200 90.400 ;
      LAYER metal3 ;
        RECT 9.200 90.300 10.000 90.400 ;
        RECT 28.400 90.300 29.200 90.400 ;
        RECT -1.900 89.700 29.200 90.300 ;
        RECT 9.200 89.600 10.000 89.700 ;
        RECT 28.400 89.600 29.200 89.700 ;
    END
  END N[7]
  PIN N[8]
    PORT
      LAYER metal1 ;
        RECT 1.200 95.600 2.000 97.200 ;
        RECT 19.600 91.600 21.200 92.400 ;
      LAYER via1 ;
        RECT 20.400 91.600 21.200 92.400 ;
      LAYER metal2 ;
        RECT 1.200 95.600 2.000 96.400 ;
        RECT 1.300 94.400 1.900 95.600 ;
        RECT 1.200 93.600 2.000 94.400 ;
        RECT 20.400 93.600 21.200 94.400 ;
        RECT 20.500 92.400 21.100 93.600 ;
        RECT 20.400 91.600 21.200 92.400 ;
      LAYER metal3 ;
        RECT 1.200 94.300 2.000 94.400 ;
        RECT 20.400 94.300 21.200 94.400 ;
        RECT -1.900 93.700 21.200 94.300 ;
        RECT 1.200 93.600 2.000 93.700 ;
        RECT 20.400 93.600 21.200 93.700 ;
    END
  END N[8]
  PIN dp[0]
    PORT
      LAYER metal1 ;
        RECT 220.400 191.800 221.200 199.800 ;
        RECT 220.600 189.600 221.200 191.800 ;
        RECT 220.400 188.300 221.200 189.600 ;
        RECT 225.200 188.300 226.000 188.400 ;
        RECT 220.400 187.700 226.000 188.300 ;
        RECT 220.400 182.200 221.200 187.700 ;
        RECT 225.200 187.600 226.000 187.700 ;
      LAYER metal2 ;
        RECT 225.200 189.600 226.000 190.400 ;
        RECT 225.300 188.400 225.900 189.600 ;
        RECT 225.200 187.600 226.000 188.400 ;
      LAYER metal3 ;
        RECT 225.200 190.300 226.000 190.400 ;
        RECT 225.200 189.700 229.100 190.300 ;
        RECT 225.200 189.600 226.000 189.700 ;
    END
  END dp[0]
  PIN dp[1]
    PORT
      LAYER metal1 ;
        RECT 215.600 71.800 216.400 79.800 ;
        RECT 215.800 69.600 216.400 71.800 ;
        RECT 215.600 62.200 216.400 69.600 ;
      LAYER via1 ;
        RECT 215.600 67.600 216.400 68.400 ;
      LAYER metal2 ;
        RECT 215.600 69.600 216.400 70.400 ;
        RECT 215.700 68.400 216.300 69.600 ;
        RECT 215.600 67.600 216.400 68.400 ;
      LAYER metal3 ;
        RECT 215.600 70.300 216.400 70.400 ;
        RECT 215.600 69.700 229.100 70.300 ;
        RECT 215.600 69.600 216.400 69.700 ;
    END
  END dp[1]
  PIN dp[2]
    PORT
      LAYER metal1 ;
        RECT 154.800 12.400 155.600 19.800 ;
        RECT 155.000 10.200 155.600 12.400 ;
        RECT 154.800 2.200 155.600 10.200 ;
      LAYER via1 ;
        RECT 154.800 3.600 155.600 4.400 ;
      LAYER metal2 ;
        RECT 154.800 3.600 155.600 4.400 ;
        RECT 154.900 -1.700 155.500 3.600 ;
        RECT 153.300 -2.300 155.500 -1.700 ;
    END
  END dp[2]
  PIN dp[3]
    PORT
      LAYER metal1 ;
        RECT 223.600 31.800 224.400 39.800 ;
        RECT 223.800 29.600 224.400 31.800 ;
        RECT 223.600 28.300 224.400 29.600 ;
        RECT 225.200 28.300 226.000 28.400 ;
        RECT 223.600 27.700 226.000 28.300 ;
        RECT 223.600 22.200 224.400 27.700 ;
        RECT 225.200 27.600 226.000 27.700 ;
      LAYER metal2 ;
        RECT 225.200 29.600 226.000 30.400 ;
        RECT 225.300 28.400 225.900 29.600 ;
        RECT 225.200 27.600 226.000 28.400 ;
      LAYER metal3 ;
        RECT 225.200 30.300 226.000 30.400 ;
        RECT 225.200 29.700 229.100 30.300 ;
        RECT 225.200 29.600 226.000 29.700 ;
    END
  END dp[3]
  PIN dp[4]
    PORT
      LAYER metal1 ;
        RECT 135.600 12.400 136.400 19.800 ;
        RECT 135.800 10.200 136.400 12.400 ;
        RECT 135.600 4.300 136.400 10.200 ;
        RECT 137.200 4.300 138.000 4.400 ;
        RECT 135.600 3.700 138.000 4.300 ;
        RECT 135.600 2.200 136.400 3.700 ;
        RECT 137.200 3.600 138.000 3.700 ;
      LAYER metal2 ;
        RECT 137.200 3.600 138.000 4.400 ;
        RECT 137.300 -1.700 137.900 3.600 ;
        RECT 135.700 -2.300 137.900 -1.700 ;
    END
  END dp[4]
  PIN dp[5]
    PORT
      LAYER metal1 ;
        RECT 220.400 74.300 221.200 79.800 ;
        RECT 225.200 74.300 226.000 74.400 ;
        RECT 220.400 73.700 226.000 74.300 ;
        RECT 220.400 71.800 221.200 73.700 ;
        RECT 225.200 73.600 226.000 73.700 ;
        RECT 220.600 69.600 221.200 71.800 ;
        RECT 220.400 62.200 221.200 69.600 ;
      LAYER metal2 ;
        RECT 225.200 73.600 226.000 74.400 ;
      LAYER metal3 ;
        RECT 225.200 74.300 226.000 74.400 ;
        RECT 225.200 73.700 229.100 74.300 ;
        RECT 225.200 73.600 226.000 73.700 ;
    END
  END dp[5]
  PIN dp[6]
    PORT
      LAYER metal1 ;
        RECT 97.200 92.400 98.000 99.800 ;
        RECT 97.200 90.200 97.800 92.400 ;
        RECT 97.200 82.200 98.000 90.200 ;
      LAYER via1 ;
        RECT 97.200 83.600 98.000 84.400 ;
      LAYER metal2 ;
        RECT 97.200 83.600 98.000 84.400 ;
        RECT 97.300 82.400 97.900 83.600 ;
        RECT 97.200 81.600 98.000 82.400 ;
        RECT 98.800 3.600 99.600 4.400 ;
        RECT 98.900 -2.300 99.500 3.600 ;
      LAYER metal3 ;
        RECT 97.200 82.300 98.000 82.400 ;
        RECT 100.400 82.300 101.200 82.400 ;
        RECT 97.200 81.700 101.200 82.300 ;
        RECT 97.200 81.600 98.000 81.700 ;
        RECT 100.400 81.600 101.200 81.700 ;
        RECT 98.800 4.300 99.600 4.400 ;
        RECT 100.400 4.300 101.200 4.400 ;
        RECT 98.800 3.700 101.200 4.300 ;
        RECT 98.800 3.600 99.600 3.700 ;
        RECT 100.400 3.600 101.200 3.700 ;
      LAYER metal4 ;
        RECT 100.200 3.400 101.400 82.600 ;
    END
  END dp[6]
  PIN dp[7]
    PORT
      LAYER metal1 ;
        RECT 223.600 151.800 224.400 159.800 ;
        RECT 223.800 149.600 224.400 151.800 ;
        RECT 223.600 148.300 224.400 149.600 ;
        RECT 225.200 148.300 226.000 148.400 ;
        RECT 223.600 147.700 226.000 148.300 ;
        RECT 223.600 142.200 224.400 147.700 ;
        RECT 225.200 147.600 226.000 147.700 ;
      LAYER metal2 ;
        RECT 225.200 149.600 226.000 150.400 ;
        RECT 225.300 148.400 225.900 149.600 ;
        RECT 225.200 147.600 226.000 148.400 ;
      LAYER metal3 ;
        RECT 225.200 150.300 226.000 150.400 ;
        RECT 225.200 149.700 229.100 150.300 ;
        RECT 225.200 149.600 226.000 149.700 ;
    END
  END dp[7]
  PIN dp[8]
    PORT
      LAYER metal1 ;
        RECT 201.200 191.800 202.000 199.800 ;
        RECT 201.400 189.600 202.000 191.800 ;
        RECT 201.200 182.200 202.000 189.600 ;
      LAYER via1 ;
        RECT 201.200 197.600 202.000 198.400 ;
      LAYER metal2 ;
        RECT 199.700 203.700 201.900 204.300 ;
        RECT 201.300 198.400 201.900 203.700 ;
        RECT 201.200 197.600 202.000 198.400 ;
    END
  END dp[8]
  PIN done
    PORT
      LAYER metal1 ;
        RECT 1.200 52.400 2.000 59.800 ;
        RECT 1.200 50.200 1.800 52.400 ;
        RECT 1.200 42.200 2.000 50.200 ;
      LAYER via1 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal2 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 1.300 48.400 1.900 49.600 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal3 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -1.900 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
    END
  END done
  PIN counter[0]
    PORT
      LAYER metal1 ;
        RECT 124.400 172.400 125.200 179.800 ;
        RECT 124.600 170.200 125.200 172.400 ;
        RECT 124.400 162.200 125.200 170.200 ;
      LAYER via1 ;
        RECT 124.400 177.600 125.200 178.400 ;
      LAYER metal2 ;
        RECT 122.900 203.700 125.100 204.300 ;
        RECT 124.500 178.400 125.100 203.700 ;
        RECT 124.400 177.600 125.200 178.400 ;
    END
  END counter[0]
  PIN counter[1]
    PORT
      LAYER metal1 ;
        RECT 110.000 191.800 110.800 199.800 ;
        RECT 110.000 189.600 110.600 191.800 ;
        RECT 110.000 182.200 110.800 189.600 ;
      LAYER via1 ;
        RECT 110.000 197.600 110.800 198.400 ;
      LAYER metal2 ;
        RECT 110.100 203.700 112.300 204.300 ;
        RECT 110.100 198.400 110.700 203.700 ;
        RECT 110.000 197.600 110.800 198.400 ;
    END
  END counter[1]
  PIN counter[2]
    PORT
      LAYER metal1 ;
        RECT 76.400 191.800 77.200 199.800 ;
        RECT 76.400 189.600 77.000 191.800 ;
        RECT 76.400 182.200 77.200 189.600 ;
      LAYER via1 ;
        RECT 76.400 197.600 77.200 198.400 ;
      LAYER metal2 ;
        RECT 76.500 203.700 78.700 204.300 ;
        RECT 76.500 198.400 77.100 203.700 ;
        RECT 76.400 197.600 77.200 198.400 ;
    END
  END counter[2]
  PIN counter[3]
    PORT
      LAYER metal1 ;
        RECT 63.600 132.400 64.400 139.800 ;
        RECT 63.600 130.200 64.200 132.400 ;
        RECT 63.600 122.200 64.400 130.200 ;
      LAYER via1 ;
        RECT 63.600 137.600 64.400 138.400 ;
      LAYER metal2 ;
        RECT 63.600 139.600 64.400 140.400 ;
        RECT 63.700 138.400 64.300 139.600 ;
        RECT 63.600 137.600 64.400 138.400 ;
      LAYER metal3 ;
        RECT 1.200 140.300 2.000 140.400 ;
        RECT 63.600 140.300 64.400 140.400 ;
        RECT 1.200 139.700 64.400 140.300 ;
        RECT 1.200 139.600 2.000 139.700 ;
        RECT 63.600 139.600 64.400 139.700 ;
        RECT 1.200 130.300 2.000 130.400 ;
        RECT -1.900 129.700 2.000 130.300 ;
        RECT 1.200 129.600 2.000 129.700 ;
      LAYER metal4 ;
        RECT 1.000 129.400 2.200 140.600 ;
    END
  END counter[3]
  PIN counter[4]
    PORT
      LAYER metal1 ;
        RECT 1.200 151.800 2.000 159.800 ;
        RECT 1.200 149.600 1.800 151.800 ;
        RECT 1.200 142.200 2.000 149.600 ;
      LAYER via1 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal2 ;
        RECT 1.200 149.600 2.000 150.400 ;
        RECT 1.300 148.400 1.900 149.600 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal3 ;
        RECT 1.200 150.300 2.000 150.400 ;
        RECT -1.900 149.700 2.000 150.300 ;
        RECT 1.200 149.600 2.000 149.700 ;
    END
  END counter[4]
  PIN counter[5]
    PORT
      LAYER metal1 ;
        RECT 1.200 111.800 2.000 119.800 ;
        RECT 1.200 109.600 1.800 111.800 ;
        RECT 1.200 102.200 2.000 109.600 ;
      LAYER via1 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal2 ;
        RECT 1.200 109.600 2.000 110.400 ;
        RECT 1.300 108.400 1.900 109.600 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal3 ;
        RECT 1.200 110.300 2.000 110.400 ;
        RECT -1.900 109.700 2.000 110.300 ;
        RECT 1.200 109.600 2.000 109.700 ;
    END
  END counter[5]
  PIN counter[6]
    PORT
      LAYER metal1 ;
        RECT 1.200 71.800 2.000 79.800 ;
        RECT 1.200 69.600 1.800 71.800 ;
        RECT 1.200 62.200 2.000 69.600 ;
      LAYER via1 ;
        RECT 1.200 67.600 2.000 68.400 ;
      LAYER metal2 ;
        RECT 1.200 69.600 2.000 70.400 ;
        RECT 1.300 68.400 1.900 69.600 ;
        RECT 1.200 67.600 2.000 68.400 ;
      LAYER metal3 ;
        RECT 1.200 70.300 2.000 70.400 ;
        RECT -1.900 69.700 2.000 70.300 ;
        RECT 1.200 69.600 2.000 69.700 ;
    END
  END counter[6]
  PIN counter[7]
    PORT
      LAYER metal1 ;
        RECT 6.000 71.800 6.800 79.800 ;
        RECT 6.000 69.600 6.600 71.800 ;
        RECT 6.000 62.200 6.800 69.600 ;
      LAYER via1 ;
        RECT 6.000 73.600 6.800 74.400 ;
      LAYER metal2 ;
        RECT 6.000 73.600 6.800 74.400 ;
      LAYER metal3 ;
        RECT 6.000 74.300 6.800 74.400 ;
        RECT -1.900 73.700 6.800 74.300 ;
        RECT 6.000 73.600 6.800 73.700 ;
    END
  END counter[7]
  PIN sr[0]
    PORT
      LAYER metal1 ;
        RECT 222.000 111.800 222.800 119.800 ;
        RECT 222.200 109.600 222.800 111.800 ;
        RECT 222.000 108.300 222.800 109.600 ;
        RECT 225.200 108.300 226.000 108.400 ;
        RECT 222.000 107.700 226.000 108.300 ;
        RECT 222.000 102.200 222.800 107.700 ;
        RECT 225.200 107.600 226.000 107.700 ;
      LAYER metal2 ;
        RECT 225.200 109.600 226.000 110.400 ;
        RECT 225.300 108.400 225.900 109.600 ;
        RECT 225.200 107.600 226.000 108.400 ;
      LAYER metal3 ;
        RECT 225.200 110.300 226.000 110.400 ;
        RECT 225.200 109.700 229.100 110.300 ;
        RECT 225.200 109.600 226.000 109.700 ;
    END
  END sr[0]
  PIN sr[1]
    PORT
      LAYER metal1 ;
        RECT 174.000 12.400 174.800 19.800 ;
        RECT 174.200 10.200 174.800 12.400 ;
        RECT 174.000 2.200 174.800 10.200 ;
      LAYER via1 ;
        RECT 174.000 3.600 174.800 4.400 ;
      LAYER metal2 ;
        RECT 174.000 3.600 174.800 4.400 ;
        RECT 174.100 -1.700 174.700 3.600 ;
        RECT 172.500 -2.300 174.700 -1.700 ;
    END
  END sr[1]
  PIN sr[2]
    PORT
      LAYER metal1 ;
        RECT 222.000 12.400 222.800 19.800 ;
        RECT 222.200 10.200 222.800 12.400 ;
        RECT 222.000 8.300 222.800 10.200 ;
        RECT 225.200 8.300 226.000 8.400 ;
        RECT 222.000 7.700 226.000 8.300 ;
        RECT 222.000 2.200 222.800 7.700 ;
        RECT 225.200 7.600 226.000 7.700 ;
      LAYER metal2 ;
        RECT 225.200 9.600 226.000 10.400 ;
        RECT 225.300 8.400 225.900 9.600 ;
        RECT 225.200 7.600 226.000 8.400 ;
      LAYER metal3 ;
        RECT 225.200 10.300 226.000 10.400 ;
        RECT 225.200 9.700 229.100 10.300 ;
        RECT 225.200 9.600 226.000 9.700 ;
    END
  END sr[2]
  PIN sr[3]
    PORT
      LAYER metal1 ;
        RECT 162.800 12.400 163.600 19.800 ;
        RECT 163.000 10.200 163.600 12.400 ;
        RECT 162.800 2.200 163.600 10.200 ;
      LAYER via1 ;
        RECT 162.800 3.600 163.600 4.400 ;
      LAYER metal2 ;
        RECT 162.800 3.600 163.600 4.400 ;
        RECT 162.900 -1.700 163.500 3.600 ;
        RECT 161.300 -2.300 163.500 -1.700 ;
    END
  END sr[3]
  PIN sr[4]
    PORT
      LAYER metal1 ;
        RECT 220.400 132.400 221.200 139.800 ;
        RECT 220.600 130.200 221.200 132.400 ;
        RECT 220.400 128.300 221.200 130.200 ;
        RECT 225.200 128.300 226.000 128.400 ;
        RECT 220.400 127.700 226.000 128.300 ;
        RECT 220.400 122.200 221.200 127.700 ;
        RECT 225.200 127.600 226.000 127.700 ;
      LAYER metal2 ;
        RECT 225.200 129.600 226.000 130.400 ;
        RECT 225.300 128.400 225.900 129.600 ;
        RECT 225.200 127.600 226.000 128.400 ;
      LAYER metal3 ;
        RECT 225.200 130.300 226.000 130.400 ;
        RECT 225.200 129.700 229.100 130.300 ;
        RECT 225.200 129.600 226.000 129.700 ;
    END
  END sr[4]
  PIN sr[5]
    PORT
      LAYER metal1 ;
        RECT 154.800 191.800 155.600 199.800 ;
        RECT 155.000 189.600 155.600 191.800 ;
        RECT 154.800 182.200 155.600 189.600 ;
      LAYER via1 ;
        RECT 154.800 197.600 155.600 198.400 ;
      LAYER metal2 ;
        RECT 153.300 203.700 155.500 204.300 ;
        RECT 154.900 198.400 155.500 203.700 ;
        RECT 154.800 197.600 155.600 198.400 ;
    END
  END sr[5]
  PIN sr[6]
    PORT
      LAYER metal1 ;
        RECT 185.200 172.400 186.000 179.800 ;
        RECT 185.400 170.200 186.000 172.400 ;
        RECT 185.200 162.200 186.000 170.200 ;
      LAYER via1 ;
        RECT 185.200 177.600 186.000 178.400 ;
      LAYER metal2 ;
        RECT 183.700 200.400 184.300 204.300 ;
        RECT 183.600 199.600 184.400 200.400 ;
        RECT 185.200 177.600 186.000 178.400 ;
      LAYER metal3 ;
        RECT 183.600 199.600 184.400 200.400 ;
        RECT 183.600 178.300 184.400 178.400 ;
        RECT 185.200 178.300 186.000 178.400 ;
        RECT 183.600 177.700 186.000 178.300 ;
        RECT 183.600 177.600 184.400 177.700 ;
        RECT 185.200 177.600 186.000 177.700 ;
      LAYER metal4 ;
        RECT 183.400 177.400 184.600 200.600 ;
    END
  END sr[6]
  PIN sr[7]
    PORT
      LAYER metal1 ;
        RECT 156.400 191.800 157.200 199.800 ;
        RECT 156.400 189.600 157.000 191.800 ;
        RECT 156.400 182.200 157.200 189.600 ;
      LAYER via1 ;
        RECT 156.400 197.600 157.200 198.400 ;
      LAYER metal2 ;
        RECT 156.500 203.700 158.700 204.300 ;
        RECT 156.500 198.400 157.100 203.700 ;
        RECT 156.400 197.600 157.200 198.400 ;
    END
  END sr[7]
  OBS
      LAYER metal1 ;
        RECT 3.800 192.400 4.600 199.800 ;
        RECT 8.200 194.400 9.000 199.800 ;
        RECT 8.200 193.600 10.000 194.400 ;
        RECT 8.200 192.600 9.000 193.600 ;
        RECT 3.800 191.800 4.800 192.400 ;
        RECT 8.200 191.800 10.000 192.600 ;
        RECT 2.800 188.800 3.600 190.400 ;
        RECT 4.200 188.400 4.800 191.800 ;
        RECT 9.200 188.400 9.800 191.800 ;
        RECT 12.400 191.600 13.200 193.200 ;
        RECT 4.200 188.300 6.800 188.400 ;
        RECT 7.600 188.300 8.400 188.400 ;
        RECT 4.200 187.700 8.400 188.300 ;
        RECT 4.200 187.600 6.800 187.700 ;
        RECT 7.600 187.600 8.400 187.700 ;
        RECT 9.200 187.600 10.000 188.400 ;
        RECT 1.400 186.200 5.000 186.600 ;
        RECT 6.000 186.200 6.600 187.600 ;
        RECT 1.200 186.000 5.200 186.200 ;
        RECT 1.200 182.200 2.000 186.000 ;
        RECT 4.400 182.200 5.200 186.000 ;
        RECT 6.000 182.200 6.800 186.200 ;
        RECT 9.200 184.200 9.800 187.600 ;
        RECT 14.000 186.200 14.800 199.800 ;
        RECT 15.600 186.800 16.400 188.400 ;
        RECT 13.000 185.600 14.800 186.200 ;
        RECT 18.800 186.300 19.600 199.800 ;
        RECT 20.400 191.800 21.200 199.800 ;
        RECT 22.000 192.400 22.800 199.800 ;
        RECT 25.200 192.400 26.000 199.800 ;
        RECT 26.800 195.800 27.600 199.800 ;
        RECT 27.000 195.600 27.600 195.800 ;
        RECT 30.000 195.800 30.800 199.800 ;
        RECT 30.000 195.600 30.600 195.800 ;
        RECT 27.000 195.000 30.600 195.600 ;
        RECT 27.000 192.400 27.600 195.000 ;
        RECT 28.400 192.800 29.200 194.400 ;
        RECT 22.000 191.800 26.000 192.400 ;
        RECT 20.600 190.400 21.200 191.800 ;
        RECT 26.800 191.600 27.600 192.400 ;
        RECT 24.400 190.400 25.200 190.800 ;
        RECT 20.400 189.800 22.800 190.400 ;
        RECT 24.400 189.800 26.000 190.400 ;
        RECT 20.400 189.600 21.200 189.800 ;
        RECT 20.400 186.300 21.200 186.400 ;
        RECT 18.800 185.700 21.200 186.300 ;
        RECT 22.200 186.200 22.800 189.800 ;
        RECT 25.200 189.600 26.000 189.800 ;
        RECT 23.600 187.600 24.400 189.200 ;
        RECT 27.000 188.400 27.600 191.600 ;
        RECT 31.600 192.300 32.400 192.400 ;
        RECT 33.200 192.300 34.000 192.400 ;
        RECT 31.600 191.700 34.000 192.300 ;
        RECT 31.600 190.800 32.400 191.700 ;
        RECT 33.200 191.600 34.000 191.700 ;
        RECT 29.200 189.600 30.800 190.400 ;
        RECT 25.200 188.300 26.000 188.400 ;
        RECT 27.000 188.300 28.600 188.400 ;
        RECT 25.200 188.200 28.600 188.300 ;
        RECT 25.200 187.700 28.800 188.200 ;
        RECT 25.200 187.600 26.000 187.700 ;
        RECT 13.000 184.400 13.800 185.600 ;
        RECT 9.200 182.200 10.000 184.200 ;
        RECT 13.000 183.600 14.800 184.400 ;
        RECT 13.000 182.200 13.800 183.600 ;
        RECT 18.800 182.200 19.600 185.700 ;
        RECT 20.400 185.600 21.200 185.700 ;
        RECT 20.600 184.800 21.400 185.600 ;
        RECT 22.000 182.200 22.800 186.200 ;
        RECT 28.000 182.200 28.800 187.700 ;
        RECT 33.200 186.800 34.000 188.400 ;
        RECT 34.800 186.200 35.600 199.800 ;
        RECT 40.200 194.300 41.000 199.800 ;
        RECT 38.100 193.700 41.000 194.300 ;
        RECT 36.400 192.300 37.200 193.200 ;
        RECT 38.100 192.300 38.700 193.700 ;
        RECT 36.400 191.700 38.700 192.300 ;
        RECT 40.200 192.600 41.000 193.700 ;
        RECT 40.200 191.800 42.000 192.600 ;
        RECT 46.600 192.400 47.400 199.800 ;
        RECT 46.400 191.800 47.400 192.400 ;
        RECT 36.400 191.600 37.200 191.700 ;
        RECT 41.200 188.400 41.800 191.800 ;
        RECT 46.400 188.400 47.000 191.800 ;
        RECT 47.600 190.300 48.400 190.400 ;
        RECT 52.400 190.300 53.200 199.800 ;
        RECT 54.000 192.400 54.800 199.800 ;
        RECT 57.200 192.400 58.000 199.800 ;
        RECT 54.000 191.800 58.000 192.400 ;
        RECT 58.800 191.800 59.600 199.800 ;
        RECT 54.800 190.400 55.600 190.800 ;
        RECT 58.800 190.400 59.400 191.800 ;
        RECT 54.000 190.300 55.600 190.400 ;
        RECT 47.600 189.800 55.600 190.300 ;
        RECT 57.200 189.800 59.600 190.400 ;
        RECT 47.600 189.700 54.800 189.800 ;
        RECT 47.600 188.800 48.400 189.700 ;
        RECT 41.200 187.600 42.000 188.400 ;
        RECT 44.400 187.600 47.000 188.400 ;
        RECT 34.800 185.600 36.600 186.200 ;
        RECT 35.800 184.300 36.600 185.600 ;
        RECT 38.000 184.300 38.800 184.400 ;
        RECT 35.800 183.700 38.800 184.300 ;
        RECT 35.800 182.200 36.600 183.700 ;
        RECT 38.000 183.600 38.800 183.700 ;
        RECT 41.200 184.200 41.800 187.600 ;
        RECT 44.600 186.200 45.200 187.600 ;
        RECT 50.800 186.800 51.600 188.400 ;
        RECT 46.200 186.200 49.800 186.600 ;
        RECT 41.200 182.200 42.000 184.200 ;
        RECT 44.400 182.200 45.200 186.200 ;
        RECT 46.000 186.000 50.000 186.200 ;
        RECT 46.000 182.200 46.800 186.000 ;
        RECT 49.200 182.200 50.000 186.000 ;
        RECT 52.400 182.200 53.200 189.700 ;
        RECT 54.000 189.600 54.800 189.700 ;
        RECT 57.200 186.200 57.800 189.800 ;
        RECT 58.800 189.600 59.600 189.800 ;
        RECT 62.000 186.400 62.800 199.800 ;
        RECT 67.800 192.600 68.600 199.800 ;
        RECT 66.800 191.800 68.600 192.600 ;
        RECT 72.600 192.400 73.400 199.800 ;
        RECT 74.000 193.600 74.800 194.400 ;
        RECT 74.200 192.400 74.800 193.600 ;
        RECT 79.600 192.400 80.400 199.800 ;
        RECT 72.600 191.800 73.600 192.400 ;
        RECT 74.200 191.800 75.600 192.400 ;
        RECT 67.000 188.400 67.600 191.800 ;
        RECT 71.600 188.800 72.400 190.400 ;
        RECT 73.000 188.400 73.600 191.800 ;
        RECT 74.800 191.600 75.600 191.800 ;
        RECT 78.200 191.800 80.400 192.400 ;
        RECT 78.200 191.200 78.800 191.800 ;
        RECT 77.600 190.400 78.800 191.200 ;
        RECT 66.800 188.300 67.600 188.400 ;
        RECT 70.000 188.300 70.800 188.400 ;
        RECT 66.800 188.200 70.800 188.300 ;
        RECT 66.800 187.700 71.600 188.200 ;
        RECT 66.800 187.600 67.600 187.700 ;
        RECT 70.000 187.600 71.600 187.700 ;
        RECT 73.000 187.600 75.600 188.400 ;
        RECT 57.200 182.200 58.000 186.200 ;
        RECT 58.800 185.600 59.600 186.400 ;
        RECT 60.400 185.600 62.800 186.400 ;
        RECT 58.600 184.800 59.400 185.600 ;
        RECT 61.000 182.200 61.800 185.600 ;
        RECT 67.000 184.200 67.600 187.600 ;
        RECT 70.800 187.200 71.600 187.600 ;
        RECT 70.200 186.200 73.800 186.600 ;
        RECT 74.800 186.200 75.400 187.600 ;
        RECT 78.200 187.400 78.800 190.400 ;
        RECT 79.600 188.800 80.400 190.400 ;
        RECT 78.200 186.800 80.400 187.400 ;
        RECT 81.200 186.800 82.000 188.400 ;
        RECT 66.800 182.200 67.600 184.200 ;
        RECT 70.000 186.000 74.000 186.200 ;
        RECT 70.000 182.200 70.800 186.000 ;
        RECT 73.200 182.200 74.000 186.000 ;
        RECT 74.800 182.200 75.600 186.200 ;
        RECT 79.600 182.200 80.400 186.800 ;
        RECT 82.800 186.200 83.600 199.800 ;
        RECT 88.400 193.600 89.200 194.400 ;
        RECT 84.400 191.600 85.200 193.200 ;
        RECT 88.400 192.400 89.000 193.600 ;
        RECT 89.800 192.400 90.600 199.800 ;
        RECT 87.600 191.800 89.000 192.400 ;
        RECT 89.600 191.800 90.600 192.400 ;
        RECT 87.600 191.600 88.400 191.800 ;
        RECT 84.500 190.300 85.100 191.600 ;
        RECT 89.600 190.300 90.200 191.800 ;
        RECT 84.500 189.700 90.200 190.300 ;
        RECT 89.600 188.400 90.200 189.700 ;
        RECT 90.800 190.300 91.600 190.400 ;
        RECT 94.000 190.300 94.800 199.800 ;
        RECT 99.800 192.600 100.600 199.800 ;
        RECT 98.800 191.800 100.600 192.600 ;
        RECT 90.800 189.700 94.800 190.300 ;
        RECT 90.800 188.800 91.600 189.700 ;
        RECT 87.600 187.600 90.200 188.400 ;
        RECT 92.400 188.200 93.200 188.400 ;
        RECT 91.600 187.600 93.200 188.200 ;
        RECT 87.800 186.200 88.400 187.600 ;
        RECT 91.600 187.200 92.400 187.600 ;
        RECT 89.400 186.200 93.000 186.600 ;
        RECT 82.800 185.600 84.600 186.200 ;
        RECT 83.800 182.200 84.600 185.600 ;
        RECT 87.600 182.200 88.400 186.200 ;
        RECT 89.200 186.000 93.200 186.200 ;
        RECT 89.200 182.200 90.000 186.000 ;
        RECT 92.400 182.200 93.200 186.000 ;
        RECT 94.000 182.200 94.800 189.700 ;
        RECT 99.000 188.400 99.600 191.800 ;
        RECT 102.000 191.600 102.800 193.200 ;
        RECT 100.400 190.300 101.200 191.200 ;
        RECT 102.100 190.300 102.700 191.600 ;
        RECT 100.400 189.700 102.700 190.300 ;
        RECT 100.400 189.600 101.200 189.700 ;
        RECT 95.600 188.300 96.400 188.400 ;
        RECT 98.800 188.300 99.600 188.400 ;
        RECT 95.600 187.700 99.600 188.300 ;
        RECT 95.600 187.600 96.400 187.700 ;
        RECT 98.800 187.600 99.600 187.700 ;
        RECT 95.600 184.800 96.400 186.400 ;
        RECT 97.200 184.800 98.000 186.400 ;
        RECT 99.000 184.200 99.600 187.600 ;
        RECT 103.600 186.200 104.400 199.800 ;
        RECT 105.200 188.300 106.000 188.400 ;
        RECT 106.800 188.300 107.600 199.800 ;
        RECT 113.200 192.400 114.000 199.800 ;
        RECT 111.800 191.800 114.000 192.400 ;
        RECT 116.400 192.000 117.200 199.800 ;
        RECT 119.600 195.200 120.400 199.800 ;
        RECT 111.800 191.200 112.400 191.800 ;
        RECT 111.200 190.400 112.400 191.200 ;
        RECT 116.200 191.200 117.200 192.000 ;
        RECT 117.800 194.600 120.400 195.200 ;
        RECT 117.800 193.000 118.400 194.600 ;
        RECT 122.800 194.400 123.600 199.800 ;
        RECT 126.000 197.000 126.800 199.800 ;
        RECT 127.600 197.000 128.400 199.800 ;
        RECT 129.200 197.000 130.000 199.800 ;
        RECT 124.200 194.400 128.400 195.200 ;
        RECT 121.000 193.600 123.600 194.400 ;
        RECT 130.800 193.600 131.600 199.800 ;
        RECT 134.000 195.000 134.800 199.800 ;
        RECT 137.200 195.000 138.000 199.800 ;
        RECT 138.800 197.000 139.600 199.800 ;
        RECT 140.400 197.000 141.200 199.800 ;
        RECT 143.600 195.200 144.400 199.800 ;
        RECT 146.800 196.400 147.600 199.800 ;
        RECT 146.800 195.800 147.800 196.400 ;
        RECT 147.200 195.200 147.800 195.800 ;
        RECT 142.400 194.400 146.600 195.200 ;
        RECT 147.200 194.600 149.200 195.200 ;
        RECT 134.000 193.600 136.600 194.400 ;
        RECT 137.200 193.800 143.000 194.400 ;
        RECT 146.000 194.000 146.600 194.400 ;
        RECT 126.000 193.000 126.800 193.200 ;
        RECT 117.800 192.400 126.800 193.000 ;
        RECT 129.200 193.000 130.000 193.200 ;
        RECT 137.200 193.000 137.800 193.800 ;
        RECT 143.600 193.200 145.000 193.800 ;
        RECT 146.000 193.200 147.600 194.000 ;
        RECT 129.200 192.400 137.800 193.000 ;
        RECT 138.800 193.000 145.000 193.200 ;
        RECT 138.800 192.600 144.200 193.000 ;
        RECT 138.800 192.400 139.600 192.600 ;
        RECT 105.200 187.700 107.600 188.300 ;
        RECT 105.200 186.800 106.000 187.700 ;
        RECT 102.600 185.600 104.400 186.200 ;
        RECT 102.600 184.400 103.400 185.600 ;
        RECT 98.800 182.200 99.600 184.200 ;
        RECT 102.000 183.600 103.400 184.400 ;
        RECT 102.600 182.200 103.400 183.600 ;
        RECT 106.800 182.200 107.600 187.700 ;
        RECT 111.800 187.400 112.400 190.400 ;
        RECT 113.200 190.300 114.000 190.400 ;
        RECT 116.200 190.300 117.000 191.200 ;
        RECT 117.800 190.600 118.400 192.400 ;
        RECT 113.200 189.700 117.000 190.300 ;
        RECT 113.200 188.800 114.000 189.700 ;
        RECT 111.800 186.800 114.000 187.400 ;
        RECT 108.400 184.800 109.200 186.400 ;
        RECT 113.200 182.200 114.000 186.800 ;
        RECT 116.200 186.800 117.000 189.700 ;
        RECT 117.600 190.000 118.400 190.600 ;
        RECT 124.400 190.000 147.800 190.600 ;
        RECT 117.600 188.000 118.200 190.000 ;
        RECT 124.400 189.400 125.200 190.000 ;
        RECT 142.000 189.600 142.800 190.000 ;
        RECT 145.200 189.600 146.000 190.000 ;
        RECT 147.000 189.800 147.800 190.000 ;
        RECT 118.800 188.600 122.600 189.400 ;
        RECT 117.600 187.400 118.800 188.000 ;
        RECT 114.800 186.300 115.600 186.400 ;
        RECT 116.200 186.300 117.200 186.800 ;
        RECT 114.800 185.700 117.200 186.300 ;
        RECT 114.800 185.600 115.600 185.700 ;
        RECT 116.400 182.200 117.200 185.700 ;
        RECT 118.000 182.200 118.800 187.400 ;
        RECT 121.800 187.400 122.600 188.600 ;
        RECT 121.800 186.800 123.600 187.400 ;
        RECT 122.800 186.200 123.600 186.800 ;
        RECT 127.600 186.400 128.400 189.200 ;
        RECT 130.800 188.600 134.000 189.400 ;
        RECT 137.800 188.600 139.800 189.400 ;
        RECT 148.400 189.000 149.200 194.600 ;
        RECT 151.600 192.400 152.400 199.800 ;
        RECT 159.600 192.400 160.400 199.800 ;
        RECT 162.800 196.400 163.600 199.800 ;
        RECT 162.600 195.800 163.600 196.400 ;
        RECT 162.600 195.200 163.200 195.800 ;
        RECT 166.000 195.200 166.800 199.800 ;
        RECT 169.200 197.000 170.000 199.800 ;
        RECT 170.800 197.000 171.600 199.800 ;
        RECT 151.600 191.800 153.800 192.400 ;
        RECT 153.200 191.200 153.800 191.800 ;
        RECT 158.200 191.800 160.400 192.400 ;
        RECT 161.200 194.600 163.200 195.200 ;
        RECT 158.200 191.200 158.800 191.800 ;
        RECT 153.200 190.400 154.400 191.200 ;
        RECT 157.600 190.400 158.800 191.200 ;
        RECT 130.400 187.800 131.200 188.000 ;
        RECT 130.400 187.200 134.800 187.800 ;
        RECT 134.000 187.000 134.800 187.200 ;
        RECT 135.600 186.800 136.400 188.400 ;
        RECT 122.800 185.400 125.200 186.200 ;
        RECT 127.600 185.600 128.600 186.400 ;
        RECT 131.600 185.600 133.200 186.400 ;
        RECT 134.000 186.200 134.800 186.400 ;
        RECT 137.800 186.200 138.600 188.600 ;
        RECT 140.400 188.200 149.200 189.000 ;
        RECT 151.600 188.800 152.400 190.400 ;
        RECT 143.800 186.800 146.800 187.600 ;
        RECT 143.800 186.200 144.600 186.800 ;
        RECT 134.000 185.600 138.600 186.200 ;
        RECT 124.400 182.200 125.200 185.400 ;
        RECT 142.000 185.400 144.600 186.200 ;
        RECT 126.000 182.200 126.800 185.000 ;
        RECT 127.600 182.200 128.400 185.000 ;
        RECT 129.200 182.200 130.000 185.000 ;
        RECT 130.800 182.200 131.600 185.000 ;
        RECT 134.000 182.200 134.800 185.000 ;
        RECT 137.200 182.200 138.000 185.000 ;
        RECT 138.800 182.200 139.600 185.000 ;
        RECT 140.400 182.200 141.200 185.000 ;
        RECT 142.000 182.200 142.800 185.400 ;
        RECT 148.400 182.200 149.200 188.200 ;
        RECT 153.200 187.400 153.800 190.400 ;
        RECT 151.600 186.800 153.800 187.400 ;
        RECT 158.200 187.400 158.800 190.400 ;
        RECT 159.600 188.800 160.400 190.400 ;
        RECT 161.200 189.000 162.000 194.600 ;
        RECT 163.800 194.400 168.000 195.200 ;
        RECT 172.400 195.000 173.200 199.800 ;
        RECT 175.600 195.000 176.400 199.800 ;
        RECT 163.800 194.000 164.400 194.400 ;
        RECT 162.800 193.200 164.400 194.000 ;
        RECT 167.400 193.800 173.200 194.400 ;
        RECT 165.400 193.200 166.800 193.800 ;
        RECT 165.400 193.000 171.600 193.200 ;
        RECT 166.200 192.600 171.600 193.000 ;
        RECT 170.800 192.400 171.600 192.600 ;
        RECT 172.600 193.000 173.200 193.800 ;
        RECT 173.800 193.600 176.400 194.400 ;
        RECT 178.800 193.600 179.600 199.800 ;
        RECT 180.400 197.000 181.200 199.800 ;
        RECT 182.000 197.000 182.800 199.800 ;
        RECT 183.600 197.000 184.400 199.800 ;
        RECT 182.000 194.400 186.200 195.200 ;
        RECT 186.800 194.400 187.600 199.800 ;
        RECT 190.000 195.200 190.800 199.800 ;
        RECT 190.000 194.600 192.600 195.200 ;
        RECT 186.800 193.600 189.400 194.400 ;
        RECT 180.400 193.000 181.200 193.200 ;
        RECT 172.600 192.400 181.200 193.000 ;
        RECT 183.600 193.000 184.400 193.200 ;
        RECT 192.000 193.000 192.600 194.600 ;
        RECT 183.600 192.400 192.600 193.000 ;
        RECT 192.000 190.600 192.600 192.400 ;
        RECT 193.200 192.000 194.000 199.800 ;
        RECT 198.000 192.400 198.800 199.800 ;
        RECT 193.200 191.200 194.200 192.000 ;
        RECT 198.000 191.800 200.200 192.400 ;
        RECT 202.800 191.800 203.600 199.800 ;
        RECT 204.400 192.400 205.200 199.800 ;
        RECT 207.600 192.400 208.400 199.800 ;
        RECT 204.400 191.800 208.400 192.400 ;
        RECT 209.800 192.600 210.600 199.800 ;
        RECT 209.800 191.800 211.600 192.600 ;
        RECT 162.600 190.000 186.000 190.600 ;
        RECT 192.000 190.000 192.800 190.600 ;
        RECT 162.600 189.800 163.600 190.000 ;
        RECT 162.800 189.600 163.600 189.800 ;
        RECT 167.600 189.600 168.400 190.000 ;
        RECT 185.200 189.400 186.000 190.000 ;
        RECT 161.200 188.200 170.000 189.000 ;
        RECT 170.600 188.600 172.600 189.400 ;
        RECT 176.400 188.600 179.600 189.400 ;
        RECT 158.200 186.800 160.400 187.400 ;
        RECT 151.600 182.200 152.400 186.800 ;
        RECT 159.600 182.200 160.400 186.800 ;
        RECT 161.200 182.200 162.000 188.200 ;
        RECT 163.600 186.800 166.600 187.600 ;
        RECT 165.800 186.200 166.600 186.800 ;
        RECT 171.800 186.200 172.600 188.600 ;
        RECT 174.000 186.800 174.800 188.400 ;
        RECT 179.200 187.800 180.000 188.000 ;
        RECT 175.600 187.200 180.000 187.800 ;
        RECT 175.600 187.000 176.400 187.200 ;
        RECT 182.000 186.400 182.800 189.200 ;
        RECT 187.800 188.600 191.600 189.400 ;
        RECT 187.800 187.400 188.600 188.600 ;
        RECT 192.200 188.000 192.800 190.000 ;
        RECT 175.600 186.200 176.400 186.400 ;
        RECT 165.800 185.400 168.400 186.200 ;
        RECT 171.800 185.600 176.400 186.200 ;
        RECT 177.200 185.600 178.800 186.400 ;
        RECT 181.800 185.600 182.800 186.400 ;
        RECT 186.800 186.800 188.600 187.400 ;
        RECT 191.600 187.400 192.800 188.000 ;
        RECT 193.400 190.300 194.200 191.200 ;
        RECT 199.600 191.200 200.200 191.800 ;
        RECT 199.600 190.400 200.800 191.200 ;
        RECT 203.000 190.400 203.600 191.800 ;
        RECT 206.800 190.400 207.600 190.800 ;
        RECT 198.000 190.300 198.800 190.400 ;
        RECT 193.400 189.700 198.800 190.300 ;
        RECT 186.800 186.200 187.600 186.800 ;
        RECT 167.600 182.200 168.400 185.400 ;
        RECT 185.200 185.400 187.600 186.200 ;
        RECT 169.200 182.200 170.000 185.000 ;
        RECT 170.800 182.200 171.600 185.000 ;
        RECT 172.400 182.200 173.200 185.000 ;
        RECT 175.600 182.200 176.400 185.000 ;
        RECT 178.800 182.200 179.600 185.000 ;
        RECT 180.400 182.200 181.200 185.000 ;
        RECT 182.000 182.200 182.800 185.000 ;
        RECT 183.600 182.200 184.400 185.000 ;
        RECT 185.200 182.200 186.000 185.400 ;
        RECT 191.600 182.200 192.400 187.400 ;
        RECT 193.400 186.800 194.200 189.700 ;
        RECT 198.000 188.800 198.800 189.700 ;
        RECT 199.600 187.400 200.200 190.400 ;
        RECT 202.800 189.800 205.200 190.400 ;
        RECT 206.800 189.800 208.400 190.400 ;
        RECT 202.800 189.600 203.600 189.800 ;
        RECT 193.200 186.000 194.200 186.800 ;
        RECT 198.000 186.800 200.200 187.400 ;
        RECT 193.200 182.200 194.000 186.000 ;
        RECT 198.000 182.200 198.800 186.800 ;
        RECT 202.800 185.600 203.600 186.400 ;
        RECT 204.600 186.200 205.200 189.800 ;
        RECT 207.600 189.600 208.400 189.800 ;
        RECT 209.200 189.600 210.000 191.200 ;
        RECT 206.000 188.300 206.800 189.200 ;
        RECT 209.300 188.300 209.900 189.600 ;
        RECT 206.000 187.700 209.900 188.300 ;
        RECT 210.800 188.400 211.400 191.800 ;
        RECT 212.400 190.300 213.200 190.400 ;
        RECT 214.000 190.300 214.800 199.800 ;
        RECT 217.200 192.400 218.000 199.800 ;
        RECT 217.200 191.800 219.400 192.400 ;
        RECT 218.800 191.200 219.400 191.800 ;
        RECT 218.800 190.400 220.000 191.200 ;
        RECT 212.400 189.700 214.800 190.300 ;
        RECT 212.400 189.600 213.200 189.700 ;
        RECT 206.000 187.600 206.800 187.700 ;
        RECT 210.800 187.600 211.600 188.400 ;
        RECT 203.000 184.800 203.800 185.600 ;
        RECT 204.400 182.200 205.200 186.200 ;
        RECT 209.200 186.300 210.000 186.400 ;
        RECT 210.800 186.300 211.400 187.600 ;
        RECT 209.200 185.700 211.500 186.300 ;
        RECT 209.200 185.600 210.000 185.700 ;
        RECT 210.800 184.200 211.400 185.700 ;
        RECT 210.800 182.200 211.600 184.200 ;
        RECT 214.000 182.200 214.800 189.700 ;
        RECT 215.600 190.300 216.400 190.400 ;
        RECT 217.200 190.300 218.000 190.400 ;
        RECT 215.600 189.700 218.000 190.300 ;
        RECT 215.600 189.600 216.400 189.700 ;
        RECT 217.200 188.800 218.000 189.700 ;
        RECT 218.800 187.400 219.400 190.400 ;
        RECT 217.200 186.800 219.400 187.400 ;
        RECT 215.600 184.800 216.400 186.400 ;
        RECT 217.200 182.200 218.000 186.800 ;
        RECT 1.200 176.000 2.000 179.800 ;
        RECT 4.400 176.000 5.200 179.800 ;
        RECT 1.200 175.800 5.200 176.000 ;
        RECT 6.000 175.800 6.800 179.800 ;
        RECT 7.600 176.000 8.400 179.800 ;
        RECT 10.800 176.000 11.600 179.800 ;
        RECT 7.600 175.800 11.600 176.000 ;
        RECT 12.400 175.800 13.200 179.800 ;
        RECT 15.600 176.000 16.400 179.800 ;
        RECT 1.400 175.400 5.000 175.800 ;
        RECT 6.000 174.400 6.600 175.800 ;
        RECT 7.800 175.400 11.400 175.800 ;
        RECT 8.400 174.400 9.200 174.800 ;
        RECT 12.400 174.400 13.000 175.800 ;
        RECT 15.400 175.200 16.400 176.000 ;
        RECT 4.200 173.600 6.800 174.400 ;
        RECT 7.600 173.800 9.200 174.400 ;
        RECT 10.600 174.300 13.200 174.400 ;
        RECT 14.000 174.300 14.800 174.400 ;
        RECT 7.600 173.600 8.400 173.800 ;
        RECT 10.600 173.700 14.800 174.300 ;
        RECT 10.600 173.600 13.200 173.700 ;
        RECT 14.000 173.600 14.800 173.700 ;
        RECT 2.800 171.600 3.600 173.200 ;
        RECT 4.200 172.300 4.800 173.600 ;
        RECT 9.200 172.300 10.000 173.200 ;
        RECT 4.200 171.700 10.000 172.300 ;
        RECT 4.200 170.200 4.800 171.700 ;
        RECT 9.200 171.600 10.000 171.700 ;
        RECT 6.000 170.200 6.800 170.400 ;
        RECT 10.600 170.200 11.200 173.600 ;
        RECT 15.400 170.800 16.200 175.200 ;
        RECT 17.200 174.600 18.000 179.800 ;
        RECT 23.600 176.600 24.400 179.800 ;
        RECT 25.200 177.000 26.000 179.800 ;
        RECT 26.800 177.000 27.600 179.800 ;
        RECT 28.400 177.000 29.200 179.800 ;
        RECT 30.000 177.000 30.800 179.800 ;
        RECT 33.200 177.000 34.000 179.800 ;
        RECT 36.400 177.000 37.200 179.800 ;
        RECT 38.000 177.000 38.800 179.800 ;
        RECT 39.600 177.000 40.400 179.800 ;
        RECT 22.000 175.800 24.400 176.600 ;
        RECT 41.200 176.600 42.000 179.800 ;
        RECT 22.000 175.200 22.800 175.800 ;
        RECT 16.800 174.000 18.000 174.600 ;
        RECT 21.000 174.600 22.800 175.200 ;
        RECT 26.800 175.600 27.800 176.400 ;
        RECT 30.800 175.600 32.400 176.400 ;
        RECT 33.200 175.800 37.800 176.400 ;
        RECT 41.200 175.800 43.800 176.600 ;
        RECT 33.200 175.600 34.000 175.800 ;
        RECT 16.800 172.000 17.400 174.000 ;
        RECT 21.000 173.400 21.800 174.600 ;
        RECT 18.000 172.600 21.800 173.400 ;
        RECT 26.800 172.800 27.600 175.600 ;
        RECT 33.200 174.800 34.000 175.000 ;
        RECT 29.600 174.200 34.000 174.800 ;
        RECT 29.600 174.000 30.400 174.200 ;
        RECT 34.800 173.600 35.600 175.200 ;
        RECT 37.000 173.400 37.800 175.800 ;
        RECT 43.000 175.200 43.800 175.800 ;
        RECT 43.000 174.400 46.000 175.200 ;
        RECT 47.600 173.800 48.400 179.800 ;
        RECT 52.000 174.200 52.800 179.800 ;
        RECT 57.200 176.000 58.000 179.800 ;
        RECT 60.400 176.000 61.200 179.800 ;
        RECT 57.200 175.800 61.200 176.000 ;
        RECT 62.000 175.800 62.800 179.800 ;
        RECT 63.600 175.800 64.400 179.800 ;
        RECT 65.200 176.000 66.000 179.800 ;
        RECT 68.400 176.000 69.200 179.800 ;
        RECT 65.200 175.800 69.200 176.000 ;
        RECT 70.000 175.800 70.800 179.800 ;
        RECT 71.600 176.000 72.400 179.800 ;
        RECT 74.800 176.000 75.600 179.800 ;
        RECT 71.600 175.800 75.600 176.000 ;
        RECT 76.400 175.800 77.200 179.800 ;
        RECT 80.800 176.200 82.400 179.800 ;
        RECT 57.400 175.400 61.000 175.800 ;
        RECT 62.000 174.400 62.600 175.800 ;
        RECT 63.800 174.400 64.400 175.800 ;
        RECT 65.400 175.400 69.000 175.800 ;
        RECT 67.600 174.400 68.400 174.800 ;
        RECT 70.200 174.400 70.800 175.800 ;
        RECT 71.800 175.400 75.400 175.800 ;
        RECT 76.400 175.200 78.800 175.800 ;
        RECT 78.000 175.000 78.800 175.200 ;
        RECT 79.400 174.800 80.200 175.600 ;
        RECT 74.000 174.400 74.800 174.800 ;
        RECT 79.400 174.400 80.000 174.800 ;
        RECT 30.000 172.600 33.200 173.400 ;
        RECT 37.000 172.600 39.000 173.400 ;
        RECT 39.600 173.000 48.400 173.800 ;
        RECT 23.600 172.000 24.400 172.600 ;
        RECT 41.200 172.000 42.000 172.400 ;
        RECT 46.200 172.000 47.000 172.200 ;
        RECT 16.800 171.400 17.600 172.000 ;
        RECT 23.600 171.400 47.000 172.000 ;
        RECT 12.400 170.200 13.200 170.400 ;
        RECT 3.800 169.600 4.800 170.200 ;
        RECT 5.400 169.600 6.800 170.200 ;
        RECT 10.200 169.600 11.200 170.200 ;
        RECT 11.800 169.600 13.200 170.200 ;
        RECT 15.400 170.000 16.400 170.800 ;
        RECT 3.800 162.200 4.600 169.600 ;
        RECT 5.400 168.400 6.000 169.600 ;
        RECT 5.200 167.600 6.000 168.400 ;
        RECT 10.200 162.200 11.000 169.600 ;
        RECT 11.800 168.400 12.400 169.600 ;
        RECT 11.600 167.600 12.400 168.400 ;
        RECT 14.000 168.300 14.800 168.400 ;
        RECT 15.600 168.300 16.400 170.000 ;
        RECT 14.000 167.700 16.400 168.300 ;
        RECT 14.000 167.600 14.800 167.700 ;
        RECT 15.600 162.200 16.400 167.700 ;
        RECT 17.000 169.600 17.600 171.400 ;
        RECT 17.000 169.000 26.000 169.600 ;
        RECT 17.000 167.400 17.600 169.000 ;
        RECT 25.200 168.800 26.000 169.000 ;
        RECT 28.400 169.000 37.000 169.600 ;
        RECT 28.400 168.800 29.200 169.000 ;
        RECT 20.200 167.600 22.800 168.400 ;
        RECT 17.000 166.800 19.600 167.400 ;
        RECT 18.800 162.200 19.600 166.800 ;
        RECT 22.000 162.200 22.800 167.600 ;
        RECT 23.400 166.800 27.600 167.600 ;
        RECT 25.200 162.200 26.000 165.000 ;
        RECT 26.800 162.200 27.600 165.000 ;
        RECT 28.400 162.200 29.200 165.000 ;
        RECT 30.000 162.200 30.800 168.400 ;
        RECT 33.200 167.600 35.800 168.400 ;
        RECT 36.400 168.200 37.000 169.000 ;
        RECT 38.000 169.400 38.800 169.600 ;
        RECT 38.000 169.000 43.400 169.400 ;
        RECT 38.000 168.800 44.200 169.000 ;
        RECT 42.800 168.200 44.200 168.800 ;
        RECT 36.400 167.600 42.200 168.200 ;
        RECT 45.200 168.000 46.800 168.800 ;
        RECT 45.200 167.600 45.800 168.000 ;
        RECT 33.200 162.200 34.000 167.000 ;
        RECT 36.400 162.200 37.200 167.000 ;
        RECT 41.600 166.800 45.800 167.600 ;
        RECT 47.600 167.400 48.400 173.000 ;
        RECT 51.000 173.800 52.800 174.200 ;
        RECT 51.000 173.600 52.600 173.800 ;
        RECT 60.200 173.600 62.800 174.400 ;
        RECT 63.600 173.600 66.200 174.400 ;
        RECT 67.600 173.800 69.200 174.400 ;
        RECT 68.400 173.600 69.200 173.800 ;
        RECT 70.000 173.600 72.600 174.400 ;
        RECT 74.000 174.300 75.600 174.400 ;
        RECT 76.400 174.300 78.000 174.400 ;
        RECT 74.000 173.800 78.000 174.300 ;
        RECT 74.800 173.700 78.000 173.800 ;
        RECT 74.800 173.600 75.600 173.700 ;
        RECT 76.400 173.600 78.000 173.700 ;
        RECT 79.200 173.600 80.000 174.400 ;
        RECT 80.800 174.200 81.400 176.200 ;
        RECT 86.000 175.800 86.800 179.800 ;
        RECT 82.000 174.800 83.600 175.600 ;
        RECT 84.200 175.200 86.800 175.800 ;
        RECT 84.200 175.000 85.000 175.200 ;
        RECT 85.200 174.200 86.800 174.400 ;
        RECT 80.800 173.600 81.800 174.200 ;
        RECT 84.600 174.000 86.800 174.200 ;
        RECT 51.000 170.400 51.600 173.600 ;
        RECT 53.200 171.600 54.800 172.400 ;
        RECT 58.800 171.600 59.600 173.200 ;
        RECT 60.200 172.300 60.800 173.600 ;
        RECT 60.200 171.700 64.300 172.300 ;
        RECT 50.800 169.600 51.600 170.400 ;
        RECT 55.600 169.600 56.400 171.200 ;
        RECT 60.200 170.200 60.800 171.700 ;
        RECT 63.700 170.400 64.300 171.700 ;
        RECT 62.000 170.200 62.800 170.400 ;
        RECT 59.800 169.600 60.800 170.200 ;
        RECT 61.400 169.600 62.800 170.200 ;
        RECT 63.600 170.200 64.400 170.400 ;
        RECT 65.600 170.200 66.200 173.600 ;
        RECT 66.800 171.600 67.600 173.200 ;
        RECT 68.400 172.300 69.200 172.400 ;
        RECT 72.000 172.300 72.600 173.600 ;
        RECT 68.400 171.700 72.600 172.300 ;
        RECT 68.400 171.600 69.200 171.700 ;
        RECT 70.000 170.200 70.800 170.400 ;
        RECT 72.000 170.200 72.600 171.700 ;
        RECT 73.200 172.300 74.000 173.200 ;
        RECT 81.200 172.400 81.800 173.600 ;
        RECT 82.400 173.600 86.800 174.000 ;
        RECT 82.400 173.400 85.200 173.600 ;
        RECT 82.400 173.200 83.200 173.400 ;
        RECT 76.400 172.300 77.200 172.400 ;
        RECT 73.200 171.700 77.200 172.300 ;
        RECT 73.200 171.600 74.000 171.700 ;
        RECT 76.400 171.600 77.200 171.700 ;
        RECT 79.600 172.300 80.400 172.400 ;
        RECT 81.200 172.300 82.000 172.400 ;
        RECT 79.600 171.700 82.000 172.300 ;
        RECT 83.800 172.200 84.600 172.400 ;
        RECT 79.600 171.600 80.400 171.700 ;
        RECT 81.200 171.600 82.000 171.700 ;
        RECT 83.000 171.600 84.600 172.200 ;
        RECT 90.800 172.300 91.600 179.800 ;
        RECT 92.400 176.000 93.200 179.800 ;
        RECT 95.600 176.000 96.400 179.800 ;
        RECT 92.400 175.800 96.400 176.000 ;
        RECT 97.200 175.800 98.000 179.800 ;
        RECT 98.800 175.800 99.600 179.800 ;
        RECT 100.400 176.000 101.200 179.800 ;
        RECT 103.600 176.000 104.400 179.800 ;
        RECT 100.400 175.800 104.400 176.000 ;
        RECT 106.800 177.800 107.600 179.800 ;
        RECT 92.600 175.400 96.200 175.800 ;
        RECT 93.200 174.400 94.000 174.800 ;
        RECT 97.200 174.400 97.800 175.800 ;
        RECT 99.000 174.400 99.600 175.800 ;
        RECT 100.600 175.400 104.200 175.800 ;
        RECT 102.800 174.400 103.600 174.800 ;
        RECT 106.800 174.400 107.400 177.800 ;
        RECT 108.400 175.600 109.200 177.200 ;
        RECT 110.600 176.800 111.400 179.800 ;
        RECT 110.000 175.800 111.400 176.800 ;
        RECT 114.800 175.800 115.600 179.800 ;
        RECT 118.000 177.800 118.800 179.800 ;
        RECT 92.400 173.800 94.000 174.400 ;
        RECT 92.400 173.600 93.200 173.800 ;
        RECT 95.400 173.600 98.000 174.400 ;
        RECT 98.800 173.600 101.400 174.400 ;
        RECT 102.800 173.800 104.400 174.400 ;
        RECT 103.600 173.600 104.400 173.800 ;
        RECT 106.800 173.600 107.600 174.400 ;
        RECT 94.000 172.300 94.800 173.200 ;
        RECT 90.800 171.700 94.800 172.300 ;
        RECT 81.200 170.200 81.800 171.600 ;
        RECT 83.000 171.400 83.800 171.600 ;
        RECT 63.600 169.600 65.000 170.200 ;
        RECT 65.600 169.600 66.600 170.200 ;
        RECT 70.000 169.600 71.400 170.200 ;
        RECT 72.000 169.600 73.000 170.200 ;
        RECT 46.400 166.800 48.400 167.400 ;
        RECT 51.000 167.000 51.600 169.600 ;
        RECT 52.400 167.600 53.200 169.200 ;
        RECT 38.000 162.200 38.800 165.000 ;
        RECT 39.600 162.200 40.400 165.000 ;
        RECT 42.800 162.200 43.600 166.800 ;
        RECT 46.400 166.200 47.000 166.800 ;
        RECT 51.000 166.400 54.600 167.000 ;
        RECT 51.000 166.200 51.600 166.400 ;
        RECT 46.000 165.600 47.000 166.200 ;
        RECT 46.000 162.200 46.800 165.600 ;
        RECT 50.800 162.200 51.600 166.200 ;
        RECT 54.000 166.200 54.600 166.400 ;
        RECT 54.000 162.200 54.800 166.200 ;
        RECT 59.800 162.200 60.600 169.600 ;
        RECT 61.400 168.400 62.000 169.600 ;
        RECT 61.200 167.600 62.000 168.400 ;
        RECT 64.400 168.400 65.000 169.600 ;
        RECT 64.400 167.600 65.200 168.400 ;
        RECT 65.800 162.200 66.600 169.600 ;
        RECT 70.800 168.400 71.400 169.600 ;
        RECT 70.800 167.600 71.600 168.400 ;
        RECT 72.200 162.200 73.000 169.600 ;
        RECT 76.400 169.600 78.800 170.200 ;
        RECT 76.400 162.200 77.200 169.600 ;
        RECT 78.000 169.400 78.800 169.600 ;
        RECT 80.800 162.200 82.400 170.200 ;
        RECT 84.200 169.600 86.800 170.200 ;
        RECT 84.200 169.400 85.000 169.600 ;
        RECT 86.000 162.200 86.800 169.600 ;
        RECT 90.800 162.200 91.600 171.700 ;
        RECT 94.000 171.600 94.800 171.700 ;
        RECT 95.400 170.200 96.000 173.600 ;
        RECT 100.800 172.300 101.400 173.600 ;
        RECT 97.300 171.700 101.400 172.300 ;
        RECT 97.300 170.400 97.900 171.700 ;
        RECT 97.200 170.200 98.000 170.400 ;
        RECT 95.000 169.600 96.000 170.200 ;
        RECT 96.600 169.600 98.000 170.200 ;
        RECT 98.800 170.200 99.600 170.400 ;
        RECT 100.800 170.200 101.400 171.700 ;
        RECT 102.000 171.600 102.800 173.200 ;
        RECT 105.200 170.800 106.000 172.400 ;
        RECT 106.800 170.200 107.400 173.600 ;
        RECT 110.000 172.400 110.600 175.800 ;
        RECT 114.800 175.600 115.400 175.800 ;
        RECT 113.600 175.200 115.400 175.600 ;
        RECT 111.200 175.000 115.400 175.200 ;
        RECT 111.200 174.600 114.200 175.000 ;
        RECT 111.200 174.400 112.000 174.600 ;
        RECT 118.000 174.400 118.600 177.800 ;
        RECT 119.600 175.600 120.400 177.200 ;
        RECT 121.200 175.200 122.000 179.800 ;
        RECT 121.200 174.600 123.400 175.200 ;
        RECT 108.400 172.300 109.200 172.400 ;
        RECT 110.000 172.300 110.800 172.400 ;
        RECT 108.400 171.700 110.800 172.300 ;
        RECT 108.400 171.600 109.200 171.700 ;
        RECT 110.000 171.600 110.800 171.700 ;
        RECT 110.000 170.200 110.600 171.600 ;
        RECT 111.400 171.000 112.000 174.400 ;
        RECT 114.800 174.300 115.600 174.400 ;
        RECT 112.800 173.800 113.600 174.000 ;
        RECT 112.800 173.200 113.800 173.800 ;
        RECT 113.200 172.400 113.800 173.200 ;
        RECT 114.800 173.700 117.100 174.300 ;
        RECT 114.800 172.800 115.600 173.700 ;
        RECT 116.500 172.400 117.100 173.700 ;
        RECT 118.000 173.600 118.800 174.400 ;
        RECT 113.200 171.600 114.000 172.400 ;
        RECT 111.400 170.400 113.800 171.000 ;
        RECT 116.400 170.800 117.200 172.400 ;
        RECT 98.800 169.600 100.200 170.200 ;
        RECT 100.800 169.600 101.800 170.200 ;
        RECT 95.000 164.400 95.800 169.600 ;
        RECT 96.600 168.400 97.200 169.600 ;
        RECT 96.400 167.600 97.200 168.400 ;
        RECT 99.600 168.400 100.200 169.600 ;
        RECT 99.600 167.600 100.400 168.400 ;
        RECT 94.000 163.600 95.800 164.400 ;
        RECT 95.000 162.200 95.800 163.600 ;
        RECT 101.000 162.200 101.800 169.600 ;
        RECT 105.800 169.400 107.600 170.200 ;
        RECT 105.800 164.400 106.600 169.400 ;
        RECT 105.800 163.600 107.600 164.400 ;
        RECT 105.800 162.200 106.600 163.600 ;
        RECT 110.000 162.200 110.800 170.200 ;
        RECT 113.200 166.200 113.800 170.400 ;
        RECT 118.000 170.200 118.600 173.600 ;
        RECT 121.200 171.600 122.000 173.200 ;
        RECT 122.800 171.600 123.400 174.600 ;
        RECT 127.600 173.800 128.400 179.800 ;
        RECT 134.000 176.600 134.800 179.800 ;
        RECT 135.600 177.000 136.400 179.800 ;
        RECT 137.200 177.000 138.000 179.800 ;
        RECT 138.800 177.000 139.600 179.800 ;
        RECT 142.000 177.000 142.800 179.800 ;
        RECT 145.200 177.000 146.000 179.800 ;
        RECT 146.800 177.000 147.600 179.800 ;
        RECT 148.400 177.000 149.200 179.800 ;
        RECT 150.000 177.000 150.800 179.800 ;
        RECT 132.200 175.800 134.800 176.600 ;
        RECT 151.600 176.600 152.400 179.800 ;
        RECT 138.200 175.800 142.800 176.400 ;
        RECT 132.200 175.200 133.000 175.800 ;
        RECT 130.000 174.400 133.000 175.200 ;
        RECT 127.600 173.000 136.400 173.800 ;
        RECT 138.200 173.400 139.000 175.800 ;
        RECT 142.000 175.600 142.800 175.800 ;
        RECT 143.600 175.600 145.200 176.400 ;
        RECT 148.200 175.600 149.200 176.400 ;
        RECT 151.600 175.800 154.000 176.600 ;
        RECT 140.400 173.600 141.200 175.200 ;
        RECT 142.000 174.800 142.800 175.000 ;
        RECT 142.000 174.200 146.400 174.800 ;
        RECT 145.600 174.000 146.400 174.200 ;
        RECT 122.800 170.800 124.000 171.600 ;
        RECT 122.800 170.200 123.400 170.800 ;
        RECT 117.000 169.400 118.800 170.200 ;
        RECT 121.200 169.600 123.400 170.200 ;
        RECT 113.200 162.200 114.000 166.200 ;
        RECT 117.000 162.200 117.800 169.400 ;
        RECT 121.200 162.200 122.000 169.600 ;
        RECT 127.600 167.400 128.400 173.000 ;
        RECT 137.000 172.600 139.000 173.400 ;
        RECT 142.800 172.600 146.000 173.400 ;
        RECT 148.400 172.800 149.200 175.600 ;
        RECT 153.200 175.200 154.000 175.800 ;
        RECT 153.200 174.600 155.000 175.200 ;
        RECT 154.200 173.400 155.000 174.600 ;
        RECT 158.000 174.600 158.800 179.800 ;
        RECT 159.600 176.000 160.400 179.800 ;
        RECT 163.000 176.400 163.800 177.200 ;
        RECT 159.600 175.200 160.600 176.000 ;
        RECT 162.800 175.600 163.600 176.400 ;
        RECT 164.400 175.800 165.200 179.800 ;
        RECT 158.000 174.000 159.200 174.600 ;
        RECT 154.200 172.600 158.000 173.400 ;
        RECT 129.000 172.000 129.800 172.200 ;
        RECT 130.800 172.000 131.600 172.400 ;
        RECT 134.000 172.000 134.800 172.400 ;
        RECT 151.600 172.000 152.400 172.600 ;
        RECT 158.600 172.000 159.200 174.000 ;
        RECT 129.000 171.400 152.400 172.000 ;
        RECT 158.400 171.400 159.200 172.000 ;
        RECT 158.400 169.600 159.000 171.400 ;
        RECT 159.800 170.800 160.600 175.200 ;
        RECT 162.800 172.200 163.600 172.400 ;
        RECT 164.600 172.200 165.200 175.800 ;
        RECT 169.200 175.600 170.000 177.200 ;
        RECT 166.000 174.300 166.800 174.400 ;
        RECT 170.800 174.300 171.600 179.800 ;
        RECT 166.000 173.700 171.600 174.300 ;
        RECT 172.400 177.000 173.200 179.000 ;
        RECT 176.600 178.400 177.400 179.000 ;
        RECT 175.600 177.600 177.400 178.400 ;
        RECT 172.400 174.800 173.000 177.000 ;
        RECT 176.600 176.000 177.400 177.600 ;
        RECT 176.600 175.400 178.200 176.000 ;
        RECT 177.400 175.000 178.200 175.400 ;
        RECT 172.400 174.200 176.600 174.800 ;
        RECT 166.000 172.800 166.800 173.700 ;
        RECT 167.600 172.200 168.400 172.400 ;
        RECT 162.800 171.600 165.200 172.200 ;
        RECT 166.800 171.600 168.400 172.200 ;
        RECT 137.200 169.400 138.000 169.600 ;
        RECT 132.600 169.000 138.000 169.400 ;
        RECT 131.800 168.800 138.000 169.000 ;
        RECT 139.000 169.000 147.600 169.600 ;
        RECT 129.200 168.000 130.800 168.800 ;
        RECT 131.800 168.200 133.200 168.800 ;
        RECT 139.000 168.200 139.600 169.000 ;
        RECT 146.800 168.800 147.600 169.000 ;
        RECT 150.000 169.000 159.000 169.600 ;
        RECT 150.000 168.800 150.800 169.000 ;
        RECT 130.200 167.600 130.800 168.000 ;
        RECT 133.800 167.600 139.600 168.200 ;
        RECT 140.200 167.600 142.800 168.400 ;
        RECT 127.600 166.800 129.600 167.400 ;
        RECT 130.200 166.800 134.400 167.600 ;
        RECT 129.000 166.200 129.600 166.800 ;
        RECT 129.000 165.600 130.000 166.200 ;
        RECT 129.200 162.200 130.000 165.600 ;
        RECT 132.400 162.200 133.200 166.800 ;
        RECT 135.600 162.200 136.400 165.000 ;
        RECT 137.200 162.200 138.000 165.000 ;
        RECT 138.800 162.200 139.600 167.000 ;
        RECT 142.000 162.200 142.800 167.000 ;
        RECT 145.200 162.200 146.000 168.400 ;
        RECT 153.200 167.600 155.800 168.400 ;
        RECT 148.400 166.800 152.600 167.600 ;
        RECT 146.800 162.200 147.600 165.000 ;
        RECT 148.400 162.200 149.200 165.000 ;
        RECT 150.000 162.200 150.800 165.000 ;
        RECT 153.200 162.200 154.000 167.600 ;
        RECT 158.400 167.400 159.000 169.000 ;
        RECT 156.400 166.800 159.000 167.400 ;
        RECT 159.600 170.000 160.600 170.800 ;
        RECT 163.000 170.200 163.600 171.600 ;
        RECT 166.800 171.200 167.600 171.600 ;
        RECT 156.400 162.200 157.200 166.800 ;
        RECT 159.600 162.200 160.400 170.000 ;
        RECT 162.800 162.200 163.600 170.200 ;
        RECT 164.400 169.600 168.400 170.200 ;
        RECT 164.400 162.200 165.200 169.600 ;
        RECT 167.600 162.200 168.400 169.600 ;
        RECT 170.800 162.200 171.600 173.700 ;
        RECT 175.600 173.800 176.600 174.200 ;
        RECT 177.600 174.400 178.200 175.000 ;
        RECT 182.000 175.200 182.800 179.800 ;
        RECT 182.000 174.600 184.200 175.200 ;
        RECT 172.400 171.600 173.200 173.200 ;
        RECT 174.000 171.600 174.800 173.200 ;
        RECT 175.600 173.000 177.000 173.800 ;
        RECT 177.600 173.600 179.600 174.400 ;
        RECT 175.600 171.000 176.200 173.000 ;
        RECT 172.400 170.400 176.200 171.000 ;
        RECT 172.400 167.000 173.000 170.400 ;
        RECT 177.600 169.800 178.200 173.600 ;
        RECT 178.800 170.800 179.600 172.400 ;
        RECT 182.000 171.600 182.800 173.200 ;
        RECT 183.600 171.600 184.200 174.600 ;
        RECT 183.600 170.800 184.800 171.600 ;
        RECT 183.600 170.200 184.200 170.800 ;
        RECT 176.600 169.200 178.200 169.800 ;
        RECT 182.000 169.600 184.200 170.200 ;
        RECT 172.400 163.000 173.200 167.000 ;
        RECT 176.600 162.200 177.400 169.200 ;
        RECT 182.000 162.200 182.800 169.600 ;
        RECT 186.800 162.200 187.600 179.800 ;
        RECT 188.400 176.300 189.200 177.200 ;
        RECT 190.000 176.300 190.800 176.400 ;
        RECT 188.400 175.700 190.800 176.300 ;
        RECT 188.400 175.600 189.200 175.700 ;
        RECT 190.000 175.600 190.800 175.700 ;
        RECT 191.600 173.800 192.400 179.800 ;
        RECT 198.000 176.600 198.800 179.800 ;
        RECT 199.600 177.000 200.400 179.800 ;
        RECT 201.200 177.000 202.000 179.800 ;
        RECT 202.800 177.000 203.600 179.800 ;
        RECT 206.000 177.000 206.800 179.800 ;
        RECT 209.200 177.000 210.000 179.800 ;
        RECT 210.800 177.000 211.600 179.800 ;
        RECT 212.400 177.000 213.200 179.800 ;
        RECT 214.000 177.000 214.800 179.800 ;
        RECT 196.200 175.800 198.800 176.600 ;
        RECT 215.600 176.600 216.400 179.800 ;
        RECT 202.200 175.800 206.800 176.400 ;
        RECT 196.200 175.200 197.000 175.800 ;
        RECT 194.000 174.400 197.000 175.200 ;
        RECT 191.600 173.000 200.400 173.800 ;
        RECT 202.200 173.400 203.000 175.800 ;
        RECT 206.000 175.600 206.800 175.800 ;
        RECT 207.600 175.600 209.200 176.400 ;
        RECT 212.200 175.600 213.200 176.400 ;
        RECT 215.600 175.800 218.000 176.600 ;
        RECT 204.400 173.600 205.200 175.200 ;
        RECT 206.000 174.800 206.800 175.000 ;
        RECT 206.000 174.200 210.400 174.800 ;
        RECT 209.600 174.000 210.400 174.200 ;
        RECT 191.600 167.400 192.400 173.000 ;
        RECT 201.000 172.600 203.000 173.400 ;
        RECT 206.800 172.600 210.000 173.400 ;
        RECT 212.400 172.800 213.200 175.600 ;
        RECT 217.200 175.200 218.000 175.800 ;
        RECT 217.200 174.600 219.000 175.200 ;
        RECT 218.200 173.400 219.000 174.600 ;
        RECT 222.000 174.600 222.800 179.800 ;
        RECT 223.600 176.000 224.400 179.800 ;
        RECT 223.600 175.200 224.600 176.000 ;
        RECT 222.000 174.000 223.200 174.600 ;
        RECT 218.200 172.600 222.000 173.400 ;
        RECT 193.000 172.000 193.800 172.200 ;
        RECT 198.000 172.000 198.800 172.400 ;
        RECT 215.600 172.000 216.400 172.600 ;
        RECT 222.600 172.000 223.200 174.000 ;
        RECT 193.000 171.400 216.400 172.000 ;
        RECT 222.400 171.400 223.200 172.000 ;
        RECT 222.400 169.600 223.000 171.400 ;
        RECT 223.800 170.800 224.600 175.200 ;
        RECT 201.200 169.400 202.000 169.600 ;
        RECT 196.600 169.000 202.000 169.400 ;
        RECT 195.800 168.800 202.000 169.000 ;
        RECT 203.000 169.000 211.600 169.600 ;
        RECT 193.200 168.000 194.800 168.800 ;
        RECT 195.800 168.200 197.200 168.800 ;
        RECT 203.000 168.200 203.600 169.000 ;
        RECT 210.800 168.800 211.600 169.000 ;
        RECT 214.000 169.000 223.000 169.600 ;
        RECT 214.000 168.800 214.800 169.000 ;
        RECT 194.200 167.600 194.800 168.000 ;
        RECT 197.800 167.600 203.600 168.200 ;
        RECT 204.200 167.600 206.800 168.400 ;
        RECT 191.600 166.800 193.600 167.400 ;
        RECT 194.200 166.800 198.400 167.600 ;
        RECT 193.000 166.200 193.600 166.800 ;
        RECT 193.000 165.600 194.000 166.200 ;
        RECT 193.200 162.200 194.000 165.600 ;
        RECT 196.400 162.200 197.200 166.800 ;
        RECT 199.600 162.200 200.400 165.000 ;
        RECT 201.200 162.200 202.000 165.000 ;
        RECT 202.800 162.200 203.600 167.000 ;
        RECT 206.000 162.200 206.800 167.000 ;
        RECT 209.200 162.200 210.000 168.400 ;
        RECT 217.200 167.600 219.800 168.400 ;
        RECT 212.400 166.800 216.600 167.600 ;
        RECT 210.800 162.200 211.600 165.000 ;
        RECT 212.400 162.200 213.200 165.000 ;
        RECT 214.000 162.200 214.800 165.000 ;
        RECT 217.200 162.200 218.000 167.600 ;
        RECT 222.400 167.400 223.000 169.000 ;
        RECT 220.400 166.800 223.000 167.400 ;
        RECT 223.600 170.000 224.600 170.800 ;
        RECT 220.400 162.200 221.200 166.800 ;
        RECT 223.600 162.200 224.400 170.000 ;
        RECT 4.400 152.400 5.200 159.800 ;
        RECT 3.000 151.800 5.200 152.400 ;
        RECT 6.600 152.600 7.400 159.800 ;
        RECT 13.400 158.400 14.200 159.800 ;
        RECT 12.400 157.600 14.200 158.400 ;
        RECT 6.600 151.800 8.400 152.600 ;
        RECT 13.400 152.400 14.200 157.600 ;
        RECT 18.800 156.400 19.600 159.800 ;
        RECT 18.600 155.800 19.600 156.400 ;
        RECT 18.600 155.200 19.200 155.800 ;
        RECT 22.000 155.200 22.800 159.800 ;
        RECT 25.200 157.000 26.000 159.800 ;
        RECT 26.800 157.000 27.600 159.800 ;
        RECT 17.200 154.600 19.200 155.200 ;
        RECT 14.800 153.600 15.600 154.400 ;
        RECT 15.000 152.400 15.600 153.600 ;
        RECT 13.400 151.800 14.400 152.400 ;
        RECT 15.000 151.800 16.400 152.400 ;
        RECT 3.000 151.200 3.600 151.800 ;
        RECT 2.400 150.400 3.600 151.200 ;
        RECT 3.000 147.400 3.600 150.400 ;
        RECT 4.400 148.800 5.200 150.400 ;
        RECT 6.000 149.600 6.800 151.200 ;
        RECT 7.600 148.400 8.200 151.800 ;
        RECT 12.400 148.800 13.200 150.400 ;
        RECT 13.800 148.400 14.400 151.800 ;
        RECT 15.600 151.600 16.400 151.800 ;
        RECT 17.200 149.000 18.000 154.600 ;
        RECT 19.800 154.400 24.000 155.200 ;
        RECT 28.400 155.000 29.200 159.800 ;
        RECT 31.600 155.000 32.400 159.800 ;
        RECT 19.800 154.000 20.400 154.400 ;
        RECT 18.800 153.200 20.400 154.000 ;
        RECT 23.400 153.800 29.200 154.400 ;
        RECT 21.400 153.200 22.800 153.800 ;
        RECT 21.400 153.000 27.600 153.200 ;
        RECT 22.200 152.600 27.600 153.000 ;
        RECT 26.800 152.400 27.600 152.600 ;
        RECT 28.600 153.000 29.200 153.800 ;
        RECT 29.800 153.600 32.400 154.400 ;
        RECT 34.800 153.600 35.600 159.800 ;
        RECT 36.400 157.000 37.200 159.800 ;
        RECT 38.000 157.000 38.800 159.800 ;
        RECT 39.600 157.000 40.400 159.800 ;
        RECT 38.000 154.400 42.200 155.200 ;
        RECT 42.800 154.400 43.600 159.800 ;
        RECT 46.000 155.200 46.800 159.800 ;
        RECT 46.000 154.600 48.600 155.200 ;
        RECT 42.800 153.600 45.400 154.400 ;
        RECT 36.400 153.000 37.200 153.200 ;
        RECT 28.600 152.400 37.200 153.000 ;
        RECT 39.600 153.000 40.400 153.200 ;
        RECT 48.000 153.000 48.600 154.600 ;
        RECT 39.600 152.400 48.600 153.000 ;
        RECT 48.000 150.600 48.600 152.400 ;
        RECT 49.200 152.000 50.000 159.800 ;
        RECT 54.800 153.600 55.600 154.400 ;
        RECT 54.800 152.400 55.400 153.600 ;
        RECT 56.200 152.400 57.000 159.800 ;
        RECT 49.200 151.200 50.200 152.000 ;
        RECT 54.000 151.800 55.400 152.400 ;
        RECT 56.000 151.800 57.000 152.400 ;
        RECT 60.400 151.800 61.200 159.800 ;
        RECT 63.600 155.800 64.400 159.800 ;
        RECT 54.000 151.600 54.800 151.800 ;
        RECT 18.600 150.000 42.000 150.600 ;
        RECT 48.000 150.000 48.800 150.600 ;
        RECT 18.600 149.800 19.400 150.000 ;
        RECT 23.600 149.600 24.400 150.000 ;
        RECT 41.200 149.400 42.000 150.000 ;
        RECT 7.600 148.300 8.400 148.400 ;
        RECT 10.800 148.300 11.600 148.400 ;
        RECT 7.600 148.200 11.600 148.300 ;
        RECT 7.600 147.700 12.400 148.200 ;
        RECT 7.600 147.600 8.400 147.700 ;
        RECT 10.800 147.600 12.400 147.700 ;
        RECT 13.800 147.600 16.400 148.400 ;
        RECT 17.200 148.200 26.000 149.000 ;
        RECT 26.600 148.600 28.600 149.400 ;
        RECT 32.400 148.600 35.600 149.400 ;
        RECT 3.000 146.800 5.200 147.400 ;
        RECT 4.400 142.200 5.200 146.800 ;
        RECT 7.600 144.200 8.200 147.600 ;
        RECT 11.600 147.200 12.400 147.600 ;
        RECT 9.200 144.800 10.000 146.400 ;
        RECT 11.000 146.200 14.600 146.600 ;
        RECT 15.600 146.200 16.200 147.600 ;
        RECT 10.800 146.000 14.800 146.200 ;
        RECT 7.600 142.200 8.400 144.200 ;
        RECT 10.800 142.200 11.600 146.000 ;
        RECT 14.000 142.200 14.800 146.000 ;
        RECT 15.600 142.200 16.400 146.200 ;
        RECT 17.200 142.200 18.000 148.200 ;
        RECT 19.600 146.800 22.600 147.600 ;
        RECT 21.800 146.200 22.600 146.800 ;
        RECT 27.800 146.200 28.600 148.600 ;
        RECT 30.000 146.800 30.800 148.400 ;
        RECT 35.200 147.800 36.000 148.000 ;
        RECT 31.600 147.200 36.000 147.800 ;
        RECT 31.600 147.000 32.400 147.200 ;
        RECT 38.000 146.400 38.800 149.200 ;
        RECT 43.800 148.600 47.600 149.400 ;
        RECT 43.800 147.400 44.600 148.600 ;
        RECT 48.200 148.000 48.800 150.000 ;
        RECT 31.600 146.200 32.400 146.400 ;
        RECT 21.800 145.400 24.400 146.200 ;
        RECT 27.800 145.600 32.400 146.200 ;
        RECT 33.200 145.600 34.800 146.400 ;
        RECT 37.800 145.600 38.800 146.400 ;
        RECT 42.800 146.800 44.600 147.400 ;
        RECT 47.600 147.400 48.800 148.000 ;
        RECT 42.800 146.200 43.600 146.800 ;
        RECT 23.600 142.200 24.400 145.400 ;
        RECT 41.200 145.400 43.600 146.200 ;
        RECT 25.200 142.200 26.000 145.000 ;
        RECT 26.800 142.200 27.600 145.000 ;
        RECT 28.400 142.200 29.200 145.000 ;
        RECT 31.600 142.200 32.400 145.000 ;
        RECT 34.800 142.200 35.600 145.000 ;
        RECT 36.400 142.200 37.200 145.000 ;
        RECT 38.000 142.200 38.800 145.000 ;
        RECT 39.600 142.200 40.400 145.000 ;
        RECT 41.200 142.200 42.000 145.400 ;
        RECT 47.600 142.200 48.400 147.400 ;
        RECT 49.400 146.800 50.200 151.200 ;
        RECT 56.000 148.400 56.600 151.800 ;
        RECT 60.400 150.400 61.000 151.800 ;
        RECT 63.600 151.600 64.200 155.800 ;
        RECT 69.400 152.600 70.200 159.800 ;
        RECT 74.800 156.400 75.600 159.800 ;
        RECT 74.600 155.800 75.600 156.400 ;
        RECT 74.600 155.200 75.200 155.800 ;
        RECT 78.000 155.200 78.800 159.800 ;
        RECT 81.200 157.000 82.000 159.800 ;
        RECT 82.800 157.000 83.600 159.800 ;
        RECT 68.400 151.800 70.200 152.600 ;
        RECT 73.200 154.600 75.200 155.200 ;
        RECT 61.800 151.000 64.200 151.600 ;
        RECT 57.200 150.300 58.000 150.400 ;
        RECT 60.400 150.300 61.200 150.400 ;
        RECT 57.200 149.700 61.200 150.300 ;
        RECT 57.200 148.800 58.000 149.700 ;
        RECT 60.400 149.600 61.200 149.700 ;
        RECT 54.000 147.600 56.600 148.400 ;
        RECT 58.800 148.200 59.600 148.400 ;
        RECT 58.000 147.600 59.600 148.200 ;
        RECT 49.200 146.000 50.200 146.800 ;
        RECT 54.200 146.200 54.800 147.600 ;
        RECT 58.000 147.200 58.800 147.600 ;
        RECT 55.800 146.200 59.400 146.600 ;
        RECT 60.400 146.200 61.000 149.600 ;
        RECT 61.800 147.600 62.400 151.000 ;
        RECT 63.600 149.600 64.400 150.400 ;
        RECT 63.600 148.800 64.200 149.600 ;
        RECT 63.200 148.000 64.400 148.800 ;
        RECT 65.200 148.300 66.000 149.200 ;
        RECT 68.600 148.400 69.200 151.800 ;
        RECT 70.000 150.300 70.800 151.200 ;
        RECT 71.600 150.300 72.400 150.400 ;
        RECT 70.000 149.700 72.400 150.300 ;
        RECT 70.000 149.600 70.800 149.700 ;
        RECT 71.600 149.600 72.400 149.700 ;
        RECT 66.800 148.300 67.600 148.400 ;
        RECT 65.200 147.700 67.600 148.300 ;
        RECT 65.200 147.600 66.000 147.700 ;
        RECT 66.800 147.600 67.600 147.700 ;
        RECT 68.400 147.600 69.200 148.400 ;
        RECT 61.600 147.400 62.400 147.600 ;
        RECT 61.600 147.000 64.600 147.400 ;
        RECT 61.600 146.800 65.800 147.000 ;
        RECT 64.000 146.400 65.800 146.800 ;
        RECT 65.200 146.200 65.800 146.400 ;
        RECT 49.200 142.200 50.000 146.000 ;
        RECT 54.000 142.200 54.800 146.200 ;
        RECT 55.600 146.000 59.600 146.200 ;
        RECT 55.600 142.200 56.400 146.000 ;
        RECT 58.800 142.200 59.600 146.000 ;
        RECT 60.400 145.200 61.800 146.200 ;
        RECT 61.000 142.200 61.800 145.200 ;
        RECT 65.200 142.200 66.000 146.200 ;
        RECT 66.800 144.800 67.600 146.400 ;
        RECT 68.600 144.400 69.200 147.600 ;
        RECT 68.400 142.200 69.200 144.400 ;
        RECT 73.200 149.000 74.000 154.600 ;
        RECT 75.800 154.400 80.000 155.200 ;
        RECT 84.400 155.000 85.200 159.800 ;
        RECT 87.600 155.000 88.400 159.800 ;
        RECT 75.800 154.000 76.400 154.400 ;
        RECT 74.800 153.200 76.400 154.000 ;
        RECT 79.400 153.800 85.200 154.400 ;
        RECT 77.400 153.200 78.800 153.800 ;
        RECT 77.400 153.000 83.600 153.200 ;
        RECT 78.200 152.600 83.600 153.000 ;
        RECT 82.800 152.400 83.600 152.600 ;
        RECT 84.600 153.000 85.200 153.800 ;
        RECT 85.800 153.600 88.400 154.400 ;
        RECT 90.800 153.600 91.600 159.800 ;
        RECT 92.400 157.000 93.200 159.800 ;
        RECT 94.000 157.000 94.800 159.800 ;
        RECT 95.600 157.000 96.400 159.800 ;
        RECT 94.000 154.400 98.200 155.200 ;
        RECT 98.800 154.400 99.600 159.800 ;
        RECT 102.000 155.200 102.800 159.800 ;
        RECT 102.000 154.600 104.600 155.200 ;
        RECT 98.800 153.600 101.400 154.400 ;
        RECT 92.400 153.000 93.200 153.200 ;
        RECT 84.600 152.400 93.200 153.000 ;
        RECT 95.600 153.000 96.400 153.200 ;
        RECT 104.000 153.000 104.600 154.600 ;
        RECT 95.600 152.400 104.600 153.000 ;
        RECT 104.000 150.600 104.600 152.400 ;
        RECT 105.200 152.000 106.000 159.800 ;
        RECT 105.200 151.200 106.200 152.000 ;
        RECT 74.600 150.000 98.000 150.600 ;
        RECT 104.000 150.000 104.800 150.600 ;
        RECT 74.600 149.800 75.400 150.000 ;
        RECT 78.000 149.600 78.800 150.000 ;
        RECT 79.600 149.600 80.400 150.000 ;
        RECT 97.200 149.400 98.000 150.000 ;
        RECT 73.200 148.200 82.000 149.000 ;
        RECT 82.600 148.600 84.600 149.400 ;
        RECT 88.400 148.600 91.600 149.400 ;
        RECT 73.200 142.200 74.000 148.200 ;
        RECT 75.600 146.800 78.600 147.600 ;
        RECT 77.800 146.200 78.600 146.800 ;
        RECT 83.800 146.200 84.600 148.600 ;
        RECT 86.000 146.800 86.800 148.400 ;
        RECT 91.200 147.800 92.000 148.000 ;
        RECT 87.600 147.200 92.000 147.800 ;
        RECT 87.600 147.000 88.400 147.200 ;
        RECT 94.000 146.400 94.800 149.200 ;
        RECT 99.800 148.600 103.600 149.400 ;
        RECT 99.800 147.400 100.600 148.600 ;
        RECT 104.200 148.000 104.800 150.000 ;
        RECT 87.600 146.200 88.400 146.400 ;
        RECT 77.800 145.400 80.400 146.200 ;
        RECT 83.800 145.600 88.400 146.200 ;
        RECT 89.200 145.600 90.800 146.400 ;
        RECT 93.800 145.600 94.800 146.400 ;
        RECT 98.800 146.800 100.600 147.400 ;
        RECT 103.600 147.400 104.800 148.000 ;
        RECT 98.800 146.200 99.600 146.800 ;
        RECT 79.600 142.200 80.400 145.400 ;
        RECT 97.200 145.400 99.600 146.200 ;
        RECT 81.200 142.200 82.000 145.000 ;
        RECT 82.800 142.200 83.600 145.000 ;
        RECT 84.400 142.200 85.200 145.000 ;
        RECT 87.600 142.200 88.400 145.000 ;
        RECT 90.800 142.200 91.600 145.000 ;
        RECT 92.400 142.200 93.200 145.000 ;
        RECT 94.000 142.200 94.800 145.000 ;
        RECT 95.600 142.200 96.400 145.000 ;
        RECT 97.200 142.200 98.000 145.400 ;
        RECT 103.600 142.200 104.400 147.400 ;
        RECT 105.400 146.800 106.200 151.200 ;
        RECT 110.000 151.200 110.800 159.800 ;
        RECT 113.200 151.200 114.000 159.800 ;
        RECT 116.400 151.200 117.200 159.800 ;
        RECT 119.600 151.200 120.400 159.800 ;
        RECT 126.000 156.400 126.800 159.800 ;
        RECT 125.800 155.800 126.800 156.400 ;
        RECT 125.800 155.200 126.400 155.800 ;
        RECT 129.200 155.200 130.000 159.800 ;
        RECT 132.400 157.000 133.200 159.800 ;
        RECT 134.000 157.000 134.800 159.800 ;
        RECT 124.400 154.600 126.400 155.200 ;
        RECT 110.000 150.400 111.800 151.200 ;
        RECT 113.200 150.400 115.400 151.200 ;
        RECT 116.400 150.400 118.600 151.200 ;
        RECT 119.600 150.400 122.000 151.200 ;
        RECT 111.000 149.000 111.800 150.400 ;
        RECT 114.600 149.000 115.400 150.400 ;
        RECT 117.800 149.000 118.600 150.400 ;
        RECT 111.000 148.200 113.600 149.000 ;
        RECT 114.600 148.200 117.000 149.000 ;
        RECT 117.800 148.200 120.400 149.000 ;
        RECT 111.000 147.600 111.800 148.200 ;
        RECT 114.600 147.600 115.400 148.200 ;
        RECT 117.800 147.600 118.600 148.200 ;
        RECT 121.200 147.600 122.000 150.400 ;
        RECT 105.200 146.000 106.200 146.800 ;
        RECT 110.000 146.800 111.800 147.600 ;
        RECT 113.200 146.800 115.400 147.600 ;
        RECT 116.400 146.800 118.600 147.600 ;
        RECT 119.600 146.800 122.000 147.600 ;
        RECT 124.400 149.000 125.200 154.600 ;
        RECT 127.000 154.400 131.200 155.200 ;
        RECT 135.600 155.000 136.400 159.800 ;
        RECT 138.800 155.000 139.600 159.800 ;
        RECT 127.000 154.000 127.600 154.400 ;
        RECT 126.000 153.200 127.600 154.000 ;
        RECT 130.600 153.800 136.400 154.400 ;
        RECT 128.600 153.200 130.000 153.800 ;
        RECT 128.600 153.000 134.800 153.200 ;
        RECT 129.400 152.600 134.800 153.000 ;
        RECT 134.000 152.400 134.800 152.600 ;
        RECT 135.800 153.000 136.400 153.800 ;
        RECT 137.000 153.600 139.600 154.400 ;
        RECT 142.000 153.600 142.800 159.800 ;
        RECT 143.600 157.000 144.400 159.800 ;
        RECT 145.200 157.000 146.000 159.800 ;
        RECT 146.800 157.000 147.600 159.800 ;
        RECT 145.200 154.400 149.400 155.200 ;
        RECT 150.000 154.400 150.800 159.800 ;
        RECT 153.200 155.200 154.000 159.800 ;
        RECT 153.200 154.600 155.800 155.200 ;
        RECT 150.000 153.600 152.600 154.400 ;
        RECT 143.600 153.000 144.400 153.200 ;
        RECT 135.800 152.400 144.400 153.000 ;
        RECT 146.800 153.000 147.600 153.200 ;
        RECT 155.200 153.000 155.800 154.600 ;
        RECT 146.800 152.400 155.800 153.000 ;
        RECT 155.200 150.600 155.800 152.400 ;
        RECT 156.400 152.000 157.200 159.800 ;
        RECT 159.600 152.400 160.400 159.800 ;
        RECT 161.000 152.400 161.800 152.600 ;
        RECT 156.400 151.200 157.400 152.000 ;
        RECT 159.600 151.800 161.800 152.400 ;
        RECT 164.000 152.400 165.600 159.800 ;
        RECT 167.600 152.400 168.400 152.600 ;
        RECT 169.200 152.400 170.000 159.800 ;
        RECT 164.000 151.800 166.000 152.400 ;
        RECT 167.600 151.800 170.000 152.400 ;
        RECT 170.800 155.000 171.600 159.000 ;
        RECT 125.800 150.000 149.200 150.600 ;
        RECT 155.200 150.000 156.000 150.600 ;
        RECT 125.800 149.800 126.600 150.000 ;
        RECT 127.600 149.600 128.400 150.000 ;
        RECT 129.200 149.600 130.000 150.000 ;
        RECT 130.800 149.600 131.600 150.000 ;
        RECT 148.400 149.400 149.200 150.000 ;
        RECT 124.400 148.200 133.200 149.000 ;
        RECT 133.800 148.600 135.800 149.400 ;
        RECT 139.600 148.600 142.800 149.400 ;
        RECT 105.200 142.200 106.000 146.000 ;
        RECT 110.000 142.200 110.800 146.800 ;
        RECT 113.200 142.200 114.000 146.800 ;
        RECT 116.400 142.200 117.200 146.800 ;
        RECT 119.600 142.200 120.400 146.800 ;
        RECT 124.400 142.200 125.200 148.200 ;
        RECT 126.800 146.800 129.800 147.600 ;
        RECT 129.000 146.200 129.800 146.800 ;
        RECT 135.000 146.200 135.800 148.600 ;
        RECT 137.200 146.800 138.000 148.400 ;
        RECT 142.400 147.800 143.200 148.000 ;
        RECT 138.800 147.200 143.200 147.800 ;
        RECT 138.800 147.000 139.600 147.200 ;
        RECT 145.200 146.400 146.000 149.200 ;
        RECT 151.000 148.600 154.800 149.400 ;
        RECT 151.000 147.400 151.800 148.600 ;
        RECT 155.400 148.000 156.000 150.000 ;
        RECT 138.800 146.200 139.600 146.400 ;
        RECT 129.000 145.400 131.600 146.200 ;
        RECT 135.000 145.600 139.600 146.200 ;
        RECT 140.400 145.600 142.000 146.400 ;
        RECT 145.000 145.600 146.000 146.400 ;
        RECT 150.000 146.800 151.800 147.400 ;
        RECT 154.800 147.400 156.000 148.000 ;
        RECT 156.600 148.300 157.400 151.200 ;
        RECT 161.200 151.200 161.800 151.800 ;
        RECT 161.200 150.600 164.600 151.200 ;
        RECT 163.800 150.400 164.600 150.600 ;
        RECT 165.400 150.400 166.000 151.800 ;
        RECT 170.800 151.600 171.400 155.000 ;
        RECT 175.000 152.800 175.800 159.800 ;
        RECT 175.000 152.200 176.600 152.800 ;
        RECT 170.800 151.000 174.600 151.600 ;
        RECT 161.600 149.800 162.400 150.000 ;
        RECT 165.400 149.800 166.800 150.400 ;
        RECT 161.600 149.200 164.200 149.800 ;
        RECT 163.600 148.600 164.200 149.200 ;
        RECT 165.000 149.600 166.800 149.800 ;
        RECT 165.000 149.200 166.000 149.600 ;
        RECT 159.600 148.300 161.200 148.400 ;
        RECT 156.600 148.200 161.200 148.300 ;
        RECT 156.600 147.700 163.000 148.200 ;
        RECT 163.600 147.800 164.400 148.600 ;
        RECT 150.000 146.200 150.800 146.800 ;
        RECT 130.800 142.200 131.600 145.400 ;
        RECT 148.400 145.400 150.800 146.200 ;
        RECT 132.400 142.200 133.200 145.000 ;
        RECT 134.000 142.200 134.800 145.000 ;
        RECT 135.600 142.200 136.400 145.000 ;
        RECT 138.800 142.200 139.600 145.000 ;
        RECT 142.000 142.200 142.800 145.000 ;
        RECT 143.600 142.200 144.400 145.000 ;
        RECT 145.200 142.200 146.000 145.000 ;
        RECT 146.800 142.200 147.600 145.000 ;
        RECT 148.400 142.200 149.200 145.400 ;
        RECT 154.800 142.200 155.600 147.400 ;
        RECT 156.600 146.800 157.400 147.700 ;
        RECT 159.600 147.600 163.000 147.700 ;
        RECT 162.400 147.200 163.000 147.600 ;
        RECT 161.000 146.800 161.800 147.000 ;
        RECT 156.400 146.300 157.400 146.800 ;
        RECT 158.000 146.300 158.800 146.400 ;
        RECT 156.400 145.700 158.800 146.300 ;
        RECT 156.400 142.200 157.200 145.700 ;
        RECT 158.000 145.600 158.800 145.700 ;
        RECT 159.600 146.200 161.800 146.800 ;
        RECT 162.400 146.600 164.400 147.200 ;
        RECT 162.800 146.400 164.400 146.600 ;
        RECT 159.600 142.200 160.400 146.200 ;
        RECT 165.000 145.800 165.600 149.200 ;
        RECT 170.800 148.800 171.600 150.400 ;
        RECT 172.400 148.800 173.200 150.400 ;
        RECT 174.000 149.000 174.600 151.000 ;
        RECT 166.400 147.600 167.200 148.400 ;
        RECT 168.400 147.600 170.000 148.400 ;
        RECT 174.000 148.200 175.400 149.000 ;
        RECT 176.000 148.400 176.600 152.200 ;
        RECT 177.200 150.300 178.000 151.200 ;
        RECT 180.400 150.300 181.200 159.800 ;
        RECT 186.800 156.400 187.600 159.800 ;
        RECT 186.600 155.800 187.600 156.400 ;
        RECT 186.600 155.200 187.200 155.800 ;
        RECT 190.000 155.200 190.800 159.800 ;
        RECT 193.200 157.000 194.000 159.800 ;
        RECT 194.800 157.000 195.600 159.800 ;
        RECT 177.200 149.700 181.200 150.300 ;
        RECT 177.200 149.600 178.000 149.700 ;
        RECT 176.000 148.300 178.000 148.400 ;
        RECT 178.800 148.300 179.600 148.400 ;
        RECT 174.000 147.800 175.000 148.200 ;
        RECT 166.400 147.200 167.000 147.600 ;
        RECT 166.200 146.400 167.000 147.200 ;
        RECT 170.800 147.200 175.000 147.800 ;
        RECT 176.000 147.700 179.600 148.300 ;
        RECT 176.000 147.600 178.000 147.700 ;
        RECT 178.800 147.600 179.600 147.700 ;
        RECT 167.600 146.800 168.400 147.000 ;
        RECT 167.600 146.200 170.000 146.800 ;
        RECT 164.000 144.400 165.600 145.800 ;
        RECT 162.800 143.600 165.600 144.400 ;
        RECT 164.000 142.200 165.600 143.600 ;
        RECT 169.200 142.200 170.000 146.200 ;
        RECT 170.800 145.000 171.400 147.200 ;
        RECT 176.000 147.000 176.600 147.600 ;
        RECT 175.800 146.600 176.600 147.000 ;
        RECT 175.000 146.000 176.600 146.600 ;
        RECT 170.800 143.000 171.600 145.000 ;
        RECT 175.000 143.000 175.800 146.000 ;
        RECT 180.400 142.200 181.200 149.700 ;
        RECT 185.200 154.600 187.200 155.200 ;
        RECT 185.200 149.000 186.000 154.600 ;
        RECT 187.800 154.400 192.000 155.200 ;
        RECT 196.400 155.000 197.200 159.800 ;
        RECT 199.600 155.000 200.400 159.800 ;
        RECT 187.800 154.000 188.400 154.400 ;
        RECT 186.800 153.200 188.400 154.000 ;
        RECT 191.400 153.800 197.200 154.400 ;
        RECT 189.400 153.200 190.800 153.800 ;
        RECT 189.400 153.000 195.600 153.200 ;
        RECT 190.200 152.600 195.600 153.000 ;
        RECT 194.800 152.400 195.600 152.600 ;
        RECT 196.600 153.000 197.200 153.800 ;
        RECT 197.800 153.600 200.400 154.400 ;
        RECT 202.800 153.600 203.600 159.800 ;
        RECT 204.400 157.000 205.200 159.800 ;
        RECT 206.000 157.000 206.800 159.800 ;
        RECT 207.600 157.000 208.400 159.800 ;
        RECT 206.000 154.400 210.200 155.200 ;
        RECT 210.800 154.400 211.600 159.800 ;
        RECT 214.000 155.200 214.800 159.800 ;
        RECT 214.000 154.600 216.600 155.200 ;
        RECT 210.800 153.600 213.400 154.400 ;
        RECT 204.400 153.000 205.200 153.200 ;
        RECT 196.600 152.400 205.200 153.000 ;
        RECT 207.600 153.000 208.400 153.200 ;
        RECT 216.000 153.000 216.600 154.600 ;
        RECT 207.600 152.400 216.600 153.000 ;
        RECT 216.000 150.600 216.600 152.400 ;
        RECT 217.200 152.000 218.000 159.800 ;
        RECT 220.400 152.400 221.200 159.800 ;
        RECT 217.200 151.200 218.200 152.000 ;
        RECT 220.400 151.800 222.600 152.400 ;
        RECT 186.600 150.000 210.000 150.600 ;
        RECT 216.000 150.000 216.800 150.600 ;
        RECT 186.600 149.800 187.400 150.000 ;
        RECT 191.600 149.600 192.400 150.000 ;
        RECT 198.000 149.600 198.800 150.000 ;
        RECT 209.200 149.400 210.000 150.000 ;
        RECT 185.200 148.200 194.000 149.000 ;
        RECT 194.600 148.600 196.600 149.400 ;
        RECT 200.400 148.600 203.600 149.400 ;
        RECT 182.000 146.300 182.800 146.400 ;
        RECT 183.600 146.300 184.400 146.400 ;
        RECT 182.000 145.700 184.400 146.300 ;
        RECT 182.000 144.800 182.800 145.700 ;
        RECT 183.600 145.600 184.400 145.700 ;
        RECT 185.200 142.200 186.000 148.200 ;
        RECT 187.600 146.800 190.600 147.600 ;
        RECT 189.800 146.200 190.600 146.800 ;
        RECT 195.800 146.200 196.600 148.600 ;
        RECT 198.000 146.800 198.800 148.400 ;
        RECT 203.200 147.800 204.000 148.000 ;
        RECT 199.600 147.200 204.000 147.800 ;
        RECT 199.600 147.000 200.400 147.200 ;
        RECT 206.000 146.400 206.800 149.200 ;
        RECT 211.800 148.600 215.600 149.400 ;
        RECT 211.800 147.400 212.600 148.600 ;
        RECT 216.200 148.000 216.800 150.000 ;
        RECT 199.600 146.200 200.400 146.400 ;
        RECT 189.800 145.400 192.400 146.200 ;
        RECT 195.800 145.600 200.400 146.200 ;
        RECT 201.200 145.600 202.800 146.400 ;
        RECT 205.800 145.600 206.800 146.400 ;
        RECT 210.800 146.800 212.600 147.400 ;
        RECT 215.600 147.400 216.800 148.000 ;
        RECT 217.400 150.300 218.200 151.200 ;
        RECT 222.000 151.200 222.600 151.800 ;
        RECT 222.000 150.400 223.200 151.200 ;
        RECT 220.400 150.300 221.200 150.400 ;
        RECT 217.400 149.700 221.200 150.300 ;
        RECT 210.800 146.200 211.600 146.800 ;
        RECT 191.600 142.200 192.400 145.400 ;
        RECT 209.200 145.400 211.600 146.200 ;
        RECT 193.200 142.200 194.000 145.000 ;
        RECT 194.800 142.200 195.600 145.000 ;
        RECT 196.400 142.200 197.200 145.000 ;
        RECT 199.600 142.200 200.400 145.000 ;
        RECT 202.800 142.200 203.600 145.000 ;
        RECT 204.400 142.200 205.200 145.000 ;
        RECT 206.000 142.200 206.800 145.000 ;
        RECT 207.600 142.200 208.400 145.000 ;
        RECT 209.200 142.200 210.000 145.400 ;
        RECT 215.600 142.200 216.400 147.400 ;
        RECT 217.400 146.800 218.200 149.700 ;
        RECT 220.400 148.800 221.200 149.700 ;
        RECT 222.000 147.400 222.600 150.400 ;
        RECT 217.200 146.000 218.200 146.800 ;
        RECT 220.400 146.800 222.600 147.400 ;
        RECT 217.200 142.200 218.000 146.000 ;
        RECT 220.400 142.200 221.200 146.800 ;
        RECT 1.200 135.800 2.000 139.800 ;
        RECT 2.800 136.000 3.600 139.800 ;
        RECT 6.000 136.000 6.800 139.800 ;
        RECT 2.800 135.800 6.800 136.000 ;
        RECT 1.400 134.400 2.000 135.800 ;
        RECT 3.000 135.400 6.600 135.800 ;
        RECT 7.600 135.600 8.400 137.200 ;
        RECT 5.200 134.400 6.000 134.800 ;
        RECT 1.200 133.600 3.800 134.400 ;
        RECT 5.200 133.800 6.800 134.400 ;
        RECT 6.000 133.600 6.800 133.800 ;
        RECT 9.200 134.300 10.000 139.800 ;
        RECT 14.000 135.800 14.800 139.800 ;
        RECT 15.400 136.400 16.200 137.200 ;
        RECT 12.400 134.300 13.200 134.400 ;
        RECT 9.200 133.700 13.200 134.300 ;
        RECT 3.200 132.400 3.800 133.600 ;
        RECT 2.800 131.600 3.800 132.400 ;
        RECT 4.400 131.600 5.200 133.200 ;
        RECT 1.200 130.200 2.000 130.400 ;
        RECT 3.200 130.200 3.800 131.600 ;
        RECT 1.200 129.600 2.600 130.200 ;
        RECT 3.200 129.600 4.200 130.200 ;
        RECT 2.000 128.400 2.600 129.600 ;
        RECT 2.000 127.600 2.800 128.400 ;
        RECT 3.400 122.200 4.200 129.600 ;
        RECT 9.200 122.200 10.000 133.700 ;
        RECT 12.400 132.800 13.200 133.700 ;
        RECT 14.000 134.300 14.600 135.800 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 19.800 135.800 21.400 139.800 ;
        RECT 28.400 138.400 29.200 139.800 ;
        RECT 28.400 137.800 29.400 138.400 ;
        RECT 28.800 137.600 29.400 137.800 ;
        RECT 31.600 137.800 32.400 139.800 ;
        RECT 31.600 137.600 32.800 137.800 ;
        RECT 28.800 137.000 32.800 137.600 ;
        RECT 25.200 136.300 26.000 136.400 ;
        RECT 26.800 136.300 28.600 136.400 ;
        RECT 18.800 134.300 19.600 134.400 ;
        RECT 14.000 133.700 19.600 134.300 ;
        RECT 10.800 132.200 11.600 132.400 ;
        RECT 14.000 132.200 14.600 133.700 ;
        RECT 18.800 133.600 19.600 133.700 ;
        RECT 19.000 133.200 19.600 133.600 ;
        RECT 19.000 132.400 19.800 133.200 ;
        RECT 20.400 132.400 21.000 135.800 ;
        RECT 25.200 135.700 28.600 136.300 ;
        RECT 25.200 135.600 26.000 135.700 ;
        RECT 26.800 135.600 28.600 135.700 ;
        RECT 22.000 132.800 22.800 134.400 ;
        RECT 28.400 133.600 30.800 134.400 ;
        RECT 15.600 132.200 16.400 132.400 ;
        RECT 10.800 131.600 12.400 132.200 ;
        RECT 14.000 131.600 16.400 132.200 ;
        RECT 11.600 131.200 12.400 131.600 ;
        RECT 15.600 130.200 16.200 131.600 ;
        RECT 17.200 130.800 18.000 132.400 ;
        RECT 20.400 131.600 21.200 132.400 ;
        RECT 23.600 132.200 24.400 132.400 ;
        RECT 22.800 131.600 24.400 132.200 ;
        RECT 30.000 131.600 31.600 132.400 ;
        RECT 20.400 131.400 21.000 131.600 ;
        RECT 19.000 130.800 21.000 131.400 ;
        RECT 22.800 131.200 23.600 131.600 ;
        RECT 19.000 130.200 19.600 130.800 ;
        RECT 32.200 130.400 32.800 137.000 ;
        RECT 39.600 135.600 40.400 137.200 ;
        RECT 41.200 136.300 42.000 139.800 ;
        RECT 44.400 137.600 45.200 139.800 ;
        RECT 42.800 136.300 43.600 137.200 ;
        RECT 41.200 135.700 43.600 136.300 ;
        RECT 41.200 132.300 42.000 135.700 ;
        RECT 42.800 135.600 43.600 135.700 ;
        RECT 44.600 134.400 45.200 137.600 ;
        RECT 44.400 133.600 45.200 134.400 ;
        RECT 51.200 134.200 52.000 139.800 ;
        RECT 57.600 134.200 58.400 139.800 ;
        RECT 51.200 133.800 53.000 134.200 ;
        RECT 57.600 133.800 59.400 134.200 ;
        RECT 51.400 133.600 53.000 133.800 ;
        RECT 57.800 133.600 59.400 133.800 ;
        RECT 42.800 132.300 43.600 132.400 ;
        RECT 41.200 131.700 43.600 132.300 ;
        RECT 10.800 129.600 14.800 130.200 ;
        RECT 10.800 122.200 11.600 129.600 ;
        RECT 14.000 122.200 14.800 129.600 ;
        RECT 15.600 122.200 16.400 130.200 ;
        RECT 17.200 122.800 18.000 130.200 ;
        RECT 18.800 123.400 19.600 130.200 ;
        RECT 20.400 129.600 24.400 130.200 ;
        RECT 32.200 129.800 35.600 130.400 ;
        RECT 20.400 122.800 21.200 129.600 ;
        RECT 17.200 122.200 21.200 122.800 ;
        RECT 23.600 122.200 24.400 129.600 ;
        RECT 34.800 129.600 35.600 129.800 ;
        RECT 25.400 128.800 29.000 129.400 ;
        RECT 25.400 128.200 26.000 128.800 ;
        RECT 25.200 122.200 26.000 128.200 ;
        RECT 28.400 128.200 29.000 128.800 ;
        RECT 30.200 129.000 33.800 129.200 ;
        RECT 34.800 129.000 35.400 129.600 ;
        RECT 30.200 128.600 34.000 129.000 ;
        RECT 30.200 128.200 30.800 128.600 ;
        RECT 28.400 122.800 29.200 128.200 ;
        RECT 30.000 123.400 30.800 128.200 ;
        RECT 31.600 122.800 32.400 128.000 ;
        RECT 33.200 123.000 34.000 128.600 ;
        RECT 34.800 123.400 35.600 129.000 ;
        RECT 28.400 122.200 32.400 122.800 ;
        RECT 33.400 122.800 34.000 123.000 ;
        RECT 36.400 123.000 37.200 129.000 ;
        RECT 36.400 122.800 37.000 123.000 ;
        RECT 33.400 122.200 37.000 122.800 ;
        RECT 41.200 122.200 42.000 131.700 ;
        RECT 42.800 131.600 43.600 131.700 ;
        RECT 44.600 130.200 45.200 133.600 ;
        RECT 46.000 130.800 46.800 132.400 ;
        RECT 49.200 131.600 50.800 132.400 ;
        RECT 44.400 129.400 46.200 130.200 ;
        RECT 47.600 129.600 48.400 131.200 ;
        RECT 52.400 130.400 53.000 133.600 ;
        RECT 55.600 131.600 57.200 132.400 ;
        RECT 52.400 129.600 53.200 130.400 ;
        RECT 54.000 129.600 54.800 131.200 ;
        RECT 58.800 130.400 59.400 133.600 ;
        RECT 58.800 129.600 59.600 130.400 ;
        RECT 45.400 122.200 46.200 129.400 ;
        RECT 50.800 127.600 51.600 129.200 ;
        RECT 52.400 127.000 53.000 129.600 ;
        RECT 55.600 128.300 56.400 128.400 ;
        RECT 57.200 128.300 58.000 129.200 ;
        RECT 55.600 127.700 58.000 128.300 ;
        RECT 55.600 127.600 56.400 127.700 ;
        RECT 57.200 127.600 58.000 127.700 ;
        RECT 58.800 127.000 59.400 129.600 ;
        RECT 49.400 126.400 53.000 127.000 ;
        RECT 49.400 126.200 50.000 126.400 ;
        RECT 49.200 122.200 50.000 126.200 ;
        RECT 52.400 126.200 53.000 126.400 ;
        RECT 55.800 126.400 59.400 127.000 ;
        RECT 55.800 126.200 56.400 126.400 ;
        RECT 52.400 122.200 53.200 126.200 ;
        RECT 55.600 122.200 56.400 126.200 ;
        RECT 58.800 126.200 59.400 126.400 ;
        RECT 58.800 122.200 59.600 126.200 ;
        RECT 60.400 122.200 61.200 139.800 ;
        RECT 62.000 135.600 62.800 137.200 ;
        RECT 66.800 135.200 67.600 139.800 ;
        RECT 70.000 136.000 70.800 139.800 ;
        RECT 65.400 134.600 67.600 135.200 ;
        RECT 69.800 135.200 70.800 136.000 ;
        RECT 65.400 131.600 66.000 134.600 ;
        RECT 66.800 132.300 67.600 133.200 ;
        RECT 69.800 132.300 70.600 135.200 ;
        RECT 71.600 134.600 72.400 139.800 ;
        RECT 78.000 136.600 78.800 139.800 ;
        RECT 79.600 137.000 80.400 139.800 ;
        RECT 81.200 137.000 82.000 139.800 ;
        RECT 82.800 137.000 83.600 139.800 ;
        RECT 84.400 137.000 85.200 139.800 ;
        RECT 87.600 137.000 88.400 139.800 ;
        RECT 90.800 137.000 91.600 139.800 ;
        RECT 92.400 137.000 93.200 139.800 ;
        RECT 94.000 137.000 94.800 139.800 ;
        RECT 76.400 135.800 78.800 136.600 ;
        RECT 95.600 136.600 96.400 139.800 ;
        RECT 76.400 135.200 77.200 135.800 ;
        RECT 66.800 131.700 70.600 132.300 ;
        RECT 66.800 131.600 67.600 131.700 ;
        RECT 64.800 130.800 66.000 131.600 ;
        RECT 65.400 130.200 66.000 130.800 ;
        RECT 69.800 130.800 70.600 131.700 ;
        RECT 71.200 134.000 72.400 134.600 ;
        RECT 75.400 134.600 77.200 135.200 ;
        RECT 81.200 135.600 82.200 136.400 ;
        RECT 85.200 135.600 86.800 136.400 ;
        RECT 87.600 135.800 92.200 136.400 ;
        RECT 95.600 135.800 98.200 136.600 ;
        RECT 87.600 135.600 88.400 135.800 ;
        RECT 71.200 132.000 71.800 134.000 ;
        RECT 75.400 133.400 76.200 134.600 ;
        RECT 72.400 132.600 76.200 133.400 ;
        RECT 81.200 132.800 82.000 135.600 ;
        RECT 87.600 134.800 88.400 135.000 ;
        RECT 84.000 134.200 88.400 134.800 ;
        RECT 84.000 134.000 84.800 134.200 ;
        RECT 89.200 133.600 90.000 135.200 ;
        RECT 91.400 133.400 92.200 135.800 ;
        RECT 97.400 135.200 98.200 135.800 ;
        RECT 97.400 134.400 100.400 135.200 ;
        RECT 102.000 133.800 102.800 139.800 ;
        RECT 106.800 135.200 107.600 139.800 ;
        RECT 110.000 135.200 110.800 139.800 ;
        RECT 113.200 135.200 114.000 139.800 ;
        RECT 116.400 135.200 117.200 139.800 ;
        RECT 84.400 132.600 87.600 133.400 ;
        RECT 91.400 132.600 93.400 133.400 ;
        RECT 94.000 133.000 102.800 133.800 ;
        RECT 78.000 132.000 78.800 132.600 ;
        RECT 95.600 132.000 96.400 132.400 ;
        RECT 100.600 132.000 101.400 132.200 ;
        RECT 71.200 131.400 72.000 132.000 ;
        RECT 78.000 131.400 101.400 132.000 ;
        RECT 65.400 129.600 67.600 130.200 ;
        RECT 69.800 130.000 70.800 130.800 ;
        RECT 66.800 122.200 67.600 129.600 ;
        RECT 70.000 122.200 70.800 130.000 ;
        RECT 71.400 129.600 72.000 131.400 ;
        RECT 71.400 129.000 80.400 129.600 ;
        RECT 71.400 127.400 72.000 129.000 ;
        RECT 79.600 128.800 80.400 129.000 ;
        RECT 82.800 129.000 91.400 129.600 ;
        RECT 82.800 128.800 83.600 129.000 ;
        RECT 74.600 127.600 77.200 128.400 ;
        RECT 71.400 126.800 74.000 127.400 ;
        RECT 73.200 122.200 74.000 126.800 ;
        RECT 76.400 122.200 77.200 127.600 ;
        RECT 77.800 126.800 82.000 127.600 ;
        RECT 79.600 122.200 80.400 125.000 ;
        RECT 81.200 122.200 82.000 125.000 ;
        RECT 82.800 122.200 83.600 125.000 ;
        RECT 84.400 122.200 85.200 128.400 ;
        RECT 87.600 127.600 90.200 128.400 ;
        RECT 90.800 128.200 91.400 129.000 ;
        RECT 92.400 129.400 93.200 129.600 ;
        RECT 92.400 129.000 97.800 129.400 ;
        RECT 92.400 128.800 98.600 129.000 ;
        RECT 97.200 128.200 98.600 128.800 ;
        RECT 90.800 127.600 96.600 128.200 ;
        RECT 99.600 128.000 101.200 128.800 ;
        RECT 99.600 127.600 100.200 128.000 ;
        RECT 87.600 122.200 88.400 127.000 ;
        RECT 90.800 122.200 91.600 127.000 ;
        RECT 96.000 126.800 100.200 127.600 ;
        RECT 102.000 127.400 102.800 133.000 ;
        RECT 105.200 134.400 107.600 135.200 ;
        RECT 108.600 134.400 110.800 135.200 ;
        RECT 111.800 134.400 114.000 135.200 ;
        RECT 115.400 134.400 117.200 135.200 ;
        RECT 121.200 135.200 122.000 139.800 ;
        RECT 124.400 135.200 125.200 139.800 ;
        RECT 127.600 135.200 128.400 139.800 ;
        RECT 130.800 135.200 131.600 139.800 ;
        RECT 134.000 135.200 134.800 139.800 ;
        RECT 137.200 136.400 138.000 139.800 ;
        RECT 137.200 135.800 138.200 136.400 ;
        RECT 121.200 134.400 123.000 135.200 ;
        RECT 124.400 134.400 126.600 135.200 ;
        RECT 127.600 134.400 129.800 135.200 ;
        RECT 130.800 134.400 133.200 135.200 ;
        RECT 134.000 134.600 136.600 135.200 ;
        RECT 105.200 131.600 106.000 134.400 ;
        RECT 108.600 133.800 109.400 134.400 ;
        RECT 111.800 133.800 112.600 134.400 ;
        RECT 115.400 133.800 116.200 134.400 ;
        RECT 106.800 133.000 109.400 133.800 ;
        RECT 110.200 133.000 112.600 133.800 ;
        RECT 113.600 133.000 116.200 133.800 ;
        RECT 108.600 131.600 109.400 133.000 ;
        RECT 111.800 131.600 112.600 133.000 ;
        RECT 115.400 131.600 116.200 133.000 ;
        RECT 122.200 133.800 123.000 134.400 ;
        RECT 125.800 133.800 126.600 134.400 ;
        RECT 129.000 133.800 129.800 134.400 ;
        RECT 122.200 133.000 124.800 133.800 ;
        RECT 125.800 133.000 128.200 133.800 ;
        RECT 129.000 133.000 131.600 133.800 ;
        RECT 122.200 131.600 123.000 133.000 ;
        RECT 125.800 131.600 126.600 133.000 ;
        RECT 129.000 131.600 129.800 133.000 ;
        RECT 132.400 131.600 133.200 134.400 ;
        RECT 134.200 132.400 135.000 133.200 ;
        RECT 134.000 131.600 135.000 132.400 ;
        RECT 136.000 133.000 136.600 134.600 ;
        RECT 137.600 134.400 138.200 135.800 ;
        RECT 145.200 135.800 146.000 139.800 ;
        RECT 146.600 136.400 147.400 137.200 ;
        RECT 137.200 133.600 138.200 134.400 ;
        RECT 136.000 132.200 137.000 133.000 ;
        RECT 105.200 130.800 107.600 131.600 ;
        RECT 108.600 130.800 110.800 131.600 ;
        RECT 111.800 130.800 114.000 131.600 ;
        RECT 115.400 130.800 117.200 131.600 ;
        RECT 100.800 126.800 102.800 127.400 ;
        RECT 92.400 122.200 93.200 125.000 ;
        RECT 94.000 122.200 94.800 125.000 ;
        RECT 97.200 122.200 98.000 126.800 ;
        RECT 100.800 126.200 101.400 126.800 ;
        RECT 100.400 125.600 101.400 126.200 ;
        RECT 100.400 122.200 101.200 125.600 ;
        RECT 106.800 122.200 107.600 130.800 ;
        RECT 110.000 122.200 110.800 130.800 ;
        RECT 113.200 122.200 114.000 130.800 ;
        RECT 116.400 122.200 117.200 130.800 ;
        RECT 121.200 130.800 123.000 131.600 ;
        RECT 124.400 130.800 126.600 131.600 ;
        RECT 127.600 130.800 129.800 131.600 ;
        RECT 130.800 130.800 133.200 131.600 ;
        RECT 121.200 122.200 122.000 130.800 ;
        RECT 124.400 122.200 125.200 130.800 ;
        RECT 127.600 122.200 128.400 130.800 ;
        RECT 130.800 122.200 131.600 130.800 ;
        RECT 136.000 130.200 136.600 132.200 ;
        RECT 137.600 130.200 138.200 133.600 ;
        RECT 143.600 132.800 144.400 134.400 ;
        RECT 142.000 132.200 142.800 132.400 ;
        RECT 145.200 132.200 145.800 135.800 ;
        RECT 146.800 135.600 147.600 136.400 ;
        RECT 146.800 134.300 147.600 134.400 ;
        RECT 148.400 134.300 149.200 139.800 ;
        RECT 150.000 135.600 150.800 137.200 ;
        RECT 151.600 135.800 152.400 139.800 ;
        RECT 153.200 136.000 154.000 139.800 ;
        RECT 156.400 136.000 157.200 139.800 ;
        RECT 153.200 135.800 157.200 136.000 ;
        RECT 158.000 136.000 158.800 139.800 ;
        RECT 161.200 136.000 162.000 139.800 ;
        RECT 158.000 135.800 162.000 136.000 ;
        RECT 151.800 134.400 152.400 135.800 ;
        RECT 153.400 135.400 157.000 135.800 ;
        RECT 158.200 135.400 161.800 135.800 ;
        RECT 162.800 135.600 163.600 139.800 ;
        RECT 164.400 135.800 165.200 139.800 ;
        RECT 166.000 136.000 166.800 139.800 ;
        RECT 169.200 136.000 170.000 139.800 ;
        RECT 171.000 136.400 171.800 137.200 ;
        RECT 166.000 135.800 170.000 136.000 ;
        RECT 155.600 134.400 156.400 134.800 ;
        RECT 158.800 134.400 159.600 134.800 ;
        RECT 162.800 134.400 163.400 135.600 ;
        RECT 164.600 134.400 165.200 135.800 ;
        RECT 166.200 135.400 169.800 135.800 ;
        RECT 170.800 135.600 171.600 136.400 ;
        RECT 172.400 135.600 173.200 139.800 ;
        RECT 168.400 134.400 169.200 134.800 ;
        RECT 146.800 133.700 149.200 134.300 ;
        RECT 146.800 133.600 147.600 133.700 ;
        RECT 146.800 132.200 147.600 132.400 ;
        RECT 142.000 131.600 143.600 132.200 ;
        RECT 145.200 131.600 147.600 132.200 ;
        RECT 142.800 131.200 143.600 131.600 ;
        RECT 146.800 130.200 147.400 131.600 ;
        RECT 134.000 129.600 136.600 130.200 ;
        RECT 134.000 122.200 134.800 129.600 ;
        RECT 137.200 129.200 138.200 130.200 ;
        RECT 142.000 129.600 146.000 130.200 ;
        RECT 137.200 122.200 138.000 129.200 ;
        RECT 142.000 122.200 142.800 129.600 ;
        RECT 145.200 122.200 146.000 129.600 ;
        RECT 146.800 122.200 147.600 130.200 ;
        RECT 148.400 122.200 149.200 133.700 ;
        RECT 150.000 134.300 150.800 134.400 ;
        RECT 151.600 134.300 154.200 134.400 ;
        RECT 150.000 133.700 154.200 134.300 ;
        RECT 155.600 133.800 157.200 134.400 ;
        RECT 150.000 133.600 150.800 133.700 ;
        RECT 151.600 133.600 154.200 133.700 ;
        RECT 156.400 133.600 157.200 133.800 ;
        RECT 158.000 133.800 159.600 134.400 ;
        RECT 158.000 133.600 158.800 133.800 ;
        RECT 161.000 133.600 163.600 134.400 ;
        RECT 164.400 133.600 167.000 134.400 ;
        RECT 168.400 133.800 170.000 134.400 ;
        RECT 169.200 133.600 170.000 133.800 ;
        RECT 151.600 130.200 152.400 130.400 ;
        RECT 153.600 130.200 154.200 133.600 ;
        RECT 154.800 132.300 155.600 133.200 ;
        RECT 159.600 132.300 160.400 133.200 ;
        RECT 154.800 131.700 160.400 132.300 ;
        RECT 154.800 131.600 155.600 131.700 ;
        RECT 159.600 131.600 160.400 131.700 ;
        RECT 161.000 130.200 161.600 133.600 ;
        RECT 162.800 130.300 163.600 130.400 ;
        RECT 164.400 130.300 165.200 130.400 ;
        RECT 162.800 130.200 165.200 130.300 ;
        RECT 166.400 130.200 167.000 133.600 ;
        RECT 167.600 131.600 168.400 133.200 ;
        RECT 170.800 132.200 171.600 132.400 ;
        RECT 172.600 132.200 173.200 135.600 ;
        RECT 174.000 134.300 174.800 134.400 ;
        RECT 177.200 134.300 178.000 139.800 ;
        RECT 178.800 136.300 179.600 137.200 ;
        RECT 182.000 136.300 182.800 136.400 ;
        RECT 183.600 136.300 184.400 139.800 ;
        RECT 178.800 135.700 184.400 136.300 ;
        RECT 178.800 135.600 179.600 135.700 ;
        RECT 182.000 135.600 182.800 135.700 ;
        RECT 174.000 133.700 178.000 134.300 ;
        RECT 174.000 132.800 174.800 133.700 ;
        RECT 175.600 132.200 176.400 132.400 ;
        RECT 170.800 131.600 173.200 132.200 ;
        RECT 174.800 131.600 176.400 132.200 ;
        RECT 171.000 130.200 171.600 131.600 ;
        RECT 174.800 131.200 175.600 131.600 ;
        RECT 151.600 129.600 153.000 130.200 ;
        RECT 153.600 129.600 154.600 130.200 ;
        RECT 152.400 128.400 153.000 129.600 ;
        RECT 152.400 127.600 153.200 128.400 ;
        RECT 153.800 122.200 154.600 129.600 ;
        RECT 160.600 129.600 161.600 130.200 ;
        RECT 162.200 129.700 165.800 130.200 ;
        RECT 162.200 129.600 163.600 129.700 ;
        RECT 164.400 129.600 165.800 129.700 ;
        RECT 166.400 129.600 167.400 130.200 ;
        RECT 160.600 122.200 161.400 129.600 ;
        RECT 162.200 128.400 162.800 129.600 ;
        RECT 162.000 127.600 162.800 128.400 ;
        RECT 165.200 128.400 165.800 129.600 ;
        RECT 165.200 127.600 166.000 128.400 ;
        RECT 166.600 122.200 167.400 129.600 ;
        RECT 170.800 122.200 171.600 130.200 ;
        RECT 172.400 129.600 176.400 130.200 ;
        RECT 172.400 122.200 173.200 129.600 ;
        RECT 175.600 122.200 176.400 129.600 ;
        RECT 177.200 122.200 178.000 133.700 ;
        RECT 183.400 135.200 184.400 135.700 ;
        RECT 183.400 130.800 184.200 135.200 ;
        RECT 185.200 134.600 186.000 139.800 ;
        RECT 191.600 136.600 192.400 139.800 ;
        RECT 193.200 137.000 194.000 139.800 ;
        RECT 194.800 137.000 195.600 139.800 ;
        RECT 196.400 137.000 197.200 139.800 ;
        RECT 198.000 137.000 198.800 139.800 ;
        RECT 201.200 137.000 202.000 139.800 ;
        RECT 204.400 137.000 205.200 139.800 ;
        RECT 206.000 137.000 206.800 139.800 ;
        RECT 207.600 137.000 208.400 139.800 ;
        RECT 190.000 135.800 192.400 136.600 ;
        RECT 209.200 136.600 210.000 139.800 ;
        RECT 190.000 135.200 190.800 135.800 ;
        RECT 184.800 134.000 186.000 134.600 ;
        RECT 189.000 134.600 190.800 135.200 ;
        RECT 194.800 135.600 195.800 136.400 ;
        RECT 198.800 135.600 200.400 136.400 ;
        RECT 201.200 135.800 205.800 136.400 ;
        RECT 209.200 135.800 211.800 136.600 ;
        RECT 201.200 135.600 202.000 135.800 ;
        RECT 184.800 132.000 185.400 134.000 ;
        RECT 189.000 133.400 189.800 134.600 ;
        RECT 186.000 132.600 189.800 133.400 ;
        RECT 194.800 132.800 195.600 135.600 ;
        RECT 201.200 134.800 202.000 135.000 ;
        RECT 197.600 134.200 202.000 134.800 ;
        RECT 197.600 134.000 198.400 134.200 ;
        RECT 202.800 133.600 203.600 135.200 ;
        RECT 205.000 133.400 205.800 135.800 ;
        RECT 211.000 135.200 211.800 135.800 ;
        RECT 211.000 134.400 214.000 135.200 ;
        RECT 215.600 133.800 216.400 139.800 ;
        RECT 217.200 135.200 218.000 139.800 ;
        RECT 217.200 134.600 219.400 135.200 ;
        RECT 198.000 132.600 201.200 133.400 ;
        RECT 205.000 132.600 207.000 133.400 ;
        RECT 207.600 133.000 216.400 133.800 ;
        RECT 191.600 132.000 192.400 132.600 ;
        RECT 202.800 132.000 203.600 132.400 ;
        RECT 209.200 132.000 210.000 132.400 ;
        RECT 214.200 132.000 215.000 132.200 ;
        RECT 184.800 131.400 185.600 132.000 ;
        RECT 191.600 131.400 215.000 132.000 ;
        RECT 183.400 130.000 184.400 130.800 ;
        RECT 183.600 122.200 184.400 130.000 ;
        RECT 185.000 129.600 185.600 131.400 ;
        RECT 185.000 129.000 194.000 129.600 ;
        RECT 185.000 127.400 185.600 129.000 ;
        RECT 193.200 128.800 194.000 129.000 ;
        RECT 196.400 129.000 205.000 129.600 ;
        RECT 196.400 128.800 197.200 129.000 ;
        RECT 188.200 127.600 190.800 128.400 ;
        RECT 185.000 126.800 187.600 127.400 ;
        RECT 186.800 122.200 187.600 126.800 ;
        RECT 190.000 122.200 190.800 127.600 ;
        RECT 191.400 126.800 195.600 127.600 ;
        RECT 193.200 122.200 194.000 125.000 ;
        RECT 194.800 122.200 195.600 125.000 ;
        RECT 196.400 122.200 197.200 125.000 ;
        RECT 198.000 122.200 198.800 128.400 ;
        RECT 201.200 127.600 203.800 128.400 ;
        RECT 204.400 128.200 205.000 129.000 ;
        RECT 206.000 129.400 206.800 129.600 ;
        RECT 206.000 129.000 211.400 129.400 ;
        RECT 206.000 128.800 212.200 129.000 ;
        RECT 210.800 128.200 212.200 128.800 ;
        RECT 204.400 127.600 210.200 128.200 ;
        RECT 213.200 128.000 214.800 128.800 ;
        RECT 213.200 127.600 213.800 128.000 ;
        RECT 201.200 122.200 202.000 127.000 ;
        RECT 204.400 122.200 205.200 127.000 ;
        RECT 209.600 126.800 213.800 127.600 ;
        RECT 215.600 127.400 216.400 133.000 ;
        RECT 217.200 131.600 218.000 133.200 ;
        RECT 218.800 131.600 219.400 134.600 ;
        RECT 218.800 130.800 220.000 131.600 ;
        RECT 218.800 130.200 219.400 130.800 ;
        RECT 214.400 126.800 216.400 127.400 ;
        RECT 217.200 129.600 219.400 130.200 ;
        RECT 206.000 122.200 206.800 125.000 ;
        RECT 207.600 122.200 208.400 125.000 ;
        RECT 210.800 122.200 211.600 126.800 ;
        RECT 214.400 126.200 215.000 126.800 ;
        RECT 214.000 125.600 215.000 126.200 ;
        RECT 214.000 122.200 214.800 125.600 ;
        RECT 217.200 122.200 218.000 129.600 ;
        RECT 4.400 112.400 5.200 119.800 ;
        RECT 3.000 111.800 5.200 112.400 ;
        RECT 7.600 112.000 8.400 119.800 ;
        RECT 10.800 115.200 11.600 119.800 ;
        RECT 3.000 111.200 3.600 111.800 ;
        RECT 2.400 110.400 3.600 111.200 ;
        RECT 7.400 111.200 8.400 112.000 ;
        RECT 9.000 114.600 11.600 115.200 ;
        RECT 9.000 113.000 9.600 114.600 ;
        RECT 14.000 114.400 14.800 119.800 ;
        RECT 17.200 117.000 18.000 119.800 ;
        RECT 18.800 117.000 19.600 119.800 ;
        RECT 20.400 117.000 21.200 119.800 ;
        RECT 15.400 114.400 19.600 115.200 ;
        RECT 12.200 113.600 14.800 114.400 ;
        RECT 22.000 113.600 22.800 119.800 ;
        RECT 25.200 115.000 26.000 119.800 ;
        RECT 28.400 115.000 29.200 119.800 ;
        RECT 30.000 117.000 30.800 119.800 ;
        RECT 31.600 117.000 32.400 119.800 ;
        RECT 34.800 115.200 35.600 119.800 ;
        RECT 38.000 116.400 38.800 119.800 ;
        RECT 38.000 115.800 39.000 116.400 ;
        RECT 38.400 115.200 39.000 115.800 ;
        RECT 33.600 114.400 37.800 115.200 ;
        RECT 38.400 114.600 40.400 115.200 ;
        RECT 25.200 113.600 27.800 114.400 ;
        RECT 28.400 113.800 34.200 114.400 ;
        RECT 37.200 114.000 37.800 114.400 ;
        RECT 17.200 113.000 18.000 113.200 ;
        RECT 9.000 112.400 18.000 113.000 ;
        RECT 20.400 113.000 21.200 113.200 ;
        RECT 28.400 113.000 29.000 113.800 ;
        RECT 34.800 113.200 36.200 113.800 ;
        RECT 37.200 113.200 38.800 114.000 ;
        RECT 20.400 112.400 29.000 113.000 ;
        RECT 30.000 113.000 36.200 113.200 ;
        RECT 30.000 112.600 35.400 113.000 ;
        RECT 30.000 112.400 30.800 112.600 ;
        RECT 3.000 107.400 3.600 110.400 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 7.400 110.300 8.200 111.200 ;
        RECT 9.000 110.600 9.600 112.400 ;
        RECT 4.400 109.700 8.200 110.300 ;
        RECT 4.400 108.800 5.200 109.700 ;
        RECT 3.000 106.800 5.200 107.400 ;
        RECT 4.400 102.200 5.200 106.800 ;
        RECT 7.400 106.800 8.200 109.700 ;
        RECT 8.800 110.000 9.600 110.600 ;
        RECT 15.600 110.000 39.000 110.600 ;
        RECT 8.800 108.000 9.400 110.000 ;
        RECT 15.600 109.400 16.400 110.000 ;
        RECT 33.200 109.600 34.000 110.000 ;
        RECT 36.400 109.600 37.200 110.000 ;
        RECT 38.200 109.800 39.000 110.000 ;
        RECT 10.000 108.600 13.800 109.400 ;
        RECT 8.800 107.400 10.000 108.000 ;
        RECT 7.400 106.000 8.400 106.800 ;
        RECT 7.600 102.200 8.400 106.000 ;
        RECT 9.200 102.200 10.000 107.400 ;
        RECT 13.000 107.400 13.800 108.600 ;
        RECT 13.000 106.800 14.800 107.400 ;
        RECT 14.000 106.200 14.800 106.800 ;
        RECT 18.800 106.400 19.600 109.200 ;
        RECT 22.000 108.600 25.200 109.400 ;
        RECT 29.000 108.600 31.000 109.400 ;
        RECT 39.600 109.000 40.400 114.600 ;
        RECT 21.600 107.800 22.400 108.000 ;
        RECT 21.600 107.200 26.000 107.800 ;
        RECT 25.200 107.000 26.000 107.200 ;
        RECT 26.800 106.800 27.600 108.400 ;
        RECT 14.000 105.400 16.400 106.200 ;
        RECT 18.800 105.600 19.800 106.400 ;
        RECT 22.800 105.600 24.400 106.400 ;
        RECT 25.200 106.200 26.000 106.400 ;
        RECT 29.000 106.200 29.800 108.600 ;
        RECT 31.600 108.200 40.400 109.000 ;
        RECT 35.000 106.800 38.000 107.600 ;
        RECT 35.000 106.200 35.800 106.800 ;
        RECT 25.200 105.600 29.800 106.200 ;
        RECT 15.600 102.200 16.400 105.400 ;
        RECT 33.200 105.400 35.800 106.200 ;
        RECT 17.200 102.200 18.000 105.000 ;
        RECT 18.800 102.200 19.600 105.000 ;
        RECT 20.400 102.200 21.200 105.000 ;
        RECT 22.000 102.200 22.800 105.000 ;
        RECT 25.200 102.200 26.000 105.000 ;
        RECT 28.400 102.200 29.200 105.000 ;
        RECT 30.000 102.200 30.800 105.000 ;
        RECT 31.600 102.200 32.400 105.000 ;
        RECT 33.200 102.200 34.000 105.400 ;
        RECT 39.600 102.200 40.400 108.200 ;
        RECT 42.800 104.800 43.600 106.400 ;
        RECT 44.400 102.200 45.200 119.800 ;
        RECT 46.000 119.200 50.000 119.800 ;
        RECT 46.000 111.800 46.800 119.200 ;
        RECT 47.600 111.800 48.400 118.600 ;
        RECT 49.200 112.400 50.000 119.200 ;
        RECT 52.400 112.400 53.200 119.800 ;
        RECT 56.600 112.600 57.400 119.800 ;
        RECT 49.200 111.800 53.200 112.400 ;
        RECT 55.600 111.800 57.400 112.600 ;
        RECT 47.800 111.200 48.400 111.800 ;
        RECT 46.000 109.600 46.800 111.200 ;
        RECT 47.800 110.600 49.800 111.200 ;
        RECT 49.200 110.400 49.800 110.600 ;
        RECT 51.600 110.400 52.400 110.800 ;
        RECT 49.200 109.600 50.000 110.400 ;
        RECT 51.600 109.800 53.200 110.400 ;
        RECT 52.400 109.600 53.200 109.800 ;
        RECT 47.800 108.800 48.600 109.600 ;
        RECT 47.800 108.400 48.400 108.800 ;
        RECT 47.600 107.600 48.400 108.400 ;
        RECT 49.200 106.200 49.800 109.600 ;
        RECT 50.800 108.300 51.600 109.200 ;
        RECT 55.800 108.400 56.400 111.800 ;
        RECT 58.800 111.600 59.600 113.200 ;
        RECT 57.200 110.300 58.000 111.200 ;
        RECT 60.400 110.300 61.200 119.800 ;
        RECT 63.600 115.800 64.400 119.800 ;
        RECT 63.800 115.600 64.400 115.800 ;
        RECT 66.800 115.800 67.600 119.800 ;
        RECT 71.600 115.800 72.400 119.800 ;
        RECT 66.800 115.600 67.400 115.800 ;
        RECT 63.800 115.000 67.400 115.600 ;
        RECT 71.800 115.600 72.400 115.800 ;
        RECT 74.800 115.800 75.600 119.800 ;
        RECT 74.800 115.600 75.400 115.800 ;
        RECT 71.800 115.000 75.400 115.600 ;
        RECT 63.800 112.400 64.400 115.000 ;
        RECT 65.200 112.800 66.000 114.400 ;
        RECT 66.800 114.300 67.600 114.400 ;
        RECT 73.200 114.300 74.000 114.400 ;
        RECT 66.800 113.700 74.000 114.300 ;
        RECT 66.800 113.600 67.600 113.700 ;
        RECT 73.200 112.800 74.000 113.700 ;
        RECT 74.800 112.400 75.400 115.000 ;
        RECT 63.600 111.600 64.400 112.400 ;
        RECT 57.200 109.700 61.200 110.300 ;
        RECT 57.200 109.600 58.000 109.700 ;
        RECT 55.600 108.300 56.400 108.400 ;
        RECT 50.800 107.700 56.400 108.300 ;
        RECT 50.800 107.600 51.600 107.700 ;
        RECT 55.600 107.600 56.400 107.700 ;
        RECT 48.600 102.200 50.200 106.200 ;
        RECT 54.000 104.800 54.800 106.400 ;
        RECT 55.800 106.300 56.400 107.600 ;
        RECT 57.200 106.300 58.000 106.400 ;
        RECT 55.700 105.700 58.000 106.300 ;
        RECT 60.400 106.200 61.200 109.700 ;
        RECT 63.800 108.400 64.400 111.600 ;
        RECT 68.400 110.800 69.200 112.400 ;
        RECT 70.000 110.800 70.800 112.400 ;
        RECT 74.800 111.600 75.600 112.400 ;
        RECT 66.000 109.600 67.600 110.400 ;
        RECT 71.600 109.600 73.200 110.400 ;
        RECT 74.800 108.400 75.400 111.600 ;
        RECT 76.400 110.300 77.200 110.400 ;
        RECT 78.000 110.300 78.800 119.800 ;
        RECT 82.800 112.800 83.600 119.800 ;
        RECT 76.400 109.700 78.800 110.300 ;
        RECT 76.400 109.600 77.200 109.700 ;
        RECT 62.000 106.800 62.800 108.400 ;
        RECT 63.800 108.200 65.400 108.400 ;
        RECT 73.800 108.200 75.400 108.400 ;
        RECT 63.800 107.800 65.600 108.200 ;
        RECT 55.800 104.200 56.400 105.700 ;
        RECT 57.200 105.600 58.000 105.700 ;
        RECT 59.400 105.600 61.200 106.200 ;
        RECT 55.600 102.200 56.400 104.200 ;
        RECT 59.400 102.200 60.200 105.600 ;
        RECT 64.800 104.400 65.600 107.800 ;
        RECT 73.600 107.800 75.400 108.200 ;
        RECT 64.800 103.600 66.000 104.400 ;
        RECT 64.800 102.200 65.600 103.600 ;
        RECT 73.600 102.200 74.400 107.800 ;
        RECT 76.400 106.800 77.200 108.400 ;
        RECT 78.000 102.200 78.800 109.700 ;
        RECT 82.600 111.800 83.600 112.800 ;
        RECT 86.000 112.400 86.800 119.800 ;
        RECT 84.200 111.800 86.800 112.400 ;
        RECT 82.600 108.400 83.200 111.800 ;
        RECT 84.200 109.800 84.800 111.800 ;
        RECT 90.800 111.200 91.600 119.800 ;
        RECT 94.000 111.200 94.800 119.800 ;
        RECT 98.800 112.800 99.600 119.800 ;
        RECT 90.800 110.400 94.800 111.200 ;
        RECT 98.600 111.800 99.600 112.800 ;
        RECT 102.000 112.400 102.800 119.800 ;
        RECT 100.200 111.800 102.800 112.400 ;
        RECT 83.800 109.000 84.800 109.800 ;
        RECT 82.600 107.600 83.600 108.400 ;
        RECT 82.600 106.200 83.200 107.600 ;
        RECT 84.200 107.400 84.800 109.000 ;
        RECT 85.800 109.600 86.800 110.400 ;
        RECT 85.800 108.800 86.600 109.600 ;
        RECT 90.800 107.600 91.600 110.400 ;
        RECT 98.600 108.400 99.200 111.800 ;
        RECT 100.200 109.800 100.800 111.800 ;
        RECT 99.800 109.000 100.800 109.800 ;
        RECT 84.200 106.800 86.800 107.400 ;
        RECT 82.600 105.600 83.600 106.200 ;
        RECT 82.800 102.200 83.600 105.600 ;
        RECT 86.000 102.200 86.800 106.800 ;
        RECT 90.800 106.800 94.800 107.600 ;
        RECT 95.600 106.800 96.400 108.400 ;
        RECT 98.600 107.600 99.600 108.400 ;
        RECT 90.800 102.200 91.600 106.800 ;
        RECT 94.000 102.200 94.800 106.800 ;
        RECT 98.600 106.200 99.200 107.600 ;
        RECT 100.200 107.400 100.800 109.000 ;
        RECT 101.800 109.600 102.800 110.400 ;
        RECT 101.800 108.800 102.600 109.600 ;
        RECT 100.200 106.800 102.800 107.400 ;
        RECT 98.600 105.600 99.600 106.200 ;
        RECT 98.800 102.200 99.600 105.600 ;
        RECT 102.000 102.200 102.800 106.800 ;
        RECT 103.600 104.800 104.400 106.400 ;
        RECT 105.200 102.200 106.000 119.800 ;
        RECT 106.800 112.400 107.600 119.800 ;
        RECT 110.000 112.800 110.800 119.800 ;
        RECT 117.000 112.800 117.800 119.800 ;
        RECT 121.200 115.000 122.000 119.000 ;
        RECT 106.800 111.800 109.400 112.400 ;
        RECT 110.000 111.800 111.000 112.800 ;
        RECT 106.800 109.600 107.800 110.400 ;
        RECT 107.000 108.800 107.800 109.600 ;
        RECT 108.800 109.800 109.400 111.800 ;
        RECT 108.800 109.000 109.800 109.800 ;
        RECT 108.800 107.400 109.400 109.000 ;
        RECT 110.400 108.400 111.000 111.800 ;
        RECT 116.200 112.200 117.800 112.800 ;
        RECT 114.800 109.600 115.600 111.200 ;
        RECT 116.200 108.400 116.800 112.200 ;
        RECT 121.400 111.600 122.000 115.000 ;
        RECT 122.800 112.400 123.600 119.800 ;
        RECT 126.000 112.800 126.800 119.800 ;
        RECT 122.800 111.800 125.400 112.400 ;
        RECT 126.000 111.800 127.000 112.800 ;
        RECT 129.200 112.400 130.000 119.800 ;
        RECT 132.400 112.800 133.200 119.800 ;
        RECT 138.800 116.400 139.600 119.800 ;
        RECT 138.600 115.800 139.600 116.400 ;
        RECT 138.600 115.200 139.200 115.800 ;
        RECT 142.000 115.200 142.800 119.800 ;
        RECT 145.200 117.000 146.000 119.800 ;
        RECT 146.800 117.000 147.600 119.800 ;
        RECT 137.200 114.600 139.200 115.200 ;
        RECT 129.200 111.800 131.800 112.400 ;
        RECT 132.400 111.800 133.400 112.800 ;
        RECT 118.200 111.000 122.000 111.600 ;
        RECT 118.200 109.000 118.800 111.000 ;
        RECT 110.000 108.300 111.000 108.400 ;
        RECT 113.200 108.300 114.000 108.400 ;
        RECT 110.000 107.700 114.000 108.300 ;
        RECT 110.000 107.600 111.000 107.700 ;
        RECT 113.200 107.600 114.000 107.700 ;
        RECT 114.800 107.600 116.800 108.400 ;
        RECT 117.400 108.200 118.800 109.000 ;
        RECT 119.600 108.800 120.400 110.400 ;
        RECT 121.200 108.800 122.000 110.400 ;
        RECT 122.800 109.600 123.800 110.400 ;
        RECT 123.000 108.800 123.800 109.600 ;
        RECT 124.800 109.800 125.400 111.800 ;
        RECT 124.800 109.000 125.800 109.800 ;
        RECT 106.800 106.800 109.400 107.400 ;
        RECT 106.800 102.200 107.600 106.800 ;
        RECT 110.400 106.200 111.000 107.600 ;
        RECT 110.000 105.600 111.000 106.200 ;
        RECT 116.200 107.000 116.800 107.600 ;
        RECT 117.800 107.800 118.800 108.200 ;
        RECT 117.800 107.200 122.000 107.800 ;
        RECT 124.800 107.400 125.400 109.000 ;
        RECT 126.400 108.400 127.000 111.800 ;
        RECT 127.600 110.300 128.400 110.400 ;
        RECT 129.200 110.300 130.200 110.400 ;
        RECT 127.600 109.700 130.200 110.300 ;
        RECT 127.600 109.600 128.400 109.700 ;
        RECT 129.200 109.600 130.200 109.700 ;
        RECT 129.400 108.800 130.200 109.600 ;
        RECT 131.200 109.800 131.800 111.800 ;
        RECT 131.200 109.000 132.200 109.800 ;
        RECT 126.000 107.600 127.000 108.400 ;
        RECT 116.200 106.600 117.000 107.000 ;
        RECT 116.200 106.000 117.800 106.600 ;
        RECT 110.000 102.200 110.800 105.600 ;
        RECT 117.000 104.400 117.800 106.000 ;
        RECT 121.400 105.000 122.000 107.200 ;
        RECT 117.000 103.600 118.800 104.400 ;
        RECT 117.000 103.000 117.800 103.600 ;
        RECT 121.200 103.000 122.000 105.000 ;
        RECT 122.800 106.800 125.400 107.400 ;
        RECT 122.800 102.200 123.600 106.800 ;
        RECT 126.400 106.200 127.000 107.600 ;
        RECT 131.200 107.400 131.800 109.000 ;
        RECT 132.800 108.400 133.400 111.800 ;
        RECT 132.400 107.600 133.400 108.400 ;
        RECT 126.000 105.600 127.000 106.200 ;
        RECT 129.200 106.800 131.800 107.400 ;
        RECT 126.000 102.200 126.800 105.600 ;
        RECT 129.200 102.200 130.000 106.800 ;
        RECT 132.800 106.200 133.400 107.600 ;
        RECT 132.400 105.600 133.400 106.200 ;
        RECT 137.200 109.000 138.000 114.600 ;
        RECT 139.800 114.400 144.000 115.200 ;
        RECT 148.400 115.000 149.200 119.800 ;
        RECT 151.600 115.000 152.400 119.800 ;
        RECT 139.800 114.000 140.400 114.400 ;
        RECT 138.800 113.200 140.400 114.000 ;
        RECT 143.400 113.800 149.200 114.400 ;
        RECT 141.400 113.200 142.800 113.800 ;
        RECT 141.400 113.000 147.600 113.200 ;
        RECT 142.200 112.600 147.600 113.000 ;
        RECT 146.800 112.400 147.600 112.600 ;
        RECT 148.600 113.000 149.200 113.800 ;
        RECT 149.800 113.600 152.400 114.400 ;
        RECT 154.800 113.600 155.600 119.800 ;
        RECT 156.400 117.000 157.200 119.800 ;
        RECT 158.000 117.000 158.800 119.800 ;
        RECT 159.600 117.000 160.400 119.800 ;
        RECT 158.000 114.400 162.200 115.200 ;
        RECT 162.800 114.400 163.600 119.800 ;
        RECT 166.000 115.200 166.800 119.800 ;
        RECT 166.000 114.600 168.600 115.200 ;
        RECT 162.800 113.600 165.400 114.400 ;
        RECT 156.400 113.000 157.200 113.200 ;
        RECT 148.600 112.400 157.200 113.000 ;
        RECT 159.600 113.000 160.400 113.200 ;
        RECT 168.000 113.000 168.600 114.600 ;
        RECT 159.600 112.400 168.600 113.000 ;
        RECT 168.000 110.600 168.600 112.400 ;
        RECT 169.200 112.000 170.000 119.800 ;
        RECT 169.200 111.200 170.200 112.000 ;
        RECT 172.400 111.800 173.200 119.800 ;
        RECT 174.000 112.400 174.800 119.800 ;
        RECT 177.200 112.400 178.000 119.800 ;
        RECT 182.000 116.400 182.800 119.800 ;
        RECT 181.800 115.800 182.800 116.400 ;
        RECT 181.800 115.200 182.400 115.800 ;
        RECT 185.200 115.200 186.000 119.800 ;
        RECT 188.400 117.000 189.200 119.800 ;
        RECT 190.000 117.000 190.800 119.800 ;
        RECT 174.000 111.800 178.000 112.400 ;
        RECT 180.400 114.600 182.400 115.200 ;
        RECT 138.600 110.000 162.000 110.600 ;
        RECT 168.000 110.000 168.800 110.600 ;
        RECT 138.600 109.800 139.400 110.000 ;
        RECT 140.400 109.600 141.200 110.000 ;
        RECT 143.600 109.600 144.400 110.000 ;
        RECT 161.200 109.400 162.000 110.000 ;
        RECT 137.200 108.200 146.000 109.000 ;
        RECT 146.600 108.600 148.600 109.400 ;
        RECT 152.400 108.600 155.600 109.400 ;
        RECT 132.400 102.200 133.200 105.600 ;
        RECT 137.200 102.200 138.000 108.200 ;
        RECT 139.600 106.800 142.600 107.600 ;
        RECT 141.800 106.200 142.600 106.800 ;
        RECT 147.800 106.200 148.600 108.600 ;
        RECT 150.000 106.800 150.800 108.400 ;
        RECT 155.200 107.800 156.000 108.000 ;
        RECT 151.600 107.200 156.000 107.800 ;
        RECT 151.600 107.000 152.400 107.200 ;
        RECT 158.000 106.400 158.800 109.200 ;
        RECT 163.800 108.600 167.600 109.400 ;
        RECT 163.800 107.400 164.600 108.600 ;
        RECT 168.200 108.000 168.800 110.000 ;
        RECT 151.600 106.200 152.400 106.400 ;
        RECT 141.800 105.400 144.400 106.200 ;
        RECT 147.800 105.600 152.400 106.200 ;
        RECT 153.200 105.600 154.800 106.400 ;
        RECT 157.800 105.600 158.800 106.400 ;
        RECT 162.800 106.800 164.600 107.400 ;
        RECT 167.600 107.400 168.800 108.000 ;
        RECT 162.800 106.200 163.600 106.800 ;
        RECT 143.600 102.200 144.400 105.400 ;
        RECT 161.200 105.400 163.600 106.200 ;
        RECT 145.200 102.200 146.000 105.000 ;
        RECT 146.800 102.200 147.600 105.000 ;
        RECT 148.400 102.200 149.200 105.000 ;
        RECT 151.600 102.200 152.400 105.000 ;
        RECT 154.800 102.200 155.600 105.000 ;
        RECT 156.400 102.200 157.200 105.000 ;
        RECT 158.000 102.200 158.800 105.000 ;
        RECT 159.600 102.200 160.400 105.000 ;
        RECT 161.200 102.200 162.000 105.400 ;
        RECT 167.600 102.200 168.400 107.400 ;
        RECT 169.400 106.800 170.200 111.200 ;
        RECT 172.600 110.400 173.200 111.800 ;
        RECT 176.400 110.400 177.200 110.800 ;
        RECT 172.400 109.800 174.800 110.400 ;
        RECT 176.400 109.800 178.000 110.400 ;
        RECT 172.400 109.600 173.200 109.800 ;
        RECT 169.200 106.000 170.200 106.800 ;
        RECT 174.200 106.400 174.800 109.800 ;
        RECT 177.200 109.600 178.000 109.800 ;
        RECT 175.600 107.600 176.400 109.200 ;
        RECT 180.400 109.000 181.200 114.600 ;
        RECT 183.000 114.400 187.200 115.200 ;
        RECT 191.600 115.000 192.400 119.800 ;
        RECT 194.800 115.000 195.600 119.800 ;
        RECT 183.000 114.000 183.600 114.400 ;
        RECT 182.000 113.200 183.600 114.000 ;
        RECT 186.600 113.800 192.400 114.400 ;
        RECT 184.600 113.200 186.000 113.800 ;
        RECT 184.600 113.000 190.800 113.200 ;
        RECT 185.400 112.600 190.800 113.000 ;
        RECT 190.000 112.400 190.800 112.600 ;
        RECT 191.800 113.000 192.400 113.800 ;
        RECT 193.000 113.600 195.600 114.400 ;
        RECT 198.000 113.600 198.800 119.800 ;
        RECT 199.600 117.000 200.400 119.800 ;
        RECT 201.200 117.000 202.000 119.800 ;
        RECT 202.800 117.000 203.600 119.800 ;
        RECT 201.200 114.400 205.400 115.200 ;
        RECT 206.000 114.400 206.800 119.800 ;
        RECT 209.200 115.200 210.000 119.800 ;
        RECT 209.200 114.600 211.800 115.200 ;
        RECT 206.000 113.600 208.600 114.400 ;
        RECT 199.600 113.000 200.400 113.200 ;
        RECT 191.800 112.400 200.400 113.000 ;
        RECT 202.800 113.000 203.600 113.200 ;
        RECT 211.200 113.000 211.800 114.600 ;
        RECT 202.800 112.400 211.800 113.000 ;
        RECT 211.200 110.600 211.800 112.400 ;
        RECT 212.400 112.000 213.200 119.800 ;
        RECT 212.400 111.200 213.400 112.000 ;
        RECT 181.800 110.000 205.200 110.600 ;
        RECT 211.200 110.000 212.000 110.600 ;
        RECT 181.800 109.800 182.600 110.000 ;
        RECT 183.600 109.600 184.400 110.000 ;
        RECT 186.800 109.600 187.600 110.000 ;
        RECT 204.400 109.400 205.200 110.000 ;
        RECT 180.400 108.200 189.200 109.000 ;
        RECT 189.800 108.600 191.800 109.400 ;
        RECT 195.600 108.600 198.800 109.400 ;
        RECT 169.200 102.200 170.000 106.000 ;
        RECT 172.400 105.600 173.200 106.400 ;
        RECT 172.600 104.800 173.400 105.600 ;
        RECT 174.000 102.200 174.800 106.400 ;
        RECT 180.400 102.200 181.200 108.200 ;
        RECT 182.800 106.800 185.800 107.600 ;
        RECT 185.000 106.200 185.800 106.800 ;
        RECT 191.000 106.200 191.800 108.600 ;
        RECT 193.200 106.800 194.000 108.400 ;
        RECT 198.400 107.800 199.200 108.000 ;
        RECT 194.800 107.200 199.200 107.800 ;
        RECT 194.800 107.000 195.600 107.200 ;
        RECT 201.200 106.400 202.000 109.200 ;
        RECT 207.000 108.600 210.800 109.400 ;
        RECT 207.000 107.400 207.800 108.600 ;
        RECT 211.400 108.000 212.000 110.000 ;
        RECT 194.800 106.200 195.600 106.400 ;
        RECT 185.000 105.400 187.600 106.200 ;
        RECT 191.000 105.600 195.600 106.200 ;
        RECT 196.400 105.600 198.000 106.400 ;
        RECT 201.000 105.600 202.000 106.400 ;
        RECT 206.000 106.800 207.800 107.400 ;
        RECT 210.800 107.400 212.000 108.000 ;
        RECT 206.000 106.200 206.800 106.800 ;
        RECT 186.800 102.200 187.600 105.400 ;
        RECT 204.400 105.400 206.800 106.200 ;
        RECT 188.400 102.200 189.200 105.000 ;
        RECT 190.000 102.200 190.800 105.000 ;
        RECT 191.600 102.200 192.400 105.000 ;
        RECT 194.800 102.200 195.600 105.000 ;
        RECT 198.000 102.200 198.800 105.000 ;
        RECT 199.600 102.200 200.400 105.000 ;
        RECT 201.200 102.200 202.000 105.000 ;
        RECT 202.800 102.200 203.600 105.000 ;
        RECT 204.400 102.200 205.200 105.400 ;
        RECT 210.800 102.200 211.600 107.400 ;
        RECT 212.600 106.800 213.400 111.200 ;
        RECT 212.400 106.000 213.400 106.800 ;
        RECT 212.400 102.200 213.200 106.000 ;
        RECT 215.600 102.200 216.400 119.800 ;
        RECT 218.800 112.400 219.600 119.800 ;
        RECT 218.800 111.800 221.000 112.400 ;
        RECT 220.400 111.200 221.000 111.800 ;
        RECT 220.400 110.400 221.600 111.200 ;
        RECT 218.800 108.800 219.600 110.400 ;
        RECT 220.400 107.400 221.000 110.400 ;
        RECT 218.800 106.800 221.000 107.400 ;
        RECT 217.200 104.800 218.000 106.400 ;
        RECT 218.800 102.200 219.600 106.800 ;
        RECT 2.800 90.300 3.600 99.800 ;
        RECT 4.400 95.800 5.200 99.800 ;
        RECT 6.000 96.000 6.800 99.800 ;
        RECT 9.200 96.000 10.000 99.800 ;
        RECT 6.000 95.800 10.000 96.000 ;
        RECT 4.600 94.400 5.200 95.800 ;
        RECT 6.200 95.400 9.800 95.800 ;
        RECT 4.400 93.600 7.000 94.400 ;
        RECT 14.400 94.200 15.200 99.800 ;
        RECT 18.400 94.200 19.200 99.800 ;
        RECT 14.400 93.800 16.200 94.200 ;
        RECT 14.600 93.600 16.200 93.800 ;
        RECT 6.400 92.400 7.000 93.600 ;
        RECT 6.000 91.600 7.000 92.400 ;
        RECT 7.600 91.600 8.400 93.200 ;
        RECT 12.400 91.600 14.000 92.400 ;
        RECT 4.400 90.300 5.200 90.400 ;
        RECT 2.800 90.200 5.200 90.300 ;
        RECT 6.400 90.200 7.000 91.600 ;
        RECT 2.800 89.700 5.800 90.200 ;
        RECT 2.800 82.200 3.600 89.700 ;
        RECT 4.400 89.600 5.800 89.700 ;
        RECT 6.400 89.600 7.400 90.200 ;
        RECT 10.800 89.600 11.600 91.200 ;
        RECT 15.600 90.400 16.200 93.600 ;
        RECT 17.400 93.800 19.200 94.200 ;
        RECT 17.400 93.600 19.000 93.800 ;
        RECT 17.400 90.400 18.000 93.600 ;
        RECT 15.600 89.600 16.400 90.400 ;
        RECT 17.200 89.600 18.000 90.400 ;
        RECT 22.000 89.600 22.800 91.200 ;
        RECT 5.200 88.400 5.800 89.600 ;
        RECT 5.200 87.600 6.000 88.400 ;
        RECT 6.600 82.200 7.400 89.600 ;
        RECT 14.000 87.600 14.800 89.200 ;
        RECT 15.600 87.000 16.200 89.600 ;
        RECT 17.400 88.400 18.000 89.600 ;
        RECT 17.200 87.600 18.000 88.400 ;
        RECT 18.800 88.300 19.600 89.200 ;
        RECT 23.600 88.300 24.400 99.800 ;
        RECT 25.200 95.600 26.000 97.200 ;
        RECT 25.200 92.300 26.000 92.400 ;
        RECT 26.800 92.300 27.600 99.800 ;
        RECT 30.000 96.000 30.800 99.800 ;
        RECT 33.200 96.000 34.000 99.800 ;
        RECT 30.000 95.800 34.000 96.000 ;
        RECT 34.800 96.300 35.600 99.800 ;
        RECT 38.000 96.300 38.800 97.200 ;
        RECT 30.200 95.400 33.800 95.800 ;
        RECT 34.800 95.700 38.800 96.300 ;
        RECT 34.800 94.400 35.400 95.700 ;
        RECT 38.000 95.600 38.800 95.700 ;
        RECT 33.000 93.600 35.600 94.400 ;
        RECT 25.200 91.700 27.600 92.300 ;
        RECT 25.200 91.600 26.000 91.700 ;
        RECT 25.200 88.300 26.000 88.400 ;
        RECT 18.800 87.700 26.000 88.300 ;
        RECT 18.800 87.600 19.600 87.700 ;
        RECT 12.600 86.400 16.200 87.000 ;
        RECT 17.400 87.000 18.000 87.600 ;
        RECT 17.400 86.400 21.000 87.000 ;
        RECT 12.600 86.200 13.200 86.400 ;
        RECT 12.400 82.200 13.200 86.200 ;
        RECT 15.600 82.200 16.400 86.400 ;
        RECT 17.400 86.200 18.000 86.400 ;
        RECT 17.200 82.200 18.000 86.200 ;
        RECT 20.400 86.200 21.000 86.400 ;
        RECT 20.400 82.200 21.200 86.200 ;
        RECT 23.600 82.200 24.400 87.700 ;
        RECT 25.200 87.600 26.000 87.700 ;
        RECT 26.800 82.200 27.600 91.700 ;
        RECT 31.600 91.600 32.400 93.200 ;
        RECT 33.000 90.200 33.600 93.600 ;
        RECT 34.800 90.200 35.600 90.400 ;
        RECT 32.600 89.600 33.600 90.200 ;
        RECT 34.200 89.600 35.600 90.200 ;
        RECT 32.600 82.200 33.400 89.600 ;
        RECT 34.200 88.400 34.800 89.600 ;
        RECT 34.000 87.600 34.800 88.400 ;
        RECT 39.600 82.200 40.400 99.800 ;
        RECT 41.200 96.000 42.000 99.800 ;
        RECT 44.400 96.000 45.200 99.800 ;
        RECT 41.200 95.800 45.200 96.000 ;
        RECT 46.000 95.800 46.800 99.800 ;
        RECT 47.600 95.800 48.400 99.800 ;
        RECT 49.200 96.000 50.000 99.800 ;
        RECT 52.400 96.000 53.200 99.800 ;
        RECT 49.200 95.800 53.200 96.000 ;
        RECT 54.000 95.800 54.800 99.800 ;
        RECT 58.200 96.800 59.000 99.800 ;
        RECT 58.200 95.800 59.600 96.800 ;
        RECT 62.000 96.000 62.800 99.800 ;
        RECT 41.400 95.400 45.000 95.800 ;
        RECT 42.000 94.400 42.800 94.800 ;
        RECT 46.000 94.400 46.600 95.800 ;
        RECT 47.800 94.400 48.400 95.800 ;
        RECT 49.400 95.400 53.000 95.800 ;
        RECT 54.200 95.600 54.800 95.800 ;
        RECT 54.200 95.200 56.000 95.600 ;
        RECT 54.200 95.000 58.400 95.200 ;
        RECT 51.600 94.400 52.400 94.800 ;
        RECT 55.400 94.600 58.400 95.000 ;
        RECT 57.600 94.400 58.400 94.600 ;
        RECT 41.200 93.800 42.800 94.400 ;
        RECT 41.200 93.600 42.000 93.800 ;
        RECT 44.200 93.600 46.800 94.400 ;
        RECT 47.600 93.600 50.200 94.400 ;
        RECT 51.600 93.800 53.200 94.400 ;
        RECT 52.400 93.600 53.200 93.800 ;
        RECT 42.800 91.600 43.600 93.200 ;
        RECT 44.200 92.300 44.800 93.600 ;
        RECT 44.200 91.700 48.300 92.300 ;
        RECT 44.200 90.200 44.800 91.700 ;
        RECT 47.700 90.400 48.300 91.700 ;
        RECT 46.000 90.200 46.800 90.400 ;
        RECT 43.800 89.600 44.800 90.200 ;
        RECT 45.400 89.600 46.800 90.200 ;
        RECT 47.600 90.200 48.400 90.400 ;
        RECT 49.600 90.200 50.200 93.600 ;
        RECT 50.800 91.600 51.600 93.200 ;
        RECT 54.000 92.800 54.800 94.400 ;
        RECT 56.000 93.800 56.800 94.000 ;
        RECT 55.800 93.200 56.800 93.800 ;
        RECT 55.800 92.400 56.400 93.200 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 57.600 91.000 58.200 94.400 ;
        RECT 59.000 92.400 59.600 95.800 ;
        RECT 61.800 95.200 62.800 96.000 ;
        RECT 58.800 92.300 59.600 92.400 ;
        RECT 60.400 92.300 61.200 92.400 ;
        RECT 58.800 91.700 61.200 92.300 ;
        RECT 58.800 91.600 59.600 91.700 ;
        RECT 60.400 91.600 61.200 91.700 ;
        RECT 55.800 90.400 58.200 91.000 ;
        RECT 47.600 89.600 49.000 90.200 ;
        RECT 49.600 89.600 50.600 90.200 ;
        RECT 43.800 82.200 44.600 89.600 ;
        RECT 45.400 88.400 46.000 89.600 ;
        RECT 45.200 87.600 46.000 88.400 ;
        RECT 48.400 88.400 49.000 89.600 ;
        RECT 48.400 87.600 49.200 88.400 ;
        RECT 49.800 82.200 50.600 89.600 ;
        RECT 55.800 86.200 56.400 90.400 ;
        RECT 59.000 90.200 59.600 91.600 ;
        RECT 55.600 82.200 56.400 86.200 ;
        RECT 58.800 82.200 59.600 90.200 ;
        RECT 61.800 90.800 62.600 95.200 ;
        RECT 63.600 94.600 64.400 99.800 ;
        RECT 70.000 96.600 70.800 99.800 ;
        RECT 71.600 97.000 72.400 99.800 ;
        RECT 73.200 97.000 74.000 99.800 ;
        RECT 74.800 97.000 75.600 99.800 ;
        RECT 76.400 97.000 77.200 99.800 ;
        RECT 79.600 97.000 80.400 99.800 ;
        RECT 82.800 97.000 83.600 99.800 ;
        RECT 84.400 97.000 85.200 99.800 ;
        RECT 86.000 97.000 86.800 99.800 ;
        RECT 68.400 95.800 70.800 96.600 ;
        RECT 87.600 96.600 88.400 99.800 ;
        RECT 68.400 95.200 69.200 95.800 ;
        RECT 63.200 94.000 64.400 94.600 ;
        RECT 67.400 94.600 69.200 95.200 ;
        RECT 73.200 95.600 74.200 96.400 ;
        RECT 77.200 95.600 78.800 96.400 ;
        RECT 79.600 95.800 84.200 96.400 ;
        RECT 87.600 95.800 90.200 96.600 ;
        RECT 79.600 95.600 80.400 95.800 ;
        RECT 63.200 92.000 63.800 94.000 ;
        RECT 67.400 93.400 68.200 94.600 ;
        RECT 64.400 92.600 68.200 93.400 ;
        RECT 73.200 92.800 74.000 95.600 ;
        RECT 79.600 94.800 80.400 95.000 ;
        RECT 76.000 94.200 80.400 94.800 ;
        RECT 76.000 94.000 76.800 94.200 ;
        RECT 81.200 93.600 82.000 95.200 ;
        RECT 83.400 93.400 84.200 95.800 ;
        RECT 89.400 95.200 90.200 95.800 ;
        RECT 89.400 94.400 92.400 95.200 ;
        RECT 94.000 93.800 94.800 99.800 ;
        RECT 100.400 95.200 101.200 99.800 ;
        RECT 103.600 96.000 104.400 99.800 ;
        RECT 76.400 92.600 79.600 93.400 ;
        RECT 83.400 92.600 85.400 93.400 ;
        RECT 86.000 93.000 94.800 93.800 ;
        RECT 70.000 92.000 70.800 92.600 ;
        RECT 87.600 92.000 88.400 92.400 ;
        RECT 89.200 92.000 90.000 92.400 ;
        RECT 92.600 92.000 93.400 92.200 ;
        RECT 63.200 91.400 64.000 92.000 ;
        RECT 70.000 91.400 93.400 92.000 ;
        RECT 61.800 90.000 62.800 90.800 ;
        RECT 62.000 82.200 62.800 90.000 ;
        RECT 63.400 89.600 64.000 91.400 ;
        RECT 63.400 89.000 72.400 89.600 ;
        RECT 63.400 87.400 64.000 89.000 ;
        RECT 71.600 88.800 72.400 89.000 ;
        RECT 74.800 89.000 83.400 89.600 ;
        RECT 74.800 88.800 75.600 89.000 ;
        RECT 66.600 87.600 69.200 88.400 ;
        RECT 63.400 86.800 66.000 87.400 ;
        RECT 65.200 82.200 66.000 86.800 ;
        RECT 68.400 82.200 69.200 87.600 ;
        RECT 69.800 86.800 74.000 87.600 ;
        RECT 71.600 82.200 72.400 85.000 ;
        RECT 73.200 82.200 74.000 85.000 ;
        RECT 74.800 82.200 75.600 85.000 ;
        RECT 76.400 82.200 77.200 88.400 ;
        RECT 79.600 87.600 82.200 88.400 ;
        RECT 82.800 88.200 83.400 89.000 ;
        RECT 84.400 89.400 85.200 89.600 ;
        RECT 84.400 89.000 89.800 89.400 ;
        RECT 84.400 88.800 90.600 89.000 ;
        RECT 89.200 88.200 90.600 88.800 ;
        RECT 82.800 87.600 88.600 88.200 ;
        RECT 91.600 88.000 93.200 88.800 ;
        RECT 91.600 87.600 92.200 88.000 ;
        RECT 79.600 82.200 80.400 87.000 ;
        RECT 82.800 82.200 83.600 87.000 ;
        RECT 88.000 86.800 92.200 87.600 ;
        RECT 94.000 87.400 94.800 93.000 ;
        RECT 99.000 94.600 101.200 95.200 ;
        RECT 103.400 95.200 104.400 96.000 ;
        RECT 99.000 91.600 99.600 94.600 ;
        RECT 100.400 92.300 101.200 93.200 ;
        RECT 103.400 92.300 104.200 95.200 ;
        RECT 105.200 94.600 106.000 99.800 ;
        RECT 111.600 96.600 112.400 99.800 ;
        RECT 113.200 97.000 114.000 99.800 ;
        RECT 114.800 97.000 115.600 99.800 ;
        RECT 116.400 97.000 117.200 99.800 ;
        RECT 118.000 97.000 118.800 99.800 ;
        RECT 121.200 97.000 122.000 99.800 ;
        RECT 124.400 97.000 125.200 99.800 ;
        RECT 126.000 97.000 126.800 99.800 ;
        RECT 127.600 97.000 128.400 99.800 ;
        RECT 110.000 95.800 112.400 96.600 ;
        RECT 129.200 96.600 130.000 99.800 ;
        RECT 110.000 95.200 110.800 95.800 ;
        RECT 100.400 91.700 104.200 92.300 ;
        RECT 100.400 91.600 101.200 91.700 ;
        RECT 98.400 90.800 99.600 91.600 ;
        RECT 99.000 90.200 99.600 90.800 ;
        RECT 103.400 90.800 104.200 91.700 ;
        RECT 104.800 94.000 106.000 94.600 ;
        RECT 109.000 94.600 110.800 95.200 ;
        RECT 114.800 95.600 115.800 96.400 ;
        RECT 118.800 95.600 120.400 96.400 ;
        RECT 121.200 95.800 125.800 96.400 ;
        RECT 129.200 95.800 131.800 96.600 ;
        RECT 121.200 95.600 122.000 95.800 ;
        RECT 104.800 92.000 105.400 94.000 ;
        RECT 109.000 93.400 109.800 94.600 ;
        RECT 106.000 92.600 109.800 93.400 ;
        RECT 114.800 92.800 115.600 95.600 ;
        RECT 121.200 94.800 122.000 95.000 ;
        RECT 117.600 94.200 122.000 94.800 ;
        RECT 117.600 94.000 118.400 94.200 ;
        RECT 122.800 93.600 123.600 95.200 ;
        RECT 125.000 93.400 125.800 95.800 ;
        RECT 131.000 95.200 131.800 95.800 ;
        RECT 131.000 94.400 134.000 95.200 ;
        RECT 135.600 93.800 136.400 99.800 ;
        RECT 138.800 95.800 139.600 99.800 ;
        RECT 140.400 96.000 141.200 99.800 ;
        RECT 143.600 96.000 144.400 99.800 ;
        RECT 145.400 96.400 146.200 97.200 ;
        RECT 140.400 95.800 144.400 96.000 ;
        RECT 139.000 94.400 139.600 95.800 ;
        RECT 140.600 95.400 144.200 95.800 ;
        RECT 145.200 95.600 146.000 96.400 ;
        RECT 146.800 95.800 147.600 99.800 ;
        RECT 142.800 94.400 143.600 94.800 ;
        RECT 118.000 92.600 121.200 93.400 ;
        RECT 125.000 92.600 127.000 93.400 ;
        RECT 127.600 93.000 136.400 93.800 ;
        RECT 138.800 93.600 141.400 94.400 ;
        RECT 142.800 94.300 144.400 94.400 ;
        RECT 145.200 94.300 146.000 94.400 ;
        RECT 142.800 93.800 146.000 94.300 ;
        RECT 143.600 93.700 146.000 93.800 ;
        RECT 143.600 93.600 144.400 93.700 ;
        RECT 145.200 93.600 146.000 93.700 ;
        RECT 111.600 92.000 112.400 92.600 ;
        RECT 129.200 92.000 130.000 92.400 ;
        RECT 130.800 92.000 131.600 92.400 ;
        RECT 134.200 92.000 135.000 92.200 ;
        RECT 104.800 91.400 105.600 92.000 ;
        RECT 111.600 91.400 135.000 92.000 ;
        RECT 99.000 89.600 101.200 90.200 ;
        RECT 103.400 90.000 104.400 90.800 ;
        RECT 92.800 86.800 94.800 87.400 ;
        RECT 84.400 82.200 85.200 85.000 ;
        RECT 86.000 82.200 86.800 85.000 ;
        RECT 89.200 82.200 90.000 86.800 ;
        RECT 92.800 86.200 93.400 86.800 ;
        RECT 92.400 85.600 93.400 86.200 ;
        RECT 92.400 82.200 93.200 85.600 ;
        RECT 100.400 82.200 101.200 89.600 ;
        RECT 103.600 82.200 104.400 90.000 ;
        RECT 105.000 89.600 105.600 91.400 ;
        RECT 105.000 89.000 114.000 89.600 ;
        RECT 105.000 87.400 105.600 89.000 ;
        RECT 113.200 88.800 114.000 89.000 ;
        RECT 116.400 89.000 125.000 89.600 ;
        RECT 116.400 88.800 117.200 89.000 ;
        RECT 108.200 87.600 110.800 88.400 ;
        RECT 105.000 86.800 107.600 87.400 ;
        RECT 106.800 82.200 107.600 86.800 ;
        RECT 110.000 82.200 110.800 87.600 ;
        RECT 111.400 86.800 115.600 87.600 ;
        RECT 113.200 82.200 114.000 85.000 ;
        RECT 114.800 82.200 115.600 85.000 ;
        RECT 116.400 82.200 117.200 85.000 ;
        RECT 118.000 82.200 118.800 88.400 ;
        RECT 121.200 87.600 123.800 88.400 ;
        RECT 124.400 88.200 125.000 89.000 ;
        RECT 126.000 89.400 126.800 89.600 ;
        RECT 126.000 89.000 131.400 89.400 ;
        RECT 126.000 88.800 132.200 89.000 ;
        RECT 130.800 88.200 132.200 88.800 ;
        RECT 124.400 87.600 130.200 88.200 ;
        RECT 133.200 88.000 134.800 88.800 ;
        RECT 133.200 87.600 133.800 88.000 ;
        RECT 121.200 82.200 122.000 87.000 ;
        RECT 124.400 82.200 125.200 87.000 ;
        RECT 129.600 86.800 133.800 87.600 ;
        RECT 135.600 87.400 136.400 93.000 ;
        RECT 138.800 90.200 139.600 90.400 ;
        RECT 140.800 90.200 141.400 93.600 ;
        RECT 142.000 92.300 142.800 93.200 ;
        RECT 143.600 92.300 144.400 92.400 ;
        RECT 142.000 91.700 144.400 92.300 ;
        RECT 142.000 91.600 142.800 91.700 ;
        RECT 143.600 91.600 144.400 91.700 ;
        RECT 145.200 92.200 146.000 92.400 ;
        RECT 147.000 92.200 147.600 95.800 ;
        RECT 153.200 97.600 154.000 99.800 ;
        RECT 153.200 94.400 153.800 97.600 ;
        RECT 154.800 95.600 155.600 97.200 ;
        RECT 156.400 95.800 157.200 99.800 ;
        RECT 160.800 96.200 162.400 99.800 ;
        RECT 156.400 95.200 158.800 95.800 ;
        RECT 158.000 95.000 158.800 95.200 ;
        RECT 159.400 94.800 160.200 95.600 ;
        RECT 159.400 94.400 160.000 94.800 ;
        RECT 148.400 92.800 149.200 94.400 ;
        RECT 153.200 93.600 154.000 94.400 ;
        RECT 156.400 93.600 158.000 94.400 ;
        RECT 159.200 93.600 160.000 94.400 ;
        RECT 150.000 92.200 150.800 92.400 ;
        RECT 145.200 91.600 147.600 92.200 ;
        RECT 149.200 91.600 150.800 92.200 ;
        RECT 145.400 90.200 146.000 91.600 ;
        RECT 149.200 91.200 150.000 91.600 ;
        RECT 151.600 90.800 152.400 92.400 ;
        RECT 153.200 90.200 153.800 93.600 ;
        RECT 160.800 92.800 161.400 96.200 ;
        RECT 166.000 95.800 166.800 99.800 ;
        RECT 167.600 96.000 168.400 99.800 ;
        RECT 170.800 96.000 171.600 99.800 ;
        RECT 167.600 95.800 171.600 96.000 ;
        RECT 172.400 95.800 173.200 99.800 ;
        RECT 174.000 96.000 174.800 99.800 ;
        RECT 177.200 96.000 178.000 99.800 ;
        RECT 174.000 95.800 178.000 96.000 ;
        RECT 178.800 95.800 179.600 99.800 ;
        RECT 162.000 95.400 163.600 95.600 ;
        RECT 162.000 94.800 164.000 95.400 ;
        RECT 164.600 95.200 166.800 95.800 ;
        RECT 167.800 95.400 171.400 95.800 ;
        RECT 164.600 95.000 165.400 95.200 ;
        RECT 163.400 94.400 164.000 94.800 ;
        RECT 168.400 94.400 169.200 94.800 ;
        RECT 172.400 94.400 173.000 95.800 ;
        RECT 174.200 95.400 177.800 95.800 ;
        RECT 174.800 94.400 175.600 94.800 ;
        RECT 178.800 94.400 179.400 95.800 ;
        RECT 163.400 94.300 166.800 94.400 ;
        RECT 167.600 94.300 169.200 94.400 ;
        RECT 162.000 93.400 162.800 94.200 ;
        RECT 163.400 93.800 169.200 94.300 ;
        RECT 165.200 93.700 168.400 93.800 ;
        RECT 165.200 93.600 166.800 93.700 ;
        RECT 167.600 93.600 168.400 93.700 ;
        RECT 170.600 93.600 173.200 94.400 ;
        RECT 174.000 93.800 175.600 94.400 ;
        RECT 174.000 93.600 174.800 93.800 ;
        RECT 177.000 93.600 179.600 94.400 ;
        RECT 182.000 93.800 182.800 99.800 ;
        RECT 188.400 96.600 189.200 99.800 ;
        RECT 190.000 97.000 190.800 99.800 ;
        RECT 191.600 97.000 192.400 99.800 ;
        RECT 193.200 97.000 194.000 99.800 ;
        RECT 196.400 97.000 197.200 99.800 ;
        RECT 199.600 97.000 200.400 99.800 ;
        RECT 201.200 97.000 202.000 99.800 ;
        RECT 202.800 97.000 203.600 99.800 ;
        RECT 204.400 97.000 205.200 99.800 ;
        RECT 186.600 95.800 189.200 96.600 ;
        RECT 206.000 96.600 206.800 99.800 ;
        RECT 192.600 95.800 197.200 96.400 ;
        RECT 186.600 95.200 187.400 95.800 ;
        RECT 184.400 94.400 187.400 95.200 ;
        RECT 160.400 92.400 161.400 92.800 ;
        RECT 159.600 92.200 161.400 92.400 ;
        RECT 162.200 92.800 162.800 93.400 ;
        RECT 162.200 92.200 164.800 92.800 ;
        RECT 159.600 91.600 161.000 92.200 ;
        RECT 164.000 92.000 164.800 92.200 ;
        RECT 166.000 92.300 166.800 92.400 ;
        RECT 169.200 92.300 170.000 93.200 ;
        RECT 166.000 91.700 170.000 92.300 ;
        RECT 166.000 91.600 166.800 91.700 ;
        RECT 169.200 91.600 170.000 91.700 ;
        RECT 160.400 90.400 161.000 91.600 ;
        RECT 161.800 91.400 162.600 91.600 ;
        RECT 161.800 90.800 165.200 91.400 ;
        RECT 159.600 90.200 161.000 90.400 ;
        RECT 164.600 90.200 165.200 90.800 ;
        RECT 170.600 90.200 171.200 93.600 ;
        RECT 175.600 91.600 176.400 93.200 ;
        RECT 172.400 90.200 173.200 90.400 ;
        RECT 177.000 90.200 177.600 93.600 ;
        RECT 182.000 93.000 190.800 93.800 ;
        RECT 192.600 93.400 193.400 95.800 ;
        RECT 196.400 95.600 197.200 95.800 ;
        RECT 198.000 95.600 199.600 96.400 ;
        RECT 202.600 95.600 203.600 96.400 ;
        RECT 206.000 95.800 208.400 96.600 ;
        RECT 194.800 93.600 195.600 95.200 ;
        RECT 196.400 94.800 197.200 95.000 ;
        RECT 196.400 94.200 200.800 94.800 ;
        RECT 200.000 94.000 200.800 94.200 ;
        RECT 178.800 90.200 179.600 90.400 ;
        RECT 138.800 89.600 140.200 90.200 ;
        RECT 140.800 89.600 141.800 90.200 ;
        RECT 139.600 88.400 140.200 89.600 ;
        RECT 139.600 87.600 140.400 88.400 ;
        RECT 134.400 86.800 136.400 87.400 ;
        RECT 126.000 82.200 126.800 85.000 ;
        RECT 127.600 82.200 128.400 85.000 ;
        RECT 130.800 82.200 131.600 86.800 ;
        RECT 134.400 86.200 135.000 86.800 ;
        RECT 134.000 85.600 135.000 86.200 ;
        RECT 134.000 82.200 134.800 85.600 ;
        RECT 141.000 82.200 141.800 89.600 ;
        RECT 145.200 82.200 146.000 90.200 ;
        RECT 146.800 89.600 150.800 90.200 ;
        RECT 146.800 82.200 147.600 89.600 ;
        RECT 150.000 82.200 150.800 89.600 ;
        RECT 152.200 89.400 154.000 90.200 ;
        RECT 156.400 89.600 158.800 90.200 ;
        RECT 159.600 89.600 162.400 90.200 ;
        RECT 152.200 82.200 153.000 89.400 ;
        RECT 156.400 82.200 157.200 89.600 ;
        RECT 158.000 89.400 158.800 89.600 ;
        RECT 160.800 82.200 162.400 89.600 ;
        RECT 164.600 89.600 166.800 90.200 ;
        RECT 164.600 89.400 165.400 89.600 ;
        RECT 166.000 82.200 166.800 89.600 ;
        RECT 170.200 89.600 171.200 90.200 ;
        RECT 171.800 89.600 173.200 90.200 ;
        RECT 176.600 89.600 177.600 90.200 ;
        RECT 178.200 89.600 179.600 90.200 ;
        RECT 170.200 82.200 171.000 89.600 ;
        RECT 171.800 88.400 172.400 89.600 ;
        RECT 171.600 87.600 172.400 88.400 ;
        RECT 176.600 82.200 177.400 89.600 ;
        RECT 178.200 88.400 178.800 89.600 ;
        RECT 178.000 87.600 178.800 88.400 ;
        RECT 182.000 87.400 182.800 93.000 ;
        RECT 191.400 92.600 193.400 93.400 ;
        RECT 197.200 92.600 200.400 93.400 ;
        RECT 202.800 92.800 203.600 95.600 ;
        RECT 207.600 95.200 208.400 95.800 ;
        RECT 207.600 94.600 209.400 95.200 ;
        RECT 208.600 93.400 209.400 94.600 ;
        RECT 212.400 94.600 213.200 99.800 ;
        RECT 214.000 96.000 214.800 99.800 ;
        RECT 217.200 97.000 218.000 99.000 ;
        RECT 214.000 95.200 215.000 96.000 ;
        RECT 212.400 94.000 213.600 94.600 ;
        RECT 208.600 92.600 212.400 93.400 ;
        RECT 183.400 92.000 184.200 92.200 ;
        RECT 185.200 92.000 186.000 92.400 ;
        RECT 188.400 92.000 189.200 92.400 ;
        RECT 206.000 92.000 206.800 92.600 ;
        RECT 213.000 92.000 213.600 94.000 ;
        RECT 183.400 91.400 206.800 92.000 ;
        RECT 212.800 91.400 213.600 92.000 ;
        RECT 212.800 89.600 213.400 91.400 ;
        RECT 214.200 90.800 215.000 95.200 ;
        RECT 217.200 94.800 217.800 97.000 ;
        RECT 221.400 96.400 222.200 99.000 ;
        RECT 220.400 96.000 222.200 96.400 ;
        RECT 220.400 95.600 223.000 96.000 ;
        RECT 221.400 95.400 223.000 95.600 ;
        RECT 222.200 95.000 223.000 95.400 ;
        RECT 217.200 94.200 221.400 94.800 ;
        RECT 220.400 93.800 221.400 94.200 ;
        RECT 222.400 94.400 223.000 95.000 ;
        RECT 217.200 91.600 218.000 93.200 ;
        RECT 218.800 91.600 219.600 93.200 ;
        RECT 220.400 93.000 221.800 93.800 ;
        RECT 222.400 93.600 224.400 94.400 ;
        RECT 220.400 91.000 221.000 93.000 ;
        RECT 191.600 89.400 192.400 89.600 ;
        RECT 187.000 89.000 192.400 89.400 ;
        RECT 186.200 88.800 192.400 89.000 ;
        RECT 193.400 89.000 202.000 89.600 ;
        RECT 183.600 88.000 185.200 88.800 ;
        RECT 186.200 88.200 187.600 88.800 ;
        RECT 193.400 88.200 194.000 89.000 ;
        RECT 201.200 88.800 202.000 89.000 ;
        RECT 204.400 89.000 213.400 89.600 ;
        RECT 204.400 88.800 205.200 89.000 ;
        RECT 184.600 87.600 185.200 88.000 ;
        RECT 188.200 87.600 194.000 88.200 ;
        RECT 194.600 87.600 197.200 88.400 ;
        RECT 182.000 86.800 184.000 87.400 ;
        RECT 184.600 86.800 188.800 87.600 ;
        RECT 183.400 86.200 184.000 86.800 ;
        RECT 183.400 85.600 184.400 86.200 ;
        RECT 183.600 82.200 184.400 85.600 ;
        RECT 186.800 82.200 187.600 86.800 ;
        RECT 190.000 82.200 190.800 85.000 ;
        RECT 191.600 82.200 192.400 85.000 ;
        RECT 193.200 82.200 194.000 87.000 ;
        RECT 196.400 82.200 197.200 87.000 ;
        RECT 199.600 82.200 200.400 88.400 ;
        RECT 207.600 87.600 210.200 88.400 ;
        RECT 202.800 86.800 207.000 87.600 ;
        RECT 201.200 82.200 202.000 85.000 ;
        RECT 202.800 82.200 203.600 85.000 ;
        RECT 204.400 82.200 205.200 85.000 ;
        RECT 207.600 82.200 208.400 87.600 ;
        RECT 212.800 87.400 213.400 89.000 ;
        RECT 210.800 86.800 213.400 87.400 ;
        RECT 214.000 90.000 215.000 90.800 ;
        RECT 217.200 90.400 221.000 91.000 ;
        RECT 210.800 82.200 211.600 86.800 ;
        RECT 214.000 82.200 214.800 90.000 ;
        RECT 217.200 87.000 217.800 90.400 ;
        RECT 222.400 89.800 223.000 93.600 ;
        RECT 223.600 90.800 224.400 92.400 ;
        RECT 221.400 89.200 223.000 89.800 ;
        RECT 217.200 83.000 218.000 87.000 ;
        RECT 221.400 82.200 222.200 89.200 ;
        RECT 4.400 72.400 5.200 79.800 ;
        RECT 9.200 72.400 10.000 79.800 ;
        RECT 3.000 71.800 5.200 72.400 ;
        RECT 7.800 71.800 10.000 72.400 ;
        RECT 12.400 72.000 13.200 79.800 ;
        RECT 15.600 75.200 16.400 79.800 ;
        RECT 3.000 71.200 3.600 71.800 ;
        RECT 7.800 71.200 8.400 71.800 ;
        RECT 2.400 70.400 3.600 71.200 ;
        RECT 7.200 70.400 8.400 71.200 ;
        RECT 12.200 71.200 13.200 72.000 ;
        RECT 13.800 74.600 16.400 75.200 ;
        RECT 13.800 73.000 14.400 74.600 ;
        RECT 18.800 74.400 19.600 79.800 ;
        RECT 22.000 77.000 22.800 79.800 ;
        RECT 23.600 77.000 24.400 79.800 ;
        RECT 25.200 77.000 26.000 79.800 ;
        RECT 20.200 74.400 24.400 75.200 ;
        RECT 17.000 73.600 19.600 74.400 ;
        RECT 26.800 73.600 27.600 79.800 ;
        RECT 30.000 75.000 30.800 79.800 ;
        RECT 33.200 75.000 34.000 79.800 ;
        RECT 34.800 77.000 35.600 79.800 ;
        RECT 36.400 77.000 37.200 79.800 ;
        RECT 39.600 75.200 40.400 79.800 ;
        RECT 42.800 76.400 43.600 79.800 ;
        RECT 42.800 75.800 43.800 76.400 ;
        RECT 43.200 75.200 43.800 75.800 ;
        RECT 38.400 74.400 42.600 75.200 ;
        RECT 43.200 74.600 45.200 75.200 ;
        RECT 30.000 73.600 32.600 74.400 ;
        RECT 33.200 73.800 39.000 74.400 ;
        RECT 42.000 74.000 42.600 74.400 ;
        RECT 22.000 73.000 22.800 73.200 ;
        RECT 13.800 72.400 22.800 73.000 ;
        RECT 25.200 73.000 26.000 73.200 ;
        RECT 33.200 73.000 33.800 73.800 ;
        RECT 39.600 73.200 41.000 73.800 ;
        RECT 42.000 73.200 43.600 74.000 ;
        RECT 25.200 72.400 33.800 73.000 ;
        RECT 34.800 73.000 41.000 73.200 ;
        RECT 34.800 72.600 40.200 73.000 ;
        RECT 34.800 72.400 35.600 72.600 ;
        RECT 3.000 67.400 3.600 70.400 ;
        RECT 4.400 68.800 5.200 70.400 ;
        RECT 7.800 67.400 8.400 70.400 ;
        RECT 9.200 68.800 10.000 70.400 ;
        RECT 3.000 66.800 5.200 67.400 ;
        RECT 7.800 66.800 10.000 67.400 ;
        RECT 4.400 62.200 5.200 66.800 ;
        RECT 9.200 62.200 10.000 66.800 ;
        RECT 12.200 66.800 13.000 71.200 ;
        RECT 13.800 70.600 14.400 72.400 ;
        RECT 13.600 70.000 14.400 70.600 ;
        RECT 20.400 70.000 43.800 70.600 ;
        RECT 13.600 68.000 14.200 70.000 ;
        RECT 20.400 69.400 21.200 70.000 ;
        RECT 38.000 69.600 38.800 70.000 ;
        RECT 43.000 69.800 43.800 70.000 ;
        RECT 14.800 68.600 18.600 69.400 ;
        RECT 13.600 67.400 14.800 68.000 ;
        RECT 12.200 66.000 13.200 66.800 ;
        RECT 12.400 62.200 13.200 66.000 ;
        RECT 14.000 62.200 14.800 67.400 ;
        RECT 17.800 67.400 18.600 68.600 ;
        RECT 17.800 66.800 19.600 67.400 ;
        RECT 18.800 66.200 19.600 66.800 ;
        RECT 23.600 66.400 24.400 69.200 ;
        RECT 26.800 68.600 30.000 69.400 ;
        RECT 33.800 68.600 35.800 69.400 ;
        RECT 44.400 69.000 45.200 74.600 ;
        RECT 26.400 67.800 27.200 68.000 ;
        RECT 26.400 67.200 30.800 67.800 ;
        RECT 30.000 67.000 30.800 67.200 ;
        RECT 31.600 66.800 32.400 68.400 ;
        RECT 18.800 65.400 21.200 66.200 ;
        RECT 23.600 65.600 24.600 66.400 ;
        RECT 27.600 65.600 29.200 66.400 ;
        RECT 30.000 66.200 30.800 66.400 ;
        RECT 33.800 66.200 34.600 68.600 ;
        RECT 36.400 68.200 45.200 69.000 ;
        RECT 39.800 66.800 42.800 67.600 ;
        RECT 39.800 66.200 40.600 66.800 ;
        RECT 30.000 65.600 34.600 66.200 ;
        RECT 20.400 62.200 21.200 65.400 ;
        RECT 38.000 65.400 40.600 66.200 ;
        RECT 22.000 62.200 22.800 65.000 ;
        RECT 23.600 62.200 24.400 65.000 ;
        RECT 25.200 62.200 26.000 65.000 ;
        RECT 26.800 62.200 27.600 65.000 ;
        RECT 30.000 62.200 30.800 65.000 ;
        RECT 33.200 62.200 34.000 65.000 ;
        RECT 34.800 62.200 35.600 65.000 ;
        RECT 36.400 62.200 37.200 65.000 ;
        RECT 38.000 62.200 38.800 65.400 ;
        RECT 44.400 62.200 45.200 68.200 ;
        RECT 47.600 64.800 48.400 66.400 ;
        RECT 49.200 62.200 50.000 79.800 ;
        RECT 50.800 75.800 51.600 79.800 ;
        RECT 51.000 75.600 51.600 75.800 ;
        RECT 54.000 75.800 54.800 79.800 ;
        RECT 58.800 75.800 59.600 79.800 ;
        RECT 54.000 75.600 54.700 75.800 ;
        RECT 51.000 75.000 54.700 75.600 ;
        RECT 59.000 75.600 59.600 75.800 ;
        RECT 62.000 75.800 62.800 79.800 ;
        RECT 62.000 75.600 62.600 75.800 ;
        RECT 59.000 75.000 62.600 75.600 ;
        RECT 51.000 72.400 51.600 75.000 ;
        RECT 52.400 72.800 53.200 74.400 ;
        RECT 54.100 74.300 54.700 75.000 ;
        RECT 60.400 74.300 61.200 74.400 ;
        RECT 54.100 73.700 61.200 74.300 ;
        RECT 50.800 71.600 51.600 72.400 ;
        RECT 51.000 68.400 51.600 71.600 ;
        RECT 55.600 70.800 56.400 72.400 ;
        RECT 57.200 70.800 58.000 72.400 ;
        RECT 60.400 71.600 61.200 73.700 ;
        RECT 62.000 72.400 62.600 75.000 ;
        RECT 65.800 74.400 66.600 79.800 ;
        RECT 64.400 73.600 65.200 74.400 ;
        RECT 65.800 73.600 67.600 74.400 ;
        RECT 64.400 72.400 65.000 73.600 ;
        RECT 65.800 72.400 66.600 73.600 ;
        RECT 62.000 71.600 62.800 72.400 ;
        RECT 63.600 71.800 65.000 72.400 ;
        RECT 65.600 71.800 66.600 72.400 ;
        RECT 72.600 72.400 73.400 79.800 ;
        RECT 74.000 73.600 74.800 74.400 ;
        RECT 74.200 72.400 74.800 73.600 ;
        RECT 72.600 71.800 73.600 72.400 ;
        RECT 74.200 71.800 75.600 72.400 ;
        RECT 63.600 71.600 64.400 71.800 ;
        RECT 53.200 69.600 54.800 70.400 ;
        RECT 58.800 69.600 60.400 70.400 ;
        RECT 62.000 68.400 62.600 71.600 ;
        RECT 65.600 68.400 66.200 71.800 ;
        RECT 66.800 70.300 67.600 70.400 ;
        RECT 71.600 70.300 72.400 70.400 ;
        RECT 66.800 69.700 72.400 70.300 ;
        RECT 66.800 68.800 67.600 69.700 ;
        RECT 71.600 68.800 72.400 69.700 ;
        RECT 73.000 70.300 73.600 71.800 ;
        RECT 74.800 71.600 75.600 71.800 ;
        RECT 76.400 71.600 77.200 73.200 ;
        RECT 76.500 70.300 77.100 71.600 ;
        RECT 73.000 69.700 77.100 70.300 ;
        RECT 78.000 70.300 78.800 79.800 ;
        RECT 82.800 72.800 83.600 79.800 ;
        RECT 82.600 71.600 83.600 72.800 ;
        RECT 86.000 72.400 86.800 79.800 ;
        RECT 90.800 76.400 91.600 79.800 ;
        RECT 90.600 75.800 91.600 76.400 ;
        RECT 90.600 75.200 91.200 75.800 ;
        RECT 94.000 75.200 94.800 79.800 ;
        RECT 97.200 77.000 98.000 79.800 ;
        RECT 98.800 77.000 99.600 79.800 ;
        RECT 84.200 71.800 86.800 72.400 ;
        RECT 89.200 74.600 91.200 75.200 ;
        RECT 81.200 70.300 82.000 70.400 ;
        RECT 78.000 69.700 82.000 70.300 ;
        RECT 73.000 68.400 73.600 69.700 ;
        RECT 51.000 68.200 52.600 68.400 ;
        RECT 61.000 68.200 62.600 68.400 ;
        RECT 51.000 67.800 52.800 68.200 ;
        RECT 52.000 62.200 52.800 67.800 ;
        RECT 60.800 67.800 62.600 68.200 ;
        RECT 60.800 62.200 61.600 67.800 ;
        RECT 63.600 67.600 66.200 68.400 ;
        RECT 68.400 68.200 69.200 68.400 ;
        RECT 67.600 67.600 69.200 68.200 ;
        RECT 70.000 68.200 70.800 68.400 ;
        RECT 70.000 67.600 71.600 68.200 ;
        RECT 73.000 67.600 75.600 68.400 ;
        RECT 63.800 66.200 64.400 67.600 ;
        RECT 67.600 67.200 68.400 67.600 ;
        RECT 70.800 67.200 71.600 67.600 ;
        RECT 65.400 66.200 69.000 66.600 ;
        RECT 70.200 66.200 73.800 66.600 ;
        RECT 74.800 66.200 75.400 67.600 ;
        RECT 78.000 66.200 78.800 69.700 ;
        RECT 81.200 69.600 82.000 69.700 ;
        RECT 82.600 68.400 83.200 71.600 ;
        RECT 84.200 69.800 84.800 71.800 ;
        RECT 83.800 69.000 84.800 69.800 ;
        RECT 79.600 66.800 80.400 68.400 ;
        RECT 82.600 67.600 83.600 68.400 ;
        RECT 63.600 62.200 64.400 66.200 ;
        RECT 65.200 66.000 69.200 66.200 ;
        RECT 65.200 62.200 66.000 66.000 ;
        RECT 68.400 62.200 69.200 66.000 ;
        RECT 70.000 66.000 74.000 66.200 ;
        RECT 70.000 62.200 70.800 66.000 ;
        RECT 73.200 62.200 74.000 66.000 ;
        RECT 74.800 62.200 75.600 66.200 ;
        RECT 77.000 65.600 78.800 66.200 ;
        RECT 82.600 66.200 83.200 67.600 ;
        RECT 84.200 67.400 84.800 69.000 ;
        RECT 85.800 69.600 86.800 70.400 ;
        RECT 85.800 68.800 86.600 69.600 ;
        RECT 89.200 69.000 90.000 74.600 ;
        RECT 91.800 74.400 96.000 75.200 ;
        RECT 100.400 75.000 101.200 79.800 ;
        RECT 103.600 75.000 104.400 79.800 ;
        RECT 91.800 74.000 92.400 74.400 ;
        RECT 90.800 73.200 92.400 74.000 ;
        RECT 95.400 73.800 101.200 74.400 ;
        RECT 93.400 73.200 94.800 73.800 ;
        RECT 93.400 73.000 99.600 73.200 ;
        RECT 94.200 72.600 99.600 73.000 ;
        RECT 98.800 72.400 99.600 72.600 ;
        RECT 100.600 73.000 101.200 73.800 ;
        RECT 101.800 73.600 104.400 74.400 ;
        RECT 106.800 73.600 107.600 79.800 ;
        RECT 108.400 77.000 109.200 79.800 ;
        RECT 110.000 77.000 110.800 79.800 ;
        RECT 111.600 77.000 112.400 79.800 ;
        RECT 110.000 74.400 114.200 75.200 ;
        RECT 114.800 74.400 115.600 79.800 ;
        RECT 118.000 75.200 118.800 79.800 ;
        RECT 118.000 74.600 120.600 75.200 ;
        RECT 114.800 73.600 117.400 74.400 ;
        RECT 108.400 73.000 109.200 73.200 ;
        RECT 100.600 72.400 109.200 73.000 ;
        RECT 111.600 73.000 112.400 73.200 ;
        RECT 120.000 73.000 120.600 74.600 ;
        RECT 111.600 72.400 120.600 73.000 ;
        RECT 120.000 70.600 120.600 72.400 ;
        RECT 121.200 72.000 122.000 79.800 ;
        RECT 127.600 76.400 128.400 79.800 ;
        RECT 127.400 75.800 128.400 76.400 ;
        RECT 127.400 75.200 128.000 75.800 ;
        RECT 130.800 75.200 131.600 79.800 ;
        RECT 134.000 77.000 134.800 79.800 ;
        RECT 135.600 77.000 136.400 79.800 ;
        RECT 126.000 74.600 128.000 75.200 ;
        RECT 121.200 71.200 122.200 72.000 ;
        RECT 90.600 70.000 114.000 70.600 ;
        RECT 120.000 70.000 120.800 70.600 ;
        RECT 90.600 69.800 91.400 70.000 ;
        RECT 92.400 69.600 93.200 70.000 ;
        RECT 94.000 69.600 94.800 70.000 ;
        RECT 95.600 69.600 96.400 70.000 ;
        RECT 113.200 69.400 114.000 70.000 ;
        RECT 89.200 68.200 98.000 69.000 ;
        RECT 98.600 68.600 100.600 69.400 ;
        RECT 104.400 68.600 107.600 69.400 ;
        RECT 84.200 66.800 86.800 67.400 ;
        RECT 82.600 65.600 83.600 66.200 ;
        RECT 77.000 62.200 77.800 65.600 ;
        RECT 82.800 62.200 83.600 65.600 ;
        RECT 86.000 62.200 86.800 66.800 ;
        RECT 89.200 62.200 90.000 68.200 ;
        RECT 91.600 66.800 94.600 67.600 ;
        RECT 93.800 66.200 94.600 66.800 ;
        RECT 99.800 66.200 100.600 68.600 ;
        RECT 102.000 66.800 102.800 68.400 ;
        RECT 107.200 67.800 108.000 68.000 ;
        RECT 103.600 67.200 108.000 67.800 ;
        RECT 103.600 67.000 104.400 67.200 ;
        RECT 110.000 66.400 110.800 69.200 ;
        RECT 115.800 68.600 119.600 69.400 ;
        RECT 115.800 67.400 116.600 68.600 ;
        RECT 120.200 68.000 120.800 70.000 ;
        RECT 103.600 66.200 104.400 66.400 ;
        RECT 93.800 65.400 96.400 66.200 ;
        RECT 99.800 65.600 104.400 66.200 ;
        RECT 105.200 65.600 106.800 66.400 ;
        RECT 109.800 65.600 110.800 66.400 ;
        RECT 114.800 66.800 116.600 67.400 ;
        RECT 119.600 67.400 120.800 68.000 ;
        RECT 114.800 66.200 115.600 66.800 ;
        RECT 95.600 62.200 96.400 65.400 ;
        RECT 113.200 65.400 115.600 66.200 ;
        RECT 97.200 62.200 98.000 65.000 ;
        RECT 98.800 62.200 99.600 65.000 ;
        RECT 100.400 62.200 101.200 65.000 ;
        RECT 103.600 62.200 104.400 65.000 ;
        RECT 106.800 62.200 107.600 65.000 ;
        RECT 108.400 62.200 109.200 65.000 ;
        RECT 110.000 62.200 110.800 65.000 ;
        RECT 111.600 62.200 112.400 65.000 ;
        RECT 113.200 62.200 114.000 65.400 ;
        RECT 119.600 62.200 120.400 67.400 ;
        RECT 121.400 66.800 122.200 71.200 ;
        RECT 121.200 66.000 122.200 66.800 ;
        RECT 126.000 69.000 126.800 74.600 ;
        RECT 128.600 74.400 132.800 75.200 ;
        RECT 137.200 75.000 138.000 79.800 ;
        RECT 140.400 75.000 141.200 79.800 ;
        RECT 128.600 74.000 129.200 74.400 ;
        RECT 127.600 73.200 129.200 74.000 ;
        RECT 132.200 73.800 138.000 74.400 ;
        RECT 130.200 73.200 131.600 73.800 ;
        RECT 130.200 73.000 136.400 73.200 ;
        RECT 131.000 72.600 136.400 73.000 ;
        RECT 135.600 72.400 136.400 72.600 ;
        RECT 137.400 73.000 138.000 73.800 ;
        RECT 138.600 73.600 141.200 74.400 ;
        RECT 143.600 73.600 144.400 79.800 ;
        RECT 145.200 77.000 146.000 79.800 ;
        RECT 146.800 77.000 147.600 79.800 ;
        RECT 148.400 77.000 149.200 79.800 ;
        RECT 146.800 74.400 151.000 75.200 ;
        RECT 151.600 74.400 152.400 79.800 ;
        RECT 154.800 75.200 155.600 79.800 ;
        RECT 154.800 74.600 157.400 75.200 ;
        RECT 151.600 73.600 154.200 74.400 ;
        RECT 145.200 73.000 146.000 73.200 ;
        RECT 137.400 72.400 146.000 73.000 ;
        RECT 148.400 73.000 149.200 73.200 ;
        RECT 156.800 73.000 157.400 74.600 ;
        RECT 148.400 72.400 157.400 73.000 ;
        RECT 156.800 70.600 157.400 72.400 ;
        RECT 158.000 72.000 158.800 79.800 ;
        RECT 162.800 76.400 163.600 79.800 ;
        RECT 162.600 75.800 163.600 76.400 ;
        RECT 162.600 75.200 163.200 75.800 ;
        RECT 166.000 75.200 166.800 79.800 ;
        RECT 169.200 77.000 170.000 79.800 ;
        RECT 170.800 77.000 171.600 79.800 ;
        RECT 161.200 74.600 163.200 75.200 ;
        RECT 158.000 71.200 159.000 72.000 ;
        RECT 127.400 70.000 150.800 70.600 ;
        RECT 156.800 70.000 157.600 70.600 ;
        RECT 127.400 69.800 128.200 70.000 ;
        RECT 130.800 69.600 131.600 70.000 ;
        RECT 132.400 69.600 133.200 70.000 ;
        RECT 150.000 69.400 150.800 70.000 ;
        RECT 126.000 68.200 134.800 69.000 ;
        RECT 135.400 68.600 137.400 69.400 ;
        RECT 141.200 68.600 144.400 69.400 ;
        RECT 121.200 62.200 122.000 66.000 ;
        RECT 126.000 62.200 126.800 68.200 ;
        RECT 128.400 66.800 131.400 67.600 ;
        RECT 130.600 66.200 131.400 66.800 ;
        RECT 136.600 66.200 137.400 68.600 ;
        RECT 138.800 66.800 139.600 68.400 ;
        RECT 144.000 67.800 144.800 68.000 ;
        RECT 140.400 67.200 144.800 67.800 ;
        RECT 140.400 67.000 141.200 67.200 ;
        RECT 146.800 66.400 147.600 69.200 ;
        RECT 152.600 68.600 156.400 69.400 ;
        RECT 152.600 67.400 153.400 68.600 ;
        RECT 157.000 68.000 157.600 70.000 ;
        RECT 140.400 66.200 141.200 66.400 ;
        RECT 130.600 65.400 133.200 66.200 ;
        RECT 136.600 65.600 141.200 66.200 ;
        RECT 142.000 65.600 143.600 66.400 ;
        RECT 146.600 65.600 147.600 66.400 ;
        RECT 151.600 66.800 153.400 67.400 ;
        RECT 156.400 67.400 157.600 68.000 ;
        RECT 151.600 66.200 152.400 66.800 ;
        RECT 132.400 62.200 133.200 65.400 ;
        RECT 150.000 65.400 152.400 66.200 ;
        RECT 134.000 62.200 134.800 65.000 ;
        RECT 135.600 62.200 136.400 65.000 ;
        RECT 137.200 62.200 138.000 65.000 ;
        RECT 140.400 62.200 141.200 65.000 ;
        RECT 143.600 62.200 144.400 65.000 ;
        RECT 145.200 62.200 146.000 65.000 ;
        RECT 146.800 62.200 147.600 65.000 ;
        RECT 148.400 62.200 149.200 65.000 ;
        RECT 150.000 62.200 150.800 65.400 ;
        RECT 156.400 62.200 157.200 67.400 ;
        RECT 158.200 66.800 159.000 71.200 ;
        RECT 158.000 66.000 159.000 66.800 ;
        RECT 161.200 69.000 162.000 74.600 ;
        RECT 163.800 74.400 168.000 75.200 ;
        RECT 172.400 75.000 173.200 79.800 ;
        RECT 175.600 75.000 176.400 79.800 ;
        RECT 163.800 74.000 164.400 74.400 ;
        RECT 162.800 73.200 164.400 74.000 ;
        RECT 167.400 73.800 173.200 74.400 ;
        RECT 165.400 73.200 166.800 73.800 ;
        RECT 165.400 73.000 171.600 73.200 ;
        RECT 166.200 72.600 171.600 73.000 ;
        RECT 170.800 72.400 171.600 72.600 ;
        RECT 172.600 73.000 173.200 73.800 ;
        RECT 173.800 73.600 176.400 74.400 ;
        RECT 178.800 73.600 179.600 79.800 ;
        RECT 180.400 77.000 181.200 79.800 ;
        RECT 182.000 77.000 182.800 79.800 ;
        RECT 183.600 77.000 184.400 79.800 ;
        RECT 182.000 74.400 186.200 75.200 ;
        RECT 186.800 74.400 187.600 79.800 ;
        RECT 190.000 75.200 190.800 79.800 ;
        RECT 190.000 74.600 192.600 75.200 ;
        RECT 186.800 73.600 189.400 74.400 ;
        RECT 180.400 73.000 181.200 73.200 ;
        RECT 172.600 72.400 181.200 73.000 ;
        RECT 183.600 73.000 184.400 73.200 ;
        RECT 192.000 73.000 192.600 74.600 ;
        RECT 183.600 72.400 192.600 73.000 ;
        RECT 192.000 70.600 192.600 72.400 ;
        RECT 193.200 72.000 194.000 79.800 ;
        RECT 193.200 71.200 194.200 72.000 ;
        RECT 162.600 70.000 186.000 70.600 ;
        RECT 192.000 70.000 192.800 70.600 ;
        RECT 162.600 69.800 163.400 70.000 ;
        RECT 164.400 69.600 165.200 70.000 ;
        RECT 167.600 69.600 168.400 70.000 ;
        RECT 185.200 69.400 186.000 70.000 ;
        RECT 161.200 68.200 170.000 69.000 ;
        RECT 170.600 68.600 172.600 69.400 ;
        RECT 176.400 68.600 179.600 69.400 ;
        RECT 158.000 62.200 158.800 66.000 ;
        RECT 161.200 62.200 162.000 68.200 ;
        RECT 163.600 66.800 166.600 67.600 ;
        RECT 165.800 66.200 166.600 66.800 ;
        RECT 171.800 66.200 172.600 68.600 ;
        RECT 174.000 66.800 174.800 68.400 ;
        RECT 179.200 67.800 180.000 68.000 ;
        RECT 175.600 67.200 180.000 67.800 ;
        RECT 175.600 67.000 176.400 67.200 ;
        RECT 182.000 66.400 182.800 69.200 ;
        RECT 187.800 68.600 191.600 69.400 ;
        RECT 187.800 67.400 188.600 68.600 ;
        RECT 192.200 68.000 192.800 70.000 ;
        RECT 175.600 66.200 176.400 66.400 ;
        RECT 165.800 65.400 168.400 66.200 ;
        RECT 171.800 65.600 176.400 66.200 ;
        RECT 177.200 65.600 178.800 66.400 ;
        RECT 181.800 65.600 182.800 66.400 ;
        RECT 186.800 66.800 188.600 67.400 ;
        RECT 191.600 67.400 192.800 68.000 ;
        RECT 186.800 66.200 187.600 66.800 ;
        RECT 167.600 62.200 168.400 65.400 ;
        RECT 185.200 65.400 187.600 66.200 ;
        RECT 169.200 62.200 170.000 65.000 ;
        RECT 170.800 62.200 171.600 65.000 ;
        RECT 172.400 62.200 173.200 65.000 ;
        RECT 175.600 62.200 176.400 65.000 ;
        RECT 178.800 62.200 179.600 65.000 ;
        RECT 180.400 62.200 181.200 65.000 ;
        RECT 182.000 62.200 182.800 65.000 ;
        RECT 183.600 62.200 184.400 65.000 ;
        RECT 185.200 62.200 186.000 65.400 ;
        RECT 191.600 62.200 192.400 67.400 ;
        RECT 193.400 66.800 194.200 71.200 ;
        RECT 193.200 66.300 194.200 66.800 ;
        RECT 199.600 70.300 200.400 79.800 ;
        RECT 201.200 72.400 202.000 79.800 ;
        RECT 204.400 72.400 205.200 79.800 ;
        RECT 201.200 71.800 205.200 72.400 ;
        RECT 206.000 71.800 206.800 79.800 ;
        RECT 210.200 72.600 211.000 79.800 ;
        RECT 209.200 71.800 211.000 72.600 ;
        RECT 212.400 72.400 213.200 79.800 ;
        RECT 217.200 72.400 218.000 79.800 ;
        RECT 212.400 71.800 214.600 72.400 ;
        RECT 217.200 71.800 219.400 72.400 ;
        RECT 202.000 70.400 202.800 70.800 ;
        RECT 206.000 70.400 206.600 71.800 ;
        RECT 201.200 70.300 202.800 70.400 ;
        RECT 199.600 69.800 202.800 70.300 ;
        RECT 204.400 69.800 206.800 70.400 ;
        RECT 199.600 69.700 202.000 69.800 ;
        RECT 198.000 66.300 198.800 66.400 ;
        RECT 193.200 65.700 198.800 66.300 ;
        RECT 193.200 62.200 194.000 65.700 ;
        RECT 198.000 64.800 198.800 65.700 ;
        RECT 199.600 62.200 200.400 69.700 ;
        RECT 201.200 69.600 202.000 69.700 ;
        RECT 202.800 67.600 203.600 69.200 ;
        RECT 204.400 66.400 205.000 69.800 ;
        RECT 206.000 69.600 206.800 69.800 ;
        RECT 209.400 68.400 210.000 71.800 ;
        RECT 214.000 71.200 214.600 71.800 ;
        RECT 218.800 71.200 219.400 71.800 ;
        RECT 210.800 69.600 211.600 71.200 ;
        RECT 214.000 70.400 215.200 71.200 ;
        RECT 218.800 70.400 220.000 71.200 ;
        RECT 212.400 68.800 213.200 70.400 ;
        RECT 209.200 68.300 210.000 68.400 ;
        RECT 206.100 67.700 210.000 68.300 ;
        RECT 206.100 66.400 206.700 67.700 ;
        RECT 209.200 67.600 210.000 67.700 ;
        RECT 204.400 62.200 205.200 66.400 ;
        RECT 206.000 65.600 206.800 66.400 ;
        RECT 205.800 64.800 206.600 65.600 ;
        RECT 207.600 64.800 208.400 66.400 ;
        RECT 209.400 64.200 210.000 67.600 ;
        RECT 214.000 67.400 214.600 70.400 ;
        RECT 217.200 68.800 218.000 70.400 ;
        RECT 218.800 67.400 219.400 70.400 ;
        RECT 209.200 62.200 210.000 64.200 ;
        RECT 212.400 66.800 214.600 67.400 ;
        RECT 217.200 66.800 219.400 67.400 ;
        RECT 212.400 62.200 213.200 66.800 ;
        RECT 217.200 62.200 218.000 66.800 ;
        RECT 4.400 55.200 5.200 59.800 ;
        RECT 7.600 56.000 8.400 59.800 ;
        RECT 3.000 54.600 5.200 55.200 ;
        RECT 7.400 55.200 8.400 56.000 ;
        RECT 3.000 51.600 3.600 54.600 ;
        RECT 4.400 52.300 5.200 53.200 ;
        RECT 7.400 52.300 8.200 55.200 ;
        RECT 9.200 54.600 10.000 59.800 ;
        RECT 15.600 56.600 16.400 59.800 ;
        RECT 17.200 57.000 18.000 59.800 ;
        RECT 18.800 57.000 19.600 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 22.000 57.000 22.800 59.800 ;
        RECT 25.200 57.000 26.000 59.800 ;
        RECT 28.400 57.000 29.200 59.800 ;
        RECT 30.000 57.000 30.800 59.800 ;
        RECT 31.600 57.000 32.400 59.800 ;
        RECT 14.000 55.800 16.400 56.600 ;
        RECT 33.200 56.600 34.000 59.800 ;
        RECT 14.000 55.200 14.800 55.800 ;
        RECT 4.400 51.700 8.200 52.300 ;
        RECT 4.400 51.600 5.200 51.700 ;
        RECT 2.400 50.800 3.600 51.600 ;
        RECT 3.000 50.200 3.600 50.800 ;
        RECT 7.400 50.800 8.200 51.700 ;
        RECT 8.800 54.000 10.000 54.600 ;
        RECT 13.000 54.600 14.800 55.200 ;
        RECT 18.800 55.600 19.800 56.400 ;
        RECT 22.800 55.600 24.400 56.400 ;
        RECT 25.200 55.800 29.800 56.400 ;
        RECT 33.200 55.800 35.800 56.600 ;
        RECT 25.200 55.600 26.000 55.800 ;
        RECT 8.800 52.000 9.400 54.000 ;
        RECT 13.000 53.400 13.800 54.600 ;
        RECT 10.000 52.600 13.800 53.400 ;
        RECT 18.800 52.800 19.600 55.600 ;
        RECT 25.200 54.800 26.000 55.000 ;
        RECT 21.600 54.200 26.000 54.800 ;
        RECT 21.600 54.000 22.400 54.200 ;
        RECT 26.800 53.600 27.600 55.200 ;
        RECT 29.000 53.400 29.800 55.800 ;
        RECT 35.000 55.200 35.800 55.800 ;
        RECT 35.000 54.400 38.000 55.200 ;
        RECT 39.600 53.800 40.400 59.800 ;
        RECT 41.200 56.300 42.000 56.400 ;
        RECT 42.800 56.300 43.600 57.200 ;
        RECT 41.200 55.700 43.600 56.300 ;
        RECT 41.200 55.600 42.000 55.700 ;
        RECT 42.800 55.600 43.600 55.700 ;
        RECT 22.000 52.600 25.200 53.400 ;
        RECT 29.000 52.600 31.000 53.400 ;
        RECT 31.600 53.000 40.400 53.800 ;
        RECT 15.600 52.000 16.400 52.600 ;
        RECT 33.200 52.000 34.000 52.400 ;
        RECT 34.800 52.000 35.600 52.400 ;
        RECT 38.000 52.200 38.800 52.400 ;
        RECT 38.000 52.000 39.000 52.200 ;
        RECT 8.800 51.400 9.600 52.000 ;
        RECT 15.600 51.400 39.000 52.000 ;
        RECT 3.000 49.600 5.200 50.200 ;
        RECT 7.400 50.000 8.400 50.800 ;
        RECT 4.400 42.200 5.200 49.600 ;
        RECT 7.600 42.200 8.400 50.000 ;
        RECT 9.000 49.600 9.600 51.400 ;
        RECT 9.000 49.000 18.000 49.600 ;
        RECT 9.000 47.400 9.600 49.000 ;
        RECT 17.200 48.800 18.000 49.000 ;
        RECT 20.400 49.000 29.000 49.600 ;
        RECT 20.400 48.800 21.200 49.000 ;
        RECT 12.200 47.600 14.800 48.400 ;
        RECT 9.000 46.800 11.600 47.400 ;
        RECT 10.800 42.200 11.600 46.800 ;
        RECT 14.000 42.200 14.800 47.600 ;
        RECT 15.400 46.800 19.600 47.600 ;
        RECT 17.200 42.200 18.000 45.000 ;
        RECT 18.800 42.200 19.600 45.000 ;
        RECT 20.400 42.200 21.200 45.000 ;
        RECT 22.000 42.200 22.800 48.400 ;
        RECT 25.200 47.600 27.800 48.400 ;
        RECT 28.400 48.200 29.000 49.000 ;
        RECT 30.000 49.400 30.800 49.600 ;
        RECT 30.000 49.000 35.400 49.400 ;
        RECT 30.000 48.800 36.200 49.000 ;
        RECT 34.800 48.200 36.200 48.800 ;
        RECT 28.400 47.600 34.200 48.200 ;
        RECT 37.200 48.000 38.800 48.800 ;
        RECT 37.200 47.600 37.800 48.000 ;
        RECT 25.200 42.200 26.000 47.000 ;
        RECT 28.400 42.200 29.200 47.000 ;
        RECT 33.600 46.800 37.800 47.600 ;
        RECT 39.600 47.400 40.400 53.000 ;
        RECT 38.400 46.800 40.400 47.400 ;
        RECT 44.400 54.300 45.200 59.800 ;
        RECT 46.200 56.400 47.000 57.200 ;
        RECT 46.000 55.600 46.800 56.400 ;
        RECT 47.600 55.800 48.400 59.800 ;
        RECT 46.000 54.300 46.800 54.400 ;
        RECT 44.400 53.700 46.800 54.300 ;
        RECT 30.000 42.200 30.800 45.000 ;
        RECT 31.600 42.200 32.400 45.000 ;
        RECT 34.800 42.200 35.600 46.800 ;
        RECT 38.400 46.200 39.000 46.800 ;
        RECT 38.000 45.600 39.000 46.200 ;
        RECT 38.000 42.200 38.800 45.600 ;
        RECT 44.400 42.200 45.200 53.700 ;
        RECT 46.000 53.600 46.800 53.700 ;
        RECT 46.000 52.200 46.800 52.400 ;
        RECT 47.800 52.200 48.400 55.800 ;
        RECT 49.200 52.800 50.000 54.400 ;
        RECT 50.800 52.200 51.600 52.400 ;
        RECT 46.000 51.600 48.400 52.200 ;
        RECT 50.000 51.600 51.600 52.200 ;
        RECT 46.200 50.200 46.800 51.600 ;
        RECT 50.000 51.200 50.800 51.600 ;
        RECT 46.000 42.200 46.800 50.200 ;
        RECT 47.600 49.600 51.600 50.200 ;
        RECT 47.600 42.200 48.400 49.600 ;
        RECT 50.800 42.200 51.600 49.600 ;
        RECT 52.400 42.200 53.200 59.800 ;
        RECT 54.000 55.600 54.800 57.200 ;
        RECT 59.200 54.200 60.000 59.800 ;
        RECT 59.200 53.800 61.000 54.200 ;
        RECT 59.400 53.600 61.000 53.800 ;
        RECT 57.200 51.600 58.800 52.400 ;
        RECT 54.000 50.300 54.800 50.400 ;
        RECT 55.600 50.300 56.400 51.200 ;
        RECT 54.000 49.700 56.400 50.300 ;
        RECT 54.000 49.600 54.800 49.700 ;
        RECT 55.600 49.600 56.400 49.700 ;
        RECT 60.400 50.400 61.000 53.600 ;
        RECT 60.400 49.600 61.200 50.400 ;
        RECT 58.800 47.600 59.600 49.200 ;
        RECT 60.400 47.000 61.000 49.600 ;
        RECT 57.400 46.400 61.000 47.000 ;
        RECT 57.200 42.200 58.000 46.400 ;
        RECT 60.400 46.200 61.000 46.400 ;
        RECT 60.400 42.200 61.200 46.200 ;
        RECT 62.000 42.200 62.800 59.800 ;
        RECT 63.600 55.600 64.400 57.200 ;
        RECT 66.800 56.000 67.600 59.800 ;
        RECT 66.600 55.200 67.600 56.000 ;
        RECT 66.600 50.800 67.400 55.200 ;
        RECT 68.400 54.600 69.200 59.800 ;
        RECT 74.800 56.600 75.600 59.800 ;
        RECT 76.400 57.000 77.200 59.800 ;
        RECT 78.000 57.000 78.800 59.800 ;
        RECT 79.600 57.000 80.400 59.800 ;
        RECT 81.200 57.000 82.000 59.800 ;
        RECT 84.400 57.000 85.200 59.800 ;
        RECT 87.600 57.000 88.400 59.800 ;
        RECT 89.200 57.000 90.000 59.800 ;
        RECT 90.800 57.000 91.600 59.800 ;
        RECT 73.200 55.800 75.600 56.600 ;
        RECT 92.400 56.600 93.200 59.800 ;
        RECT 73.200 55.200 74.000 55.800 ;
        RECT 68.000 54.000 69.200 54.600 ;
        RECT 72.200 54.600 74.000 55.200 ;
        RECT 78.000 55.600 79.000 56.400 ;
        RECT 82.000 55.600 83.600 56.400 ;
        RECT 84.400 55.800 89.000 56.400 ;
        RECT 92.400 55.800 95.000 56.600 ;
        RECT 84.400 55.600 85.200 55.800 ;
        RECT 68.000 52.000 68.600 54.000 ;
        RECT 72.200 53.400 73.000 54.600 ;
        RECT 69.200 52.600 73.000 53.400 ;
        RECT 78.000 52.800 78.800 55.600 ;
        RECT 84.400 54.800 85.200 55.000 ;
        RECT 80.800 54.200 85.200 54.800 ;
        RECT 80.800 54.000 81.600 54.200 ;
        RECT 86.000 53.600 86.800 55.200 ;
        RECT 88.200 53.400 89.000 55.800 ;
        RECT 94.200 55.200 95.000 55.800 ;
        RECT 94.200 54.400 97.200 55.200 ;
        RECT 98.800 53.800 99.600 59.800 ;
        RECT 102.000 55.600 102.800 57.200 ;
        RECT 81.200 52.600 84.400 53.400 ;
        RECT 88.200 52.600 90.200 53.400 ;
        RECT 90.800 53.000 99.600 53.800 ;
        RECT 74.800 52.000 75.600 52.600 ;
        RECT 92.400 52.000 93.200 52.400 ;
        RECT 94.000 52.000 94.800 52.400 ;
        RECT 97.400 52.000 98.200 52.200 ;
        RECT 68.000 51.400 68.800 52.000 ;
        RECT 74.800 51.400 98.200 52.000 ;
        RECT 66.600 50.000 67.600 50.800 ;
        RECT 66.800 42.200 67.600 50.000 ;
        RECT 68.200 49.600 68.800 51.400 ;
        RECT 68.200 49.000 77.200 49.600 ;
        RECT 68.200 47.400 68.800 49.000 ;
        RECT 76.400 48.800 77.200 49.000 ;
        RECT 79.600 49.000 88.200 49.600 ;
        RECT 79.600 48.800 80.400 49.000 ;
        RECT 71.400 47.600 74.000 48.400 ;
        RECT 68.200 46.800 70.800 47.400 ;
        RECT 70.000 42.200 70.800 46.800 ;
        RECT 73.200 42.200 74.000 47.600 ;
        RECT 74.600 46.800 78.800 47.600 ;
        RECT 76.400 42.200 77.200 45.000 ;
        RECT 78.000 42.200 78.800 45.000 ;
        RECT 79.600 42.200 80.400 45.000 ;
        RECT 81.200 42.200 82.000 48.400 ;
        RECT 84.400 47.600 87.000 48.400 ;
        RECT 87.600 48.200 88.200 49.000 ;
        RECT 89.200 49.400 90.000 49.600 ;
        RECT 89.200 49.000 94.600 49.400 ;
        RECT 89.200 48.800 95.400 49.000 ;
        RECT 94.000 48.200 95.400 48.800 ;
        RECT 87.600 47.600 93.400 48.200 ;
        RECT 96.400 48.000 98.000 48.800 ;
        RECT 96.400 47.600 97.000 48.000 ;
        RECT 84.400 42.200 85.200 47.000 ;
        RECT 87.600 42.200 88.400 47.000 ;
        RECT 92.800 46.800 97.000 47.600 ;
        RECT 98.800 47.400 99.600 53.000 ;
        RECT 97.600 46.800 99.600 47.400 ;
        RECT 89.200 42.200 90.000 45.000 ;
        RECT 90.800 42.200 91.600 45.000 ;
        RECT 94.000 42.200 94.800 46.800 ;
        RECT 97.600 46.200 98.200 46.800 ;
        RECT 97.200 45.600 98.200 46.200 ;
        RECT 97.200 42.200 98.000 45.600 ;
        RECT 103.600 42.200 104.400 59.800 ;
        RECT 106.800 55.200 107.600 59.800 ;
        RECT 110.000 55.200 110.800 59.800 ;
        RECT 113.200 55.200 114.000 59.800 ;
        RECT 116.400 55.200 117.200 59.800 ;
        RECT 120.800 58.400 121.600 59.800 ;
        RECT 120.800 57.600 122.000 58.400 ;
        RECT 106.800 54.400 108.600 55.200 ;
        RECT 110.000 54.400 112.200 55.200 ;
        RECT 113.200 54.400 115.400 55.200 ;
        RECT 116.400 54.400 118.800 55.200 ;
        RECT 107.800 53.800 108.600 54.400 ;
        RECT 111.400 53.800 112.200 54.400 ;
        RECT 114.600 53.800 115.400 54.400 ;
        RECT 107.800 53.000 110.400 53.800 ;
        RECT 111.400 53.000 113.800 53.800 ;
        RECT 114.600 53.000 117.200 53.800 ;
        RECT 107.800 51.600 108.600 53.000 ;
        RECT 111.400 51.600 112.200 53.000 ;
        RECT 114.600 51.600 115.400 53.000 ;
        RECT 118.000 51.600 118.800 54.400 ;
        RECT 120.800 54.200 121.600 57.600 ;
        RECT 129.200 56.000 130.000 59.800 ;
        RECT 106.800 50.800 108.600 51.600 ;
        RECT 110.000 50.800 112.200 51.600 ;
        RECT 113.200 50.800 115.400 51.600 ;
        RECT 116.400 50.800 118.800 51.600 ;
        RECT 119.800 53.800 121.600 54.200 ;
        RECT 129.000 55.200 130.000 56.000 ;
        RECT 119.800 53.600 121.400 53.800 ;
        RECT 106.800 42.200 107.600 50.800 ;
        RECT 110.000 42.200 110.800 50.800 ;
        RECT 113.200 42.200 114.000 50.800 ;
        RECT 116.400 42.200 117.200 50.800 ;
        RECT 119.800 50.400 120.400 53.600 ;
        RECT 122.000 51.600 123.600 52.400 ;
        RECT 119.600 49.600 120.400 50.400 ;
        RECT 122.800 50.300 123.600 50.400 ;
        RECT 124.400 50.300 125.200 51.200 ;
        RECT 129.000 50.800 129.800 55.200 ;
        RECT 130.800 54.600 131.600 59.800 ;
        RECT 137.200 56.600 138.000 59.800 ;
        RECT 138.800 57.000 139.600 59.800 ;
        RECT 140.400 57.000 141.200 59.800 ;
        RECT 142.000 57.000 142.800 59.800 ;
        RECT 143.600 57.000 144.400 59.800 ;
        RECT 146.800 57.000 147.600 59.800 ;
        RECT 150.000 57.000 150.800 59.800 ;
        RECT 151.600 57.000 152.400 59.800 ;
        RECT 153.200 57.000 154.000 59.800 ;
        RECT 135.600 55.800 138.000 56.600 ;
        RECT 154.800 56.600 155.600 59.800 ;
        RECT 135.600 55.200 136.400 55.800 ;
        RECT 130.400 54.000 131.600 54.600 ;
        RECT 134.600 54.600 136.400 55.200 ;
        RECT 140.400 55.600 141.400 56.400 ;
        RECT 144.400 55.600 146.000 56.400 ;
        RECT 146.800 55.800 151.400 56.400 ;
        RECT 154.800 55.800 157.400 56.600 ;
        RECT 146.800 55.600 147.600 55.800 ;
        RECT 130.400 52.000 131.000 54.000 ;
        RECT 134.600 53.400 135.400 54.600 ;
        RECT 131.600 52.600 135.400 53.400 ;
        RECT 140.400 52.800 141.200 55.600 ;
        RECT 146.800 54.800 147.600 55.000 ;
        RECT 143.200 54.200 147.600 54.800 ;
        RECT 143.200 54.000 144.000 54.200 ;
        RECT 148.400 53.600 149.200 55.200 ;
        RECT 150.600 53.400 151.400 55.800 ;
        RECT 156.600 55.200 157.400 55.800 ;
        RECT 156.600 54.400 159.600 55.200 ;
        RECT 161.200 53.800 162.000 59.800 ;
        RECT 162.800 55.600 163.600 57.200 ;
        RECT 143.600 52.600 146.800 53.400 ;
        RECT 150.600 52.600 152.600 53.400 ;
        RECT 153.200 53.000 162.000 53.800 ;
        RECT 137.200 52.000 138.000 52.600 ;
        RECT 154.800 52.000 155.600 52.400 ;
        RECT 159.600 52.200 160.400 52.400 ;
        RECT 159.600 52.000 160.600 52.200 ;
        RECT 130.400 51.400 131.200 52.000 ;
        RECT 137.200 51.400 160.600 52.000 ;
        RECT 129.000 50.300 130.000 50.800 ;
        RECT 122.800 49.700 130.000 50.300 ;
        RECT 122.800 49.600 123.600 49.700 ;
        RECT 124.400 49.600 125.200 49.700 ;
        RECT 119.800 47.000 120.400 49.600 ;
        RECT 121.200 48.300 122.000 49.200 ;
        RECT 124.400 48.300 125.200 48.400 ;
        RECT 121.200 47.700 125.200 48.300 ;
        RECT 121.200 47.600 122.000 47.700 ;
        RECT 124.400 47.600 125.200 47.700 ;
        RECT 119.800 46.400 123.400 47.000 ;
        RECT 119.800 46.200 120.400 46.400 ;
        RECT 119.600 42.200 120.400 46.200 ;
        RECT 122.800 46.200 123.400 46.400 ;
        RECT 122.800 42.200 123.600 46.200 ;
        RECT 129.200 42.200 130.000 49.700 ;
        RECT 130.600 49.600 131.200 51.400 ;
        RECT 130.600 49.000 139.600 49.600 ;
        RECT 130.600 47.400 131.200 49.000 ;
        RECT 138.800 48.800 139.600 49.000 ;
        RECT 142.000 49.000 150.600 49.600 ;
        RECT 142.000 48.800 142.800 49.000 ;
        RECT 133.800 47.600 136.400 48.400 ;
        RECT 130.600 46.800 133.200 47.400 ;
        RECT 132.400 42.200 133.200 46.800 ;
        RECT 135.600 42.200 136.400 47.600 ;
        RECT 137.000 46.800 141.200 47.600 ;
        RECT 138.800 42.200 139.600 45.000 ;
        RECT 140.400 42.200 141.200 45.000 ;
        RECT 142.000 42.200 142.800 45.000 ;
        RECT 143.600 42.200 144.400 48.400 ;
        RECT 146.800 47.600 149.400 48.400 ;
        RECT 150.000 48.200 150.600 49.000 ;
        RECT 151.600 49.400 152.400 49.600 ;
        RECT 151.600 49.000 157.000 49.400 ;
        RECT 151.600 48.800 157.800 49.000 ;
        RECT 156.400 48.200 157.800 48.800 ;
        RECT 150.000 47.600 155.800 48.200 ;
        RECT 158.800 48.000 160.400 48.800 ;
        RECT 158.800 47.600 159.400 48.000 ;
        RECT 146.800 42.200 147.600 47.000 ;
        RECT 150.000 42.200 150.800 47.000 ;
        RECT 155.200 46.800 159.400 47.600 ;
        RECT 161.200 47.400 162.000 53.000 ;
        RECT 160.000 46.800 162.000 47.400 ;
        RECT 164.400 54.300 165.200 59.800 ;
        RECT 169.200 55.800 170.000 59.800 ;
        RECT 170.600 56.400 171.400 57.200 ;
        RECT 170.800 56.300 171.600 56.400 ;
        RECT 172.400 56.300 173.200 59.800 ;
        RECT 167.600 54.300 168.400 54.400 ;
        RECT 164.400 53.700 168.400 54.300 ;
        RECT 151.600 42.200 152.400 45.000 ;
        RECT 153.200 42.200 154.000 45.000 ;
        RECT 156.400 42.200 157.200 46.800 ;
        RECT 160.000 46.200 160.600 46.800 ;
        RECT 159.600 45.600 160.600 46.200 ;
        RECT 159.600 42.200 160.400 45.600 ;
        RECT 164.400 42.200 165.200 53.700 ;
        RECT 167.600 52.800 168.400 53.700 ;
        RECT 166.000 52.200 166.800 52.400 ;
        RECT 169.200 52.200 169.800 55.800 ;
        RECT 170.800 55.700 173.200 56.300 ;
        RECT 174.000 56.000 174.800 59.800 ;
        RECT 177.200 56.000 178.000 59.800 ;
        RECT 174.000 55.800 178.000 56.000 ;
        RECT 178.800 56.000 179.600 59.800 ;
        RECT 182.000 56.000 182.800 59.800 ;
        RECT 178.800 55.800 182.800 56.000 ;
        RECT 183.600 55.800 184.400 59.800 ;
        RECT 170.800 55.600 171.600 55.700 ;
        RECT 172.600 54.400 173.200 55.700 ;
        RECT 174.200 55.400 177.800 55.800 ;
        RECT 179.000 55.400 182.600 55.800 ;
        RECT 176.400 54.400 177.200 54.800 ;
        RECT 179.600 54.400 180.400 54.800 ;
        RECT 183.600 54.400 184.200 55.800 ;
        RECT 172.400 53.600 175.000 54.400 ;
        RECT 176.400 53.800 178.000 54.400 ;
        RECT 177.200 53.600 178.000 53.800 ;
        RECT 178.800 53.800 180.400 54.400 ;
        RECT 178.800 53.600 179.600 53.800 ;
        RECT 181.800 53.600 184.400 54.400 ;
        RECT 186.800 53.800 187.600 59.800 ;
        RECT 193.200 56.600 194.000 59.800 ;
        RECT 194.800 57.000 195.600 59.800 ;
        RECT 196.400 57.000 197.200 59.800 ;
        RECT 198.000 57.000 198.800 59.800 ;
        RECT 201.200 57.000 202.000 59.800 ;
        RECT 204.400 57.000 205.200 59.800 ;
        RECT 206.000 57.000 206.800 59.800 ;
        RECT 207.600 57.000 208.400 59.800 ;
        RECT 209.200 57.000 210.000 59.800 ;
        RECT 191.400 55.800 194.000 56.600 ;
        RECT 210.800 56.600 211.600 59.800 ;
        RECT 197.400 55.800 202.000 56.400 ;
        RECT 191.400 55.200 192.200 55.800 ;
        RECT 189.200 54.400 192.200 55.200 ;
        RECT 170.800 52.200 171.600 52.400 ;
        RECT 166.000 51.600 167.600 52.200 ;
        RECT 169.200 51.600 171.600 52.200 ;
        RECT 166.800 51.200 167.600 51.600 ;
        RECT 170.800 50.200 171.400 51.600 ;
        RECT 172.400 50.200 173.200 50.400 ;
        RECT 174.400 50.200 175.000 53.600 ;
        RECT 175.600 52.300 176.400 53.200 ;
        RECT 180.400 52.300 181.200 53.200 ;
        RECT 175.600 51.700 181.200 52.300 ;
        RECT 175.600 51.600 176.400 51.700 ;
        RECT 180.400 51.600 181.200 51.700 ;
        RECT 181.800 50.200 182.400 53.600 ;
        RECT 186.800 53.000 195.600 53.800 ;
        RECT 197.400 53.400 198.200 55.800 ;
        RECT 201.200 55.600 202.000 55.800 ;
        RECT 202.800 55.600 204.400 56.400 ;
        RECT 207.400 55.600 208.400 56.400 ;
        RECT 210.800 55.800 213.200 56.600 ;
        RECT 199.600 53.600 200.400 55.200 ;
        RECT 201.200 54.800 202.000 55.000 ;
        RECT 201.200 54.200 205.600 54.800 ;
        RECT 204.800 54.000 205.600 54.200 ;
        RECT 183.600 50.200 184.400 50.400 ;
        RECT 166.000 49.600 170.000 50.200 ;
        RECT 166.000 42.200 166.800 49.600 ;
        RECT 169.200 42.200 170.000 49.600 ;
        RECT 170.800 42.200 171.600 50.200 ;
        RECT 172.400 49.600 173.800 50.200 ;
        RECT 174.400 49.600 175.400 50.200 ;
        RECT 173.200 48.400 173.800 49.600 ;
        RECT 173.200 47.600 174.000 48.400 ;
        RECT 174.600 42.200 175.400 49.600 ;
        RECT 181.400 49.600 182.400 50.200 ;
        RECT 183.000 49.600 184.400 50.200 ;
        RECT 181.400 44.400 182.200 49.600 ;
        RECT 183.000 48.400 183.600 49.600 ;
        RECT 182.800 47.600 183.600 48.400 ;
        RECT 186.800 47.400 187.600 53.000 ;
        RECT 196.200 52.600 198.200 53.400 ;
        RECT 202.000 52.600 205.200 53.400 ;
        RECT 207.600 52.800 208.400 55.600 ;
        RECT 212.400 55.200 213.200 55.800 ;
        RECT 212.400 54.600 214.200 55.200 ;
        RECT 213.400 53.400 214.200 54.600 ;
        RECT 217.200 54.600 218.000 59.800 ;
        RECT 218.800 56.000 219.600 59.800 ;
        RECT 220.400 56.300 221.200 56.400 ;
        RECT 222.000 56.300 222.800 57.200 ;
        RECT 218.800 55.200 219.800 56.000 ;
        RECT 220.400 55.700 222.800 56.300 ;
        RECT 220.400 55.600 221.200 55.700 ;
        RECT 222.000 55.600 222.800 55.700 ;
        RECT 217.200 54.000 218.400 54.600 ;
        RECT 213.400 52.600 217.200 53.400 ;
        RECT 188.200 52.000 189.000 52.200 ;
        RECT 193.200 52.000 194.000 52.400 ;
        RECT 210.800 52.000 211.600 52.600 ;
        RECT 217.800 52.000 218.400 54.000 ;
        RECT 188.200 51.400 211.600 52.000 ;
        RECT 217.600 51.400 218.400 52.000 ;
        RECT 217.600 49.600 218.200 51.400 ;
        RECT 219.000 50.800 219.800 55.200 ;
        RECT 196.400 49.400 197.200 49.600 ;
        RECT 191.800 49.000 197.200 49.400 ;
        RECT 191.000 48.800 197.200 49.000 ;
        RECT 198.200 49.000 206.800 49.600 ;
        RECT 188.400 48.000 190.000 48.800 ;
        RECT 191.000 48.200 192.400 48.800 ;
        RECT 198.200 48.200 198.800 49.000 ;
        RECT 206.000 48.800 206.800 49.000 ;
        RECT 209.200 49.000 218.200 49.600 ;
        RECT 209.200 48.800 210.000 49.000 ;
        RECT 189.400 47.600 190.000 48.000 ;
        RECT 193.000 47.600 198.800 48.200 ;
        RECT 199.400 47.600 202.000 48.400 ;
        RECT 186.800 46.800 188.800 47.400 ;
        RECT 189.400 46.800 193.600 47.600 ;
        RECT 188.200 46.200 188.800 46.800 ;
        RECT 188.200 45.600 189.200 46.200 ;
        RECT 180.400 43.600 182.200 44.400 ;
        RECT 181.400 42.200 182.200 43.600 ;
        RECT 188.400 42.200 189.200 45.600 ;
        RECT 191.600 42.200 192.400 46.800 ;
        RECT 194.800 42.200 195.600 45.000 ;
        RECT 196.400 42.200 197.200 45.000 ;
        RECT 198.000 42.200 198.800 47.000 ;
        RECT 201.200 42.200 202.000 47.000 ;
        RECT 204.400 42.200 205.200 48.400 ;
        RECT 212.400 47.600 215.000 48.400 ;
        RECT 207.600 46.800 211.800 47.600 ;
        RECT 206.000 42.200 206.800 45.000 ;
        RECT 207.600 42.200 208.400 45.000 ;
        RECT 209.200 42.200 210.000 45.000 ;
        RECT 212.400 42.200 213.200 47.600 ;
        RECT 217.600 47.400 218.200 49.000 ;
        RECT 215.600 46.800 218.200 47.400 ;
        RECT 218.800 50.000 219.800 50.800 ;
        RECT 215.600 42.200 216.400 46.800 ;
        RECT 218.800 42.200 219.600 50.000 ;
        RECT 223.600 42.200 224.400 59.800 ;
        RECT 2.800 32.000 3.600 39.800 ;
        RECT 6.000 35.200 6.800 39.800 ;
        RECT 2.600 31.200 3.600 32.000 ;
        RECT 4.200 34.600 6.800 35.200 ;
        RECT 4.200 33.000 4.800 34.600 ;
        RECT 9.200 34.400 10.000 39.800 ;
        RECT 12.400 37.000 13.200 39.800 ;
        RECT 14.000 37.000 14.800 39.800 ;
        RECT 15.600 37.000 16.400 39.800 ;
        RECT 10.600 34.400 14.800 35.200 ;
        RECT 7.400 33.600 10.000 34.400 ;
        RECT 17.200 33.600 18.000 39.800 ;
        RECT 20.400 35.000 21.200 39.800 ;
        RECT 23.600 35.000 24.400 39.800 ;
        RECT 25.200 37.000 26.000 39.800 ;
        RECT 26.800 37.000 27.600 39.800 ;
        RECT 30.000 35.200 30.800 39.800 ;
        RECT 33.200 36.400 34.000 39.800 ;
        RECT 33.200 35.800 34.200 36.400 ;
        RECT 33.600 35.200 34.200 35.800 ;
        RECT 28.800 34.400 33.000 35.200 ;
        RECT 33.600 34.600 35.600 35.200 ;
        RECT 20.400 33.600 23.000 34.400 ;
        RECT 23.600 33.800 29.400 34.400 ;
        RECT 32.400 34.000 33.000 34.400 ;
        RECT 12.400 33.000 13.200 33.200 ;
        RECT 4.200 32.400 13.200 33.000 ;
        RECT 15.600 33.000 16.400 33.200 ;
        RECT 23.600 33.000 24.200 33.800 ;
        RECT 30.000 33.200 31.400 33.800 ;
        RECT 32.400 33.200 34.000 34.000 ;
        RECT 15.600 32.400 24.200 33.000 ;
        RECT 25.200 33.000 31.400 33.200 ;
        RECT 25.200 32.600 30.600 33.000 ;
        RECT 25.200 32.400 26.000 32.600 ;
        RECT 2.600 26.800 3.400 31.200 ;
        RECT 4.200 30.600 4.800 32.400 ;
        RECT 28.200 31.800 29.000 32.000 ;
        RECT 31.600 31.800 32.400 32.400 ;
        RECT 5.400 31.200 32.400 31.800 ;
        RECT 5.400 31.000 6.200 31.200 ;
        RECT 4.000 30.000 4.800 30.600 ;
        RECT 4.000 28.000 4.600 30.000 ;
        RECT 5.200 28.600 9.000 29.400 ;
        RECT 4.000 27.400 5.200 28.000 ;
        RECT 2.600 26.000 3.600 26.800 ;
        RECT 2.800 22.200 3.600 26.000 ;
        RECT 4.400 22.200 5.200 27.400 ;
        RECT 8.200 27.400 9.000 28.600 ;
        RECT 8.200 26.800 10.000 27.400 ;
        RECT 9.200 26.200 10.000 26.800 ;
        RECT 14.000 26.400 14.800 29.200 ;
        RECT 17.200 28.600 20.400 29.400 ;
        RECT 24.200 28.600 26.200 29.400 ;
        RECT 34.800 29.000 35.600 34.600 ;
        RECT 38.000 31.800 38.800 39.800 ;
        RECT 41.200 35.800 42.000 39.800 ;
        RECT 38.000 30.400 38.600 31.800 ;
        RECT 41.200 31.600 41.800 35.800 ;
        RECT 39.400 31.000 41.800 31.600 ;
        RECT 36.400 30.300 37.200 30.400 ;
        RECT 38.000 30.300 38.800 30.400 ;
        RECT 36.400 29.700 38.800 30.300 ;
        RECT 36.400 29.600 37.200 29.700 ;
        RECT 38.000 29.600 38.800 29.700 ;
        RECT 16.800 27.800 17.600 28.000 ;
        RECT 16.800 27.200 21.200 27.800 ;
        RECT 20.400 27.000 21.200 27.200 ;
        RECT 22.000 26.800 22.800 28.400 ;
        RECT 9.200 25.400 11.600 26.200 ;
        RECT 14.000 25.600 15.000 26.400 ;
        RECT 18.000 25.600 19.600 26.400 ;
        RECT 20.400 26.200 21.200 26.400 ;
        RECT 24.200 26.200 25.000 28.600 ;
        RECT 26.800 28.200 35.600 29.000 ;
        RECT 30.200 26.800 33.200 27.600 ;
        RECT 30.200 26.200 31.000 26.800 ;
        RECT 20.400 25.600 25.000 26.200 ;
        RECT 10.800 22.200 11.600 25.400 ;
        RECT 28.400 25.400 31.000 26.200 ;
        RECT 12.400 22.200 13.200 25.000 ;
        RECT 14.000 22.200 14.800 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 17.200 22.200 18.000 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 26.800 22.200 27.600 25.000 ;
        RECT 28.400 22.200 29.200 25.400 ;
        RECT 34.800 22.200 35.600 28.200 ;
        RECT 38.000 26.200 38.600 29.600 ;
        RECT 39.400 27.600 40.000 31.000 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 41.200 28.800 41.800 29.600 ;
        RECT 40.800 28.200 41.800 28.800 ;
        RECT 40.800 28.000 41.600 28.200 ;
        RECT 42.800 27.600 43.600 29.200 ;
        RECT 46.000 28.300 46.800 39.800 ;
        RECT 50.200 32.400 51.000 39.800 ;
        RECT 51.600 33.600 52.400 34.400 ;
        RECT 51.800 32.400 52.400 33.600 ;
        RECT 50.200 31.800 51.200 32.400 ;
        RECT 51.800 31.800 53.200 32.400 ;
        RECT 55.600 32.000 56.400 39.800 ;
        RECT 58.800 35.200 59.600 39.800 ;
        RECT 49.200 28.800 50.000 30.400 ;
        RECT 50.600 28.400 51.200 31.800 ;
        RECT 52.400 31.600 53.200 31.800 ;
        RECT 55.400 31.200 56.400 32.000 ;
        RECT 57.000 34.600 59.600 35.200 ;
        RECT 57.000 33.000 57.600 34.600 ;
        RECT 62.000 34.400 62.800 39.800 ;
        RECT 65.200 37.000 66.000 39.800 ;
        RECT 66.800 37.000 67.600 39.800 ;
        RECT 68.400 37.000 69.200 39.800 ;
        RECT 63.400 34.400 67.600 35.200 ;
        RECT 60.200 33.600 62.800 34.400 ;
        RECT 70.000 33.600 70.800 39.800 ;
        RECT 73.200 35.000 74.000 39.800 ;
        RECT 76.400 35.000 77.200 39.800 ;
        RECT 78.000 37.000 78.800 39.800 ;
        RECT 79.600 37.000 80.400 39.800 ;
        RECT 82.800 35.200 83.600 39.800 ;
        RECT 86.000 36.400 86.800 39.800 ;
        RECT 86.000 35.800 87.000 36.400 ;
        RECT 86.400 35.200 87.000 35.800 ;
        RECT 81.600 34.400 85.800 35.200 ;
        RECT 86.400 34.600 88.400 35.200 ;
        RECT 73.200 33.600 75.800 34.400 ;
        RECT 76.400 33.800 82.200 34.400 ;
        RECT 85.200 34.000 85.800 34.400 ;
        RECT 65.200 33.000 66.000 33.200 ;
        RECT 57.000 32.400 66.000 33.000 ;
        RECT 68.400 33.000 69.200 33.200 ;
        RECT 76.400 33.000 77.000 33.800 ;
        RECT 82.800 33.200 84.200 33.800 ;
        RECT 85.200 33.200 86.800 34.000 ;
        RECT 68.400 32.400 77.000 33.000 ;
        RECT 78.000 33.000 84.200 33.200 ;
        RECT 78.000 32.600 83.400 33.000 ;
        RECT 78.000 32.400 78.800 32.600 ;
        RECT 47.600 28.300 48.400 28.400 ;
        RECT 46.000 28.200 48.400 28.300 ;
        RECT 46.000 27.700 49.200 28.200 ;
        RECT 39.200 27.400 40.000 27.600 ;
        RECT 39.200 27.000 42.200 27.400 ;
        RECT 39.200 26.800 43.400 27.000 ;
        RECT 41.600 26.400 43.400 26.800 ;
        RECT 42.800 26.200 43.400 26.400 ;
        RECT 38.000 25.200 39.400 26.200 ;
        RECT 38.600 22.200 39.400 25.200 ;
        RECT 42.800 22.200 43.600 26.200 ;
        RECT 44.400 24.800 45.200 26.400 ;
        RECT 46.000 22.200 46.800 27.700 ;
        RECT 47.600 27.600 49.200 27.700 ;
        RECT 50.600 27.600 53.200 28.400 ;
        RECT 48.400 27.200 49.200 27.600 ;
        RECT 47.800 26.200 51.400 26.600 ;
        RECT 52.400 26.200 53.000 27.600 ;
        RECT 55.400 26.800 56.200 31.200 ;
        RECT 57.000 30.600 57.600 32.400 ;
        RECT 56.800 30.000 57.600 30.600 ;
        RECT 63.600 30.000 87.000 30.600 ;
        RECT 56.800 28.000 57.400 30.000 ;
        RECT 63.600 29.400 64.400 30.000 ;
        RECT 81.200 29.600 82.000 30.000 ;
        RECT 84.400 29.600 85.200 30.000 ;
        RECT 86.200 29.800 87.000 30.000 ;
        RECT 58.000 28.600 61.800 29.400 ;
        RECT 56.800 27.400 58.000 28.000 ;
        RECT 47.600 26.000 51.600 26.200 ;
        RECT 47.600 22.200 48.400 26.000 ;
        RECT 50.800 22.200 51.600 26.000 ;
        RECT 52.400 22.200 53.200 26.200 ;
        RECT 55.400 26.000 56.400 26.800 ;
        RECT 55.600 22.200 56.400 26.000 ;
        RECT 57.200 22.200 58.000 27.400 ;
        RECT 61.000 27.400 61.800 28.600 ;
        RECT 61.000 26.800 62.800 27.400 ;
        RECT 62.000 26.200 62.800 26.800 ;
        RECT 66.800 26.400 67.600 29.200 ;
        RECT 70.000 28.600 73.200 29.400 ;
        RECT 77.000 28.600 79.000 29.400 ;
        RECT 87.600 29.000 88.400 34.600 ;
        RECT 92.400 32.800 93.200 39.800 ;
        RECT 69.600 27.800 70.400 28.000 ;
        RECT 69.600 27.200 74.000 27.800 ;
        RECT 73.200 27.000 74.000 27.200 ;
        RECT 74.800 26.800 75.600 28.400 ;
        RECT 62.000 25.400 64.400 26.200 ;
        RECT 66.800 25.600 67.800 26.400 ;
        RECT 70.800 25.600 72.400 26.400 ;
        RECT 73.200 26.200 74.000 26.400 ;
        RECT 77.000 26.200 77.800 28.600 ;
        RECT 79.600 28.200 88.400 29.000 ;
        RECT 92.200 31.800 93.200 32.800 ;
        RECT 95.600 32.400 96.400 39.800 ;
        RECT 93.800 31.800 96.400 32.400 ;
        RECT 97.200 32.400 98.000 39.800 ;
        RECT 100.400 32.800 101.200 39.800 ;
        RECT 97.200 31.800 99.800 32.400 ;
        RECT 100.400 31.800 101.400 32.800 ;
        RECT 92.200 28.400 92.800 31.800 ;
        RECT 93.800 29.800 94.400 31.800 ;
        RECT 93.400 29.000 94.400 29.800 ;
        RECT 83.000 26.800 86.000 27.600 ;
        RECT 83.000 26.200 83.800 26.800 ;
        RECT 73.200 25.600 77.800 26.200 ;
        RECT 63.600 22.200 64.400 25.400 ;
        RECT 81.200 25.400 83.800 26.200 ;
        RECT 65.200 22.200 66.000 25.000 ;
        RECT 66.800 22.200 67.600 25.000 ;
        RECT 68.400 22.200 69.200 25.000 ;
        RECT 70.000 22.200 70.800 25.000 ;
        RECT 73.200 22.200 74.000 25.000 ;
        RECT 76.400 22.200 77.200 25.000 ;
        RECT 78.000 22.200 78.800 25.000 ;
        RECT 79.600 22.200 80.400 25.000 ;
        RECT 81.200 22.200 82.000 25.400 ;
        RECT 87.600 22.200 88.400 28.200 ;
        RECT 89.200 28.300 90.000 28.400 ;
        RECT 92.200 28.300 93.200 28.400 ;
        RECT 89.200 27.700 93.200 28.300 ;
        RECT 89.200 27.600 90.000 27.700 ;
        RECT 92.200 27.600 93.200 27.700 ;
        RECT 92.200 26.200 92.800 27.600 ;
        RECT 93.800 27.400 94.400 29.000 ;
        RECT 95.400 30.300 96.400 30.400 ;
        RECT 97.200 30.300 98.200 30.400 ;
        RECT 95.400 29.700 98.200 30.300 ;
        RECT 95.400 29.600 96.400 29.700 ;
        RECT 97.200 29.600 98.200 29.700 ;
        RECT 95.400 28.800 96.200 29.600 ;
        RECT 97.400 28.800 98.200 29.600 ;
        RECT 99.200 29.800 99.800 31.800 ;
        RECT 99.200 29.000 100.200 29.800 ;
        RECT 99.200 27.400 99.800 29.000 ;
        RECT 100.800 28.400 101.400 31.800 ;
        RECT 105.200 31.200 106.000 39.800 ;
        RECT 108.400 31.200 109.200 39.800 ;
        RECT 113.200 36.400 114.000 39.800 ;
        RECT 113.000 35.800 114.000 36.400 ;
        RECT 113.000 35.200 113.600 35.800 ;
        RECT 116.400 35.200 117.200 39.800 ;
        RECT 119.600 37.000 120.400 39.800 ;
        RECT 121.200 37.000 122.000 39.800 ;
        RECT 105.200 30.400 109.200 31.200 ;
        RECT 100.400 27.600 101.400 28.400 ;
        RECT 108.400 27.600 109.200 30.400 ;
        RECT 93.800 26.800 96.400 27.400 ;
        RECT 92.200 25.600 93.200 26.200 ;
        RECT 92.400 22.200 93.200 25.600 ;
        RECT 95.600 22.200 96.400 26.800 ;
        RECT 97.200 26.800 99.800 27.400 ;
        RECT 97.200 22.200 98.000 26.800 ;
        RECT 100.800 26.200 101.400 27.600 ;
        RECT 100.400 25.600 101.400 26.200 ;
        RECT 105.200 26.800 109.200 27.600 ;
        RECT 100.400 22.200 101.200 25.600 ;
        RECT 105.200 22.200 106.000 26.800 ;
        RECT 108.400 22.200 109.200 26.800 ;
        RECT 111.600 34.600 113.600 35.200 ;
        RECT 111.600 29.000 112.400 34.600 ;
        RECT 114.200 34.400 118.400 35.200 ;
        RECT 122.800 35.000 123.600 39.800 ;
        RECT 126.000 35.000 126.800 39.800 ;
        RECT 114.200 34.000 114.800 34.400 ;
        RECT 113.200 33.200 114.800 34.000 ;
        RECT 117.800 33.800 123.600 34.400 ;
        RECT 115.800 33.200 117.200 33.800 ;
        RECT 115.800 33.000 122.000 33.200 ;
        RECT 116.600 32.600 122.000 33.000 ;
        RECT 121.200 32.400 122.000 32.600 ;
        RECT 123.000 33.000 123.600 33.800 ;
        RECT 124.200 33.600 126.800 34.400 ;
        RECT 129.200 33.600 130.000 39.800 ;
        RECT 130.800 37.000 131.600 39.800 ;
        RECT 132.400 37.000 133.200 39.800 ;
        RECT 134.000 37.000 134.800 39.800 ;
        RECT 132.400 34.400 136.600 35.200 ;
        RECT 137.200 34.400 138.000 39.800 ;
        RECT 140.400 35.200 141.200 39.800 ;
        RECT 140.400 34.600 143.000 35.200 ;
        RECT 137.200 33.600 139.800 34.400 ;
        RECT 130.800 33.000 131.600 33.200 ;
        RECT 123.000 32.400 131.600 33.000 ;
        RECT 134.000 33.000 134.800 33.200 ;
        RECT 142.400 33.000 143.000 34.600 ;
        RECT 134.000 32.400 143.000 33.000 ;
        RECT 142.400 30.600 143.000 32.400 ;
        RECT 143.600 32.000 144.400 39.800 ;
        RECT 143.600 31.200 144.600 32.000 ;
        RECT 113.000 30.000 136.400 30.600 ;
        RECT 142.400 30.000 143.200 30.600 ;
        RECT 113.000 29.800 113.800 30.000 ;
        RECT 114.800 29.600 115.600 30.000 ;
        RECT 118.000 29.600 118.800 30.000 ;
        RECT 135.600 29.400 136.400 30.000 ;
        RECT 111.600 28.200 120.400 29.000 ;
        RECT 121.000 28.600 123.000 29.400 ;
        RECT 126.800 28.600 130.000 29.400 ;
        RECT 111.600 22.200 112.400 28.200 ;
        RECT 114.000 26.800 117.000 27.600 ;
        RECT 116.200 26.200 117.000 26.800 ;
        RECT 122.200 26.200 123.000 28.600 ;
        RECT 124.400 26.800 125.200 28.400 ;
        RECT 129.600 27.800 130.400 28.000 ;
        RECT 126.000 27.200 130.400 27.800 ;
        RECT 126.000 27.000 126.800 27.200 ;
        RECT 132.400 26.400 133.200 29.200 ;
        RECT 138.200 28.600 142.000 29.400 ;
        RECT 138.200 27.400 139.000 28.600 ;
        RECT 142.600 28.000 143.200 30.000 ;
        RECT 126.000 26.200 126.800 26.400 ;
        RECT 116.200 25.400 118.800 26.200 ;
        RECT 122.200 25.600 126.800 26.200 ;
        RECT 127.600 25.600 129.200 26.400 ;
        RECT 132.200 25.600 133.200 26.400 ;
        RECT 137.200 26.800 139.000 27.400 ;
        RECT 142.000 27.400 143.200 28.000 ;
        RECT 137.200 26.200 138.000 26.800 ;
        RECT 118.000 22.200 118.800 25.400 ;
        RECT 135.600 25.400 138.000 26.200 ;
        RECT 119.600 22.200 120.400 25.000 ;
        RECT 121.200 22.200 122.000 25.000 ;
        RECT 122.800 22.200 123.600 25.000 ;
        RECT 126.000 22.200 126.800 25.000 ;
        RECT 129.200 22.200 130.000 25.000 ;
        RECT 130.800 22.200 131.600 25.000 ;
        RECT 132.400 22.200 133.200 25.000 ;
        RECT 134.000 22.200 134.800 25.000 ;
        RECT 135.600 22.200 136.400 25.400 ;
        RECT 142.000 22.200 142.800 27.400 ;
        RECT 143.800 26.800 144.600 31.200 ;
        RECT 143.600 26.300 144.600 26.800 ;
        RECT 150.000 30.300 150.800 39.800 ;
        RECT 155.400 32.800 156.200 39.800 ;
        RECT 159.600 35.000 160.400 39.000 ;
        RECT 154.600 32.200 156.200 32.800 ;
        RECT 153.200 30.300 154.000 31.200 ;
        RECT 150.000 29.700 154.000 30.300 ;
        RECT 148.400 26.300 149.200 26.400 ;
        RECT 143.600 25.700 149.200 26.300 ;
        RECT 143.600 22.200 144.400 25.700 ;
        RECT 148.400 24.800 149.200 25.700 ;
        RECT 150.000 22.200 150.800 29.700 ;
        RECT 153.200 29.600 154.000 29.700 ;
        RECT 154.600 28.400 155.200 32.200 ;
        RECT 159.800 31.600 160.400 35.000 ;
        RECT 161.200 34.300 162.000 34.400 ;
        RECT 162.800 34.300 163.600 39.800 ;
        RECT 166.000 35.200 166.800 39.800 ;
        RECT 161.200 33.700 163.600 34.300 ;
        RECT 161.200 33.600 162.000 33.700 ;
        RECT 162.800 32.000 163.600 33.700 ;
        RECT 156.600 31.000 160.400 31.600 ;
        RECT 162.600 31.200 163.600 32.000 ;
        RECT 164.200 34.600 166.800 35.200 ;
        RECT 164.200 33.000 164.800 34.600 ;
        RECT 169.200 34.400 170.000 39.800 ;
        RECT 172.400 37.000 173.200 39.800 ;
        RECT 174.000 37.000 174.800 39.800 ;
        RECT 175.600 37.000 176.400 39.800 ;
        RECT 170.600 34.400 174.800 35.200 ;
        RECT 167.400 33.600 170.000 34.400 ;
        RECT 177.200 33.600 178.000 39.800 ;
        RECT 180.400 35.000 181.200 39.800 ;
        RECT 183.600 35.000 184.400 39.800 ;
        RECT 185.200 37.000 186.000 39.800 ;
        RECT 186.800 37.000 187.600 39.800 ;
        RECT 190.000 35.200 190.800 39.800 ;
        RECT 193.200 36.400 194.000 39.800 ;
        RECT 193.200 35.800 194.200 36.400 ;
        RECT 193.600 35.200 194.200 35.800 ;
        RECT 188.800 34.400 193.000 35.200 ;
        RECT 193.600 34.600 195.600 35.200 ;
        RECT 180.400 33.600 183.000 34.400 ;
        RECT 183.600 33.800 189.400 34.400 ;
        RECT 192.400 34.000 193.000 34.400 ;
        RECT 172.400 33.000 173.200 33.200 ;
        RECT 164.200 32.400 173.200 33.000 ;
        RECT 175.600 33.000 176.400 33.200 ;
        RECT 183.600 33.000 184.200 33.800 ;
        RECT 190.000 33.200 191.400 33.800 ;
        RECT 192.400 33.200 194.000 34.000 ;
        RECT 175.600 32.400 184.200 33.000 ;
        RECT 185.200 33.000 191.400 33.200 ;
        RECT 185.200 32.600 190.600 33.000 ;
        RECT 185.200 32.400 186.000 32.600 ;
        RECT 156.600 29.000 157.200 31.000 ;
        RECT 151.600 28.300 152.400 28.400 ;
        RECT 153.200 28.300 155.200 28.400 ;
        RECT 151.600 27.700 155.200 28.300 ;
        RECT 155.800 28.200 157.200 29.000 ;
        RECT 158.000 28.800 158.800 30.400 ;
        RECT 159.600 28.800 160.400 30.400 ;
        RECT 151.600 27.600 152.400 27.700 ;
        RECT 153.200 27.600 155.200 27.700 ;
        RECT 154.600 27.000 155.200 27.600 ;
        RECT 156.200 27.800 157.200 28.200 ;
        RECT 156.200 27.200 160.400 27.800 ;
        RECT 154.600 26.600 155.400 27.000 ;
        RECT 154.600 26.000 156.200 26.600 ;
        RECT 155.400 23.000 156.200 26.000 ;
        RECT 159.800 25.000 160.400 27.200 ;
        RECT 162.600 26.800 163.400 31.200 ;
        RECT 164.200 30.600 164.800 32.400 ;
        RECT 164.000 30.000 164.800 30.600 ;
        RECT 170.800 30.000 194.200 30.600 ;
        RECT 164.000 28.000 164.600 30.000 ;
        RECT 170.800 29.400 171.600 30.000 ;
        RECT 188.400 29.600 189.200 30.000 ;
        RECT 190.000 29.600 190.800 30.000 ;
        RECT 193.200 29.800 194.200 30.000 ;
        RECT 193.200 29.600 194.000 29.800 ;
        RECT 165.200 28.600 169.000 29.400 ;
        RECT 164.000 27.400 165.200 28.000 ;
        RECT 162.600 26.000 163.600 26.800 ;
        RECT 159.600 23.000 160.400 25.000 ;
        RECT 162.800 22.200 163.600 26.000 ;
        RECT 164.400 22.200 165.200 27.400 ;
        RECT 168.200 27.400 169.000 28.600 ;
        RECT 168.200 26.800 170.000 27.400 ;
        RECT 169.200 26.200 170.000 26.800 ;
        RECT 174.000 26.400 174.800 29.200 ;
        RECT 177.200 28.600 180.400 29.400 ;
        RECT 184.200 28.600 186.200 29.400 ;
        RECT 194.800 29.000 195.600 34.600 ;
        RECT 198.000 31.800 198.800 39.800 ;
        RECT 199.600 32.400 200.400 39.800 ;
        RECT 202.800 32.400 203.600 39.800 ;
        RECT 199.600 31.800 203.600 32.400 ;
        RECT 198.200 30.400 198.800 31.800 ;
        RECT 202.000 30.400 202.800 30.800 ;
        RECT 198.000 29.800 200.400 30.400 ;
        RECT 202.000 29.800 203.600 30.400 ;
        RECT 198.000 29.600 198.800 29.800 ;
        RECT 176.800 27.800 177.600 28.000 ;
        RECT 176.800 27.200 181.200 27.800 ;
        RECT 180.400 27.000 181.200 27.200 ;
        RECT 182.000 26.800 182.800 28.400 ;
        RECT 169.200 25.400 171.600 26.200 ;
        RECT 174.000 25.600 175.000 26.400 ;
        RECT 178.000 25.600 179.600 26.400 ;
        RECT 180.400 26.200 181.200 26.400 ;
        RECT 184.200 26.200 185.000 28.600 ;
        RECT 186.800 28.200 195.600 29.000 ;
        RECT 190.200 26.800 193.200 27.600 ;
        RECT 190.200 26.200 191.000 26.800 ;
        RECT 180.400 25.600 185.000 26.200 ;
        RECT 170.800 22.200 171.600 25.400 ;
        RECT 188.400 25.400 191.000 26.200 ;
        RECT 172.400 22.200 173.200 25.000 ;
        RECT 174.000 22.200 174.800 25.000 ;
        RECT 175.600 22.200 176.400 25.000 ;
        RECT 177.200 22.200 178.000 25.000 ;
        RECT 180.400 22.200 181.200 25.000 ;
        RECT 183.600 22.200 184.400 25.000 ;
        RECT 185.200 22.200 186.000 25.000 ;
        RECT 186.800 22.200 187.600 25.000 ;
        RECT 188.400 22.200 189.200 25.400 ;
        RECT 194.800 22.200 195.600 28.200 ;
        RECT 196.400 28.300 197.200 28.400 ;
        RECT 199.800 28.300 200.400 29.800 ;
        RECT 202.800 29.600 203.600 29.800 ;
        RECT 196.400 27.700 200.400 28.300 ;
        RECT 196.400 27.600 197.200 27.700 ;
        RECT 198.000 25.600 198.800 26.400 ;
        RECT 199.800 26.200 200.400 27.700 ;
        RECT 201.200 28.300 202.000 29.200 ;
        RECT 204.400 28.300 205.200 39.800 ;
        RECT 207.600 35.000 208.400 39.000 ;
        RECT 211.800 38.400 212.600 39.800 ;
        RECT 211.800 37.600 213.200 38.400 ;
        RECT 207.600 31.600 208.200 35.000 ;
        RECT 211.800 32.800 212.600 37.600 ;
        RECT 211.800 32.200 213.400 32.800 ;
        RECT 207.600 31.000 211.400 31.600 ;
        RECT 207.600 28.800 208.400 30.400 ;
        RECT 209.200 28.800 210.000 30.400 ;
        RECT 210.800 29.000 211.400 31.000 ;
        RECT 206.000 28.300 206.800 28.400 ;
        RECT 201.200 27.700 206.800 28.300 ;
        RECT 210.800 28.200 212.200 29.000 ;
        RECT 212.800 28.400 213.400 32.200 ;
        RECT 214.000 30.300 214.800 31.200 ;
        RECT 217.200 30.300 218.000 39.800 ;
        RECT 220.400 32.400 221.200 39.800 ;
        RECT 220.400 31.800 222.600 32.400 ;
        RECT 222.000 31.200 222.600 31.800 ;
        RECT 222.000 30.400 223.200 31.200 ;
        RECT 214.000 29.700 218.000 30.300 ;
        RECT 214.000 29.600 214.800 29.700 ;
        RECT 210.800 27.800 211.800 28.200 ;
        RECT 201.200 27.600 202.000 27.700 ;
        RECT 198.200 24.800 199.000 25.600 ;
        RECT 199.600 22.200 200.400 26.200 ;
        RECT 204.400 22.200 205.200 27.700 ;
        RECT 206.000 27.600 206.800 27.700 ;
        RECT 207.600 27.200 211.800 27.800 ;
        RECT 212.800 27.600 214.800 28.400 ;
        RECT 206.000 24.800 206.800 26.400 ;
        RECT 207.600 25.000 208.200 27.200 ;
        RECT 212.800 27.000 213.400 27.600 ;
        RECT 212.600 26.600 213.400 27.000 ;
        RECT 211.800 26.000 213.400 26.600 ;
        RECT 207.600 23.000 208.400 25.000 ;
        RECT 211.800 23.000 212.600 26.000 ;
        RECT 217.200 22.200 218.000 29.700 ;
        RECT 218.800 30.300 219.600 30.400 ;
        RECT 220.400 30.300 221.200 30.400 ;
        RECT 218.800 29.700 221.200 30.300 ;
        RECT 218.800 29.600 219.600 29.700 ;
        RECT 220.400 28.800 221.200 29.700 ;
        RECT 222.000 27.400 222.600 30.400 ;
        RECT 220.400 26.800 222.600 27.400 ;
        RECT 218.800 24.800 219.600 26.400 ;
        RECT 220.400 22.200 221.200 26.800 ;
        RECT 2.800 16.000 3.600 19.800 ;
        RECT 2.600 15.200 3.600 16.000 ;
        RECT 2.600 10.800 3.400 15.200 ;
        RECT 4.400 14.600 5.200 19.800 ;
        RECT 10.800 16.600 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 14.000 17.000 14.800 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 17.200 17.000 18.000 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 26.800 17.000 27.600 19.800 ;
        RECT 9.200 15.800 11.600 16.600 ;
        RECT 28.400 16.600 29.200 19.800 ;
        RECT 9.200 15.200 10.000 15.800 ;
        RECT 4.000 14.000 5.200 14.600 ;
        RECT 8.200 14.600 10.000 15.200 ;
        RECT 14.000 15.600 15.000 16.400 ;
        RECT 18.000 15.600 19.600 16.400 ;
        RECT 20.400 15.800 25.000 16.400 ;
        RECT 28.400 15.800 31.000 16.600 ;
        RECT 20.400 15.600 21.200 15.800 ;
        RECT 4.000 12.000 4.600 14.000 ;
        RECT 8.200 13.400 9.000 14.600 ;
        RECT 5.200 12.600 9.000 13.400 ;
        RECT 14.000 12.800 14.800 15.600 ;
        RECT 20.400 14.800 21.200 15.000 ;
        RECT 16.800 14.200 21.200 14.800 ;
        RECT 16.800 14.000 17.600 14.200 ;
        RECT 22.000 13.600 22.800 15.200 ;
        RECT 24.200 13.400 25.000 15.800 ;
        RECT 30.200 15.200 31.000 15.800 ;
        RECT 30.200 14.400 33.200 15.200 ;
        RECT 34.800 13.800 35.600 19.800 ;
        RECT 39.600 17.800 40.400 19.800 ;
        RECT 36.400 16.300 37.200 16.400 ;
        RECT 38.000 16.300 38.800 17.200 ;
        RECT 39.800 16.300 40.400 17.800 ;
        RECT 41.200 16.300 42.000 16.400 ;
        RECT 36.400 15.700 38.800 16.300 ;
        RECT 39.700 15.700 42.000 16.300 ;
        RECT 36.400 15.600 37.200 15.700 ;
        RECT 38.000 15.600 38.800 15.700 ;
        RECT 39.800 14.400 40.400 15.700 ;
        RECT 41.200 15.600 42.000 15.700 ;
        RECT 17.200 12.600 20.400 13.400 ;
        RECT 24.200 12.600 26.200 13.400 ;
        RECT 26.800 13.000 35.600 13.800 ;
        RECT 39.600 13.600 40.400 14.400 ;
        RECT 10.800 12.000 11.600 12.600 ;
        RECT 28.400 12.000 29.200 12.400 ;
        RECT 31.600 12.000 32.400 12.400 ;
        RECT 33.400 12.000 34.200 12.200 ;
        RECT 4.000 11.400 4.800 12.000 ;
        RECT 10.800 11.400 34.200 12.000 ;
        RECT 2.600 10.000 3.600 10.800 ;
        RECT 2.800 2.200 3.600 10.000 ;
        RECT 4.200 9.600 4.800 11.400 ;
        RECT 4.200 9.000 13.200 9.600 ;
        RECT 4.200 7.400 4.800 9.000 ;
        RECT 12.400 8.800 13.200 9.000 ;
        RECT 15.600 9.000 24.200 9.600 ;
        RECT 15.600 8.800 16.400 9.000 ;
        RECT 7.400 7.600 10.000 8.400 ;
        RECT 4.200 6.800 6.800 7.400 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 7.600 ;
        RECT 10.600 6.800 14.800 7.600 ;
        RECT 12.400 2.200 13.200 5.000 ;
        RECT 14.000 2.200 14.800 5.000 ;
        RECT 15.600 2.200 16.400 5.000 ;
        RECT 17.200 2.200 18.000 8.400 ;
        RECT 20.400 7.600 23.000 8.400 ;
        RECT 23.600 8.200 24.200 9.000 ;
        RECT 25.200 9.400 26.000 9.600 ;
        RECT 25.200 9.000 30.600 9.400 ;
        RECT 25.200 8.800 31.400 9.000 ;
        RECT 30.000 8.200 31.400 8.800 ;
        RECT 23.600 7.600 29.400 8.200 ;
        RECT 32.400 8.000 34.000 8.800 ;
        RECT 32.400 7.600 33.000 8.000 ;
        RECT 20.400 2.200 21.200 7.000 ;
        RECT 23.600 2.200 24.400 7.000 ;
        RECT 28.800 6.800 33.000 7.600 ;
        RECT 34.800 7.400 35.600 13.000 ;
        RECT 39.800 10.200 40.400 13.600 ;
        RECT 41.200 12.300 42.000 12.400 ;
        RECT 42.800 12.300 43.600 19.800 ;
        RECT 44.400 16.300 45.200 17.200 ;
        RECT 47.600 16.300 48.400 19.800 ;
        RECT 44.400 15.700 48.400 16.300 ;
        RECT 44.400 15.600 45.200 15.700 ;
        RECT 41.200 11.700 43.600 12.300 ;
        RECT 41.200 10.800 42.000 11.700 ;
        RECT 39.600 9.400 41.400 10.200 ;
        RECT 33.600 6.800 35.600 7.400 ;
        RECT 25.200 2.200 26.000 5.000 ;
        RECT 26.800 2.200 27.600 5.000 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.600 6.200 34.200 6.800 ;
        RECT 33.200 5.600 34.200 6.200 ;
        RECT 33.200 2.200 34.000 5.600 ;
        RECT 40.600 2.200 41.400 9.400 ;
        RECT 42.800 2.200 43.600 11.700 ;
        RECT 47.400 15.200 48.400 15.700 ;
        RECT 47.400 10.800 48.200 15.200 ;
        RECT 49.200 14.600 50.000 19.800 ;
        RECT 55.600 16.600 56.400 19.800 ;
        RECT 57.200 17.000 58.000 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 60.400 17.000 61.200 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 65.200 17.000 66.000 19.800 ;
        RECT 68.400 17.000 69.200 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 71.600 17.000 72.400 19.800 ;
        RECT 54.000 15.800 56.400 16.600 ;
        RECT 73.200 16.600 74.000 19.800 ;
        RECT 54.000 15.200 54.800 15.800 ;
        RECT 48.800 14.000 50.000 14.600 ;
        RECT 53.000 14.600 54.800 15.200 ;
        RECT 58.800 15.600 59.800 16.400 ;
        RECT 62.800 15.600 64.400 16.400 ;
        RECT 65.200 15.800 69.800 16.400 ;
        RECT 73.200 15.800 75.800 16.600 ;
        RECT 65.200 15.600 66.000 15.800 ;
        RECT 48.800 12.000 49.400 14.000 ;
        RECT 53.000 13.400 53.800 14.600 ;
        RECT 50.000 12.600 53.800 13.400 ;
        RECT 58.800 12.800 59.600 15.600 ;
        RECT 65.200 14.800 66.000 15.000 ;
        RECT 61.600 14.200 66.000 14.800 ;
        RECT 61.600 14.000 62.400 14.200 ;
        RECT 69.000 13.400 69.800 15.800 ;
        RECT 75.000 15.200 75.800 15.800 ;
        RECT 75.000 14.400 78.000 15.200 ;
        RECT 79.600 13.800 80.400 19.800 ;
        RECT 84.400 15.200 85.200 19.800 ;
        RECT 87.600 15.200 88.400 19.800 ;
        RECT 90.800 15.200 91.600 19.800 ;
        RECT 94.000 15.200 94.800 19.800 ;
        RECT 62.000 12.600 65.200 13.400 ;
        RECT 69.000 12.600 71.000 13.400 ;
        RECT 71.600 13.000 80.400 13.800 ;
        RECT 55.600 12.000 56.400 12.600 ;
        RECT 73.200 12.000 74.000 12.400 ;
        RECT 76.400 12.000 77.200 12.400 ;
        RECT 78.200 12.000 79.000 12.200 ;
        RECT 48.800 11.400 49.600 12.000 ;
        RECT 55.600 11.400 79.000 12.000 ;
        RECT 47.400 10.000 48.400 10.800 ;
        RECT 47.600 2.200 48.400 10.000 ;
        RECT 49.000 9.600 49.600 11.400 ;
        RECT 49.000 9.000 58.000 9.600 ;
        RECT 49.000 7.400 49.600 9.000 ;
        RECT 57.200 8.800 58.000 9.000 ;
        RECT 60.400 9.000 69.000 9.600 ;
        RECT 60.400 8.800 61.200 9.000 ;
        RECT 52.200 7.600 54.800 8.400 ;
        RECT 49.000 6.800 51.600 7.400 ;
        RECT 50.800 2.200 51.600 6.800 ;
        RECT 54.000 2.200 54.800 7.600 ;
        RECT 55.400 6.800 59.600 7.600 ;
        RECT 57.200 2.200 58.000 5.000 ;
        RECT 58.800 2.200 59.600 5.000 ;
        RECT 60.400 2.200 61.200 5.000 ;
        RECT 62.000 2.200 62.800 8.400 ;
        RECT 65.200 7.600 67.800 8.400 ;
        RECT 68.400 8.200 69.000 9.000 ;
        RECT 70.000 9.400 70.800 9.600 ;
        RECT 70.000 9.000 75.400 9.400 ;
        RECT 70.000 8.800 76.200 9.000 ;
        RECT 74.800 8.200 76.200 8.800 ;
        RECT 68.400 7.600 74.200 8.200 ;
        RECT 77.200 8.000 78.800 8.800 ;
        RECT 77.200 7.600 77.800 8.000 ;
        RECT 65.200 2.200 66.000 7.000 ;
        RECT 68.400 2.200 69.200 7.000 ;
        RECT 73.600 6.800 77.800 7.600 ;
        RECT 79.600 7.400 80.400 13.000 ;
        RECT 82.800 14.400 85.200 15.200 ;
        RECT 86.200 14.400 88.400 15.200 ;
        RECT 89.400 14.400 91.600 15.200 ;
        RECT 93.000 14.400 94.800 15.200 ;
        RECT 82.800 11.600 83.600 14.400 ;
        RECT 86.200 13.800 87.000 14.400 ;
        RECT 89.400 13.800 90.200 14.400 ;
        RECT 93.000 13.800 93.800 14.400 ;
        RECT 84.400 13.000 87.000 13.800 ;
        RECT 87.800 13.000 90.200 13.800 ;
        RECT 91.200 13.000 93.800 13.800 ;
        RECT 86.200 11.600 87.000 13.000 ;
        RECT 89.400 11.600 90.200 13.000 ;
        RECT 93.000 11.600 93.800 13.000 ;
        RECT 97.200 13.800 98.000 19.800 ;
        RECT 103.600 16.600 104.400 19.800 ;
        RECT 105.200 17.000 106.000 19.800 ;
        RECT 106.800 17.000 107.600 19.800 ;
        RECT 108.400 17.000 109.200 19.800 ;
        RECT 111.600 17.000 112.400 19.800 ;
        RECT 114.800 17.000 115.600 19.800 ;
        RECT 116.400 17.000 117.200 19.800 ;
        RECT 118.000 17.000 118.800 19.800 ;
        RECT 119.600 17.000 120.400 19.800 ;
        RECT 101.800 15.800 104.400 16.600 ;
        RECT 121.200 16.600 122.000 19.800 ;
        RECT 107.800 15.800 112.400 16.400 ;
        RECT 101.800 15.200 102.600 15.800 ;
        RECT 99.600 14.400 102.600 15.200 ;
        RECT 97.200 13.000 106.000 13.800 ;
        RECT 107.800 13.400 108.600 15.800 ;
        RECT 111.600 15.600 112.400 15.800 ;
        RECT 113.200 15.600 114.800 16.400 ;
        RECT 117.800 15.600 118.800 16.400 ;
        RECT 121.200 15.800 123.600 16.600 ;
        RECT 110.000 13.600 110.800 15.200 ;
        RECT 111.600 14.800 112.400 15.000 ;
        RECT 111.600 14.200 116.000 14.800 ;
        RECT 115.200 14.000 116.000 14.200 ;
        RECT 82.800 10.800 85.200 11.600 ;
        RECT 86.200 10.800 88.400 11.600 ;
        RECT 89.400 10.800 91.600 11.600 ;
        RECT 93.000 10.800 94.800 11.600 ;
        RECT 78.400 6.800 80.400 7.400 ;
        RECT 70.000 2.200 70.800 5.000 ;
        RECT 71.600 2.200 72.400 5.000 ;
        RECT 74.800 2.200 75.600 6.800 ;
        RECT 78.400 6.200 79.000 6.800 ;
        RECT 78.000 5.600 79.000 6.200 ;
        RECT 78.000 2.200 78.800 5.600 ;
        RECT 84.400 2.200 85.200 10.800 ;
        RECT 87.600 2.200 88.400 10.800 ;
        RECT 90.800 2.200 91.600 10.800 ;
        RECT 94.000 2.200 94.800 10.800 ;
        RECT 97.200 7.400 98.000 13.000 ;
        RECT 106.600 12.600 108.600 13.400 ;
        RECT 112.400 12.600 115.600 13.400 ;
        RECT 118.000 12.800 118.800 15.600 ;
        RECT 122.800 15.200 123.600 15.800 ;
        RECT 122.800 14.600 124.600 15.200 ;
        RECT 123.800 13.400 124.600 14.600 ;
        RECT 127.600 14.600 128.400 19.800 ;
        RECT 129.200 16.000 130.000 19.800 ;
        RECT 129.200 15.200 130.200 16.000 ;
        RECT 127.600 14.000 128.800 14.600 ;
        RECT 123.800 12.600 127.600 13.400 ;
        RECT 98.600 12.000 99.400 12.200 ;
        RECT 100.400 12.000 101.200 12.400 ;
        RECT 103.600 12.000 104.400 12.400 ;
        RECT 121.200 12.000 122.000 12.600 ;
        RECT 128.200 12.000 128.800 14.000 ;
        RECT 98.600 11.400 122.000 12.000 ;
        RECT 128.000 11.400 128.800 12.000 ;
        RECT 129.400 12.300 130.200 15.200 ;
        RECT 132.400 15.200 133.200 19.800 ;
        RECT 138.800 15.600 139.600 17.200 ;
        RECT 132.400 14.600 134.600 15.200 ;
        RECT 132.400 12.300 133.200 13.200 ;
        RECT 129.400 11.700 133.200 12.300 ;
        RECT 128.000 9.600 128.600 11.400 ;
        RECT 129.400 10.800 130.200 11.700 ;
        RECT 132.400 11.600 133.200 11.700 ;
        RECT 134.000 11.600 134.600 14.600 ;
        RECT 140.400 12.300 141.200 19.800 ;
        RECT 145.800 16.000 146.600 19.000 ;
        RECT 150.000 17.000 150.800 19.000 ;
        RECT 145.000 15.400 146.600 16.000 ;
        RECT 145.000 15.000 145.800 15.400 ;
        RECT 145.000 14.400 145.600 15.000 ;
        RECT 150.200 14.800 150.800 17.000 ;
        RECT 142.000 14.300 142.800 14.400 ;
        RECT 143.600 14.300 145.600 14.400 ;
        RECT 142.000 13.700 145.600 14.300 ;
        RECT 146.600 14.200 150.800 14.800 ;
        RECT 151.600 15.200 152.400 19.800 ;
        RECT 151.600 14.600 153.800 15.200 ;
        RECT 146.600 13.800 147.600 14.200 ;
        RECT 142.000 13.600 142.800 13.700 ;
        RECT 143.600 13.600 145.600 13.700 ;
        RECT 143.600 12.300 144.400 12.400 ;
        RECT 140.400 11.700 144.400 12.300 ;
        RECT 106.800 9.400 107.600 9.600 ;
        RECT 102.200 9.000 107.600 9.400 ;
        RECT 101.400 8.800 107.600 9.000 ;
        RECT 108.600 9.000 117.200 9.600 ;
        RECT 98.800 8.000 100.400 8.800 ;
        RECT 101.400 8.200 102.800 8.800 ;
        RECT 108.600 8.200 109.200 9.000 ;
        RECT 116.400 8.800 117.200 9.000 ;
        RECT 119.600 9.000 128.600 9.600 ;
        RECT 119.600 8.800 120.400 9.000 ;
        RECT 99.800 7.600 100.400 8.000 ;
        RECT 103.400 7.600 109.200 8.200 ;
        RECT 109.800 7.600 112.400 8.400 ;
        RECT 97.200 6.800 99.200 7.400 ;
        RECT 99.800 6.800 104.000 7.600 ;
        RECT 98.600 6.200 99.200 6.800 ;
        RECT 98.600 5.600 99.600 6.200 ;
        RECT 98.800 2.200 99.600 5.600 ;
        RECT 102.000 2.200 102.800 6.800 ;
        RECT 105.200 2.200 106.000 5.000 ;
        RECT 106.800 2.200 107.600 5.000 ;
        RECT 108.400 2.200 109.200 7.000 ;
        RECT 111.600 2.200 112.400 7.000 ;
        RECT 114.800 2.200 115.600 8.400 ;
        RECT 122.800 7.600 125.400 8.400 ;
        RECT 118.000 6.800 122.200 7.600 ;
        RECT 116.400 2.200 117.200 5.000 ;
        RECT 118.000 2.200 118.800 5.000 ;
        RECT 119.600 2.200 120.400 5.000 ;
        RECT 122.800 2.200 123.600 7.600 ;
        RECT 128.000 7.400 128.600 9.000 ;
        RECT 126.000 6.800 128.600 7.400 ;
        RECT 129.200 10.000 130.200 10.800 ;
        RECT 134.000 10.800 135.200 11.600 ;
        RECT 134.000 10.200 134.600 10.800 ;
        RECT 126.000 2.200 126.800 6.800 ;
        RECT 129.200 2.200 130.000 10.000 ;
        RECT 132.400 9.600 134.600 10.200 ;
        RECT 132.400 2.200 133.200 9.600 ;
        RECT 140.400 2.200 141.200 11.700 ;
        RECT 143.600 10.800 144.400 11.700 ;
        RECT 145.000 9.800 145.600 13.600 ;
        RECT 146.200 13.000 147.600 13.800 ;
        RECT 147.000 11.000 147.600 13.000 ;
        RECT 148.400 11.600 149.200 13.200 ;
        RECT 150.000 11.600 150.800 13.200 ;
        RECT 151.600 11.600 152.400 13.200 ;
        RECT 153.200 11.600 153.800 14.600 ;
        RECT 147.000 10.400 150.800 11.000 ;
        RECT 145.000 9.200 146.600 9.800 ;
        RECT 145.800 2.200 146.600 9.200 ;
        RECT 150.200 7.000 150.800 10.400 ;
        RECT 153.200 10.800 154.400 11.600 ;
        RECT 153.200 10.200 153.800 10.800 ;
        RECT 150.000 3.000 150.800 7.000 ;
        RECT 151.600 9.600 153.800 10.200 ;
        RECT 151.600 2.200 152.400 9.600 ;
        RECT 156.400 2.200 157.200 19.800 ;
        RECT 158.000 15.600 158.800 17.200 ;
        RECT 159.600 15.200 160.400 19.800 ;
        RECT 167.600 15.800 168.400 19.800 ;
        RECT 169.000 16.400 169.800 17.200 ;
        RECT 159.600 14.600 161.800 15.200 ;
        RECT 158.000 12.300 158.800 12.400 ;
        RECT 159.600 12.300 160.400 13.200 ;
        RECT 158.000 11.700 160.400 12.300 ;
        RECT 158.000 11.600 158.800 11.700 ;
        RECT 159.600 11.600 160.400 11.700 ;
        RECT 161.200 11.600 161.800 14.600 ;
        RECT 166.000 12.800 166.800 14.400 ;
        RECT 164.400 12.200 165.200 12.400 ;
        RECT 167.600 12.200 168.200 15.800 ;
        RECT 169.200 15.600 170.000 16.400 ;
        RECT 170.800 15.200 171.600 19.800 ;
        RECT 175.600 15.600 176.400 19.800 ;
        RECT 177.200 16.000 178.000 19.800 ;
        RECT 180.400 16.000 181.200 19.800 ;
        RECT 177.200 15.800 181.200 16.000 ;
        RECT 170.800 14.600 173.000 15.200 ;
        RECT 169.200 12.200 170.000 12.400 ;
        RECT 164.400 11.600 166.000 12.200 ;
        RECT 167.600 11.600 170.000 12.200 ;
        RECT 170.800 11.600 171.600 13.200 ;
        RECT 172.400 11.600 173.000 14.600 ;
        RECT 175.800 14.400 176.400 15.600 ;
        RECT 177.400 15.400 181.000 15.800 ;
        RECT 179.600 14.400 180.400 14.800 ;
        RECT 175.600 13.600 178.200 14.400 ;
        RECT 179.600 13.800 181.200 14.400 ;
        RECT 180.400 13.600 181.200 13.800 ;
        RECT 183.600 13.800 184.400 19.800 ;
        RECT 190.000 16.600 190.800 19.800 ;
        RECT 191.600 17.000 192.400 19.800 ;
        RECT 193.200 17.000 194.000 19.800 ;
        RECT 194.800 17.000 195.600 19.800 ;
        RECT 198.000 17.000 198.800 19.800 ;
        RECT 201.200 17.000 202.000 19.800 ;
        RECT 202.800 17.000 203.600 19.800 ;
        RECT 204.400 17.000 205.200 19.800 ;
        RECT 206.000 17.000 206.800 19.800 ;
        RECT 188.200 15.800 190.800 16.600 ;
        RECT 207.600 16.600 208.400 19.800 ;
        RECT 194.200 15.800 198.800 16.400 ;
        RECT 188.200 15.200 189.000 15.800 ;
        RECT 186.000 14.400 189.000 15.200 ;
        RECT 161.200 10.800 162.400 11.600 ;
        RECT 165.200 11.200 166.000 11.600 ;
        RECT 161.200 10.200 161.800 10.800 ;
        RECT 169.200 10.200 169.800 11.600 ;
        RECT 172.400 10.800 173.600 11.600 ;
        RECT 172.400 10.200 173.000 10.800 ;
        RECT 159.600 9.600 161.800 10.200 ;
        RECT 164.400 9.600 168.400 10.200 ;
        RECT 159.600 2.200 160.400 9.600 ;
        RECT 164.400 2.200 165.200 9.600 ;
        RECT 167.600 2.200 168.400 9.600 ;
        RECT 169.200 2.200 170.000 10.200 ;
        RECT 170.800 9.600 173.000 10.200 ;
        RECT 175.600 10.200 176.400 10.400 ;
        RECT 177.600 10.200 178.200 13.600 ;
        RECT 178.800 11.600 179.600 13.200 ;
        RECT 183.600 13.000 192.400 13.800 ;
        RECT 194.200 13.400 195.000 15.800 ;
        RECT 198.000 15.600 198.800 15.800 ;
        RECT 199.600 15.600 201.200 16.400 ;
        RECT 204.200 15.600 205.200 16.400 ;
        RECT 207.600 15.800 210.000 16.600 ;
        RECT 196.400 13.600 197.200 15.200 ;
        RECT 198.000 14.800 198.800 15.000 ;
        RECT 198.000 14.200 202.400 14.800 ;
        RECT 201.600 14.000 202.400 14.200 ;
        RECT 175.600 9.600 177.000 10.200 ;
        RECT 177.600 9.600 178.600 10.200 ;
        RECT 170.800 2.200 171.600 9.600 ;
        RECT 176.400 8.400 177.000 9.600 ;
        RECT 176.400 7.600 177.200 8.400 ;
        RECT 177.800 2.200 178.600 9.600 ;
        RECT 183.600 7.400 184.400 13.000 ;
        RECT 193.000 12.600 195.000 13.400 ;
        RECT 198.800 12.600 202.000 13.400 ;
        RECT 204.400 12.800 205.200 15.600 ;
        RECT 209.200 15.200 210.000 15.800 ;
        RECT 209.200 14.600 211.000 15.200 ;
        RECT 210.200 13.400 211.000 14.600 ;
        RECT 214.000 14.600 214.800 19.800 ;
        RECT 215.600 16.000 216.400 19.800 ;
        RECT 215.600 15.200 216.600 16.000 ;
        RECT 214.000 14.000 215.200 14.600 ;
        RECT 210.200 12.600 214.000 13.400 ;
        RECT 185.000 12.000 185.800 12.200 ;
        RECT 190.000 12.000 190.800 12.400 ;
        RECT 207.600 12.000 208.400 12.600 ;
        RECT 214.600 12.000 215.200 14.000 ;
        RECT 185.000 11.400 208.400 12.000 ;
        RECT 214.400 11.400 215.200 12.000 ;
        RECT 215.800 12.300 216.600 15.200 ;
        RECT 218.800 15.200 219.600 19.800 ;
        RECT 218.800 14.600 221.000 15.200 ;
        RECT 218.800 12.300 219.600 13.200 ;
        RECT 215.800 11.700 219.600 12.300 ;
        RECT 214.400 9.600 215.000 11.400 ;
        RECT 215.800 10.800 216.600 11.700 ;
        RECT 218.800 11.600 219.600 11.700 ;
        RECT 220.400 11.600 221.000 14.600 ;
        RECT 193.200 9.400 194.000 9.600 ;
        RECT 188.600 9.000 194.000 9.400 ;
        RECT 187.800 8.800 194.000 9.000 ;
        RECT 195.000 9.000 203.600 9.600 ;
        RECT 185.200 8.000 186.800 8.800 ;
        RECT 187.800 8.200 189.200 8.800 ;
        RECT 195.000 8.200 195.600 9.000 ;
        RECT 202.800 8.800 203.600 9.000 ;
        RECT 206.000 9.000 215.000 9.600 ;
        RECT 206.000 8.800 206.800 9.000 ;
        RECT 186.200 7.600 186.800 8.000 ;
        RECT 189.800 7.600 195.600 8.200 ;
        RECT 196.200 7.600 198.800 8.400 ;
        RECT 183.600 6.800 185.600 7.400 ;
        RECT 186.200 6.800 190.400 7.600 ;
        RECT 185.000 6.200 185.600 6.800 ;
        RECT 185.000 5.600 186.000 6.200 ;
        RECT 185.200 2.200 186.000 5.600 ;
        RECT 188.400 2.200 189.200 6.800 ;
        RECT 191.600 2.200 192.400 5.000 ;
        RECT 193.200 2.200 194.000 5.000 ;
        RECT 194.800 2.200 195.600 7.000 ;
        RECT 198.000 2.200 198.800 7.000 ;
        RECT 201.200 2.200 202.000 8.400 ;
        RECT 209.200 7.600 211.800 8.400 ;
        RECT 204.400 6.800 208.600 7.600 ;
        RECT 202.800 2.200 203.600 5.000 ;
        RECT 204.400 2.200 205.200 5.000 ;
        RECT 206.000 2.200 206.800 5.000 ;
        RECT 209.200 2.200 210.000 7.600 ;
        RECT 214.400 7.400 215.000 9.000 ;
        RECT 212.400 6.800 215.000 7.400 ;
        RECT 215.600 10.000 216.600 10.800 ;
        RECT 220.400 10.800 221.600 11.600 ;
        RECT 220.400 10.200 221.000 10.800 ;
        RECT 212.400 2.200 213.200 6.800 ;
        RECT 215.600 2.200 216.400 10.000 ;
        RECT 218.800 9.600 221.000 10.200 ;
        RECT 218.800 2.200 219.600 9.600 ;
      LAYER via1 ;
        RECT 9.200 193.600 10.000 194.400 ;
        RECT 2.800 189.600 3.600 190.400 ;
        RECT 15.600 187.600 16.400 188.400 ;
        RECT 28.400 193.600 29.200 194.400 ;
        RECT 30.000 189.600 30.800 190.400 ;
        RECT 14.000 183.600 14.800 184.400 ;
        RECT 22.000 183.600 22.800 184.400 ;
        RECT 33.200 187.600 34.000 188.400 ;
        RECT 50.800 187.600 51.600 188.400 ;
        RECT 44.400 183.600 45.200 184.400 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 71.600 189.600 72.400 190.400 ;
        RECT 74.800 187.600 75.600 188.400 ;
        RECT 57.200 183.600 58.000 184.400 ;
        RECT 79.600 189.600 80.400 190.400 ;
        RECT 82.800 189.600 83.600 190.400 ;
        RECT 81.200 187.600 82.000 188.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 95.600 185.600 96.400 186.400 ;
        RECT 97.200 185.600 98.000 186.400 ;
        RECT 105.200 187.600 106.000 188.400 ;
        RECT 127.600 194.400 128.400 195.200 ;
        RECT 130.800 195.000 131.600 195.800 ;
        RECT 126.000 192.400 126.800 193.200 ;
        RECT 108.400 185.600 109.200 186.400 ;
        RECT 135.600 187.600 136.400 188.400 ;
        RECT 132.400 185.600 133.200 186.400 ;
        RECT 151.600 189.600 152.400 190.400 ;
        RECT 126.000 184.200 126.800 185.000 ;
        RECT 127.600 184.200 128.400 185.000 ;
        RECT 129.200 184.200 130.000 185.000 ;
        RECT 130.800 184.200 131.600 185.000 ;
        RECT 134.000 184.200 134.800 185.000 ;
        RECT 137.200 184.200 138.000 185.000 ;
        RECT 138.800 184.200 139.600 185.000 ;
        RECT 140.400 184.200 141.200 185.000 ;
        RECT 159.600 189.600 160.400 190.400 ;
        RECT 178.800 195.000 179.600 195.800 ;
        RECT 175.600 193.600 176.400 194.400 ;
        RECT 180.400 192.400 181.200 193.200 ;
        RECT 185.200 189.600 186.000 190.400 ;
        RECT 169.200 188.200 170.000 189.000 ;
        RECT 178.800 188.600 179.600 189.400 ;
        RECT 174.000 187.600 174.800 188.400 ;
        RECT 169.200 184.200 170.000 185.000 ;
        RECT 170.800 184.200 171.600 185.000 ;
        RECT 172.400 184.200 173.200 185.000 ;
        RECT 175.600 184.200 176.400 185.000 ;
        RECT 178.800 184.200 179.600 185.000 ;
        RECT 180.400 184.200 181.200 185.000 ;
        RECT 182.000 184.200 182.800 185.000 ;
        RECT 183.600 184.200 184.400 185.000 ;
        RECT 193.200 183.600 194.000 184.400 ;
        RECT 204.400 183.600 205.200 184.400 ;
        RECT 215.600 185.600 216.400 186.400 ;
        RECT 6.000 169.600 6.800 170.400 ;
        RECT 31.600 175.600 32.400 176.400 ;
        RECT 33.200 174.200 34.000 175.000 ;
        RECT 23.600 171.600 24.400 172.400 ;
        RECT 12.400 169.600 13.200 170.400 ;
        RECT 26.800 166.800 27.600 167.600 ;
        RECT 30.000 166.200 30.800 167.000 ;
        RECT 25.200 164.200 26.000 165.000 ;
        RECT 26.800 164.200 27.600 165.000 ;
        RECT 28.400 164.200 29.200 165.000 ;
        RECT 33.200 166.200 34.000 167.000 ;
        RECT 36.400 166.200 37.200 167.000 ;
        RECT 82.800 174.800 83.600 175.600 ;
        RECT 54.000 171.600 54.800 172.400 ;
        RECT 38.000 164.200 38.800 165.000 ;
        RECT 39.600 164.200 40.400 165.000 ;
        RECT 54.000 163.600 54.800 164.400 ;
        RECT 62.000 169.600 62.800 170.400 ;
        RECT 86.000 173.600 86.800 174.400 ;
        RECT 105.200 171.600 106.000 172.400 ;
        RECT 116.400 171.600 117.200 172.400 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 135.600 173.000 136.400 173.800 ;
        RECT 145.200 172.600 146.000 173.400 ;
        RECT 164.400 177.600 165.200 178.400 ;
        RECT 130.800 171.600 131.600 172.400 ;
        RECT 159.800 173.600 160.600 174.400 ;
        RECT 170.800 173.600 171.600 174.400 ;
        RECT 137.200 168.800 138.000 169.600 ;
        RECT 142.000 167.600 142.800 168.400 ;
        RECT 138.800 166.200 139.600 167.000 ;
        RECT 135.600 164.200 136.400 165.000 ;
        RECT 137.200 164.200 138.000 165.000 ;
        RECT 142.000 166.200 142.800 167.000 ;
        RECT 145.200 166.200 146.000 167.000 ;
        RECT 146.800 164.200 147.600 165.000 ;
        RECT 148.400 164.200 149.200 165.000 ;
        RECT 150.000 164.200 150.800 165.000 ;
        RECT 167.600 171.600 168.400 172.400 ;
        RECT 178.800 171.600 179.600 172.400 ;
        RECT 186.800 171.600 187.600 172.400 ;
        RECT 199.600 173.000 200.400 173.800 ;
        RECT 209.200 172.600 210.000 173.400 ;
        RECT 223.600 177.600 224.400 178.400 ;
        RECT 198.000 171.600 198.800 172.400 ;
        RECT 201.200 168.800 202.000 169.600 ;
        RECT 206.000 167.600 206.800 168.400 ;
        RECT 202.800 166.200 203.600 167.000 ;
        RECT 199.600 164.200 200.400 165.000 ;
        RECT 201.200 164.200 202.000 165.000 ;
        RECT 206.000 166.200 206.800 167.000 ;
        RECT 209.200 166.200 210.000 167.000 ;
        RECT 210.800 164.200 211.600 165.000 ;
        RECT 212.400 164.200 213.200 165.000 ;
        RECT 214.000 164.200 214.800 165.000 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 12.400 149.600 13.200 150.400 ;
        RECT 34.800 155.000 35.600 155.800 ;
        RECT 31.600 153.600 32.400 154.400 ;
        RECT 49.200 155.600 50.000 156.400 ;
        RECT 36.400 152.400 37.200 153.200 ;
        RECT 41.200 149.600 42.000 150.400 ;
        RECT 25.200 148.200 26.000 149.000 ;
        RECT 34.800 148.600 35.600 149.400 ;
        RECT 9.200 145.600 10.000 146.400 ;
        RECT 30.000 147.600 30.800 148.400 ;
        RECT 25.200 144.200 26.000 145.000 ;
        RECT 26.800 144.200 27.600 145.000 ;
        RECT 28.400 144.200 29.200 145.000 ;
        RECT 31.600 144.200 32.400 145.000 ;
        RECT 34.800 144.200 35.600 145.000 ;
        RECT 36.400 144.200 37.200 145.000 ;
        RECT 38.000 144.200 38.800 145.000 ;
        RECT 39.600 144.200 40.400 145.000 ;
        RECT 58.800 147.600 59.600 148.400 ;
        RECT 63.600 148.000 64.400 148.800 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 66.800 145.600 67.600 146.400 ;
        RECT 68.400 143.600 69.200 144.400 ;
        RECT 90.800 155.000 91.600 155.800 ;
        RECT 87.600 153.600 88.400 154.400 ;
        RECT 105.200 157.600 106.000 158.400 ;
        RECT 92.400 152.400 93.200 153.200 ;
        RECT 97.200 149.600 98.000 150.400 ;
        RECT 81.200 148.200 82.000 149.000 ;
        RECT 90.800 148.600 91.600 149.400 ;
        RECT 86.000 147.600 86.800 148.400 ;
        RECT 81.200 144.200 82.000 145.000 ;
        RECT 82.800 144.200 83.600 145.000 ;
        RECT 84.400 144.200 85.200 145.000 ;
        RECT 87.600 144.200 88.400 145.000 ;
        RECT 90.800 144.200 91.600 145.000 ;
        RECT 92.400 144.200 93.200 145.000 ;
        RECT 94.000 144.200 94.800 145.000 ;
        RECT 95.600 144.200 96.400 145.000 ;
        RECT 142.000 155.000 142.800 155.800 ;
        RECT 138.800 153.600 139.600 154.400 ;
        RECT 143.600 152.400 144.400 153.200 ;
        RECT 161.000 151.800 161.800 152.600 ;
        RECT 132.400 148.200 133.200 149.000 ;
        RECT 142.000 148.600 142.800 149.400 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 137.200 147.600 138.000 148.400 ;
        RECT 170.800 149.600 171.600 150.400 ;
        RECT 132.400 144.200 133.200 145.000 ;
        RECT 134.000 144.200 134.800 145.000 ;
        RECT 135.600 144.200 136.400 145.000 ;
        RECT 138.800 144.200 139.600 145.000 ;
        RECT 142.000 144.200 142.800 145.000 ;
        RECT 143.600 144.200 144.400 145.000 ;
        RECT 145.200 144.200 146.000 145.000 ;
        RECT 146.800 144.200 147.600 145.000 ;
        RECT 161.000 146.200 161.800 147.000 ;
        RECT 172.400 149.600 173.200 150.400 ;
        RECT 169.200 147.600 170.000 148.400 ;
        RECT 202.800 155.000 203.600 155.800 ;
        RECT 199.600 153.600 200.400 154.400 ;
        RECT 204.400 152.400 205.200 153.200 ;
        RECT 209.200 149.600 210.000 150.400 ;
        RECT 193.200 148.200 194.000 149.000 ;
        RECT 202.800 148.600 203.600 149.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 193.200 144.200 194.000 145.000 ;
        RECT 194.800 144.200 195.600 145.000 ;
        RECT 196.400 144.200 197.200 145.000 ;
        RECT 199.600 144.200 200.400 145.000 ;
        RECT 202.800 144.200 203.600 145.000 ;
        RECT 204.400 144.200 205.200 145.000 ;
        RECT 206.000 144.200 206.800 145.000 ;
        RECT 207.600 144.200 208.400 145.000 ;
        RECT 217.200 145.600 218.000 146.400 ;
        RECT 12.400 133.600 13.200 134.400 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 30.000 133.600 30.800 134.400 ;
        RECT 17.200 131.600 18.000 132.400 ;
        RECT 23.600 131.600 24.400 132.400 ;
        RECT 18.800 123.600 19.600 124.400 ;
        RECT 34.800 123.600 35.600 124.400 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 49.200 123.600 50.000 124.400 ;
        RECT 55.600 123.600 56.400 124.400 ;
        RECT 70.000 137.600 70.800 138.400 ;
        RECT 86.000 135.600 86.800 136.400 ;
        RECT 87.600 134.200 88.400 135.000 ;
        RECT 78.000 131.600 78.800 132.400 ;
        RECT 60.400 127.600 61.200 128.400 ;
        RECT 81.200 126.800 82.000 127.600 ;
        RECT 84.400 126.200 85.200 127.000 ;
        RECT 79.600 124.200 80.400 125.000 ;
        RECT 81.200 124.200 82.000 125.000 ;
        RECT 82.800 124.200 83.600 125.000 ;
        RECT 87.600 126.200 88.400 127.000 ;
        RECT 90.800 126.200 91.600 127.000 ;
        RECT 137.200 137.600 138.000 138.400 ;
        RECT 145.200 137.600 146.000 138.400 ;
        RECT 105.200 133.600 106.000 134.400 ;
        RECT 92.400 124.200 93.200 125.000 ;
        RECT 94.000 124.200 94.800 125.000 ;
        RECT 143.600 133.600 144.400 134.400 ;
        RECT 164.400 137.600 165.200 138.400 ;
        RECT 130.800 123.600 131.600 124.400 ;
        RECT 174.000 133.600 174.800 134.400 ;
        RECT 175.600 131.600 176.400 132.400 ;
        RECT 199.600 135.600 200.400 136.400 ;
        RECT 201.200 134.200 202.000 135.000 ;
        RECT 202.800 131.600 203.600 132.400 ;
        RECT 209.200 131.600 210.000 132.400 ;
        RECT 194.800 126.800 195.600 127.600 ;
        RECT 198.000 126.200 198.800 127.000 ;
        RECT 193.200 124.200 194.000 125.000 ;
        RECT 194.800 124.200 195.600 125.000 ;
        RECT 196.400 124.200 197.200 125.000 ;
        RECT 201.200 126.200 202.000 127.000 ;
        RECT 204.400 126.200 205.200 127.000 ;
        RECT 206.000 124.200 206.800 125.000 ;
        RECT 207.600 124.200 208.400 125.000 ;
        RECT 7.600 117.600 8.400 118.400 ;
        RECT 18.800 114.400 19.600 115.200 ;
        RECT 22.000 115.000 22.800 115.800 ;
        RECT 44.400 117.600 45.200 118.400 ;
        RECT 17.200 112.400 18.000 113.200 ;
        RECT 26.800 107.600 27.600 108.400 ;
        RECT 23.600 105.600 24.400 106.400 ;
        RECT 17.200 104.200 18.000 105.000 ;
        RECT 18.800 104.200 19.600 105.000 ;
        RECT 20.400 104.200 21.200 105.000 ;
        RECT 22.000 104.200 22.800 105.000 ;
        RECT 25.200 104.200 26.000 105.000 ;
        RECT 28.400 104.200 29.200 105.000 ;
        RECT 30.000 104.200 30.800 105.000 ;
        RECT 31.600 104.200 32.400 105.000 ;
        RECT 42.800 105.600 43.600 106.400 ;
        RECT 71.600 117.600 72.400 118.400 ;
        RECT 65.200 113.600 66.000 114.400 ;
        RECT 73.200 113.600 74.000 114.400 ;
        RECT 54.000 105.600 54.800 106.400 ;
        RECT 49.200 103.600 50.000 104.400 ;
        RECT 68.400 111.600 69.200 112.400 ;
        RECT 70.000 111.600 70.800 112.400 ;
        RECT 66.800 109.600 67.600 110.400 ;
        RECT 82.800 117.600 83.600 118.400 ;
        RECT 62.000 107.600 62.800 108.400 ;
        RECT 65.200 103.600 66.000 104.400 ;
        RECT 76.400 107.600 77.200 108.400 ;
        RECT 94.000 113.600 94.800 114.400 ;
        RECT 86.000 109.600 86.800 110.400 ;
        RECT 95.600 107.600 96.400 108.400 ;
        RECT 78.000 103.600 78.800 104.400 ;
        RECT 102.000 109.600 102.800 110.400 ;
        RECT 105.200 107.600 106.000 108.400 ;
        RECT 98.800 103.600 99.600 104.400 ;
        RECT 103.600 105.600 104.400 106.400 ;
        RECT 126.000 117.600 126.800 118.400 ;
        RECT 119.600 109.600 120.400 110.400 ;
        RECT 121.200 109.600 122.000 110.400 ;
        RECT 118.000 103.600 118.800 104.400 ;
        RECT 154.800 115.000 155.600 115.800 ;
        RECT 151.600 113.600 152.400 114.400 ;
        RECT 156.400 112.400 157.200 113.200 ;
        RECT 161.200 109.600 162.000 110.400 ;
        RECT 145.200 108.200 146.000 109.000 ;
        RECT 154.800 108.600 155.600 109.400 ;
        RECT 132.400 103.600 133.200 104.400 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 145.200 104.200 146.000 105.000 ;
        RECT 146.800 104.200 147.600 105.000 ;
        RECT 148.400 104.200 149.200 105.000 ;
        RECT 151.600 104.200 152.400 105.000 ;
        RECT 154.800 104.200 155.600 105.000 ;
        RECT 156.400 104.200 157.200 105.000 ;
        RECT 158.000 104.200 158.800 105.000 ;
        RECT 159.600 104.200 160.400 105.000 ;
        RECT 198.000 115.000 198.800 115.800 ;
        RECT 194.800 113.600 195.600 114.400 ;
        RECT 199.600 112.400 200.400 113.200 ;
        RECT 204.400 109.600 205.200 110.400 ;
        RECT 188.400 108.200 189.200 109.000 ;
        RECT 198.000 108.600 198.800 109.400 ;
        RECT 174.000 105.600 174.800 106.400 ;
        RECT 169.200 103.600 170.000 104.400 ;
        RECT 193.200 107.600 194.000 108.400 ;
        RECT 188.400 104.200 189.200 105.000 ;
        RECT 190.000 104.200 190.800 105.000 ;
        RECT 191.600 104.200 192.400 105.000 ;
        RECT 194.800 104.200 195.600 105.000 ;
        RECT 198.000 104.200 198.800 105.000 ;
        RECT 199.600 104.200 200.400 105.000 ;
        RECT 201.200 104.200 202.000 105.000 ;
        RECT 202.800 104.200 203.600 105.000 ;
        RECT 212.400 105.600 213.200 106.400 ;
        RECT 218.800 109.600 219.600 110.400 ;
        RECT 217.200 105.600 218.000 106.400 ;
        RECT 215.600 103.600 216.400 104.400 ;
        RECT 15.600 85.600 16.400 86.400 ;
        RECT 54.000 93.600 54.800 94.400 ;
        RECT 34.800 89.600 35.600 90.400 ;
        RECT 39.600 89.600 40.400 90.400 ;
        RECT 46.000 89.600 46.800 90.400 ;
        RECT 78.000 95.600 78.800 96.400 ;
        RECT 79.600 94.200 80.400 95.000 ;
        RECT 103.600 97.600 104.400 98.400 ;
        RECT 89.200 91.600 90.000 92.400 ;
        RECT 62.000 83.600 62.800 84.400 ;
        RECT 73.200 86.800 74.000 87.600 ;
        RECT 76.400 86.200 77.200 87.000 ;
        RECT 71.600 84.200 72.400 85.000 ;
        RECT 73.200 84.200 74.000 85.000 ;
        RECT 74.800 84.200 75.600 85.000 ;
        RECT 79.600 86.200 80.400 87.000 ;
        RECT 82.800 86.200 83.600 87.000 ;
        RECT 119.600 95.600 120.400 96.400 ;
        RECT 121.200 94.200 122.000 95.000 ;
        RECT 140.400 93.600 141.200 94.400 ;
        RECT 111.600 91.600 112.400 92.400 ;
        RECT 130.800 91.600 131.600 92.400 ;
        RECT 84.400 84.200 85.200 85.000 ;
        RECT 86.000 84.200 86.800 85.000 ;
        RECT 114.800 86.800 115.600 87.600 ;
        RECT 118.000 86.200 118.800 87.000 ;
        RECT 113.200 84.200 114.000 85.000 ;
        RECT 114.800 84.200 115.600 85.000 ;
        RECT 116.400 84.200 117.200 85.000 ;
        RECT 121.200 86.200 122.000 87.000 ;
        RECT 124.400 86.200 125.200 87.000 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 151.600 91.600 152.400 92.400 ;
        RECT 172.400 97.600 173.200 98.400 ;
        RECT 178.800 97.600 179.600 98.400 ;
        RECT 162.800 94.800 163.600 95.600 ;
        RECT 126.000 84.200 126.800 85.000 ;
        RECT 127.600 84.200 128.400 85.000 ;
        RECT 145.200 87.600 146.000 88.400 ;
        RECT 172.400 89.600 173.200 90.400 ;
        RECT 190.000 93.000 190.800 93.800 ;
        RECT 178.800 89.600 179.600 90.400 ;
        RECT 199.600 92.600 200.400 93.400 ;
        RECT 185.200 91.600 186.000 92.400 ;
        RECT 191.600 88.800 192.400 89.600 ;
        RECT 196.400 87.600 197.200 88.400 ;
        RECT 193.200 86.200 194.000 87.000 ;
        RECT 190.000 84.200 190.800 85.000 ;
        RECT 191.600 84.200 192.400 85.000 ;
        RECT 196.400 86.200 197.200 87.000 ;
        RECT 199.600 86.200 200.400 87.000 ;
        RECT 201.200 84.200 202.000 85.000 ;
        RECT 202.800 84.200 203.600 85.000 ;
        RECT 204.400 84.200 205.200 85.000 ;
        RECT 214.000 83.600 214.800 84.400 ;
        RECT 223.600 91.600 224.400 92.400 ;
        RECT 12.400 77.600 13.200 78.400 ;
        RECT 23.600 74.400 24.400 75.200 ;
        RECT 26.800 75.000 27.600 75.800 ;
        RECT 22.000 72.400 22.800 73.200 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 28.400 65.600 29.200 66.400 ;
        RECT 22.000 64.200 22.800 65.000 ;
        RECT 23.600 64.200 24.400 65.000 ;
        RECT 25.200 64.200 26.000 65.000 ;
        RECT 26.800 64.200 27.600 65.000 ;
        RECT 30.000 64.200 30.800 65.000 ;
        RECT 33.200 64.200 34.000 65.000 ;
        RECT 34.800 64.200 35.600 65.000 ;
        RECT 36.400 64.200 37.200 65.000 ;
        RECT 58.800 77.600 59.600 78.400 ;
        RECT 52.400 73.600 53.200 74.400 ;
        RECT 49.200 69.600 50.000 70.400 ;
        RECT 47.600 65.600 48.400 66.400 ;
        RECT 55.600 71.600 56.400 72.400 ;
        RECT 57.200 71.600 58.000 72.400 ;
        RECT 66.800 73.600 67.600 74.400 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 66.800 69.600 67.600 70.400 ;
        RECT 82.800 71.600 83.600 72.400 ;
        RECT 68.400 67.600 69.200 68.400 ;
        RECT 79.600 67.600 80.400 68.400 ;
        RECT 86.000 69.600 86.800 70.400 ;
        RECT 106.800 75.000 107.600 75.800 ;
        RECT 103.600 73.600 104.400 74.400 ;
        RECT 108.400 72.400 109.200 73.200 ;
        RECT 121.200 73.600 122.000 74.400 ;
        RECT 97.200 68.200 98.000 69.000 ;
        RECT 106.800 68.600 107.600 69.400 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 97.200 64.200 98.000 65.000 ;
        RECT 98.800 64.200 99.600 65.000 ;
        RECT 100.400 64.200 101.200 65.000 ;
        RECT 103.600 64.200 104.400 65.000 ;
        RECT 106.800 64.200 107.600 65.000 ;
        RECT 108.400 64.200 109.200 65.000 ;
        RECT 110.000 64.200 110.800 65.000 ;
        RECT 111.600 64.200 112.400 65.000 ;
        RECT 143.600 75.000 144.400 75.800 ;
        RECT 140.400 73.600 141.200 74.400 ;
        RECT 145.200 72.400 146.000 73.200 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 134.000 68.200 134.800 69.000 ;
        RECT 143.600 68.600 144.400 69.400 ;
        RECT 138.800 67.600 139.600 68.400 ;
        RECT 134.000 64.200 134.800 65.000 ;
        RECT 135.600 64.200 136.400 65.000 ;
        RECT 137.200 64.200 138.000 65.000 ;
        RECT 140.400 64.200 141.200 65.000 ;
        RECT 143.600 64.200 144.400 65.000 ;
        RECT 145.200 64.200 146.000 65.000 ;
        RECT 146.800 64.200 147.600 65.000 ;
        RECT 148.400 64.200 149.200 65.000 ;
        RECT 178.800 75.000 179.600 75.800 ;
        RECT 175.600 73.600 176.400 74.400 ;
        RECT 180.400 72.400 181.200 73.200 ;
        RECT 185.200 69.600 186.000 70.400 ;
        RECT 169.200 68.200 170.000 69.000 ;
        RECT 178.800 68.600 179.600 69.400 ;
        RECT 158.000 63.600 158.800 64.400 ;
        RECT 174.000 67.600 174.800 68.400 ;
        RECT 169.200 64.200 170.000 65.000 ;
        RECT 170.800 64.200 171.600 65.000 ;
        RECT 172.400 64.200 173.200 65.000 ;
        RECT 175.600 64.200 176.400 65.000 ;
        RECT 178.800 64.200 179.600 65.000 ;
        RECT 180.400 64.200 181.200 65.000 ;
        RECT 182.000 64.200 182.800 65.000 ;
        RECT 183.600 64.200 184.400 65.000 ;
        RECT 198.000 65.600 198.800 66.400 ;
        RECT 212.400 69.600 213.200 70.400 ;
        RECT 204.400 65.600 205.200 66.400 ;
        RECT 207.600 65.600 208.400 66.400 ;
        RECT 217.200 69.600 218.000 70.400 ;
        RECT 7.600 55.600 8.400 56.400 ;
        RECT 23.600 55.600 24.400 56.400 ;
        RECT 25.200 54.200 26.000 55.000 ;
        RECT 34.800 51.600 35.600 52.400 ;
        RECT 38.000 51.600 38.800 52.400 ;
        RECT 18.800 46.800 19.600 47.600 ;
        RECT 22.000 46.200 22.800 47.000 ;
        RECT 17.200 44.200 18.000 45.000 ;
        RECT 18.800 44.200 19.600 45.000 ;
        RECT 20.400 44.200 21.200 45.000 ;
        RECT 25.200 46.200 26.000 47.000 ;
        RECT 28.400 46.200 29.200 47.000 ;
        RECT 30.000 44.200 30.800 45.000 ;
        RECT 31.600 44.200 32.400 45.000 ;
        RECT 49.200 53.600 50.000 54.400 ;
        RECT 50.800 51.600 51.600 52.400 ;
        RECT 52.400 43.600 53.200 44.400 ;
        RECT 57.200 45.600 58.000 46.400 ;
        RECT 66.600 51.600 67.400 52.400 ;
        RECT 82.800 55.600 83.600 56.400 ;
        RECT 84.400 54.200 85.200 55.000 ;
        RECT 103.600 55.600 104.400 56.400 ;
        RECT 94.000 51.600 94.800 52.400 ;
        RECT 62.000 47.600 62.800 48.400 ;
        RECT 78.000 46.800 78.800 47.600 ;
        RECT 81.200 46.200 82.000 47.000 ;
        RECT 76.400 44.200 77.200 45.000 ;
        RECT 78.000 44.200 78.800 45.000 ;
        RECT 79.600 44.200 80.400 45.000 ;
        RECT 84.400 46.200 85.200 47.000 ;
        RECT 87.600 46.200 88.400 47.000 ;
        RECT 89.200 44.200 90.000 45.000 ;
        RECT 90.800 44.200 91.600 45.000 ;
        RECT 121.200 57.600 122.000 58.400 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 145.200 55.600 146.000 56.400 ;
        RECT 146.800 54.200 147.600 55.000 ;
        RECT 137.200 51.600 138.000 52.400 ;
        RECT 159.600 51.600 160.400 52.400 ;
        RECT 116.400 43.600 117.200 44.400 ;
        RECT 122.800 43.600 123.600 44.400 ;
        RECT 140.400 46.800 141.200 47.600 ;
        RECT 143.600 46.200 144.400 47.000 ;
        RECT 138.800 44.200 139.600 45.000 ;
        RECT 140.400 44.200 141.200 45.000 ;
        RECT 142.000 44.200 142.800 45.000 ;
        RECT 146.800 46.200 147.600 47.000 ;
        RECT 150.000 46.200 150.800 47.000 ;
        RECT 169.200 57.600 170.000 58.400 ;
        RECT 151.600 44.200 152.400 45.000 ;
        RECT 153.200 44.200 154.000 45.000 ;
        RECT 164.400 43.600 165.200 44.400 ;
        RECT 194.800 53.000 195.600 53.800 ;
        RECT 183.600 49.600 184.400 50.400 ;
        RECT 204.400 52.600 205.200 53.400 ;
        RECT 223.600 57.600 224.400 58.400 ;
        RECT 193.200 51.600 194.000 52.400 ;
        RECT 196.400 48.800 197.200 49.600 ;
        RECT 201.200 47.600 202.000 48.400 ;
        RECT 198.000 46.200 198.800 47.000 ;
        RECT 194.800 44.200 195.600 45.000 ;
        RECT 196.400 44.200 197.200 45.000 ;
        RECT 201.200 46.200 202.000 47.000 ;
        RECT 204.400 46.200 205.200 47.000 ;
        RECT 206.000 44.200 206.800 45.000 ;
        RECT 207.600 44.200 208.400 45.000 ;
        RECT 209.200 44.200 210.000 45.000 ;
        RECT 218.800 43.600 219.600 44.400 ;
        RECT 2.800 37.600 3.600 38.400 ;
        RECT 14.000 34.400 14.800 35.200 ;
        RECT 17.200 35.000 18.000 35.800 ;
        RECT 12.400 32.400 13.200 33.200 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 18.800 25.600 19.600 26.400 ;
        RECT 12.400 24.200 13.200 25.000 ;
        RECT 14.000 24.200 14.800 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 17.200 24.200 18.000 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 26.800 24.200 27.600 25.000 ;
        RECT 49.200 29.600 50.000 30.400 ;
        RECT 66.800 34.400 67.600 35.200 ;
        RECT 70.000 35.000 70.800 35.800 ;
        RECT 65.200 32.400 66.000 33.200 ;
        RECT 55.400 29.600 56.200 30.400 ;
        RECT 44.400 25.600 45.200 26.400 ;
        RECT 52.400 27.600 53.200 28.400 ;
        RECT 74.800 27.600 75.600 28.400 ;
        RECT 71.600 25.600 72.400 26.400 ;
        RECT 105.200 33.600 106.000 34.400 ;
        RECT 65.200 24.200 66.000 25.000 ;
        RECT 66.800 24.200 67.600 25.000 ;
        RECT 68.400 24.200 69.200 25.000 ;
        RECT 70.000 24.200 70.800 25.000 ;
        RECT 73.200 24.200 74.000 25.000 ;
        RECT 76.400 24.200 77.200 25.000 ;
        RECT 78.000 24.200 78.800 25.000 ;
        RECT 79.600 24.200 80.400 25.000 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 100.400 23.600 101.200 24.400 ;
        RECT 129.200 35.000 130.000 35.800 ;
        RECT 126.000 33.600 126.800 34.400 ;
        RECT 130.800 32.400 131.600 33.200 ;
        RECT 135.600 29.600 136.400 30.400 ;
        RECT 119.600 28.200 120.400 29.000 ;
        RECT 129.200 28.600 130.000 29.400 ;
        RECT 124.400 27.600 125.200 28.400 ;
        RECT 119.600 24.200 120.400 25.000 ;
        RECT 121.200 24.200 122.000 25.000 ;
        RECT 122.800 24.200 123.600 25.000 ;
        RECT 126.000 24.200 126.800 25.000 ;
        RECT 129.200 24.200 130.000 25.000 ;
        RECT 130.800 24.200 131.600 25.000 ;
        RECT 132.400 24.200 133.200 25.000 ;
        RECT 134.000 24.200 134.800 25.000 ;
        RECT 148.400 25.600 149.200 26.400 ;
        RECT 174.000 34.400 174.800 35.200 ;
        RECT 177.200 35.000 178.000 35.800 ;
        RECT 172.400 32.400 173.200 33.200 ;
        RECT 158.000 29.600 158.800 30.400 ;
        RECT 159.600 29.600 160.400 30.400 ;
        RECT 170.800 29.600 171.600 30.400 ;
        RECT 162.800 23.600 163.600 24.400 ;
        RECT 182.000 27.600 182.800 28.400 ;
        RECT 178.800 25.600 179.600 26.400 ;
        RECT 172.400 24.200 173.200 25.000 ;
        RECT 174.000 24.200 174.800 25.000 ;
        RECT 175.600 24.200 176.400 25.000 ;
        RECT 177.200 24.200 178.000 25.000 ;
        RECT 180.400 24.200 181.200 25.000 ;
        RECT 183.600 24.200 184.400 25.000 ;
        RECT 185.200 24.200 186.000 25.000 ;
        RECT 186.800 24.200 187.600 25.000 ;
        RECT 212.400 37.600 213.200 38.400 ;
        RECT 207.600 29.600 208.400 30.400 ;
        RECT 209.200 29.600 210.000 30.400 ;
        RECT 206.000 25.600 206.800 26.400 ;
        RECT 218.800 25.600 219.600 26.400 ;
        RECT 2.800 15.600 3.600 16.400 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 20.400 14.200 21.200 15.000 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 14.000 6.800 14.800 7.600 ;
        RECT 17.200 6.200 18.000 7.000 ;
        RECT 12.400 4.200 13.200 5.000 ;
        RECT 14.000 4.200 14.800 5.000 ;
        RECT 15.600 4.200 16.400 5.000 ;
        RECT 20.400 6.200 21.200 7.000 ;
        RECT 23.600 6.200 24.400 7.000 ;
        RECT 25.200 4.200 26.000 5.000 ;
        RECT 26.800 4.200 27.600 5.000 ;
        RECT 63.600 15.600 64.400 16.400 ;
        RECT 65.200 14.200 66.000 15.000 ;
        RECT 55.600 11.600 56.400 12.400 ;
        RECT 76.400 11.600 77.200 12.400 ;
        RECT 58.800 6.800 59.600 7.600 ;
        RECT 62.000 6.200 62.800 7.000 ;
        RECT 57.200 4.200 58.000 5.000 ;
        RECT 58.800 4.200 59.600 5.000 ;
        RECT 60.400 4.200 61.200 5.000 ;
        RECT 65.200 6.200 66.000 7.000 ;
        RECT 68.400 6.200 69.200 7.000 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 105.200 13.000 106.000 13.800 ;
        RECT 70.000 4.200 70.800 5.000 ;
        RECT 71.600 4.200 72.400 5.000 ;
        RECT 114.800 12.600 115.600 13.400 ;
        RECT 100.400 11.600 101.200 12.400 ;
        RECT 106.800 8.800 107.600 9.600 ;
        RECT 111.600 7.600 112.400 8.400 ;
        RECT 108.400 6.200 109.200 7.000 ;
        RECT 105.200 4.200 106.000 5.000 ;
        RECT 106.800 4.200 107.600 5.000 ;
        RECT 111.600 6.200 112.400 7.000 ;
        RECT 114.800 6.200 115.600 7.000 ;
        RECT 116.400 4.200 117.200 5.000 ;
        RECT 118.000 4.200 118.800 5.000 ;
        RECT 119.600 4.200 120.400 5.000 ;
        RECT 167.600 17.600 168.400 18.400 ;
        RECT 156.400 11.600 157.200 12.400 ;
        RECT 166.000 13.600 166.800 14.400 ;
        RECT 191.600 13.000 192.400 13.800 ;
        RECT 201.200 12.600 202.000 13.400 ;
        RECT 215.600 17.600 216.400 18.400 ;
        RECT 190.000 11.600 190.800 12.400 ;
        RECT 193.200 8.800 194.000 9.600 ;
        RECT 198.000 7.600 198.800 8.400 ;
        RECT 194.800 6.200 195.600 7.000 ;
        RECT 191.600 4.200 192.400 5.000 ;
        RECT 193.200 4.200 194.000 5.000 ;
        RECT 198.000 6.200 198.800 7.000 ;
        RECT 201.200 6.200 202.000 7.000 ;
        RECT 202.800 4.200 203.600 5.000 ;
        RECT 204.400 4.200 205.200 5.000 ;
        RECT 206.000 4.200 206.800 5.000 ;
      LAYER metal2 ;
        RECT 9.200 193.600 10.000 194.400 ;
        RECT 28.400 193.600 29.200 194.400 ;
        RECT 12.400 191.600 13.200 192.400 ;
        RECT 33.200 191.600 34.000 192.400 ;
        RECT 36.400 191.600 37.200 192.400 ;
        RECT 74.800 192.300 75.600 192.400 ;
        RECT 73.300 191.700 75.600 192.300 ;
        RECT 12.500 190.400 13.100 191.600 ;
        RECT 2.800 189.600 3.600 190.400 ;
        RECT 7.600 189.600 8.400 190.400 ;
        RECT 12.400 189.600 13.200 190.400 ;
        RECT 25.200 189.600 26.000 190.400 ;
        RECT 30.000 189.600 30.800 190.400 ;
        RECT 2.900 180.400 3.500 189.600 ;
        RECT 7.700 188.400 8.300 189.600 ;
        RECT 33.300 188.400 33.900 191.600 ;
        RECT 36.500 190.400 37.100 191.600 ;
        RECT 36.400 189.600 37.200 190.400 ;
        RECT 71.600 189.600 72.400 190.400 ;
        RECT 7.600 187.600 8.400 188.400 ;
        RECT 15.600 187.600 16.400 188.400 ;
        RECT 23.600 187.600 24.400 188.400 ;
        RECT 25.200 187.600 26.000 188.400 ;
        RECT 33.200 187.600 34.000 188.400 ;
        RECT 50.800 187.600 51.600 188.400 ;
        RECT 23.700 186.400 24.300 187.600 ;
        RECT 33.300 186.400 33.900 187.600 ;
        RECT 50.900 186.400 51.500 187.600 ;
        RECT 23.600 185.600 24.400 186.400 ;
        RECT 33.200 185.600 34.000 186.400 ;
        RECT 50.800 185.600 51.600 186.400 ;
        RECT 58.800 185.600 59.600 186.400 ;
        RECT 60.400 185.600 61.200 186.400 ;
        RECT 58.900 184.400 59.500 185.600 ;
        RECT 14.000 183.600 14.800 184.400 ;
        RECT 22.000 183.600 22.800 184.400 ;
        RECT 38.000 183.600 38.800 184.400 ;
        RECT 44.400 183.600 45.200 184.400 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 57.200 183.600 58.000 184.400 ;
        RECT 58.800 183.600 59.600 184.400 ;
        RECT 2.800 179.600 3.600 180.400 ;
        RECT 2.900 172.400 3.500 179.600 ;
        RECT 7.600 177.600 8.400 178.400 ;
        RECT 7.700 174.400 8.300 177.600 ;
        RECT 14.100 176.400 14.700 183.600 ;
        RECT 22.100 178.400 22.700 183.600 ;
        RECT 38.100 180.400 38.700 183.600 ;
        RECT 38.000 179.600 38.800 180.400 ;
        RECT 22.000 177.600 22.800 178.400 ;
        RECT 14.000 175.600 14.800 176.400 ;
        RECT 22.000 175.600 22.800 176.400 ;
        RECT 7.600 173.600 8.400 174.400 ;
        RECT 14.000 173.600 14.800 174.400 ;
        RECT 2.800 171.600 3.600 172.400 ;
        RECT 6.000 169.600 6.800 170.400 ;
        RECT 12.400 169.600 13.200 170.400 ;
        RECT 12.500 158.400 13.100 169.600 ;
        RECT 14.000 167.600 14.800 168.400 ;
        RECT 12.400 157.600 13.200 158.400 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 6.000 149.600 6.800 150.400 ;
        RECT 12.400 149.600 13.200 150.400 ;
        RECT 4.500 136.300 5.100 149.600 ;
        RECT 12.500 148.400 13.100 149.600 ;
        RECT 10.800 147.600 11.600 148.400 ;
        RECT 12.400 147.600 13.200 148.400 ;
        RECT 9.200 145.600 10.000 146.400 ;
        RECT 9.300 136.400 9.900 145.600 ;
        RECT 6.000 136.300 6.800 136.400 ;
        RECT 4.500 135.700 6.800 136.300 ;
        RECT 6.000 135.600 6.800 135.700 ;
        RECT 7.600 135.600 8.400 136.400 ;
        RECT 9.200 135.600 10.000 136.400 ;
        RECT 6.100 134.400 6.700 135.600 ;
        RECT 4.400 133.600 5.200 134.400 ;
        RECT 6.000 133.600 6.800 134.400 ;
        RECT 4.500 132.400 5.100 133.600 ;
        RECT 2.800 131.600 3.600 132.400 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 1.200 129.600 2.000 130.400 ;
        RECT 1.300 118.400 1.900 129.600 ;
        RECT 7.700 118.400 8.300 135.600 ;
        RECT 10.900 132.400 11.500 147.600 ;
        RECT 14.100 136.400 14.700 167.600 ;
        RECT 15.600 151.600 16.400 152.400 ;
        RECT 14.000 135.600 14.800 136.400 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 12.400 133.600 13.200 134.400 ;
        RECT 10.800 131.600 11.600 132.400 ;
        RECT 12.500 130.400 13.100 133.600 ;
        RECT 12.400 129.600 13.200 130.400 ;
        RECT 15.700 128.400 16.300 135.600 ;
        RECT 22.100 134.400 22.700 175.600 ;
        RECT 23.600 171.600 24.400 172.400 ;
        RECT 23.700 150.400 24.300 171.600 ;
        RECT 25.200 164.200 26.000 177.800 ;
        RECT 26.800 164.200 27.600 177.800 ;
        RECT 28.400 164.200 29.200 177.800 ;
        RECT 30.000 166.200 30.800 177.800 ;
        RECT 31.600 175.600 32.400 176.400 ;
        RECT 31.700 164.300 32.300 175.600 ;
        RECT 33.200 166.200 34.000 177.800 ;
        RECT 34.800 173.600 35.600 174.400 ;
        RECT 36.400 166.200 37.200 177.800 ;
        RECT 31.700 163.700 33.900 164.300 ;
        RECT 38.000 164.200 38.800 177.800 ;
        RECT 39.600 164.200 40.400 177.800 ;
        RECT 44.500 172.400 45.100 183.600 ;
        RECT 52.500 176.400 53.100 183.600 ;
        RECT 54.000 179.600 54.800 180.400 ;
        RECT 52.400 175.600 53.200 176.400 ;
        RECT 54.100 172.400 54.700 179.600 ;
        RECT 57.300 178.400 57.900 183.600 ;
        RECT 71.700 180.400 72.300 189.600 ;
        RECT 58.800 179.600 59.600 180.400 ;
        RECT 71.600 179.600 72.400 180.400 ;
        RECT 57.200 177.600 58.000 178.400 ;
        RECT 58.900 176.400 59.500 179.600 ;
        RECT 62.000 177.600 62.800 178.400 ;
        RECT 58.800 175.600 59.600 176.400 ;
        RECT 55.600 173.600 56.400 174.400 ;
        RECT 44.400 171.600 45.200 172.400 ;
        RECT 52.400 171.600 53.200 172.400 ;
        RECT 54.000 171.600 54.800 172.400 ;
        RECT 52.500 168.400 53.100 171.600 ;
        RECT 55.700 170.400 56.300 173.600 ;
        RECT 58.900 172.400 59.500 175.600 ;
        RECT 58.800 171.600 59.600 172.400 ;
        RECT 62.100 170.400 62.700 177.600 ;
        RECT 73.300 174.400 73.900 191.700 ;
        RECT 74.800 191.600 75.600 191.700 ;
        RECT 87.600 191.600 88.400 192.400 ;
        RECT 79.600 189.600 80.400 190.400 ;
        RECT 82.800 189.600 83.600 190.400 ;
        RECT 74.800 187.600 75.600 188.400 ;
        RECT 79.700 186.400 80.300 189.600 ;
        RECT 81.200 187.600 82.000 188.400 ;
        RECT 87.700 186.400 88.300 191.600 ;
        RECT 100.400 189.600 101.200 190.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 95.600 187.600 96.400 188.400 ;
        RECT 74.800 185.600 75.600 186.400 ;
        RECT 79.600 185.600 80.400 186.400 ;
        RECT 87.600 185.600 88.400 186.400 ;
        RECT 92.400 185.600 93.200 186.400 ;
        RECT 95.600 185.600 96.400 186.400 ;
        RECT 97.200 185.600 98.000 186.400 ;
        RECT 74.900 174.400 75.500 185.600 ;
        RECT 78.000 175.000 78.800 175.800 ;
        RECT 84.200 175.600 85.000 175.800 ;
        RECT 79.400 175.000 85.000 175.600 ;
        RECT 63.600 173.600 64.400 174.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 73.200 173.600 74.000 174.400 ;
        RECT 74.800 173.600 75.600 174.400 ;
        RECT 76.400 173.600 77.200 174.400 ;
        RECT 78.000 174.200 78.600 175.000 ;
        RECT 79.400 174.800 80.200 175.000 ;
        RECT 82.800 174.800 83.600 175.000 ;
        RECT 78.000 173.600 83.600 174.200 ;
        RECT 55.600 169.600 56.400 170.400 ;
        RECT 58.800 169.600 59.600 170.400 ;
        RECT 62.000 169.600 62.800 170.400 ;
        RECT 52.400 167.600 53.200 168.400 ;
        RECT 23.600 149.600 24.400 150.400 ;
        RECT 25.200 144.200 26.000 157.800 ;
        RECT 26.800 144.200 27.600 157.800 ;
        RECT 28.400 144.200 29.200 155.800 ;
        RECT 30.000 153.600 30.800 154.400 ;
        RECT 30.100 148.400 30.700 153.600 ;
        RECT 30.000 147.600 30.800 148.400 ;
        RECT 31.600 144.200 32.400 155.800 ;
        RECT 33.300 146.400 33.900 163.700 ;
        RECT 54.000 163.600 54.800 164.400 ;
        RECT 33.200 145.600 34.000 146.400 ;
        RECT 25.200 135.600 26.000 136.400 ;
        RECT 30.000 135.600 30.800 136.400 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 17.200 131.600 18.000 132.400 ;
        RECT 23.600 131.600 24.400 132.400 ;
        RECT 23.700 128.400 24.300 131.600 ;
        RECT 15.600 127.600 16.400 128.400 ;
        RECT 23.600 127.600 24.400 128.400 ;
        RECT 1.200 117.600 2.000 118.400 ;
        RECT 7.600 117.600 8.400 118.400 ;
        RECT 14.000 105.600 14.800 106.400 ;
        RECT 10.800 99.600 11.600 100.400 ;
        RECT 7.600 95.600 8.400 96.400 ;
        RECT 7.700 92.400 8.300 95.600 ;
        RECT 6.000 91.600 6.800 92.400 ;
        RECT 7.600 91.600 8.400 92.400 ;
        RECT 10.900 90.400 11.500 99.600 ;
        RECT 12.400 91.600 13.200 92.400 ;
        RECT 10.800 89.600 11.600 90.400 ;
        RECT 14.100 90.300 14.700 105.600 ;
        RECT 15.700 100.400 16.300 127.600 ;
        RECT 18.800 123.600 19.600 124.400 ;
        RECT 18.900 120.400 19.500 123.600 ;
        RECT 18.800 119.600 19.600 120.400 ;
        RECT 25.300 118.400 25.900 135.600 ;
        RECT 30.100 134.400 30.700 135.600 ;
        RECT 30.000 133.600 30.800 134.400 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 30.100 124.400 30.700 131.600 ;
        RECT 30.000 123.600 30.800 124.400 ;
        RECT 26.800 119.600 27.600 120.400 ;
        RECT 17.200 104.200 18.000 117.800 ;
        RECT 18.800 104.200 19.600 117.800 ;
        RECT 20.400 104.200 21.200 117.800 ;
        RECT 25.200 117.600 26.000 118.400 ;
        RECT 22.000 104.200 22.800 115.800 ;
        RECT 23.600 107.600 24.400 108.400 ;
        RECT 23.700 106.400 24.300 107.600 ;
        RECT 23.600 105.600 24.400 106.400 ;
        RECT 25.200 104.200 26.000 115.800 ;
        RECT 26.900 108.400 27.500 119.600 ;
        RECT 26.800 107.600 27.600 108.400 ;
        RECT 28.400 104.200 29.200 115.800 ;
        RECT 30.000 104.200 30.800 117.800 ;
        RECT 31.600 104.200 32.400 117.800 ;
        RECT 33.300 108.400 33.900 145.600 ;
        RECT 34.800 144.200 35.600 155.800 ;
        RECT 36.400 144.200 37.200 157.800 ;
        RECT 38.000 144.200 38.800 157.800 ;
        RECT 39.600 144.200 40.400 157.800 ;
        RECT 49.200 155.600 50.000 156.400 ;
        RECT 54.100 152.400 54.700 163.600 ;
        RECT 54.000 151.600 54.800 152.400 ;
        RECT 41.200 149.600 42.000 150.400 ;
        RECT 58.900 148.400 59.500 169.600 ;
        RECT 63.700 154.400 64.300 173.600 ;
        RECT 66.800 171.600 67.600 172.400 ;
        RECT 68.400 171.600 69.200 172.400 ;
        RECT 63.600 153.600 64.400 154.400 ;
        RECT 44.400 147.600 45.200 148.400 ;
        RECT 58.800 147.600 59.600 148.400 ;
        RECT 63.600 148.300 64.400 148.800 ;
        RECT 62.100 148.000 64.400 148.300 ;
        RECT 66.800 148.300 67.600 148.400 ;
        RECT 68.500 148.300 69.100 171.600 ;
        RECT 70.000 169.600 70.800 170.400 ;
        RECT 62.100 147.700 64.300 148.000 ;
        RECT 66.800 147.700 69.100 148.300 ;
        RECT 44.500 138.400 45.100 147.600 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 54.100 138.400 54.700 143.600 ;
        RECT 44.400 137.600 45.200 138.400 ;
        RECT 54.000 137.600 54.800 138.400 ;
        RECT 39.600 135.600 40.400 136.400 ;
        RECT 42.800 131.600 43.600 132.400 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 55.600 131.600 56.400 132.400 ;
        RECT 46.100 128.400 46.700 131.600 ;
        RECT 47.600 129.600 48.400 130.400 ;
        RECT 54.000 129.600 54.800 130.400 ;
        RECT 46.000 127.600 46.800 128.400 ;
        RECT 50.800 127.600 51.600 128.400 ;
        RECT 55.600 127.600 56.400 128.400 ;
        RECT 55.700 126.400 56.300 127.600 ;
        RECT 44.400 125.600 45.200 126.400 ;
        RECT 55.600 125.600 56.400 126.400 ;
        RECT 58.900 126.300 59.500 147.600 ;
        RECT 62.100 136.400 62.700 147.700 ;
        RECT 66.800 147.600 67.600 147.700 ;
        RECT 66.800 145.600 67.600 146.400 ;
        RECT 62.000 135.600 62.800 136.400 ;
        RECT 62.100 134.400 62.700 135.600 ;
        RECT 62.000 133.600 62.800 134.400 ;
        RECT 62.100 130.400 62.700 133.600 ;
        RECT 66.900 132.400 67.500 145.600 ;
        RECT 68.400 143.600 69.200 144.400 ;
        RECT 66.800 131.600 67.600 132.400 ;
        RECT 62.000 129.600 62.800 130.400 ;
        RECT 60.400 127.600 61.200 128.400 ;
        RECT 58.900 125.700 61.100 126.300 ;
        RECT 34.800 123.600 35.600 124.400 ;
        RECT 34.900 116.400 35.500 123.600 ;
        RECT 44.500 118.400 45.100 125.600 ;
        RECT 46.000 123.600 46.800 124.400 ;
        RECT 49.200 123.600 50.000 124.400 ;
        RECT 55.600 123.600 56.400 124.400 ;
        RECT 44.400 117.600 45.200 118.400 ;
        RECT 34.800 115.600 35.600 116.400 ;
        RECT 46.100 110.400 46.700 123.600 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 46.000 109.600 46.800 110.400 ;
        RECT 33.200 107.600 34.000 108.400 ;
        RECT 46.100 106.400 46.700 109.600 ;
        RECT 47.600 108.300 48.400 108.400 ;
        RECT 49.300 108.300 49.900 123.600 ;
        RECT 52.400 109.600 53.200 110.400 ;
        RECT 52.500 108.400 53.100 109.600 ;
        RECT 47.600 107.700 49.900 108.300 ;
        RECT 47.600 107.600 48.400 107.700 ;
        RECT 52.400 107.600 53.200 108.400 ;
        RECT 42.800 105.600 43.600 106.400 ;
        RECT 46.000 105.600 46.800 106.400 ;
        RECT 54.000 106.300 54.800 106.400 ;
        RECT 55.700 106.300 56.300 123.600 ;
        RECT 58.800 113.600 59.600 114.400 ;
        RECT 58.900 112.400 59.500 113.600 ;
        RECT 58.800 111.600 59.600 112.400 ;
        RECT 54.000 105.700 56.300 106.300 ;
        RECT 54.000 105.600 54.800 105.700 ;
        RECT 57.200 105.600 58.000 106.400 ;
        RECT 49.200 103.600 50.000 104.400 ;
        RECT 15.600 99.600 16.400 100.400 ;
        RECT 34.800 99.600 35.600 100.400 ;
        RECT 25.200 95.600 26.000 96.400 ;
        RECT 31.600 93.600 32.400 94.400 ;
        RECT 31.700 92.400 32.300 93.600 ;
        RECT 22.000 91.600 22.800 92.400 ;
        RECT 25.200 91.600 26.000 92.400 ;
        RECT 31.600 91.600 32.400 92.400 ;
        RECT 22.100 90.400 22.700 91.600 ;
        RECT 34.900 90.400 35.500 99.600 ;
        RECT 41.200 93.600 42.000 94.400 ;
        RECT 47.600 93.600 48.400 94.400 ;
        RECT 41.300 92.400 41.900 93.600 ;
        RECT 41.200 91.600 42.000 92.400 ;
        RECT 42.800 91.600 43.600 92.400 ;
        RECT 12.500 89.700 14.700 90.300 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 9.300 66.400 9.900 69.600 ;
        RECT 9.200 65.600 10.000 66.400 ;
        RECT 7.600 55.600 8.400 56.400 ;
        RECT 10.900 38.400 11.500 89.600 ;
        RECT 12.500 78.400 13.100 89.700 ;
        RECT 22.000 89.600 22.800 90.400 ;
        RECT 34.800 89.600 35.600 90.400 ;
        RECT 39.600 89.600 40.400 90.400 ;
        RECT 42.900 88.400 43.500 91.600 ;
        RECT 46.000 89.600 46.800 90.400 ;
        RECT 14.000 87.600 14.800 88.400 ;
        RECT 17.200 87.600 18.000 88.400 ;
        RECT 25.200 87.600 26.000 88.400 ;
        RECT 42.800 87.600 43.600 88.400 ;
        RECT 15.600 85.600 16.400 86.400 ;
        RECT 12.400 77.600 13.200 78.400 ;
        RECT 12.500 70.400 13.100 77.600 ;
        RECT 12.400 69.600 13.200 70.400 ;
        RECT 22.000 64.200 22.800 77.800 ;
        RECT 23.600 64.200 24.400 77.800 ;
        RECT 25.200 64.200 26.000 77.800 ;
        RECT 26.800 64.200 27.600 75.800 ;
        RECT 28.400 65.600 29.200 66.400 ;
        RECT 28.500 62.400 29.100 65.600 ;
        RECT 30.000 64.200 30.800 75.800 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 31.700 68.400 32.300 71.600 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 33.200 64.200 34.000 75.800 ;
        RECT 34.800 64.200 35.600 77.800 ;
        RECT 36.400 64.200 37.200 77.800 ;
        RECT 46.000 75.600 46.800 76.400 ;
        RECT 38.000 69.600 38.800 70.400 ;
        RECT 23.600 61.600 24.400 62.400 ;
        RECT 28.400 61.600 29.200 62.400 ;
        RECT 17.200 44.200 18.000 57.800 ;
        RECT 18.800 44.200 19.600 57.800 ;
        RECT 20.400 44.200 21.200 57.800 ;
        RECT 22.000 46.200 22.800 57.800 ;
        RECT 23.700 56.400 24.300 61.600 ;
        RECT 23.600 55.600 24.400 56.400 ;
        RECT 23.700 42.400 24.300 55.600 ;
        RECT 25.200 46.200 26.000 57.800 ;
        RECT 26.800 53.600 27.600 54.400 ;
        RECT 26.900 52.400 27.500 53.600 ;
        RECT 26.800 51.600 27.600 52.400 ;
        RECT 28.400 46.200 29.200 57.800 ;
        RECT 30.000 44.200 30.800 57.800 ;
        RECT 31.600 44.200 32.400 57.800 ;
        RECT 38.100 52.400 38.700 69.600 ;
        RECT 46.100 56.400 46.700 75.600 ;
        RECT 47.700 72.400 48.300 93.600 ;
        RECT 49.300 92.300 49.900 103.600 ;
        RECT 52.400 99.600 53.200 100.400 ;
        RECT 52.500 94.400 53.100 99.600 ;
        RECT 52.400 93.600 53.200 94.400 ;
        RECT 54.000 93.600 54.800 94.400 ;
        RECT 50.800 92.300 51.600 92.400 ;
        RECT 49.300 91.700 51.600 92.300 ;
        RECT 50.800 91.600 51.600 91.700 ;
        RECT 52.500 76.400 53.100 93.600 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 55.700 86.400 56.300 91.600 ;
        RECT 55.600 85.600 56.400 86.400 ;
        RECT 52.400 75.600 53.200 76.400 ;
        RECT 57.300 74.400 57.900 105.600 ;
        RECT 60.500 100.400 61.100 125.700 ;
        RECT 65.200 115.600 66.000 116.400 ;
        RECT 65.300 114.400 65.900 115.600 ;
        RECT 65.200 113.600 66.000 114.400 ;
        RECT 66.800 113.600 67.600 114.400 ;
        RECT 66.900 110.400 67.500 113.600 ;
        RECT 68.500 112.400 69.100 143.600 ;
        RECT 70.100 138.400 70.700 169.600 ;
        RECT 74.900 168.400 75.500 173.600 ;
        RECT 76.500 172.400 77.100 173.600 ;
        RECT 76.400 171.600 77.200 172.400 ;
        RECT 76.400 169.600 77.200 170.400 ;
        RECT 78.000 170.200 78.600 173.600 ;
        RECT 79.600 171.600 80.400 172.400 ;
        RECT 83.000 172.200 83.600 173.600 ;
        RECT 83.000 171.400 83.800 172.200 ;
        RECT 84.400 170.200 85.000 175.000 ;
        RECT 92.500 174.400 93.100 185.600 ;
        RECT 95.700 184.400 96.300 185.600 ;
        RECT 95.600 183.600 96.400 184.400 ;
        RECT 95.700 174.400 96.300 183.600 ;
        RECT 100.500 174.400 101.100 189.600 ;
        RECT 105.200 187.600 106.000 188.400 ;
        RECT 105.300 186.400 105.900 187.600 ;
        RECT 105.200 185.600 106.000 186.400 ;
        RECT 108.400 185.600 109.200 186.400 ;
        RECT 114.800 185.600 115.600 186.400 ;
        RECT 102.000 183.600 102.800 184.400 ;
        RECT 108.500 176.400 109.100 185.600 ;
        RECT 126.000 184.200 126.800 197.800 ;
        RECT 127.600 184.200 128.400 197.800 ;
        RECT 129.200 184.200 130.000 197.800 ;
        RECT 130.800 184.200 131.600 195.800 ;
        RECT 132.400 185.600 133.200 186.400 ;
        RECT 108.400 175.600 109.200 176.400 ;
        RECT 119.600 175.600 120.400 176.400 ;
        RECT 86.000 173.600 86.800 174.400 ;
        RECT 92.400 173.600 93.200 174.400 ;
        RECT 95.600 173.600 96.400 174.400 ;
        RECT 100.400 173.600 101.200 174.400 ;
        RECT 103.600 173.600 104.400 174.400 ;
        RECT 118.000 173.600 118.800 174.400 ;
        RECT 92.500 170.400 93.100 173.600 ;
        RECT 102.000 171.600 102.800 172.400 ;
        RECT 105.200 171.600 106.000 172.400 ;
        RECT 108.400 171.600 109.200 172.400 ;
        RECT 113.200 171.600 114.000 172.400 ;
        RECT 116.400 171.600 117.200 172.400 ;
        RECT 119.700 172.300 120.300 175.600 ;
        RECT 132.500 172.400 133.100 185.600 ;
        RECT 134.000 184.200 134.800 195.800 ;
        RECT 135.600 189.600 136.400 190.400 ;
        RECT 135.700 188.400 136.300 189.600 ;
        RECT 135.600 187.600 136.400 188.400 ;
        RECT 137.200 184.200 138.000 195.800 ;
        RECT 138.800 184.200 139.600 197.800 ;
        RECT 140.400 184.200 141.200 197.800 ;
        RECT 145.200 189.600 146.000 190.400 ;
        RECT 151.600 189.600 152.400 190.400 ;
        RECT 159.600 189.600 160.400 190.400 ;
        RECT 162.800 189.600 163.600 190.400 ;
        RECT 121.200 172.300 122.000 172.400 ;
        RECT 130.800 172.300 131.600 172.400 ;
        RECT 119.700 171.700 122.000 172.300 ;
        RECT 121.200 171.600 122.000 171.700 ;
        RECT 129.300 171.700 131.600 172.300 ;
        RECT 105.300 170.400 105.900 171.600 ;
        RECT 113.300 170.400 113.900 171.600 ;
        RECT 71.600 167.600 72.400 168.400 ;
        RECT 74.800 167.600 75.600 168.400 ;
        RECT 71.700 156.400 72.300 167.600 ;
        RECT 71.600 155.600 72.400 156.400 ;
        RECT 71.700 150.400 72.300 155.600 ;
        RECT 76.500 152.400 77.100 169.600 ;
        RECT 78.000 169.400 78.800 170.200 ;
        RECT 84.200 169.400 85.000 170.200 ;
        RECT 92.400 169.600 93.200 170.400 ;
        RECT 98.800 169.600 99.600 170.400 ;
        RECT 105.200 169.600 106.000 170.400 ;
        RECT 113.200 169.600 114.000 170.400 ;
        RECT 94.000 163.600 94.800 164.400 ;
        RECT 94.100 160.400 94.700 163.600 ;
        RECT 86.000 159.600 86.800 160.400 ;
        RECT 94.000 159.600 94.800 160.400 ;
        RECT 76.400 151.600 77.200 152.400 ;
        RECT 71.600 149.600 72.400 150.400 ;
        RECT 70.000 137.600 70.800 138.400 ;
        RECT 71.600 129.600 72.400 130.400 ;
        RECT 71.700 118.400 72.300 129.600 ;
        RECT 71.600 117.600 72.400 118.400 ;
        RECT 73.200 113.600 74.000 114.400 ;
        RECT 68.400 111.600 69.200 112.400 ;
        RECT 70.000 111.600 70.800 112.400 ;
        RECT 68.500 110.400 69.100 111.600 ;
        RECT 62.000 109.600 62.800 110.400 ;
        RECT 66.800 109.600 67.600 110.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 62.100 108.400 62.700 109.600 ;
        RECT 70.100 108.400 70.700 111.600 ;
        RECT 76.500 110.400 77.100 151.600 ;
        RECT 78.000 149.600 78.800 150.400 ;
        RECT 78.100 132.400 78.700 149.600 ;
        RECT 81.200 144.200 82.000 157.800 ;
        RECT 82.800 144.200 83.600 157.800 ;
        RECT 84.400 144.200 85.200 155.800 ;
        RECT 86.100 148.400 86.700 159.600 ;
        RECT 105.300 158.400 105.900 169.600 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 86.000 147.600 86.800 148.400 ;
        RECT 87.600 144.200 88.400 155.800 ;
        RECT 89.200 145.600 90.000 146.400 ;
        RECT 90.800 144.200 91.600 155.800 ;
        RECT 92.400 144.200 93.200 157.800 ;
        RECT 94.000 144.200 94.800 157.800 ;
        RECT 95.600 144.200 96.400 157.800 ;
        RECT 105.200 157.600 106.000 158.400 ;
        RECT 97.200 149.600 98.000 150.400 ;
        RECT 97.300 148.400 97.900 149.600 ;
        RECT 97.200 147.600 98.000 148.400 ;
        RECT 78.000 131.600 78.800 132.400 ;
        RECT 78.100 122.400 78.700 131.600 ;
        RECT 79.600 124.200 80.400 137.800 ;
        RECT 81.200 124.200 82.000 137.800 ;
        RECT 82.800 124.200 83.600 137.800 ;
        RECT 84.400 126.200 85.200 137.800 ;
        RECT 86.000 135.600 86.800 136.400 ;
        RECT 87.600 126.200 88.400 137.800 ;
        RECT 89.200 137.600 90.000 138.400 ;
        RECT 89.300 134.400 89.900 137.600 ;
        RECT 89.200 133.600 90.000 134.400 ;
        RECT 90.800 126.200 91.600 137.800 ;
        RECT 92.400 124.200 93.200 137.800 ;
        RECT 94.000 124.200 94.800 137.800 ;
        RECT 105.200 135.600 106.000 136.400 ;
        RECT 105.300 134.400 105.900 135.600 ;
        RECT 105.200 133.600 106.000 134.400 ;
        RECT 78.000 121.600 78.800 122.400 ;
        RECT 82.800 121.600 83.600 122.400 ;
        RECT 82.900 118.400 83.500 121.600 ;
        RECT 82.800 117.600 83.600 118.400 ;
        RECT 106.900 114.400 107.500 163.600 ;
        RECT 116.500 138.400 117.100 171.600 ;
        RECT 121.300 170.400 121.900 171.600 ;
        RECT 121.200 169.600 122.000 170.400 ;
        RECT 129.300 150.400 129.900 171.700 ;
        RECT 130.800 171.600 131.600 171.700 ;
        RECT 132.400 171.600 133.200 172.400 ;
        RECT 135.600 164.200 136.400 177.800 ;
        RECT 137.200 164.200 138.000 177.800 ;
        RECT 138.800 166.200 139.600 177.800 ;
        RECT 140.400 177.600 141.200 178.400 ;
        RECT 140.500 174.400 141.100 177.600 ;
        RECT 140.400 173.600 141.200 174.400 ;
        RECT 140.400 171.600 141.200 172.400 ;
        RECT 121.200 149.600 122.000 150.400 ;
        RECT 127.600 149.600 128.400 150.400 ;
        RECT 129.200 149.600 130.000 150.400 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 116.400 137.600 117.200 138.400 ;
        RECT 119.600 133.600 120.400 134.400 ;
        RECT 94.000 113.600 94.800 114.400 ;
        RECT 106.800 113.600 107.600 114.400 ;
        RECT 94.100 112.400 94.700 113.600 ;
        RECT 94.000 111.600 94.800 112.400 ;
        RECT 102.000 111.600 102.800 112.400 ;
        RECT 102.100 110.400 102.700 111.600 ;
        RECT 119.700 110.400 120.300 133.600 ;
        RECT 121.300 110.400 121.900 149.600 ;
        RECT 127.700 148.400 128.300 149.600 ;
        RECT 127.600 147.600 128.400 148.400 ;
        RECT 132.400 144.200 133.200 157.800 ;
        RECT 134.000 144.200 134.800 157.800 ;
        RECT 135.600 144.200 136.400 155.800 ;
        RECT 137.200 147.600 138.000 148.400 ;
        RECT 137.300 142.400 137.900 147.600 ;
        RECT 138.800 144.200 139.600 155.800 ;
        RECT 140.500 146.400 141.100 171.600 ;
        RECT 142.000 166.200 142.800 177.800 ;
        RECT 143.600 175.600 144.400 176.400 ;
        RECT 143.700 172.400 144.300 175.600 ;
        RECT 143.600 171.600 144.400 172.400 ;
        RECT 145.200 166.200 146.000 177.800 ;
        RECT 146.800 164.200 147.600 177.800 ;
        RECT 148.400 164.200 149.200 177.800 ;
        RECT 150.000 164.200 150.800 177.800 ;
        RECT 140.400 145.600 141.200 146.400 ;
        RECT 142.000 144.200 142.800 155.800 ;
        RECT 143.600 144.200 144.400 157.800 ;
        RECT 145.200 144.200 146.000 157.800 ;
        RECT 146.800 144.200 147.600 157.800 ;
        RECT 137.200 141.600 138.000 142.400 ;
        RECT 145.200 141.600 146.000 142.400 ;
        RECT 145.300 138.400 145.900 141.600 ;
        RECT 137.200 137.600 138.000 138.400 ;
        RECT 145.200 137.600 146.000 138.400 ;
        RECT 151.700 136.400 152.300 189.600 ;
        RECT 159.700 174.400 160.300 189.600 ;
        RECT 169.200 184.200 170.000 197.800 ;
        RECT 170.800 184.200 171.600 197.800 ;
        RECT 172.400 184.200 173.200 195.800 ;
        RECT 174.000 187.600 174.800 188.400 ;
        RECT 172.400 181.600 173.200 182.400 ;
        RECT 174.100 182.300 174.700 187.600 ;
        RECT 175.600 184.200 176.400 195.800 ;
        RECT 177.200 185.600 178.000 186.400 ;
        RECT 174.100 181.700 176.300 182.300 ;
        RECT 164.400 177.600 165.200 178.400 ;
        RECT 162.800 175.600 163.600 176.400 ;
        RECT 169.200 175.600 170.000 176.400 ;
        RECT 169.300 174.400 169.900 175.600 ;
        RECT 159.600 173.600 160.600 174.400 ;
        RECT 169.200 173.600 170.000 174.400 ;
        RECT 170.800 173.600 171.600 174.400 ;
        RECT 167.600 171.600 168.400 172.400 ;
        RECT 167.700 158.400 168.300 171.600 ;
        RECT 167.600 157.600 168.400 158.400 ;
        RECT 161.000 151.800 161.800 152.600 ;
        RECT 167.600 151.800 168.400 152.600 ;
        RECT 161.000 147.000 161.600 151.800 ;
        RECT 163.600 148.400 164.400 148.600 ;
        RECT 167.800 148.400 168.400 151.800 ;
        RECT 169.300 148.400 169.900 173.600 ;
        RECT 172.500 172.400 173.100 181.600 ;
        RECT 175.700 178.400 176.300 181.700 ;
        RECT 175.600 177.600 176.400 178.400 ;
        RECT 177.300 176.400 177.900 185.600 ;
        RECT 178.800 184.200 179.600 195.800 ;
        RECT 180.400 184.200 181.200 197.800 ;
        RECT 182.000 184.200 182.800 197.800 ;
        RECT 183.600 184.200 184.400 197.800 ;
        RECT 185.200 189.600 186.000 190.400 ;
        RECT 207.600 189.600 208.400 190.400 ;
        RECT 212.400 189.600 213.200 190.400 ;
        RECT 215.600 189.600 216.400 190.400 ;
        RECT 185.300 186.400 185.900 189.600 ;
        RECT 206.000 187.600 206.800 188.400 ;
        RECT 185.200 185.600 186.000 186.400 ;
        RECT 198.000 185.600 198.800 186.400 ;
        RECT 202.800 185.600 203.600 186.400 ;
        RECT 193.200 183.600 194.000 184.400 ;
        RECT 193.300 182.400 193.900 183.600 ;
        RECT 190.000 181.600 190.800 182.400 ;
        RECT 193.200 181.600 194.000 182.400 ;
        RECT 190.100 176.400 190.700 181.600 ;
        RECT 177.200 175.600 178.000 176.400 ;
        RECT 190.000 175.600 190.800 176.400 ;
        RECT 174.000 173.600 174.800 174.400 ;
        RECT 174.100 172.400 174.700 173.600 ;
        RECT 177.300 172.400 177.900 175.600 ;
        RECT 198.100 172.400 198.700 185.600 ;
        RECT 206.100 184.400 206.700 187.600 ;
        RECT 215.700 186.400 216.300 189.600 ;
        RECT 209.200 185.600 210.000 186.400 ;
        RECT 215.600 185.600 216.400 186.400 ;
        RECT 204.400 183.600 205.200 184.400 ;
        RECT 206.000 183.600 206.800 184.400 ;
        RECT 172.400 172.300 173.200 172.400 ;
        RECT 170.900 171.700 173.200 172.300 ;
        RECT 170.900 150.400 171.500 171.700 ;
        RECT 172.400 171.600 173.200 171.700 ;
        RECT 174.000 171.600 174.800 172.400 ;
        RECT 177.200 171.600 178.000 172.400 ;
        RECT 178.800 171.600 179.600 172.400 ;
        RECT 182.000 171.600 182.800 172.400 ;
        RECT 186.800 171.600 187.600 172.400 ;
        RECT 198.000 171.600 198.800 172.400 ;
        RECT 170.800 149.600 171.600 150.400 ;
        RECT 172.400 150.300 173.200 150.400 ;
        RECT 172.400 149.700 174.700 150.300 ;
        RECT 172.400 149.600 173.200 149.700 ;
        RECT 163.600 147.800 168.400 148.400 ;
        RECT 162.800 147.000 163.600 147.200 ;
        RECT 166.200 147.000 167.000 147.200 ;
        RECT 167.800 147.000 168.400 147.800 ;
        RECT 169.200 147.600 170.000 148.400 ;
        RECT 158.000 145.600 158.800 146.400 ;
        RECT 161.000 146.200 161.800 147.000 ;
        RECT 162.800 146.400 167.000 147.000 ;
        RECT 167.600 146.200 168.400 147.000 ;
        RECT 158.100 136.400 158.700 145.600 ;
        RECT 162.800 143.600 163.600 144.400 ;
        RECT 164.400 141.600 165.200 142.400 ;
        RECT 164.500 138.400 165.100 141.600 ;
        RECT 164.400 137.600 165.200 138.400 ;
        RECT 167.600 137.600 168.400 138.400 ;
        RECT 146.800 136.300 147.600 136.400 ;
        RECT 146.800 135.700 149.100 136.300 ;
        RECT 146.800 135.600 147.600 135.700 ;
        RECT 143.600 133.600 144.400 134.400 ;
        RECT 146.800 133.600 147.600 134.400 ;
        RECT 148.500 134.300 149.100 135.700 ;
        RECT 150.000 135.600 150.800 136.400 ;
        RECT 151.600 135.600 152.400 136.400 ;
        RECT 158.000 135.600 158.800 136.400 ;
        RECT 162.800 135.600 163.600 136.400 ;
        RECT 158.100 134.400 158.700 135.600 ;
        RECT 150.000 134.300 150.800 134.400 ;
        RECT 148.500 133.700 150.800 134.300 ;
        RECT 150.000 133.600 150.800 133.700 ;
        RECT 156.400 133.600 157.200 134.400 ;
        RECT 158.000 133.600 158.800 134.400 ;
        RECT 156.500 132.400 157.100 133.600 ;
        RECT 167.700 132.400 168.300 137.600 ;
        RECT 170.800 135.600 171.600 136.400 ;
        RECT 172.400 135.600 173.200 136.400 ;
        RECT 174.100 134.400 174.700 149.700 ;
        RECT 178.800 147.600 179.600 148.400 ;
        RECT 182.100 136.400 182.700 171.600 ;
        RECT 183.600 145.600 184.400 146.400 ;
        RECT 193.200 144.200 194.000 157.800 ;
        RECT 194.800 144.200 195.600 157.800 ;
        RECT 196.400 144.200 197.200 155.800 ;
        RECT 198.100 150.400 198.700 171.600 ;
        RECT 199.600 164.200 200.400 177.800 ;
        RECT 201.200 164.200 202.000 177.800 ;
        RECT 202.800 166.200 203.600 177.800 ;
        RECT 204.500 174.400 205.100 183.600 ;
        RECT 215.700 178.400 216.300 185.600 ;
        RECT 204.400 173.600 205.200 174.400 ;
        RECT 206.000 166.200 206.800 177.800 ;
        RECT 207.600 175.600 208.400 176.400 ;
        RECT 207.700 160.400 208.300 175.600 ;
        RECT 209.200 166.200 210.000 177.800 ;
        RECT 210.800 164.200 211.600 177.800 ;
        RECT 212.400 164.200 213.200 177.800 ;
        RECT 214.000 164.200 214.800 177.800 ;
        RECT 215.600 177.600 216.400 178.400 ;
        RECT 223.600 177.600 224.400 178.400 ;
        RECT 201.200 159.600 202.000 160.400 ;
        RECT 207.600 159.600 208.400 160.400 ;
        RECT 198.000 149.600 198.800 150.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 199.600 144.200 200.400 155.800 ;
        RECT 201.300 146.400 201.900 159.600 ;
        RECT 201.200 145.600 202.000 146.400 ;
        RECT 201.300 140.300 201.900 145.600 ;
        RECT 202.800 144.200 203.600 155.800 ;
        RECT 204.400 144.200 205.200 157.800 ;
        RECT 206.000 144.200 206.800 157.800 ;
        RECT 207.600 144.200 208.400 157.800 ;
        RECT 209.200 149.600 210.000 150.400 ;
        RECT 199.700 139.700 201.900 140.300 ;
        RECT 178.800 135.600 179.600 136.400 ;
        RECT 182.000 135.600 182.800 136.400 ;
        RECT 178.900 134.400 179.500 135.600 ;
        RECT 169.200 133.600 170.000 134.400 ;
        RECT 174.000 133.600 174.800 134.400 ;
        RECT 178.800 133.600 179.600 134.400 ;
        RECT 127.600 131.600 128.400 132.400 ;
        RECT 134.000 131.600 134.800 132.400 ;
        RECT 142.000 131.600 142.800 132.400 ;
        RECT 154.800 131.600 155.600 132.400 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 167.600 131.600 168.400 132.400 ;
        RECT 175.600 131.600 176.400 132.400 ;
        RECT 126.000 127.600 126.800 128.400 ;
        RECT 126.100 118.400 126.700 127.600 ;
        RECT 126.000 117.600 126.800 118.400 ;
        RECT 127.700 112.400 128.300 131.600 ;
        RECT 142.100 128.400 142.700 131.600 ;
        RECT 151.600 129.600 152.400 130.400 ;
        RECT 154.900 128.400 155.500 131.600 ;
        RECT 164.400 129.600 165.200 130.400 ;
        RECT 142.000 127.600 142.800 128.400 ;
        RECT 154.800 127.600 155.600 128.400 ;
        RECT 130.800 123.600 131.600 124.400 ;
        RECT 122.800 111.600 123.600 112.400 ;
        RECT 127.600 111.600 128.400 112.400 ;
        RECT 122.900 110.400 123.500 111.600 ;
        RECT 127.700 110.400 128.300 111.600 ;
        RECT 71.600 109.600 72.400 110.400 ;
        RECT 76.400 109.600 77.200 110.400 ;
        RECT 86.000 109.600 86.800 110.400 ;
        RECT 102.000 109.600 102.800 110.400 ;
        RECT 106.800 109.600 107.600 110.400 ;
        RECT 113.200 109.600 114.000 110.400 ;
        RECT 114.800 109.600 115.600 110.400 ;
        RECT 119.600 109.600 120.400 110.400 ;
        RECT 121.200 109.600 122.000 110.400 ;
        RECT 122.800 109.600 123.600 110.400 ;
        RECT 127.600 109.600 128.400 110.400 ;
        RECT 113.300 108.400 113.900 109.600 ;
        RECT 114.900 108.400 115.500 109.600 ;
        RECT 62.000 107.600 62.800 108.400 ;
        RECT 70.000 107.600 70.800 108.400 ;
        RECT 76.400 107.600 77.200 108.400 ;
        RECT 95.600 107.600 96.400 108.400 ;
        RECT 105.200 107.600 106.000 108.400 ;
        RECT 113.200 107.600 114.000 108.400 ;
        RECT 114.800 107.600 115.600 108.400 ;
        RECT 65.200 103.600 66.000 104.400 ;
        RECT 60.400 99.600 61.200 100.400 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 60.400 93.600 61.200 94.400 ;
        RECT 58.900 78.400 59.500 93.600 ;
        RECT 60.500 92.400 61.100 93.600 ;
        RECT 60.400 91.600 61.200 92.400 ;
        RECT 62.000 83.600 62.800 84.400 ;
        RECT 58.800 77.600 59.600 78.400 ;
        RECT 52.400 73.600 53.200 74.400 ;
        RECT 57.200 73.600 58.000 74.400 ;
        RECT 58.800 73.600 59.600 74.400 ;
        RECT 47.600 71.600 48.400 72.400 ;
        RECT 55.600 71.600 56.400 72.400 ;
        RECT 57.200 71.600 58.000 72.400 ;
        RECT 49.200 69.600 50.000 70.400 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 57.300 68.400 57.900 71.600 ;
        RECT 58.900 70.400 59.500 73.600 ;
        RECT 60.400 71.600 61.200 72.400 ;
        RECT 58.800 69.600 59.600 70.400 ;
        RECT 57.200 67.600 58.000 68.400 ;
        RECT 47.600 65.600 48.400 66.400 ;
        RECT 60.500 56.400 61.100 71.600 ;
        RECT 62.100 70.300 62.700 83.600 ;
        RECT 63.600 71.600 64.400 72.400 ;
        RECT 63.700 70.400 64.300 71.600 ;
        RECT 63.600 70.300 64.400 70.400 ;
        RECT 62.100 69.700 64.400 70.300 ;
        RECT 65.300 70.300 65.900 103.600 ;
        RECT 68.400 79.600 69.200 80.400 ;
        RECT 66.800 73.600 67.600 74.400 ;
        RECT 66.800 70.300 67.600 70.400 ;
        RECT 65.300 69.700 67.600 70.300 ;
        RECT 62.100 66.400 62.700 69.700 ;
        RECT 63.600 69.600 64.400 69.700 ;
        RECT 66.800 69.600 67.600 69.700 ;
        RECT 68.500 68.400 69.100 79.600 ;
        RECT 70.100 72.400 70.700 107.600 ;
        RECT 76.500 100.400 77.100 107.600 ;
        RECT 103.600 105.600 104.400 106.400 ;
        RECT 78.000 103.600 78.800 104.400 ;
        RECT 98.800 103.600 99.600 104.400 ;
        RECT 76.400 99.600 77.200 100.400 ;
        RECT 78.100 98.400 78.700 103.600 ;
        RECT 71.600 84.200 72.400 97.800 ;
        RECT 73.200 84.200 74.000 97.800 ;
        RECT 74.800 84.200 75.600 97.800 ;
        RECT 76.400 86.200 77.200 97.800 ;
        RECT 78.000 97.600 78.800 98.400 ;
        RECT 78.000 95.600 78.800 96.400 ;
        RECT 79.600 86.200 80.400 97.800 ;
        RECT 81.200 93.600 82.000 94.400 ;
        RECT 82.800 86.200 83.600 97.800 ;
        RECT 84.400 84.200 85.200 97.800 ;
        RECT 86.000 84.200 86.800 97.800 ;
        RECT 89.200 91.600 90.000 92.400 ;
        RECT 79.600 81.600 80.400 82.400 ;
        RECT 70.000 71.600 70.800 72.400 ;
        RECT 74.800 71.600 75.600 72.400 ;
        RECT 70.000 69.600 70.800 70.400 ;
        RECT 70.100 68.400 70.700 69.600 ;
        RECT 79.700 68.400 80.300 81.600 ;
        RECT 89.300 72.400 89.900 91.600 ;
        RECT 98.900 80.400 99.500 103.600 ;
        RECT 103.700 98.400 104.300 105.600 ;
        RECT 121.300 104.400 121.900 109.600 ;
        RECT 130.900 106.400 131.500 123.600 ;
        RECT 140.400 109.600 141.200 110.400 ;
        RECT 130.800 105.600 131.600 106.400 ;
        RECT 142.000 105.600 142.800 106.400 ;
        RECT 118.000 103.600 118.800 104.400 ;
        RECT 121.200 103.600 122.000 104.400 ;
        RECT 118.100 100.400 118.700 103.600 ;
        RECT 118.000 99.600 118.800 100.400 ;
        RECT 122.800 99.600 123.600 100.400 ;
        RECT 103.600 97.600 104.400 98.400 ;
        RECT 105.200 95.600 106.000 96.400 ;
        RECT 98.800 79.600 99.600 80.400 ;
        RECT 82.800 71.600 83.600 72.400 ;
        RECT 89.200 71.600 90.000 72.400 ;
        RECT 92.400 71.600 93.200 72.400 ;
        RECT 92.500 70.400 93.100 71.600 ;
        RECT 81.200 69.600 82.000 70.400 ;
        RECT 86.000 69.600 86.800 70.400 ;
        RECT 92.400 69.600 93.200 70.400 ;
        RECT 94.000 69.600 94.800 70.400 ;
        RECT 81.300 68.400 81.900 69.600 ;
        RECT 68.400 67.600 69.200 68.400 ;
        RECT 70.000 67.600 70.800 68.400 ;
        RECT 79.600 67.600 80.400 68.400 ;
        RECT 81.200 67.600 82.000 68.400 ;
        RECT 62.000 65.600 62.800 66.400 ;
        RECT 41.200 55.600 42.000 56.400 ;
        RECT 46.000 55.600 46.800 56.400 ;
        RECT 54.000 55.600 54.800 56.400 ;
        RECT 60.400 55.600 61.200 56.400 ;
        RECT 63.600 55.600 64.400 56.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 49.200 53.600 50.000 54.400 ;
        RECT 54.100 52.400 54.700 55.600 ;
        RECT 57.200 53.600 58.000 54.400 ;
        RECT 57.300 52.400 57.900 53.600 ;
        RECT 34.800 51.600 35.600 52.400 ;
        RECT 38.000 51.600 38.800 52.400 ;
        RECT 46.000 51.600 46.800 52.400 ;
        RECT 50.800 51.600 51.600 52.400 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 57.200 51.600 58.000 52.400 ;
        RECT 34.900 42.400 35.500 51.600 ;
        RECT 50.900 48.400 51.500 51.600 ;
        RECT 54.100 50.400 54.700 51.600 ;
        RECT 63.700 50.400 64.300 55.600 ;
        RECT 68.500 54.400 69.100 67.600 ;
        RECT 79.700 64.400 80.300 67.600 ;
        RECT 79.600 63.600 80.400 64.400 ;
        RECT 68.400 53.600 69.200 54.400 ;
        RECT 66.600 51.600 67.600 52.400 ;
        RECT 54.000 49.600 54.800 50.400 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 50.800 47.600 51.600 48.400 ;
        RECT 57.200 47.600 58.000 48.400 ;
        RECT 58.800 47.600 59.600 48.400 ;
        RECT 62.000 47.600 62.800 48.400 ;
        RECT 57.300 46.400 57.900 47.600 ;
        RECT 57.200 45.600 58.000 46.400 ;
        RECT 52.400 43.600 53.200 44.400 ;
        RECT 76.400 44.200 77.200 57.800 ;
        RECT 78.000 44.200 78.800 57.800 ;
        RECT 79.600 44.200 80.400 57.800 ;
        RECT 81.200 46.200 82.000 57.800 ;
        RECT 82.800 55.600 83.600 56.400 ;
        RECT 18.800 41.600 19.600 42.400 ;
        RECT 23.600 41.600 24.400 42.400 ;
        RECT 31.600 41.600 32.400 42.400 ;
        RECT 34.800 41.600 35.600 42.400 ;
        RECT 2.800 37.600 3.600 38.400 ;
        RECT 10.800 37.600 11.600 38.400 ;
        RECT 12.400 24.200 13.200 37.800 ;
        RECT 14.000 24.200 14.800 37.800 ;
        RECT 15.600 24.200 16.400 37.800 ;
        RECT 17.200 24.200 18.000 35.800 ;
        RECT 18.900 26.400 19.500 41.600 ;
        RECT 18.800 25.600 19.600 26.400 ;
        RECT 2.800 15.600 3.600 16.400 ;
        RECT 12.400 4.200 13.200 17.800 ;
        RECT 14.000 4.200 14.800 17.800 ;
        RECT 15.600 4.200 16.400 17.800 ;
        RECT 17.200 6.200 18.000 17.800 ;
        RECT 18.900 16.400 19.500 25.600 ;
        RECT 20.400 24.200 21.200 35.800 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 23.600 24.200 24.400 35.800 ;
        RECT 25.200 24.200 26.000 37.800 ;
        RECT 26.800 24.200 27.600 37.800 ;
        RECT 31.700 32.400 32.300 41.600 ;
        RECT 52.500 32.400 53.100 43.600 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 20.400 6.200 21.200 17.800 ;
        RECT 22.000 13.600 22.800 14.400 ;
        RECT 23.600 6.200 24.400 17.800 ;
        RECT 25.200 4.200 26.000 17.800 ;
        RECT 26.800 4.200 27.600 17.800 ;
        RECT 31.700 12.400 32.300 31.600 ;
        RECT 36.400 29.600 37.200 30.400 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 44.400 29.600 45.200 30.400 ;
        RECT 49.200 29.600 50.000 30.400 ;
        RECT 55.400 29.600 56.400 30.400 ;
        RECT 36.500 28.400 37.100 29.600 ;
        RECT 36.400 27.600 37.200 28.400 ;
        RECT 42.800 28.300 43.600 28.400 ;
        RECT 41.300 27.700 43.600 28.300 ;
        RECT 41.300 16.400 41.900 27.700 ;
        RECT 42.800 27.600 43.600 27.700 ;
        RECT 44.500 26.400 45.100 29.600 ;
        RECT 49.300 28.400 49.900 29.600 ;
        RECT 49.200 27.600 50.000 28.400 ;
        RECT 52.400 27.600 53.200 28.400 ;
        RECT 44.400 25.600 45.200 26.400 ;
        RECT 63.600 25.600 64.400 26.400 ;
        RECT 36.400 15.600 37.200 16.400 ;
        RECT 41.200 15.600 42.000 16.400 ;
        RECT 44.400 15.600 45.200 16.400 ;
        RECT 44.500 14.400 45.100 15.600 ;
        RECT 44.400 13.600 45.200 14.400 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 55.600 11.600 56.400 12.400 ;
        RECT 57.200 4.200 58.000 17.800 ;
        RECT 58.800 4.200 59.600 17.800 ;
        RECT 60.400 4.200 61.200 17.800 ;
        RECT 62.000 6.200 62.800 17.800 ;
        RECT 63.700 16.400 64.300 25.600 ;
        RECT 65.200 24.200 66.000 37.800 ;
        RECT 66.800 24.200 67.600 37.800 ;
        RECT 68.400 24.200 69.200 37.800 ;
        RECT 70.000 24.200 70.800 35.800 ;
        RECT 71.600 25.600 72.400 26.400 ;
        RECT 73.200 24.200 74.000 35.800 ;
        RECT 74.800 27.600 75.600 28.400 ;
        RECT 76.400 24.200 77.200 35.800 ;
        RECT 78.000 24.200 78.800 37.800 ;
        RECT 79.600 24.200 80.400 37.800 ;
        RECT 82.900 26.400 83.500 55.600 ;
        RECT 84.400 46.200 85.200 57.800 ;
        RECT 86.000 53.600 86.800 54.400 ;
        RECT 86.100 50.400 86.700 53.600 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 87.600 46.200 88.400 57.800 ;
        RECT 89.200 44.200 90.000 57.800 ;
        RECT 90.800 44.200 91.600 57.800 ;
        RECT 94.100 52.400 94.700 69.600 ;
        RECT 97.200 64.200 98.000 77.800 ;
        RECT 98.800 64.200 99.600 77.800 ;
        RECT 100.400 64.200 101.200 75.800 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 103.600 64.200 104.400 75.800 ;
        RECT 105.300 66.400 105.900 95.600 ;
        RECT 111.600 91.600 112.400 92.400 ;
        RECT 113.200 84.200 114.000 97.800 ;
        RECT 114.800 84.200 115.600 97.800 ;
        RECT 116.400 84.200 117.200 97.800 ;
        RECT 118.000 86.200 118.800 97.800 ;
        RECT 119.600 95.600 120.400 96.400 ;
        RECT 121.200 86.200 122.000 97.800 ;
        RECT 122.900 94.400 123.500 99.600 ;
        RECT 122.800 93.600 123.600 94.400 ;
        RECT 124.400 86.200 125.200 97.800 ;
        RECT 126.000 84.200 126.800 97.800 ;
        RECT 127.600 84.200 128.400 97.800 ;
        RECT 130.900 96.400 131.500 105.600 ;
        RECT 132.400 103.600 133.200 104.400 ;
        RECT 130.800 95.600 131.600 96.400 ;
        RECT 130.800 91.600 131.600 92.400 ;
        RECT 124.400 79.600 125.200 80.400 ;
        RECT 105.200 65.600 106.000 66.400 ;
        RECT 106.800 64.200 107.600 75.800 ;
        RECT 108.400 64.200 109.200 77.800 ;
        RECT 110.000 64.200 110.800 77.800 ;
        RECT 111.600 64.200 112.400 77.800 ;
        RECT 121.200 73.600 122.000 74.400 ;
        RECT 121.200 67.600 122.000 68.400 ;
        RECT 121.300 58.400 121.900 67.600 ;
        RECT 122.800 63.600 123.600 64.400 ;
        RECT 122.900 58.400 123.500 63.600 ;
        RECT 121.200 57.600 122.000 58.400 ;
        RECT 122.800 57.600 123.600 58.400 ;
        RECT 102.000 55.600 102.800 56.400 ;
        RECT 103.600 55.600 104.400 56.400 ;
        RECT 122.900 52.400 123.500 57.600 ;
        RECT 94.000 51.600 94.800 52.400 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 124.500 50.400 125.100 79.600 ;
        RECT 130.900 70.400 131.500 91.600 ;
        RECT 132.500 84.400 133.100 103.600 ;
        RECT 140.400 95.600 141.200 96.400 ;
        RECT 140.500 94.400 141.100 95.600 ;
        RECT 138.800 93.600 139.600 94.400 ;
        RECT 140.400 93.600 141.200 94.400 ;
        RECT 138.900 90.400 139.500 93.600 ;
        RECT 138.800 89.600 139.600 90.400 ;
        RECT 132.400 83.600 133.200 84.400 ;
        RECT 130.800 69.600 131.600 70.400 ;
        RECT 134.000 64.200 134.800 77.800 ;
        RECT 135.600 64.200 136.400 77.800 ;
        RECT 137.200 64.200 138.000 75.800 ;
        RECT 138.900 74.400 139.500 89.600 ;
        RECT 138.800 73.600 139.600 74.400 ;
        RECT 138.800 67.600 139.600 68.400 ;
        RECT 138.900 62.400 139.500 67.600 ;
        RECT 140.400 64.200 141.200 75.800 ;
        RECT 142.100 68.400 142.700 105.600 ;
        RECT 145.200 104.200 146.000 117.800 ;
        RECT 146.800 104.200 147.600 117.800 ;
        RECT 148.400 104.200 149.200 115.800 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 150.100 104.400 150.700 107.600 ;
        RECT 150.000 103.600 150.800 104.400 ;
        RECT 151.600 104.200 152.400 115.800 ;
        RECT 153.200 105.600 154.000 106.400 ;
        RECT 153.200 103.600 154.000 104.400 ;
        RECT 154.800 104.200 155.600 115.800 ;
        RECT 156.400 104.200 157.200 117.800 ;
        RECT 158.000 104.200 158.800 117.800 ;
        RECT 159.600 104.200 160.400 117.800 ;
        RECT 161.200 109.600 162.000 110.400 ;
        RECT 153.300 98.400 153.900 103.600 ;
        RECT 164.500 100.400 165.100 129.600 ;
        RECT 175.700 128.400 176.300 131.600 ;
        RECT 175.600 128.300 176.400 128.400 ;
        RECT 175.600 127.700 177.900 128.300 ;
        RECT 175.600 127.600 176.400 127.700 ;
        RECT 177.300 110.400 177.900 127.700 ;
        RECT 193.200 124.200 194.000 137.800 ;
        RECT 194.800 124.200 195.600 137.800 ;
        RECT 196.400 124.200 197.200 137.800 ;
        RECT 198.000 126.200 198.800 137.800 ;
        RECT 199.700 136.400 200.300 139.700 ;
        RECT 199.600 135.600 200.400 136.400 ;
        RECT 201.200 126.200 202.000 137.800 ;
        RECT 202.800 135.600 203.600 136.400 ;
        RECT 202.900 134.400 203.500 135.600 ;
        RECT 202.800 133.600 203.600 134.400 ;
        RECT 202.800 131.600 203.600 132.400 ;
        RECT 202.900 124.300 203.500 131.600 ;
        RECT 204.400 126.200 205.200 137.800 ;
        RECT 202.900 123.700 205.100 124.300 ;
        RECT 206.000 124.200 206.800 137.800 ;
        RECT 207.600 124.200 208.400 137.800 ;
        RECT 209.300 132.400 209.900 149.600 ;
        RECT 217.200 145.600 218.000 146.400 ;
        RECT 209.200 131.600 210.000 132.400 ;
        RECT 217.200 131.600 218.000 132.400 ;
        RECT 177.200 109.600 178.000 110.400 ;
        RECT 183.600 109.600 184.400 110.400 ;
        RECT 175.600 107.600 176.400 108.400 ;
        RECT 172.400 105.600 173.200 106.400 ;
        RECT 174.000 105.600 174.800 106.400 ;
        RECT 169.200 103.600 170.000 104.400 ;
        RECT 164.400 99.600 165.200 100.400 ;
        RECT 153.200 97.600 154.000 98.400 ;
        RECT 154.800 97.600 155.600 98.400 ;
        RECT 154.900 96.400 155.500 97.600 ;
        RECT 145.200 95.600 146.000 96.400 ;
        RECT 154.800 95.600 155.600 96.400 ;
        RECT 156.400 95.600 157.200 96.400 ;
        RECT 156.500 94.400 157.100 95.600 ;
        RECT 158.000 95.000 158.800 95.800 ;
        RECT 159.400 95.000 163.600 95.600 ;
        RECT 164.600 95.000 165.400 95.800 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 156.400 93.600 157.200 94.400 ;
        RECT 158.000 94.200 158.600 95.000 ;
        RECT 159.400 94.800 160.200 95.000 ;
        RECT 162.800 94.800 163.600 95.000 ;
        RECT 158.000 93.600 162.800 94.200 ;
        RECT 145.300 92.400 145.900 93.600 ;
        RECT 143.600 91.600 144.400 92.400 ;
        RECT 145.200 91.600 146.000 92.400 ;
        RECT 143.700 90.400 144.300 91.600 ;
        RECT 148.500 90.400 149.100 93.600 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 151.600 91.600 152.400 92.400 ;
        RECT 143.600 89.600 144.400 90.400 ;
        RECT 148.400 89.600 149.200 90.400 ;
        RECT 151.700 88.400 152.300 91.600 ;
        RECT 158.000 90.200 158.600 93.600 ;
        RECT 162.000 93.400 162.800 93.600 ;
        RECT 161.200 91.600 162.000 92.400 ;
        RECT 158.000 89.400 158.800 90.200 ;
        RECT 159.600 89.600 160.400 90.400 ;
        RECT 145.200 87.600 146.000 88.400 ;
        RECT 151.600 87.600 152.400 88.400 ;
        RECT 142.000 67.600 142.800 68.400 ;
        RECT 142.100 66.400 142.700 67.600 ;
        RECT 142.000 65.600 142.800 66.400 ;
        RECT 143.600 64.200 144.400 75.800 ;
        RECT 145.200 64.200 146.000 77.800 ;
        RECT 146.800 64.200 147.600 77.800 ;
        RECT 148.400 64.200 149.200 77.800 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 158.000 63.600 158.800 64.400 ;
        RECT 138.800 61.600 139.600 62.400 ;
        RECT 137.200 51.600 138.000 52.400 ;
        RECT 122.800 49.600 123.600 50.400 ;
        RECT 124.400 49.600 125.200 50.400 ;
        RECT 124.500 48.400 125.100 49.600 ;
        RECT 124.400 47.600 125.200 48.400 ;
        RECT 116.400 43.600 117.200 44.400 ;
        RECT 122.800 43.600 123.600 44.400 ;
        RECT 105.200 33.600 106.000 34.400 ;
        RECT 105.300 30.400 105.900 33.600 ;
        RECT 84.400 29.600 85.200 30.400 ;
        RECT 89.200 29.600 90.000 30.400 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 105.200 29.600 106.000 30.400 ;
        RECT 114.800 29.600 115.600 30.400 ;
        RECT 82.800 25.600 83.600 26.400 ;
        RECT 63.600 15.600 64.400 16.400 ;
        RECT 65.200 6.200 66.000 17.800 ;
        RECT 68.400 6.200 69.200 17.800 ;
        RECT 70.000 4.200 70.800 17.800 ;
        RECT 71.600 4.200 72.400 17.800 ;
        RECT 82.900 14.400 83.500 25.600 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 84.500 12.400 85.100 29.600 ;
        RECT 89.300 28.400 89.900 29.600 ;
        RECT 114.900 28.400 115.500 29.600 ;
        RECT 89.200 27.600 90.000 28.400 ;
        RECT 100.400 27.600 101.200 28.400 ;
        RECT 114.800 27.600 115.600 28.400 ;
        RECT 100.500 24.400 101.100 27.600 ;
        RECT 116.500 26.400 117.100 43.600 ;
        RECT 122.900 38.400 123.500 43.600 ;
        RECT 113.200 25.600 114.000 26.400 ;
        RECT 116.400 25.600 117.200 26.400 ;
        RECT 100.400 23.600 101.200 24.400 ;
        RECT 100.500 12.400 101.100 23.600 ;
        RECT 76.400 11.600 77.200 12.400 ;
        RECT 84.400 11.600 85.200 12.400 ;
        RECT 100.400 11.600 101.200 12.400 ;
        RECT 105.200 4.200 106.000 17.800 ;
        RECT 106.800 4.200 107.600 17.800 ;
        RECT 108.400 6.200 109.200 17.800 ;
        RECT 110.000 13.600 110.800 14.400 ;
        RECT 111.600 6.200 112.400 17.800 ;
        RECT 113.300 16.400 113.900 25.600 ;
        RECT 119.600 24.200 120.400 37.800 ;
        RECT 121.200 24.200 122.000 37.800 ;
        RECT 122.800 37.600 123.600 38.400 ;
        RECT 137.300 38.300 137.900 51.600 ;
        RECT 138.800 44.200 139.600 57.800 ;
        RECT 140.400 44.200 141.200 57.800 ;
        RECT 142.000 44.200 142.800 57.800 ;
        RECT 143.600 46.200 144.400 57.800 ;
        RECT 145.200 55.600 146.000 56.400 ;
        RECT 122.800 24.200 123.600 35.800 ;
        RECT 124.400 27.600 125.200 28.400 ;
        RECT 126.000 24.200 126.800 35.800 ;
        RECT 127.600 25.600 128.400 26.400 ;
        RECT 129.200 24.200 130.000 35.800 ;
        RECT 130.800 24.200 131.600 37.800 ;
        RECT 132.400 24.200 133.200 37.800 ;
        RECT 134.000 24.200 134.800 37.800 ;
        RECT 135.700 37.700 137.900 38.300 ;
        RECT 135.700 30.400 136.300 37.700 ;
        RECT 135.600 29.600 136.400 30.400 ;
        RECT 145.300 26.400 145.900 55.600 ;
        RECT 146.800 46.200 147.600 57.800 ;
        RECT 148.400 55.600 149.200 56.400 ;
        RECT 148.500 54.400 149.100 55.600 ;
        RECT 148.400 53.600 149.200 54.400 ;
        RECT 150.000 46.200 150.800 57.800 ;
        RECT 151.600 44.200 152.400 57.800 ;
        RECT 153.200 44.200 154.000 57.800 ;
        RECT 159.600 51.600 160.400 52.400 ;
        RECT 159.700 40.400 160.300 51.600 ;
        RECT 159.600 39.600 160.400 40.400 ;
        RECT 150.000 37.600 150.800 38.400 ;
        RECT 159.600 37.600 160.400 38.400 ;
        RECT 145.200 25.600 146.000 26.400 ;
        RECT 148.400 25.600 149.200 26.400 ;
        RECT 113.200 15.600 114.000 16.400 ;
        RECT 114.800 6.200 115.600 17.800 ;
        RECT 116.400 4.200 117.200 17.800 ;
        RECT 118.000 4.200 118.800 17.800 ;
        RECT 119.600 4.200 120.400 17.800 ;
        RECT 138.800 15.600 139.600 16.400 ;
        RECT 138.900 12.400 139.500 15.600 ;
        RECT 148.500 14.400 149.100 25.600 ;
        RECT 142.000 13.600 142.800 14.400 ;
        RECT 148.400 13.600 149.200 14.400 ;
        RECT 150.100 12.400 150.700 37.600 ;
        RECT 158.000 31.600 158.800 32.400 ;
        RECT 158.100 30.400 158.700 31.600 ;
        RECT 159.700 30.400 160.300 37.600 ;
        RECT 161.300 34.400 161.900 91.600 ;
        RECT 164.800 90.200 165.400 95.000 ;
        RECT 167.600 93.600 168.400 94.400 ;
        RECT 167.700 92.400 168.300 93.600 ;
        RECT 166.000 91.600 166.800 92.400 ;
        RECT 167.600 91.600 168.400 92.400 ;
        RECT 164.600 89.400 165.400 90.200 ;
        RECT 164.400 69.600 165.200 70.400 ;
        RECT 162.800 63.600 163.600 64.400 ;
        RECT 162.900 56.400 163.500 63.600 ;
        RECT 162.800 55.600 163.600 56.400 ;
        RECT 162.900 54.400 163.500 55.600 ;
        RECT 162.800 53.600 163.600 54.400 ;
        RECT 166.100 52.400 166.700 91.600 ;
        RECT 169.300 84.400 169.900 103.600 ;
        RECT 172.500 98.400 173.100 105.600 ;
        RECT 188.400 104.200 189.200 117.800 ;
        RECT 190.000 104.200 190.800 117.800 ;
        RECT 191.600 104.200 192.400 115.800 ;
        RECT 193.200 107.600 194.000 108.400 ;
        RECT 193.300 106.400 193.900 107.600 ;
        RECT 193.200 105.600 194.000 106.400 ;
        RECT 194.800 104.200 195.600 115.800 ;
        RECT 196.400 105.600 197.200 106.400 ;
        RECT 196.500 102.300 197.100 105.600 ;
        RECT 198.000 104.200 198.800 115.800 ;
        RECT 199.600 104.200 200.400 117.800 ;
        RECT 201.200 104.200 202.000 117.800 ;
        RECT 202.800 104.200 203.600 117.800 ;
        RECT 204.500 110.400 205.100 123.700 ;
        RECT 204.400 109.600 205.200 110.400 ;
        RECT 207.600 109.600 208.400 110.400 ;
        RECT 196.500 101.700 198.700 102.300 ;
        RECT 172.400 97.600 173.200 98.400 ;
        RECT 178.800 97.600 179.600 98.400 ;
        RECT 174.000 93.600 174.800 94.400 ;
        RECT 175.600 91.600 176.400 92.400 ;
        RECT 185.200 91.600 186.000 92.400 ;
        RECT 172.400 89.600 173.200 90.400 ;
        RECT 172.500 86.400 173.100 89.600 ;
        RECT 172.400 85.600 173.200 86.400 ;
        RECT 175.700 84.400 176.300 91.600 ;
        RECT 178.800 89.600 179.600 90.400 ;
        RECT 177.200 87.600 178.000 88.400 ;
        RECT 169.200 83.600 170.000 84.400 ;
        RECT 175.600 83.600 176.400 84.400 ;
        RECT 169.200 64.200 170.000 77.800 ;
        RECT 170.800 64.200 171.600 77.800 ;
        RECT 172.400 64.200 173.200 75.800 ;
        RECT 174.000 67.600 174.800 68.400 ;
        RECT 174.100 66.400 174.700 67.600 ;
        RECT 174.000 65.600 174.800 66.400 ;
        RECT 175.600 64.200 176.400 75.800 ;
        RECT 177.300 68.400 177.900 87.600 ;
        RECT 178.900 86.400 179.500 89.600 ;
        RECT 178.800 85.600 179.600 86.400 ;
        RECT 177.200 67.600 178.000 68.400 ;
        RECT 177.300 66.400 177.900 67.600 ;
        RECT 177.200 65.600 178.000 66.400 ;
        RECT 177.200 63.600 178.000 64.400 ;
        RECT 178.800 64.200 179.600 75.800 ;
        RECT 180.400 64.200 181.200 77.800 ;
        RECT 182.000 64.200 182.800 77.800 ;
        RECT 183.600 64.200 184.400 77.800 ;
        RECT 185.300 70.400 185.900 91.600 ;
        RECT 190.000 84.200 190.800 97.800 ;
        RECT 191.600 84.200 192.400 97.800 ;
        RECT 193.200 86.200 194.000 97.800 ;
        RECT 194.800 93.600 195.600 94.400 ;
        RECT 196.400 86.200 197.200 97.800 ;
        RECT 198.100 96.400 198.700 101.700 ;
        RECT 198.000 95.600 198.800 96.400 ;
        RECT 198.100 88.400 198.700 95.600 ;
        RECT 198.000 87.600 198.800 88.400 ;
        RECT 199.600 86.200 200.400 97.800 ;
        RECT 201.200 84.200 202.000 97.800 ;
        RECT 202.800 84.200 203.600 97.800 ;
        RECT 204.400 84.200 205.200 97.800 ;
        RECT 185.200 69.600 186.000 70.400 ;
        RECT 198.000 69.600 198.800 70.400 ;
        RECT 198.100 66.400 198.700 69.600 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 207.700 66.400 208.300 109.600 ;
        RECT 215.600 107.600 216.400 108.400 ;
        RECT 212.400 105.600 213.200 106.400 ;
        RECT 215.700 104.400 216.300 107.600 ;
        RECT 217.300 106.400 217.900 131.600 ;
        RECT 218.800 109.600 219.600 110.400 ;
        RECT 217.200 105.600 218.000 106.400 ;
        RECT 215.600 103.600 216.400 104.400 ;
        RECT 215.700 92.400 216.300 103.600 ;
        RECT 220.400 95.600 221.200 96.400 ;
        RECT 220.500 94.400 221.100 95.600 ;
        RECT 220.400 93.600 221.200 94.400 ;
        RECT 215.600 91.600 216.400 92.400 ;
        RECT 217.200 91.600 218.000 92.400 ;
        RECT 218.800 91.600 219.600 92.400 ;
        RECT 223.600 91.600 224.400 92.400 ;
        RECT 217.300 84.400 217.900 91.600 ;
        RECT 210.800 83.600 211.600 84.400 ;
        RECT 214.000 83.600 214.800 84.400 ;
        RECT 217.200 83.600 218.000 84.400 ;
        RECT 210.900 70.400 211.500 83.600 ;
        RECT 210.800 69.600 211.600 70.400 ;
        RECT 212.400 69.600 213.200 70.400 ;
        RECT 210.900 68.400 211.500 69.600 ;
        RECT 214.100 68.400 214.700 83.600 ;
        RECT 217.200 69.600 218.000 70.400 ;
        RECT 217.300 68.400 217.900 69.600 ;
        RECT 210.800 67.600 211.600 68.400 ;
        RECT 214.000 67.600 214.800 68.400 ;
        RECT 217.200 67.600 218.000 68.400 ;
        RECT 220.400 67.600 221.200 68.400 ;
        RECT 198.000 65.600 198.800 66.400 ;
        RECT 204.400 65.600 205.200 66.400 ;
        RECT 207.600 65.600 208.400 66.400 ;
        RECT 207.700 64.400 208.300 65.600 ;
        RECT 207.600 63.600 208.400 64.400 ;
        RECT 169.200 61.600 170.000 62.400 ;
        RECT 169.300 58.400 169.900 61.600 ;
        RECT 169.200 57.600 170.000 58.400 ;
        RECT 172.400 57.600 173.200 58.400 ;
        RECT 169.200 53.600 170.000 54.400 ;
        RECT 162.800 51.600 163.600 52.400 ;
        RECT 166.000 51.600 166.800 52.400 ;
        RECT 161.200 33.600 162.000 34.400 ;
        RECT 158.000 29.600 158.800 30.400 ;
        RECT 159.600 29.600 160.400 30.400 ;
        RECT 151.600 27.600 152.400 28.400 ;
        RECT 162.900 26.300 163.500 51.600 ;
        RECT 166.100 50.400 166.700 51.600 ;
        RECT 166.000 49.600 166.800 50.400 ;
        RECT 164.400 43.600 165.200 44.400 ;
        RECT 164.500 32.400 165.100 43.600 ;
        RECT 164.400 31.600 165.200 32.400 ;
        RECT 167.600 27.600 168.400 28.400 ;
        RECT 162.900 25.700 165.100 26.300 ;
        RECT 158.000 23.600 158.800 24.400 ;
        RECT 162.800 23.600 163.600 24.400 ;
        RECT 158.100 16.400 158.700 23.600 ;
        RECT 158.000 15.600 158.800 16.400 ;
        RECT 151.600 13.600 152.400 14.400 ;
        RECT 151.700 12.400 152.300 13.600 ;
        RECT 158.100 12.400 158.700 15.600 ;
        RECT 164.500 12.400 165.100 25.700 ;
        RECT 167.700 18.400 168.300 27.600 ;
        RECT 169.300 20.300 169.900 53.600 ;
        RECT 172.500 50.400 173.100 57.600 ;
        RECT 177.300 54.400 177.900 63.600 ;
        RECT 183.600 57.600 184.400 58.400 ;
        RECT 177.200 53.600 178.000 54.400 ;
        RECT 178.800 53.600 179.600 54.400 ;
        RECT 175.600 51.600 176.400 52.400 ;
        RECT 183.700 50.400 184.300 57.600 ;
        RECT 193.200 51.600 194.000 52.400 ;
        RECT 172.400 49.600 173.200 50.400 ;
        RECT 183.600 49.600 184.400 50.400 ;
        RECT 180.400 43.600 181.200 44.400 ;
        RECT 170.800 39.600 171.600 40.400 ;
        RECT 170.900 30.400 171.500 39.600 ;
        RECT 180.500 38.400 181.100 43.600 ;
        RECT 170.800 29.600 171.600 30.400 ;
        RECT 172.400 24.200 173.200 37.800 ;
        RECT 174.000 24.200 174.800 37.800 ;
        RECT 175.600 24.200 176.400 37.800 ;
        RECT 180.400 37.600 181.200 38.400 ;
        RECT 177.200 24.200 178.000 35.800 ;
        RECT 178.800 25.600 179.600 26.400 ;
        RECT 178.800 23.600 179.600 24.400 ;
        RECT 180.400 24.200 181.200 35.800 ;
        RECT 182.000 27.600 182.800 28.400 ;
        RECT 183.600 24.200 184.400 35.800 ;
        RECT 185.200 24.200 186.000 37.800 ;
        RECT 186.800 24.200 187.600 37.800 ;
        RECT 193.300 30.400 193.900 51.600 ;
        RECT 194.800 44.200 195.600 57.800 ;
        RECT 196.400 44.200 197.200 57.800 ;
        RECT 198.000 46.200 198.800 57.800 ;
        RECT 199.600 53.600 200.400 54.400 ;
        RECT 201.200 46.200 202.000 57.800 ;
        RECT 202.800 55.600 203.600 56.400 ;
        RECT 202.900 40.400 203.500 55.600 ;
        RECT 204.400 46.200 205.200 57.800 ;
        RECT 206.000 44.200 206.800 57.800 ;
        RECT 207.600 44.200 208.400 57.800 ;
        RECT 209.200 44.200 210.000 57.800 ;
        RECT 199.600 39.600 200.400 40.400 ;
        RECT 202.800 39.600 203.600 40.400 ;
        RECT 198.000 37.600 198.800 38.400 ;
        RECT 190.000 29.600 190.800 30.400 ;
        RECT 193.200 29.600 194.000 30.400 ;
        RECT 169.300 19.700 171.500 20.300 ;
        RECT 167.600 17.600 168.400 18.400 ;
        RECT 169.200 15.600 170.000 16.400 ;
        RECT 166.000 13.600 166.800 14.400 ;
        RECT 170.900 12.400 171.500 19.700 ;
        RECT 175.600 15.600 176.400 16.400 ;
        RECT 175.600 13.600 176.400 14.400 ;
        RECT 132.400 11.600 133.200 12.400 ;
        RECT 138.800 11.600 139.600 12.400 ;
        RECT 148.400 11.600 149.200 12.400 ;
        RECT 150.000 11.600 150.800 12.400 ;
        RECT 151.600 11.600 152.400 12.400 ;
        RECT 156.400 11.600 157.200 12.400 ;
        RECT 158.000 11.600 158.800 12.400 ;
        RECT 164.400 11.600 165.200 12.400 ;
        RECT 170.800 11.600 171.600 12.400 ;
        RECT 175.700 10.400 176.300 13.600 ;
        RECT 178.900 12.400 179.500 23.600 ;
        RECT 180.400 17.600 181.200 18.400 ;
        RECT 180.500 14.400 181.100 17.600 ;
        RECT 180.400 13.600 181.200 14.400 ;
        RECT 190.100 12.400 190.700 29.600 ;
        RECT 196.400 27.600 197.200 28.400 ;
        RECT 178.800 11.600 179.600 12.400 ;
        RECT 190.000 11.600 190.800 12.400 ;
        RECT 175.600 9.600 176.400 10.400 ;
        RECT 191.600 4.200 192.400 17.800 ;
        RECT 193.200 4.200 194.000 17.800 ;
        RECT 194.800 6.200 195.600 17.800 ;
        RECT 196.500 14.400 197.100 27.600 ;
        RECT 198.100 26.400 198.700 37.600 ;
        RECT 199.700 26.400 200.300 39.600 ;
        RECT 210.900 30.400 211.500 67.600 ;
        RECT 220.500 56.400 221.100 67.600 ;
        RECT 223.700 58.400 224.300 91.600 ;
        RECT 223.600 57.600 224.400 58.400 ;
        RECT 220.400 55.600 221.200 56.400 ;
        RECT 212.400 53.600 213.200 54.400 ;
        RECT 212.500 38.400 213.100 53.600 ;
        RECT 218.800 43.600 219.600 44.400 ;
        RECT 212.400 37.600 213.200 38.400 ;
        RECT 218.900 30.400 219.500 43.600 ;
        RECT 202.800 29.600 203.600 30.400 ;
        RECT 207.600 29.600 208.400 30.400 ;
        RECT 209.200 29.600 210.000 30.400 ;
        RECT 210.800 29.600 211.600 30.400 ;
        RECT 218.800 29.600 219.600 30.400 ;
        RECT 198.000 25.600 198.800 26.400 ;
        RECT 199.600 25.600 200.400 26.400 ;
        RECT 196.400 13.600 197.200 14.400 ;
        RECT 198.000 6.200 198.800 17.800 ;
        RECT 199.700 16.400 200.300 25.600 ;
        RECT 202.900 24.400 203.500 29.600 ;
        RECT 209.300 28.400 209.900 29.600 ;
        RECT 206.000 27.600 206.800 28.400 ;
        RECT 209.200 27.600 210.000 28.400 ;
        RECT 218.900 26.400 219.500 29.600 ;
        RECT 206.000 25.600 206.800 26.400 ;
        RECT 218.800 25.600 219.600 26.400 ;
        RECT 202.800 23.600 203.600 24.400 ;
        RECT 206.100 20.400 206.700 25.600 ;
        RECT 206.000 19.600 206.800 20.400 ;
        RECT 215.600 19.600 216.400 20.400 ;
        RECT 215.700 18.400 216.300 19.600 ;
        RECT 199.600 15.600 200.400 16.400 ;
        RECT 201.200 6.200 202.000 17.800 ;
        RECT 202.800 4.200 203.600 17.800 ;
        RECT 204.400 4.200 205.200 17.800 ;
        RECT 206.000 4.200 206.800 17.800 ;
        RECT 215.600 17.600 216.400 18.400 ;
      LAYER via2 ;
        RECT 159.600 173.600 160.400 174.400 ;
        RECT 66.800 51.600 67.600 52.400 ;
        RECT 55.600 29.600 56.400 30.400 ;
      LAYER metal3 ;
        RECT 9.200 194.300 10.000 194.400 ;
        RECT 28.400 194.300 29.200 194.400 ;
        RECT 9.200 193.700 29.200 194.300 ;
        RECT 9.200 193.600 10.000 193.700 ;
        RECT 28.400 193.600 29.200 193.700 ;
        RECT 7.600 190.300 8.400 190.400 ;
        RECT 12.400 190.300 13.200 190.400 ;
        RECT 7.600 189.700 13.200 190.300 ;
        RECT 7.600 189.600 8.400 189.700 ;
        RECT 12.400 189.600 13.200 189.700 ;
        RECT 25.200 190.300 26.000 190.400 ;
        RECT 30.000 190.300 30.800 190.400 ;
        RECT 36.400 190.300 37.200 190.400 ;
        RECT 25.200 189.700 37.200 190.300 ;
        RECT 25.200 189.600 26.000 189.700 ;
        RECT 30.000 189.600 30.800 189.700 ;
        RECT 36.400 189.600 37.200 189.700 ;
        RECT 82.800 190.300 83.600 190.400 ;
        RECT 135.600 190.300 136.400 190.400 ;
        RECT 82.800 189.700 136.400 190.300 ;
        RECT 82.800 189.600 83.600 189.700 ;
        RECT 135.600 189.600 136.400 189.700 ;
        RECT 145.200 190.300 146.000 190.400 ;
        RECT 162.800 190.300 163.600 190.400 ;
        RECT 145.200 189.700 163.600 190.300 ;
        RECT 145.200 189.600 146.000 189.700 ;
        RECT 162.800 189.600 163.600 189.700 ;
        RECT 207.600 190.300 208.400 190.400 ;
        RECT 212.400 190.300 213.200 190.400 ;
        RECT 207.600 189.700 213.200 190.300 ;
        RECT 207.600 189.600 208.400 189.700 ;
        RECT 212.400 189.600 213.200 189.700 ;
        RECT 15.600 188.300 16.400 188.400 ;
        RECT 20.400 188.300 21.200 188.400 ;
        RECT 25.200 188.300 26.000 188.400 ;
        RECT 15.600 187.700 26.000 188.300 ;
        RECT 15.600 187.600 16.400 187.700 ;
        RECT 20.400 187.600 21.200 187.700 ;
        RECT 25.200 187.600 26.000 187.700 ;
        RECT 74.800 188.300 75.600 188.400 ;
        RECT 81.200 188.300 82.000 188.400 ;
        RECT 74.800 187.700 82.000 188.300 ;
        RECT 74.800 187.600 75.600 187.700 ;
        RECT 81.200 187.600 82.000 187.700 ;
        RECT 92.400 188.300 93.200 188.400 ;
        RECT 95.600 188.300 96.400 188.400 ;
        RECT 92.400 187.700 96.400 188.300 ;
        RECT 92.400 187.600 93.200 187.700 ;
        RECT 95.600 187.600 96.400 187.700 ;
        RECT 23.600 186.300 24.400 186.400 ;
        RECT 33.200 186.300 34.000 186.400 ;
        RECT 50.800 186.300 51.600 186.400 ;
        RECT 60.400 186.300 61.200 186.400 ;
        RECT 23.600 185.700 61.200 186.300 ;
        RECT 23.600 185.600 24.400 185.700 ;
        RECT 33.200 185.600 34.000 185.700 ;
        RECT 50.800 185.600 51.600 185.700 ;
        RECT 60.400 185.600 61.200 185.700 ;
        RECT 74.800 186.300 75.600 186.400 ;
        RECT 79.600 186.300 80.400 186.400 ;
        RECT 74.800 185.700 80.400 186.300 ;
        RECT 74.800 185.600 75.600 185.700 ;
        RECT 79.600 185.600 80.400 185.700 ;
        RECT 87.600 186.300 88.400 186.400 ;
        RECT 92.400 186.300 93.200 186.400 ;
        RECT 87.600 185.700 93.200 186.300 ;
        RECT 87.600 185.600 88.400 185.700 ;
        RECT 92.400 185.600 93.200 185.700 ;
        RECT 97.200 186.300 98.000 186.400 ;
        RECT 105.200 186.300 106.000 186.400 ;
        RECT 97.200 185.700 106.000 186.300 ;
        RECT 97.200 185.600 98.000 185.700 ;
        RECT 105.200 185.600 106.000 185.700 ;
        RECT 108.400 186.300 109.200 186.400 ;
        RECT 114.800 186.300 115.600 186.400 ;
        RECT 108.400 185.700 115.600 186.300 ;
        RECT 108.400 185.600 109.200 185.700 ;
        RECT 114.800 185.600 115.600 185.700 ;
        RECT 185.200 186.300 186.000 186.400 ;
        RECT 198.000 186.300 198.800 186.400 ;
        RECT 185.200 185.700 198.800 186.300 ;
        RECT 185.200 185.600 186.000 185.700 ;
        RECT 198.000 185.600 198.800 185.700 ;
        RECT 202.800 186.300 203.600 186.400 ;
        RECT 209.200 186.300 210.000 186.400 ;
        RECT 202.800 185.700 210.000 186.300 ;
        RECT 202.800 185.600 203.600 185.700 ;
        RECT 209.200 185.600 210.000 185.700 ;
        RECT 58.800 184.300 59.600 184.400 ;
        RECT 87.700 184.300 88.300 185.600 ;
        RECT 58.800 183.700 88.300 184.300 ;
        RECT 95.600 184.300 96.400 184.400 ;
        RECT 102.000 184.300 102.800 184.400 ;
        RECT 206.000 184.300 206.800 184.400 ;
        RECT 95.600 183.700 102.800 184.300 ;
        RECT 58.800 183.600 59.600 183.700 ;
        RECT 95.600 183.600 96.400 183.700 ;
        RECT 102.000 183.600 102.800 183.700 ;
        RECT 177.300 183.700 206.800 184.300 ;
        RECT 172.400 182.300 173.200 182.400 ;
        RECT 177.300 182.300 177.900 183.700 ;
        RECT 206.000 183.600 206.800 183.700 ;
        RECT 172.400 181.700 177.900 182.300 ;
        RECT 190.000 182.300 190.800 182.400 ;
        RECT 193.200 182.300 194.000 182.400 ;
        RECT 190.000 181.700 194.000 182.300 ;
        RECT 172.400 181.600 173.200 181.700 ;
        RECT 190.000 181.600 190.800 181.700 ;
        RECT 193.200 181.600 194.000 181.700 ;
        RECT 2.800 180.300 3.600 180.400 ;
        RECT 38.000 180.300 38.800 180.400 ;
        RECT 54.000 180.300 54.800 180.400 ;
        RECT 2.800 179.700 54.800 180.300 ;
        RECT 2.800 179.600 3.600 179.700 ;
        RECT 38.000 179.600 38.800 179.700 ;
        RECT 54.000 179.600 54.800 179.700 ;
        RECT 58.800 180.300 59.600 180.400 ;
        RECT 71.600 180.300 72.400 180.400 ;
        RECT 58.800 179.700 72.400 180.300 ;
        RECT 58.800 179.600 59.600 179.700 ;
        RECT 71.600 179.600 72.400 179.700 ;
        RECT 7.600 178.300 8.400 178.400 ;
        RECT 22.000 178.300 22.800 178.400 ;
        RECT 7.600 177.700 22.800 178.300 ;
        RECT 7.600 177.600 8.400 177.700 ;
        RECT 22.000 177.600 22.800 177.700 ;
        RECT 57.200 178.300 58.000 178.400 ;
        RECT 62.000 178.300 62.800 178.400 ;
        RECT 57.200 177.700 62.800 178.300 ;
        RECT 57.200 177.600 58.000 177.700 ;
        RECT 62.000 177.600 62.800 177.700 ;
        RECT 140.400 178.300 141.200 178.400 ;
        RECT 164.400 178.300 165.200 178.400 ;
        RECT 140.400 177.700 165.200 178.300 ;
        RECT 140.400 177.600 141.200 177.700 ;
        RECT 164.400 177.600 165.200 177.700 ;
        RECT 215.600 178.300 216.400 178.400 ;
        RECT 223.600 178.300 224.400 178.400 ;
        RECT 215.600 177.700 224.400 178.300 ;
        RECT 215.600 177.600 216.400 177.700 ;
        RECT 223.600 177.600 224.400 177.700 ;
        RECT 14.000 176.300 14.800 176.400 ;
        RECT 22.000 176.300 22.800 176.400 ;
        RECT 14.000 175.700 22.800 176.300 ;
        RECT 14.000 175.600 14.800 175.700 ;
        RECT 22.000 175.600 22.800 175.700 ;
        RECT 52.400 176.300 53.200 176.400 ;
        RECT 58.800 176.300 59.600 176.400 ;
        RECT 52.400 175.700 59.600 176.300 ;
        RECT 52.400 175.600 53.200 175.700 ;
        RECT 58.800 175.600 59.600 175.700 ;
        RECT 161.200 176.300 162.000 176.400 ;
        RECT 162.800 176.300 163.600 176.400 ;
        RECT 161.200 175.700 163.600 176.300 ;
        RECT 161.200 175.600 162.000 175.700 ;
        RECT 162.800 175.600 163.600 175.700 ;
        RECT 177.200 176.300 178.000 176.400 ;
        RECT 207.600 176.300 208.400 176.400 ;
        RECT 177.200 175.700 208.400 176.300 ;
        RECT 177.200 175.600 178.000 175.700 ;
        RECT 207.600 175.600 208.400 175.700 ;
        RECT 14.000 174.300 14.800 174.400 ;
        RECT 34.800 174.300 35.600 174.400 ;
        RECT 14.000 173.700 35.600 174.300 ;
        RECT 14.000 173.600 14.800 173.700 ;
        RECT 34.800 173.600 35.600 173.700 ;
        RECT 55.600 174.300 56.400 174.400 ;
        RECT 68.400 174.300 69.200 174.400 ;
        RECT 73.200 174.300 74.000 174.400 ;
        RECT 55.600 173.700 74.000 174.300 ;
        RECT 55.600 173.600 56.400 173.700 ;
        RECT 68.400 173.600 69.200 173.700 ;
        RECT 73.200 173.600 74.000 173.700 ;
        RECT 76.400 174.300 77.200 174.400 ;
        RECT 86.000 174.300 86.800 174.400 ;
        RECT 95.600 174.300 96.400 174.400 ;
        RECT 76.400 173.700 96.400 174.300 ;
        RECT 76.400 173.600 77.200 173.700 ;
        RECT 86.000 173.600 86.800 173.700 ;
        RECT 95.600 173.600 96.400 173.700 ;
        RECT 100.400 174.300 101.200 174.400 ;
        RECT 103.600 174.300 104.400 174.400 ;
        RECT 118.000 174.300 118.800 174.400 ;
        RECT 100.400 173.700 118.800 174.300 ;
        RECT 100.400 173.600 101.200 173.700 ;
        RECT 103.600 173.600 104.400 173.700 ;
        RECT 118.000 173.600 118.800 173.700 ;
        RECT 159.600 174.300 160.400 174.400 ;
        RECT 169.200 174.300 170.000 174.400 ;
        RECT 159.600 173.700 170.000 174.300 ;
        RECT 159.600 173.600 160.400 173.700 ;
        RECT 169.200 173.600 170.000 173.700 ;
        RECT 170.800 174.300 171.600 174.400 ;
        RECT 174.000 174.300 174.800 174.400 ;
        RECT 170.800 173.700 174.800 174.300 ;
        RECT 170.800 173.600 171.600 173.700 ;
        RECT 174.000 173.600 174.800 173.700 ;
        RECT 44.400 172.300 45.200 172.400 ;
        RECT 52.400 172.300 53.200 172.400 ;
        RECT 44.400 171.700 53.200 172.300 ;
        RECT 44.400 171.600 45.200 171.700 ;
        RECT 52.400 171.600 53.200 171.700 ;
        RECT 66.800 172.300 67.600 172.400 ;
        RECT 79.600 172.300 80.400 172.400 ;
        RECT 66.800 171.700 80.400 172.300 ;
        RECT 66.800 171.600 67.600 171.700 ;
        RECT 79.600 171.600 80.400 171.700 ;
        RECT 102.000 172.300 102.800 172.400 ;
        RECT 108.400 172.300 109.200 172.400 ;
        RECT 102.000 171.700 109.200 172.300 ;
        RECT 102.000 171.600 102.800 171.700 ;
        RECT 108.400 171.600 109.200 171.700 ;
        RECT 132.400 172.300 133.200 172.400 ;
        RECT 140.400 172.300 141.200 172.400 ;
        RECT 143.600 172.300 144.400 172.400 ;
        RECT 177.200 172.300 178.000 172.400 ;
        RECT 132.400 171.700 178.000 172.300 ;
        RECT 132.400 171.600 133.200 171.700 ;
        RECT 140.400 171.600 141.200 171.700 ;
        RECT 143.600 171.600 144.400 171.700 ;
        RECT 177.200 171.600 178.000 171.700 ;
        RECT 178.800 172.300 179.600 172.400 ;
        RECT 186.800 172.300 187.600 172.400 ;
        RECT 178.800 171.700 187.600 172.300 ;
        RECT 178.800 171.600 179.600 171.700 ;
        RECT 186.800 171.600 187.600 171.700 ;
        RECT 6.000 170.300 6.800 170.400 ;
        RECT 55.600 170.300 56.400 170.400 ;
        RECT 58.800 170.300 59.600 170.400 ;
        RECT 6.000 169.700 59.600 170.300 ;
        RECT 6.000 169.600 6.800 169.700 ;
        RECT 55.600 169.600 56.400 169.700 ;
        RECT 58.800 169.600 59.600 169.700 ;
        RECT 76.400 170.300 77.200 170.400 ;
        RECT 92.400 170.300 93.200 170.400 ;
        RECT 98.800 170.300 99.600 170.400 ;
        RECT 76.400 169.700 99.600 170.300 ;
        RECT 76.400 169.600 77.200 169.700 ;
        RECT 92.400 169.600 93.200 169.700 ;
        RECT 98.800 169.600 99.600 169.700 ;
        RECT 105.200 170.300 106.000 170.400 ;
        RECT 113.200 170.300 114.000 170.400 ;
        RECT 121.200 170.300 122.000 170.400 ;
        RECT 105.200 169.700 122.000 170.300 ;
        RECT 105.200 169.600 106.000 169.700 ;
        RECT 113.200 169.600 114.000 169.700 ;
        RECT 121.200 169.600 122.000 169.700 ;
        RECT 71.600 168.300 72.400 168.400 ;
        RECT 74.800 168.300 75.600 168.400 ;
        RECT 71.600 167.700 75.600 168.300 ;
        RECT 71.600 167.600 72.400 167.700 ;
        RECT 74.800 167.600 75.600 167.700 ;
        RECT 86.000 160.300 86.800 160.400 ;
        RECT 94.000 160.300 94.800 160.400 ;
        RECT 86.000 159.700 94.800 160.300 ;
        RECT 86.000 159.600 86.800 159.700 ;
        RECT 94.000 159.600 94.800 159.700 ;
        RECT 201.200 160.300 202.000 160.400 ;
        RECT 207.600 160.300 208.400 160.400 ;
        RECT 201.200 159.700 208.400 160.300 ;
        RECT 201.200 159.600 202.000 159.700 ;
        RECT 207.600 159.600 208.400 159.700 ;
        RECT 167.600 157.600 168.400 158.400 ;
        RECT 49.200 156.300 50.000 156.400 ;
        RECT 71.600 156.300 72.400 156.400 ;
        RECT 49.200 155.700 72.400 156.300 ;
        RECT 49.200 155.600 50.000 155.700 ;
        RECT 71.600 155.600 72.400 155.700 ;
        RECT 30.000 154.300 30.800 154.400 ;
        RECT 63.600 154.300 64.400 154.400 ;
        RECT 30.000 153.700 64.400 154.300 ;
        RECT 30.000 153.600 30.800 153.700 ;
        RECT 63.600 153.600 64.400 153.700 ;
        RECT 15.600 152.300 16.400 152.400 ;
        RECT 76.400 152.300 77.200 152.400 ;
        RECT 15.600 151.700 77.200 152.300 ;
        RECT 15.600 151.600 16.400 151.700 ;
        RECT 76.400 151.600 77.200 151.700 ;
        RECT 6.000 150.300 6.800 150.400 ;
        RECT 7.600 150.300 8.400 150.400 ;
        RECT 6.000 149.700 8.400 150.300 ;
        RECT 6.000 149.600 6.800 149.700 ;
        RECT 7.600 149.600 8.400 149.700 ;
        RECT 36.400 150.300 37.200 150.400 ;
        RECT 41.200 150.300 42.000 150.400 ;
        RECT 78.000 150.300 78.800 150.400 ;
        RECT 36.400 149.700 78.800 150.300 ;
        RECT 36.400 149.600 37.200 149.700 ;
        RECT 41.200 149.600 42.000 149.700 ;
        RECT 78.000 149.600 78.800 149.700 ;
        RECT 121.200 150.300 122.000 150.400 ;
        RECT 170.800 150.300 171.600 150.400 ;
        RECT 121.200 149.700 171.600 150.300 ;
        RECT 121.200 149.600 122.000 149.700 ;
        RECT 170.800 149.600 171.600 149.700 ;
        RECT 12.400 148.300 13.200 148.400 ;
        RECT 44.400 148.300 45.200 148.400 ;
        RECT 12.400 147.700 45.200 148.300 ;
        RECT 12.400 147.600 13.200 147.700 ;
        RECT 44.400 147.600 45.200 147.700 ;
        RECT 97.200 148.300 98.000 148.400 ;
        RECT 127.600 148.300 128.400 148.400 ;
        RECT 97.200 147.700 128.400 148.300 ;
        RECT 97.200 147.600 98.000 147.700 ;
        RECT 127.600 147.600 128.400 147.700 ;
        RECT 178.800 148.300 179.600 148.400 ;
        RECT 198.000 148.300 198.800 148.400 ;
        RECT 178.800 147.700 198.800 148.300 ;
        RECT 178.800 147.600 179.600 147.700 ;
        RECT 198.000 147.600 198.800 147.700 ;
        RECT 33.200 146.300 34.000 146.400 ;
        RECT 71.600 146.300 72.400 146.400 ;
        RECT 89.200 146.300 90.000 146.400 ;
        RECT 90.800 146.300 91.600 146.400 ;
        RECT 33.200 145.700 91.600 146.300 ;
        RECT 33.200 145.600 34.000 145.700 ;
        RECT 71.600 145.600 72.400 145.700 ;
        RECT 89.200 145.600 90.000 145.700 ;
        RECT 90.800 145.600 91.600 145.700 ;
        RECT 119.600 146.300 120.400 146.400 ;
        RECT 140.400 146.300 141.200 146.400 ;
        RECT 119.600 145.700 141.200 146.300 ;
        RECT 119.600 145.600 120.400 145.700 ;
        RECT 140.400 145.600 141.200 145.700 ;
        RECT 183.600 146.300 184.400 146.400 ;
        RECT 217.200 146.300 218.000 146.400 ;
        RECT 183.600 145.700 218.000 146.300 ;
        RECT 183.600 145.600 184.400 145.700 ;
        RECT 217.200 145.600 218.000 145.700 ;
        RECT 154.800 144.300 155.600 144.400 ;
        RECT 162.800 144.300 163.600 144.400 ;
        RECT 154.800 143.700 163.600 144.300 ;
        RECT 154.800 143.600 155.600 143.700 ;
        RECT 162.800 143.600 163.600 143.700 ;
        RECT 137.200 142.300 138.000 142.400 ;
        RECT 145.200 142.300 146.000 142.400 ;
        RECT 137.200 141.700 146.000 142.300 ;
        RECT 137.200 141.600 138.000 141.700 ;
        RECT 145.200 141.600 146.000 141.700 ;
        RECT 161.200 142.300 162.000 142.400 ;
        RECT 164.400 142.300 165.200 142.400 ;
        RECT 161.200 141.700 165.200 142.300 ;
        RECT 161.200 141.600 162.000 141.700 ;
        RECT 164.400 141.600 165.200 141.700 ;
        RECT 54.000 138.300 54.800 138.400 ;
        RECT 89.200 138.300 90.000 138.400 ;
        RECT 54.000 137.700 90.000 138.300 ;
        RECT 54.000 137.600 54.800 137.700 ;
        RECT 89.200 137.600 90.000 137.700 ;
        RECT 116.400 138.300 117.200 138.400 ;
        RECT 137.200 138.300 138.000 138.400 ;
        RECT 167.600 138.300 168.400 138.400 ;
        RECT 116.400 137.700 168.400 138.300 ;
        RECT 116.400 137.600 117.200 137.700 ;
        RECT 137.200 137.600 138.000 137.700 ;
        RECT 167.600 137.600 168.400 137.700 ;
        RECT 6.000 136.300 6.800 136.400 ;
        RECT 9.200 136.300 10.000 136.400 ;
        RECT 14.000 136.300 14.800 136.400 ;
        RECT 30.000 136.300 30.800 136.400 ;
        RECT 39.600 136.300 40.400 136.400 ;
        RECT 6.000 135.700 40.400 136.300 ;
        RECT 6.000 135.600 6.800 135.700 ;
        RECT 9.200 135.600 10.000 135.700 ;
        RECT 14.000 135.600 14.800 135.700 ;
        RECT 30.000 135.600 30.800 135.700 ;
        RECT 39.600 135.600 40.400 135.700 ;
        RECT 86.000 136.300 86.800 136.400 ;
        RECT 90.800 136.300 91.600 136.400 ;
        RECT 105.200 136.300 106.000 136.400 ;
        RECT 86.000 135.700 106.000 136.300 ;
        RECT 86.000 135.600 86.800 135.700 ;
        RECT 90.800 135.600 91.600 135.700 ;
        RECT 105.200 135.600 106.000 135.700 ;
        RECT 150.000 136.300 150.800 136.400 ;
        RECT 151.600 136.300 152.400 136.400 ;
        RECT 158.000 136.300 158.800 136.400 ;
        RECT 150.000 135.700 158.800 136.300 ;
        RECT 150.000 135.600 150.800 135.700 ;
        RECT 151.600 135.600 152.400 135.700 ;
        RECT 158.000 135.600 158.800 135.700 ;
        RECT 162.800 136.300 163.600 136.400 ;
        RECT 170.800 136.300 171.600 136.400 ;
        RECT 162.800 135.700 171.600 136.300 ;
        RECT 162.800 135.600 163.600 135.700 ;
        RECT 170.800 135.600 171.600 135.700 ;
        RECT 172.400 136.300 173.200 136.400 ;
        RECT 202.800 136.300 203.600 136.400 ;
        RECT 172.400 135.700 203.600 136.300 ;
        RECT 172.400 135.600 173.200 135.700 ;
        RECT 202.800 135.600 203.600 135.700 ;
        RECT 4.400 134.300 5.200 134.400 ;
        RECT 7.600 134.300 8.400 134.400 ;
        RECT 62.000 134.300 62.800 134.400 ;
        RECT 4.400 133.700 62.800 134.300 ;
        RECT 4.400 133.600 5.200 133.700 ;
        RECT 7.600 133.600 8.400 133.700 ;
        RECT 62.000 133.600 62.800 133.700 ;
        RECT 119.600 134.300 120.400 134.400 ;
        RECT 143.600 134.300 144.400 134.400 ;
        RECT 146.800 134.300 147.600 134.400 ;
        RECT 119.600 133.700 147.600 134.300 ;
        RECT 119.600 133.600 120.400 133.700 ;
        RECT 143.600 133.600 144.400 133.700 ;
        RECT 146.800 133.600 147.600 133.700 ;
        RECT 169.200 134.300 170.000 134.400 ;
        RECT 178.800 134.300 179.600 134.400 ;
        RECT 169.200 133.700 179.600 134.300 ;
        RECT 169.200 133.600 170.000 133.700 ;
        RECT 178.800 133.600 179.600 133.700 ;
        RECT 2.800 132.300 3.600 132.400 ;
        RECT 17.200 132.300 18.000 132.400 ;
        RECT 2.800 131.700 18.000 132.300 ;
        RECT 2.800 131.600 3.600 131.700 ;
        RECT 17.200 131.600 18.000 131.700 ;
        RECT 42.800 132.300 43.600 132.400 ;
        RECT 49.200 132.300 50.000 132.400 ;
        RECT 55.600 132.300 56.400 132.400 ;
        RECT 42.800 131.700 56.400 132.300 ;
        RECT 42.800 131.600 43.600 131.700 ;
        RECT 49.200 131.600 50.000 131.700 ;
        RECT 55.600 131.600 56.400 131.700 ;
        RECT 127.600 132.300 128.400 132.400 ;
        RECT 134.000 132.300 134.800 132.400 ;
        RECT 127.600 131.700 134.800 132.300 ;
        RECT 127.600 131.600 128.400 131.700 ;
        RECT 134.000 131.600 134.800 131.700 ;
        RECT 156.400 132.300 157.200 132.400 ;
        RECT 158.000 132.300 158.800 132.400 ;
        RECT 217.200 132.300 218.000 132.400 ;
        RECT 156.400 131.700 218.000 132.300 ;
        RECT 156.400 131.600 157.200 131.700 ;
        RECT 158.000 131.600 158.800 131.700 ;
        RECT 217.200 131.600 218.000 131.700 ;
        RECT 12.400 130.300 13.200 130.400 ;
        RECT 47.600 130.300 48.400 130.400 ;
        RECT 54.000 130.300 54.800 130.400 ;
        RECT 12.400 129.700 54.800 130.300 ;
        RECT 12.400 129.600 13.200 129.700 ;
        RECT 47.600 129.600 48.400 129.700 ;
        RECT 54.000 129.600 54.800 129.700 ;
        RECT 62.000 130.300 62.800 130.400 ;
        RECT 71.600 130.300 72.400 130.400 ;
        RECT 62.000 129.700 72.400 130.300 ;
        RECT 62.000 129.600 62.800 129.700 ;
        RECT 71.600 129.600 72.400 129.700 ;
        RECT 151.600 130.300 152.400 130.400 ;
        RECT 164.400 130.300 165.200 130.400 ;
        RECT 151.600 129.700 165.200 130.300 ;
        RECT 151.600 129.600 152.400 129.700 ;
        RECT 164.400 129.600 165.200 129.700 ;
        RECT 15.600 128.300 16.400 128.400 ;
        RECT 23.600 128.300 24.400 128.400 ;
        RECT 15.600 127.700 24.400 128.300 ;
        RECT 15.600 127.600 16.400 127.700 ;
        RECT 23.600 127.600 24.400 127.700 ;
        RECT 46.000 128.300 46.800 128.400 ;
        RECT 50.800 128.300 51.600 128.400 ;
        RECT 60.400 128.300 61.200 128.400 ;
        RECT 46.000 127.700 61.200 128.300 ;
        RECT 46.000 127.600 46.800 127.700 ;
        RECT 50.800 127.600 51.600 127.700 ;
        RECT 60.400 127.600 61.200 127.700 ;
        RECT 126.000 128.300 126.800 128.400 ;
        RECT 142.000 128.300 142.800 128.400 ;
        RECT 154.800 128.300 155.600 128.400 ;
        RECT 175.600 128.300 176.400 128.400 ;
        RECT 126.000 127.700 176.400 128.300 ;
        RECT 126.000 127.600 126.800 127.700 ;
        RECT 142.000 127.600 142.800 127.700 ;
        RECT 154.800 127.600 155.600 127.700 ;
        RECT 175.600 127.600 176.400 127.700 ;
        RECT 44.400 126.300 45.200 126.400 ;
        RECT 55.600 126.300 56.400 126.400 ;
        RECT 44.400 125.700 56.400 126.300 ;
        RECT 44.400 125.600 45.200 125.700 ;
        RECT 55.600 125.600 56.400 125.700 ;
        RECT 30.000 124.300 30.800 124.400 ;
        RECT 46.000 124.300 46.800 124.400 ;
        RECT 30.000 123.700 46.800 124.300 ;
        RECT 30.000 123.600 30.800 123.700 ;
        RECT 46.000 123.600 46.800 123.700 ;
        RECT 78.000 122.300 78.800 122.400 ;
        RECT 82.800 122.300 83.600 122.400 ;
        RECT 78.000 121.700 83.600 122.300 ;
        RECT 78.000 121.600 78.800 121.700 ;
        RECT 82.800 121.600 83.600 121.700 ;
        RECT 18.800 120.300 19.600 120.400 ;
        RECT 26.800 120.300 27.600 120.400 ;
        RECT 18.800 119.700 27.600 120.300 ;
        RECT 18.800 119.600 19.600 119.700 ;
        RECT 26.800 119.600 27.600 119.700 ;
        RECT 1.200 118.300 2.000 118.400 ;
        RECT 7.600 118.300 8.400 118.400 ;
        RECT 25.200 118.300 26.000 118.400 ;
        RECT 1.200 117.700 26.000 118.300 ;
        RECT 1.200 117.600 2.000 117.700 ;
        RECT 7.600 117.600 8.400 117.700 ;
        RECT 25.200 117.600 26.000 117.700 ;
        RECT 34.800 116.300 35.600 116.400 ;
        RECT 65.200 116.300 66.000 116.400 ;
        RECT 34.800 115.700 66.000 116.300 ;
        RECT 34.800 115.600 35.600 115.700 ;
        RECT 65.200 115.600 66.000 115.700 ;
        RECT 58.800 114.300 59.600 114.400 ;
        RECT 73.200 114.300 74.000 114.400 ;
        RECT 106.800 114.300 107.600 114.400 ;
        RECT 58.800 113.700 107.600 114.300 ;
        RECT 58.800 113.600 59.600 113.700 ;
        RECT 73.200 113.600 74.000 113.700 ;
        RECT 106.800 113.600 107.600 113.700 ;
        RECT 94.000 112.300 94.800 112.400 ;
        RECT 102.000 112.300 102.800 112.400 ;
        RECT 122.800 112.300 123.600 112.400 ;
        RECT 127.600 112.300 128.400 112.400 ;
        RECT 94.000 111.700 128.400 112.300 ;
        RECT 94.000 111.600 94.800 111.700 ;
        RECT 102.000 111.600 102.800 111.700 ;
        RECT 122.800 111.600 123.600 111.700 ;
        RECT 127.600 111.600 128.400 111.700 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 62.000 110.300 62.800 110.400 ;
        RECT 68.400 110.300 69.200 110.400 ;
        RECT 71.600 110.300 72.400 110.400 ;
        RECT 62.000 109.700 72.400 110.300 ;
        RECT 62.000 109.600 62.800 109.700 ;
        RECT 68.400 109.600 69.200 109.700 ;
        RECT 71.600 109.600 72.400 109.700 ;
        RECT 86.000 110.300 86.800 110.400 ;
        RECT 90.800 110.300 91.600 110.400 ;
        RECT 106.800 110.300 107.600 110.400 ;
        RECT 86.000 109.700 107.600 110.300 ;
        RECT 86.000 109.600 86.800 109.700 ;
        RECT 90.800 109.600 91.600 109.700 ;
        RECT 106.800 109.600 107.600 109.700 ;
        RECT 113.200 110.300 114.000 110.400 ;
        RECT 140.400 110.300 141.200 110.400 ;
        RECT 113.200 109.700 141.200 110.300 ;
        RECT 113.200 109.600 114.000 109.700 ;
        RECT 140.400 109.600 141.200 109.700 ;
        RECT 161.200 110.300 162.000 110.400 ;
        RECT 183.600 110.300 184.400 110.400 ;
        RECT 161.200 109.700 184.400 110.300 ;
        RECT 161.200 109.600 162.000 109.700 ;
        RECT 183.600 109.600 184.400 109.700 ;
        RECT 207.600 110.300 208.400 110.400 ;
        RECT 218.800 110.300 219.600 110.400 ;
        RECT 207.600 109.700 219.600 110.300 ;
        RECT 207.600 109.600 208.400 109.700 ;
        RECT 218.800 109.600 219.600 109.700 ;
        RECT 23.600 108.300 24.400 108.400 ;
        RECT 33.200 108.300 34.000 108.400 ;
        RECT 23.600 107.700 34.000 108.300 ;
        RECT 23.600 107.600 24.400 107.700 ;
        RECT 33.200 107.600 34.000 107.700 ;
        RECT 52.400 108.300 53.200 108.400 ;
        RECT 70.000 108.300 70.800 108.400 ;
        RECT 95.600 108.300 96.400 108.400 ;
        RECT 52.400 107.700 96.400 108.300 ;
        RECT 52.400 107.600 53.200 107.700 ;
        RECT 70.000 107.600 70.800 107.700 ;
        RECT 95.600 107.600 96.400 107.700 ;
        RECT 105.200 108.300 106.000 108.400 ;
        RECT 114.800 108.300 115.600 108.400 ;
        RECT 105.200 107.700 115.600 108.300 ;
        RECT 105.200 107.600 106.000 107.700 ;
        RECT 114.800 107.600 115.600 107.700 ;
        RECT 175.600 108.300 176.400 108.400 ;
        RECT 215.600 108.300 216.400 108.400 ;
        RECT 175.600 107.700 216.400 108.300 ;
        RECT 175.600 107.600 176.400 107.700 ;
        RECT 215.600 107.600 216.400 107.700 ;
        RECT 14.000 106.300 14.800 106.400 ;
        RECT 42.800 106.300 43.600 106.400 ;
        RECT 46.000 106.300 46.800 106.400 ;
        RECT 14.000 105.700 46.800 106.300 ;
        RECT 14.000 105.600 14.800 105.700 ;
        RECT 42.800 105.600 43.600 105.700 ;
        RECT 46.000 105.600 46.800 105.700 ;
        RECT 130.800 106.300 131.600 106.400 ;
        RECT 142.000 106.300 142.800 106.400 ;
        RECT 153.200 106.300 154.000 106.400 ;
        RECT 130.800 105.700 154.000 106.300 ;
        RECT 130.800 105.600 131.600 105.700 ;
        RECT 142.000 105.600 142.800 105.700 ;
        RECT 153.200 105.600 154.000 105.700 ;
        RECT 174.000 106.300 174.800 106.400 ;
        RECT 193.200 106.300 194.000 106.400 ;
        RECT 174.000 105.700 194.000 106.300 ;
        RECT 174.000 105.600 174.800 105.700 ;
        RECT 193.200 105.600 194.000 105.700 ;
        RECT 212.400 106.300 213.200 106.400 ;
        RECT 217.200 106.300 218.000 106.400 ;
        RECT 212.400 105.700 218.000 106.300 ;
        RECT 212.400 105.600 213.200 105.700 ;
        RECT 217.200 105.600 218.000 105.700 ;
        RECT 121.200 104.300 122.000 104.400 ;
        RECT 122.800 104.300 123.600 104.400 ;
        RECT 121.200 103.700 123.600 104.300 ;
        RECT 121.200 103.600 122.000 103.700 ;
        RECT 122.800 103.600 123.600 103.700 ;
        RECT 150.000 104.300 150.800 104.400 ;
        RECT 153.200 104.300 154.000 104.400 ;
        RECT 150.000 103.700 154.000 104.300 ;
        RECT 150.000 103.600 150.800 103.700 ;
        RECT 153.200 103.600 154.000 103.700 ;
        RECT 10.800 100.300 11.600 100.400 ;
        RECT 15.600 100.300 16.400 100.400 ;
        RECT 34.800 100.300 35.600 100.400 ;
        RECT 52.400 100.300 53.200 100.400 ;
        RECT 60.400 100.300 61.200 100.400 ;
        RECT 76.400 100.300 77.200 100.400 ;
        RECT 10.800 99.700 77.200 100.300 ;
        RECT 10.800 99.600 11.600 99.700 ;
        RECT 15.600 99.600 16.400 99.700 ;
        RECT 34.800 99.600 35.600 99.700 ;
        RECT 52.400 99.600 53.200 99.700 ;
        RECT 60.400 99.600 61.200 99.700 ;
        RECT 76.400 99.600 77.200 99.700 ;
        RECT 118.000 100.300 118.800 100.400 ;
        RECT 122.800 100.300 123.600 100.400 ;
        RECT 118.000 99.700 123.600 100.300 ;
        RECT 118.000 99.600 118.800 99.700 ;
        RECT 122.800 99.600 123.600 99.700 ;
        RECT 164.400 100.300 165.200 100.400 ;
        RECT 170.800 100.300 171.600 100.400 ;
        RECT 164.400 99.700 171.600 100.300 ;
        RECT 164.400 99.600 165.200 99.700 ;
        RECT 170.800 99.600 171.600 99.700 ;
        RECT 78.000 97.600 78.800 98.400 ;
        RECT 154.800 98.300 155.600 98.400 ;
        RECT 178.800 98.300 179.600 98.400 ;
        RECT 154.800 97.700 179.600 98.300 ;
        RECT 154.800 97.600 155.600 97.700 ;
        RECT 178.800 97.600 179.600 97.700 ;
        RECT 7.600 96.300 8.400 96.400 ;
        RECT 20.400 96.300 21.200 96.400 ;
        RECT 25.200 96.300 26.000 96.400 ;
        RECT 7.600 95.700 26.000 96.300 ;
        RECT 7.600 95.600 8.400 95.700 ;
        RECT 20.400 95.600 21.200 95.700 ;
        RECT 25.200 95.600 26.000 95.700 ;
        RECT 71.600 96.300 72.400 96.400 ;
        RECT 78.000 96.300 78.800 96.400 ;
        RECT 71.600 95.700 78.800 96.300 ;
        RECT 71.600 95.600 72.400 95.700 ;
        RECT 78.000 95.600 78.800 95.700 ;
        RECT 105.200 96.300 106.000 96.400 ;
        RECT 119.600 96.300 120.400 96.400 ;
        RECT 130.800 96.300 131.600 96.400 ;
        RECT 105.200 95.700 131.600 96.300 ;
        RECT 105.200 95.600 106.000 95.700 ;
        RECT 119.600 95.600 120.400 95.700 ;
        RECT 130.800 95.600 131.600 95.700 ;
        RECT 140.400 96.300 141.200 96.400 ;
        RECT 145.200 96.300 146.000 96.400 ;
        RECT 140.400 95.700 146.000 96.300 ;
        RECT 140.400 95.600 141.200 95.700 ;
        RECT 145.200 95.600 146.000 95.700 ;
        RECT 156.400 96.300 157.200 96.400 ;
        RECT 158.000 96.300 158.800 96.400 ;
        RECT 156.400 95.700 158.800 96.300 ;
        RECT 156.400 95.600 157.200 95.700 ;
        RECT 158.000 95.600 158.800 95.700 ;
        RECT 25.300 94.300 25.900 95.600 ;
        RECT 31.600 94.300 32.400 94.400 ;
        RECT 25.300 93.700 32.400 94.300 ;
        RECT 31.600 93.600 32.400 93.700 ;
        RECT 54.000 94.300 54.800 94.400 ;
        RECT 58.800 94.300 59.600 94.400 ;
        RECT 54.000 93.700 59.600 94.300 ;
        RECT 54.000 93.600 54.800 93.700 ;
        RECT 58.800 93.600 59.600 93.700 ;
        RECT 60.400 94.300 61.200 94.400 ;
        RECT 81.200 94.300 82.000 94.400 ;
        RECT 60.400 93.700 82.000 94.300 ;
        RECT 60.400 93.600 61.200 93.700 ;
        RECT 81.200 93.600 82.000 93.700 ;
        RECT 138.800 94.300 139.600 94.400 ;
        RECT 174.000 94.300 174.800 94.400 ;
        RECT 138.800 93.700 174.800 94.300 ;
        RECT 138.800 93.600 139.600 93.700 ;
        RECT 174.000 93.600 174.800 93.700 ;
        RECT 194.800 94.300 195.600 94.400 ;
        RECT 220.400 94.300 221.200 94.400 ;
        RECT 194.800 93.700 221.200 94.300 ;
        RECT 194.800 93.600 195.600 93.700 ;
        RECT 220.400 93.600 221.200 93.700 ;
        RECT 6.000 92.300 6.800 92.400 ;
        RECT 12.400 92.300 13.200 92.400 ;
        RECT 6.000 91.700 13.200 92.300 ;
        RECT 6.000 91.600 6.800 91.700 ;
        RECT 12.400 91.600 13.200 91.700 ;
        RECT 22.000 92.300 22.800 92.400 ;
        RECT 25.200 92.300 26.000 92.400 ;
        RECT 41.200 92.300 42.000 92.400 ;
        RECT 22.000 91.700 42.000 92.300 ;
        RECT 22.000 91.600 22.800 91.700 ;
        RECT 25.200 91.600 26.000 91.700 ;
        RECT 41.200 91.600 42.000 91.700 ;
        RECT 89.200 92.300 90.000 92.400 ;
        RECT 111.600 92.300 112.400 92.400 ;
        RECT 89.200 91.700 112.400 92.300 ;
        RECT 89.200 91.600 90.000 91.700 ;
        RECT 111.600 91.600 112.400 91.700 ;
        RECT 145.200 92.300 146.000 92.400 ;
        RECT 150.000 92.300 150.800 92.400 ;
        RECT 154.800 92.300 155.600 92.400 ;
        RECT 145.200 91.700 155.600 92.300 ;
        RECT 145.200 91.600 146.000 91.700 ;
        RECT 150.000 91.600 150.800 91.700 ;
        RECT 154.800 91.600 155.600 91.700 ;
        RECT 161.200 92.300 162.000 92.400 ;
        RECT 167.600 92.300 168.400 92.400 ;
        RECT 161.200 91.700 168.400 92.300 ;
        RECT 161.200 91.600 162.000 91.700 ;
        RECT 167.600 91.600 168.400 91.700 ;
        RECT 215.600 92.300 216.400 92.400 ;
        RECT 218.800 92.300 219.600 92.400 ;
        RECT 215.600 91.700 219.600 92.300 ;
        RECT 215.600 91.600 216.400 91.700 ;
        RECT 218.800 91.600 219.600 91.700 ;
        RECT 39.600 90.300 40.400 90.400 ;
        RECT 46.000 90.300 46.800 90.400 ;
        RECT 39.600 89.700 46.800 90.300 ;
        RECT 39.600 89.600 40.400 89.700 ;
        RECT 46.000 89.600 46.800 89.700 ;
        RECT 143.600 90.300 144.400 90.400 ;
        RECT 148.400 90.300 149.200 90.400 ;
        RECT 159.600 90.300 160.400 90.400 ;
        RECT 143.600 89.700 160.400 90.300 ;
        RECT 143.600 89.600 144.400 89.700 ;
        RECT 148.400 89.600 149.200 89.700 ;
        RECT 159.600 89.600 160.400 89.700 ;
        RECT 14.000 88.300 14.800 88.400 ;
        RECT 17.200 88.300 18.000 88.400 ;
        RECT 14.000 87.700 18.000 88.300 ;
        RECT 14.000 87.600 14.800 87.700 ;
        RECT 17.200 87.600 18.000 87.700 ;
        RECT 25.200 88.300 26.000 88.400 ;
        RECT 42.800 88.300 43.600 88.400 ;
        RECT 25.200 87.700 43.600 88.300 ;
        RECT 25.200 87.600 26.000 87.700 ;
        RECT 42.800 87.600 43.600 87.700 ;
        RECT 145.200 88.300 146.000 88.400 ;
        RECT 151.600 88.300 152.400 88.400 ;
        RECT 145.200 87.700 152.400 88.300 ;
        RECT 145.200 87.600 146.000 87.700 ;
        RECT 151.600 87.600 152.400 87.700 ;
        RECT 177.200 88.300 178.000 88.400 ;
        RECT 198.000 88.300 198.800 88.400 ;
        RECT 177.200 87.700 198.800 88.300 ;
        RECT 177.200 87.600 178.000 87.700 ;
        RECT 198.000 87.600 198.800 87.700 ;
        RECT 15.600 86.300 16.400 86.400 ;
        RECT 55.600 86.300 56.400 86.400 ;
        RECT 15.600 85.700 56.400 86.300 ;
        RECT 15.600 85.600 16.400 85.700 ;
        RECT 55.600 85.600 56.400 85.700 ;
        RECT 170.800 86.300 171.600 86.400 ;
        RECT 172.400 86.300 173.200 86.400 ;
        RECT 178.800 86.300 179.600 86.400 ;
        RECT 170.800 85.700 179.600 86.300 ;
        RECT 170.800 85.600 171.600 85.700 ;
        RECT 172.400 85.600 173.200 85.700 ;
        RECT 178.800 85.600 179.600 85.700 ;
        RECT 132.400 84.300 133.200 84.400 ;
        RECT 138.800 84.300 139.600 84.400 ;
        RECT 132.400 83.700 139.600 84.300 ;
        RECT 132.400 83.600 133.200 83.700 ;
        RECT 138.800 83.600 139.600 83.700 ;
        RECT 169.200 84.300 170.000 84.400 ;
        RECT 175.600 84.300 176.400 84.400 ;
        RECT 177.200 84.300 178.000 84.400 ;
        RECT 169.200 83.700 178.000 84.300 ;
        RECT 169.200 83.600 170.000 83.700 ;
        RECT 175.600 83.600 176.400 83.700 ;
        RECT 177.200 83.600 178.000 83.700 ;
        RECT 210.800 84.300 211.600 84.400 ;
        RECT 217.200 84.300 218.000 84.400 ;
        RECT 210.800 83.700 218.000 84.300 ;
        RECT 210.800 83.600 211.600 83.700 ;
        RECT 217.200 83.600 218.000 83.700 ;
        RECT 78.000 82.300 78.800 82.400 ;
        RECT 79.600 82.300 80.400 82.400 ;
        RECT 78.000 81.700 80.400 82.300 ;
        RECT 78.000 81.600 78.800 81.700 ;
        RECT 79.600 81.600 80.400 81.700 ;
        RECT 68.400 80.300 69.200 80.400 ;
        RECT 98.800 80.300 99.600 80.400 ;
        RECT 124.400 80.300 125.200 80.400 ;
        RECT 68.400 79.700 125.200 80.300 ;
        RECT 68.400 79.600 69.200 79.700 ;
        RECT 98.800 79.600 99.600 79.700 ;
        RECT 124.400 79.600 125.200 79.700 ;
        RECT 46.000 76.300 46.800 76.400 ;
        RECT 52.400 76.300 53.200 76.400 ;
        RECT 46.000 75.700 53.200 76.300 ;
        RECT 46.000 75.600 46.800 75.700 ;
        RECT 52.400 75.600 53.200 75.700 ;
        RECT 52.400 74.300 53.200 74.400 ;
        RECT 57.200 74.300 58.000 74.400 ;
        RECT 52.400 73.700 58.000 74.300 ;
        RECT 52.400 73.600 53.200 73.700 ;
        RECT 57.200 73.600 58.000 73.700 ;
        RECT 58.800 74.300 59.600 74.400 ;
        RECT 66.800 74.300 67.600 74.400 ;
        RECT 121.200 74.300 122.000 74.400 ;
        RECT 138.800 74.300 139.600 74.400 ;
        RECT 58.800 73.700 67.600 74.300 ;
        RECT 58.800 73.600 59.600 73.700 ;
        RECT 66.800 73.600 67.600 73.700 ;
        RECT 74.900 73.700 139.600 74.300 ;
        RECT 74.900 72.400 75.500 73.700 ;
        RECT 121.200 73.600 122.000 73.700 ;
        RECT 138.800 73.600 139.600 73.700 ;
        RECT 31.600 72.300 32.400 72.400 ;
        RECT 47.600 72.300 48.400 72.400 ;
        RECT 31.600 71.700 48.400 72.300 ;
        RECT 31.600 71.600 32.400 71.700 ;
        RECT 47.600 71.600 48.400 71.700 ;
        RECT 55.600 72.300 56.400 72.400 ;
        RECT 70.000 72.300 70.800 72.400 ;
        RECT 74.800 72.300 75.600 72.400 ;
        RECT 55.600 71.700 75.600 72.300 ;
        RECT 55.600 71.600 56.400 71.700 ;
        RECT 70.000 71.600 70.800 71.700 ;
        RECT 74.800 71.600 75.600 71.700 ;
        RECT 82.800 72.300 83.600 72.400 ;
        RECT 89.200 72.300 90.000 72.400 ;
        RECT 92.400 72.300 93.200 72.400 ;
        RECT 82.800 71.700 93.200 72.300 ;
        RECT 82.800 71.600 83.600 71.700 ;
        RECT 89.200 71.600 90.000 71.700 ;
        RECT 92.400 71.600 93.200 71.700 ;
        RECT 4.400 70.300 5.200 70.400 ;
        RECT 12.400 70.300 13.200 70.400 ;
        RECT 4.400 69.700 13.200 70.300 ;
        RECT 4.400 69.600 5.200 69.700 ;
        RECT 12.400 69.600 13.200 69.700 ;
        RECT 49.200 70.300 50.000 70.400 ;
        RECT 54.000 70.300 54.800 70.400 ;
        RECT 63.600 70.300 64.400 70.400 ;
        RECT 70.000 70.300 70.800 70.400 ;
        RECT 49.200 69.700 54.800 70.300 ;
        RECT 62.100 69.700 70.800 70.300 ;
        RECT 49.200 69.600 50.000 69.700 ;
        RECT 54.000 69.600 54.800 69.700 ;
        RECT 63.600 69.600 64.400 69.700 ;
        RECT 70.000 69.600 70.800 69.700 ;
        RECT 86.000 70.300 86.800 70.400 ;
        RECT 90.800 70.300 91.600 70.400 ;
        RECT 86.000 69.700 91.600 70.300 ;
        RECT 86.000 69.600 86.800 69.700 ;
        RECT 90.800 69.600 91.600 69.700 ;
        RECT 150.000 70.300 150.800 70.400 ;
        RECT 164.400 70.300 165.200 70.400 ;
        RECT 150.000 69.700 165.200 70.300 ;
        RECT 150.000 69.600 150.800 69.700 ;
        RECT 164.400 69.600 165.200 69.700 ;
        RECT 198.000 70.300 198.800 70.400 ;
        RECT 212.400 70.300 213.200 70.400 ;
        RECT 198.000 69.700 213.200 70.300 ;
        RECT 198.000 69.600 198.800 69.700 ;
        RECT 212.400 69.600 213.200 69.700 ;
        RECT 57.200 68.300 58.000 68.400 ;
        RECT 79.600 68.300 80.400 68.400 ;
        RECT 57.200 67.700 80.400 68.300 ;
        RECT 57.200 67.600 58.000 67.700 ;
        RECT 79.600 67.600 80.400 67.700 ;
        RECT 81.200 68.300 82.000 68.400 ;
        RECT 102.000 68.300 102.800 68.400 ;
        RECT 81.200 67.700 102.800 68.300 ;
        RECT 81.200 67.600 82.000 67.700 ;
        RECT 102.000 67.600 102.800 67.700 ;
        RECT 121.200 68.300 122.000 68.400 ;
        RECT 122.800 68.300 123.600 68.400 ;
        RECT 121.200 67.700 123.600 68.300 ;
        RECT 121.200 67.600 122.000 67.700 ;
        RECT 122.800 67.600 123.600 67.700 ;
        RECT 142.000 68.300 142.800 68.400 ;
        RECT 177.200 68.300 178.000 68.400 ;
        RECT 142.000 67.700 178.000 68.300 ;
        RECT 142.000 67.600 142.800 67.700 ;
        RECT 177.200 67.600 178.000 67.700 ;
        RECT 202.800 68.300 203.600 68.400 ;
        RECT 210.800 68.300 211.600 68.400 ;
        RECT 202.800 67.700 211.600 68.300 ;
        RECT 202.800 67.600 203.600 67.700 ;
        RECT 210.800 67.600 211.600 67.700 ;
        RECT 214.000 68.300 214.800 68.400 ;
        RECT 217.200 68.300 218.000 68.400 ;
        RECT 220.400 68.300 221.200 68.400 ;
        RECT 214.000 67.700 221.200 68.300 ;
        RECT 214.000 67.600 214.800 67.700 ;
        RECT 217.200 67.600 218.000 67.700 ;
        RECT 220.400 67.600 221.200 67.700 ;
        RECT 9.200 66.300 10.000 66.400 ;
        RECT 47.600 66.300 48.400 66.400 ;
        RECT 62.000 66.300 62.800 66.400 ;
        RECT 9.200 65.700 62.800 66.300 ;
        RECT 9.200 65.600 10.000 65.700 ;
        RECT 47.600 65.600 48.400 65.700 ;
        RECT 62.000 65.600 62.800 65.700 ;
        RECT 174.000 66.300 174.800 66.400 ;
        RECT 204.400 66.300 205.200 66.400 ;
        RECT 174.000 65.700 205.200 66.300 ;
        RECT 174.000 65.600 174.800 65.700 ;
        RECT 204.400 65.600 205.200 65.700 ;
        RECT 79.600 64.300 80.400 64.400 ;
        RECT 122.800 64.300 123.600 64.400 ;
        RECT 79.600 63.700 123.600 64.300 ;
        RECT 79.600 63.600 80.400 63.700 ;
        RECT 122.800 63.600 123.600 63.700 ;
        RECT 158.000 64.300 158.800 64.400 ;
        RECT 162.800 64.300 163.600 64.400 ;
        RECT 158.000 63.700 163.600 64.300 ;
        RECT 158.000 63.600 158.800 63.700 ;
        RECT 162.800 63.600 163.600 63.700 ;
        RECT 177.200 64.300 178.000 64.400 ;
        RECT 207.600 64.300 208.400 64.400 ;
        RECT 177.200 63.700 208.400 64.300 ;
        RECT 177.200 63.600 178.000 63.700 ;
        RECT 207.600 63.600 208.400 63.700 ;
        RECT 23.600 62.300 24.400 62.400 ;
        RECT 28.400 62.300 29.200 62.400 ;
        RECT 23.600 61.700 29.200 62.300 ;
        RECT 23.600 61.600 24.400 61.700 ;
        RECT 28.400 61.600 29.200 61.700 ;
        RECT 138.800 62.300 139.600 62.400 ;
        RECT 169.200 62.300 170.000 62.400 ;
        RECT 138.800 61.700 170.000 62.300 ;
        RECT 138.800 61.600 139.600 61.700 ;
        RECT 169.200 61.600 170.000 61.700 ;
        RECT 122.800 58.300 123.600 58.400 ;
        RECT 170.800 58.300 171.600 58.400 ;
        RECT 172.400 58.300 173.200 58.400 ;
        RECT 183.600 58.300 184.400 58.400 ;
        RECT 122.800 57.700 184.400 58.300 ;
        RECT 122.800 57.600 123.600 57.700 ;
        RECT 170.800 57.600 171.600 57.700 ;
        RECT 172.400 57.600 173.200 57.700 ;
        RECT 183.600 57.600 184.400 57.700 ;
        RECT 7.600 56.300 8.400 56.400 ;
        RECT 41.200 56.300 42.000 56.400 ;
        RECT 7.600 55.700 42.000 56.300 ;
        RECT 7.600 55.600 8.400 55.700 ;
        RECT 41.200 55.600 42.000 55.700 ;
        RECT 60.400 56.300 61.200 56.400 ;
        RECT 102.000 56.300 102.800 56.400 ;
        RECT 60.400 55.700 102.800 56.300 ;
        RECT 60.400 55.600 61.200 55.700 ;
        RECT 102.000 55.600 102.800 55.700 ;
        RECT 103.600 56.300 104.400 56.400 ;
        RECT 148.400 56.300 149.200 56.400 ;
        RECT 103.600 55.700 149.200 56.300 ;
        RECT 103.600 55.600 104.400 55.700 ;
        RECT 148.400 55.600 149.200 55.700 ;
        RECT 46.000 54.300 46.800 54.400 ;
        RECT 49.200 54.300 50.000 54.400 ;
        RECT 46.000 53.700 50.000 54.300 ;
        RECT 46.000 53.600 46.800 53.700 ;
        RECT 49.200 53.600 50.000 53.700 ;
        RECT 57.200 54.300 58.000 54.400 ;
        RECT 68.400 54.300 69.200 54.400 ;
        RECT 57.200 53.700 69.200 54.300 ;
        RECT 57.200 53.600 58.000 53.700 ;
        RECT 68.400 53.600 69.200 53.700 ;
        RECT 162.800 54.300 163.600 54.400 ;
        RECT 169.200 54.300 170.000 54.400 ;
        RECT 178.800 54.300 179.600 54.400 ;
        RECT 162.800 53.700 179.600 54.300 ;
        RECT 162.800 53.600 163.600 53.700 ;
        RECT 169.200 53.600 170.000 53.700 ;
        RECT 178.800 53.600 179.600 53.700 ;
        RECT 199.600 54.300 200.400 54.400 ;
        RECT 212.400 54.300 213.200 54.400 ;
        RECT 199.600 53.700 213.200 54.300 ;
        RECT 199.600 53.600 200.400 53.700 ;
        RECT 212.400 53.600 213.200 53.700 ;
        RECT 26.800 52.300 27.600 52.400 ;
        RECT 46.000 52.300 46.800 52.400 ;
        RECT 26.800 51.700 46.800 52.300 ;
        RECT 26.800 51.600 27.600 51.700 ;
        RECT 46.000 51.600 46.800 51.700 ;
        RECT 54.000 52.300 54.800 52.400 ;
        RECT 66.800 52.300 67.600 52.400 ;
        RECT 54.000 51.700 67.600 52.300 ;
        RECT 54.000 51.600 54.800 51.700 ;
        RECT 66.800 51.600 67.600 51.700 ;
        RECT 138.800 52.300 139.600 52.400 ;
        RECT 162.800 52.300 163.600 52.400 ;
        RECT 175.600 52.300 176.400 52.400 ;
        RECT 138.800 51.700 176.400 52.300 ;
        RECT 138.800 51.600 139.600 51.700 ;
        RECT 162.800 51.600 163.600 51.700 ;
        RECT 175.600 51.600 176.400 51.700 ;
        RECT 63.600 50.300 64.400 50.400 ;
        RECT 86.000 50.300 86.800 50.400 ;
        RECT 122.800 50.300 123.600 50.400 ;
        RECT 63.600 49.700 123.600 50.300 ;
        RECT 63.600 49.600 64.400 49.700 ;
        RECT 86.000 49.600 86.800 49.700 ;
        RECT 122.800 49.600 123.600 49.700 ;
        RECT 124.400 50.300 125.200 50.400 ;
        RECT 166.000 50.300 166.800 50.400 ;
        RECT 124.400 49.700 166.800 50.300 ;
        RECT 124.400 49.600 125.200 49.700 ;
        RECT 166.000 49.600 166.800 49.700 ;
        RECT 50.800 48.300 51.600 48.400 ;
        RECT 57.200 48.300 58.000 48.400 ;
        RECT 50.800 47.700 58.000 48.300 ;
        RECT 50.800 47.600 51.600 47.700 ;
        RECT 57.200 47.600 58.000 47.700 ;
        RECT 58.800 48.300 59.600 48.400 ;
        RECT 62.000 48.300 62.800 48.400 ;
        RECT 58.800 47.700 62.800 48.300 ;
        RECT 58.800 47.600 59.600 47.700 ;
        RECT 62.000 47.600 62.800 47.700 ;
        RECT 18.800 42.300 19.600 42.400 ;
        RECT 23.600 42.300 24.400 42.400 ;
        RECT 18.800 41.700 24.400 42.300 ;
        RECT 18.800 41.600 19.600 41.700 ;
        RECT 23.600 41.600 24.400 41.700 ;
        RECT 31.600 42.300 32.400 42.400 ;
        RECT 34.800 42.300 35.600 42.400 ;
        RECT 31.600 41.700 35.600 42.300 ;
        RECT 31.600 41.600 32.400 41.700 ;
        RECT 34.800 41.600 35.600 41.700 ;
        RECT 159.600 40.300 160.400 40.400 ;
        RECT 170.800 40.300 171.600 40.400 ;
        RECT 159.600 39.700 171.600 40.300 ;
        RECT 159.600 39.600 160.400 39.700 ;
        RECT 170.800 39.600 171.600 39.700 ;
        RECT 199.600 40.300 200.400 40.400 ;
        RECT 202.800 40.300 203.600 40.400 ;
        RECT 199.600 39.700 203.600 40.300 ;
        RECT 199.600 39.600 200.400 39.700 ;
        RECT 202.800 39.600 203.600 39.700 ;
        RECT 2.800 38.300 3.600 38.400 ;
        RECT 10.800 38.300 11.600 38.400 ;
        RECT 2.800 37.700 11.600 38.300 ;
        RECT 2.800 37.600 3.600 37.700 ;
        RECT 10.800 37.600 11.600 37.700 ;
        RECT 122.800 38.300 123.600 38.400 ;
        RECT 150.000 38.300 150.800 38.400 ;
        RECT 159.600 38.300 160.400 38.400 ;
        RECT 122.800 37.700 160.400 38.300 ;
        RECT 122.800 37.600 123.600 37.700 ;
        RECT 150.000 37.600 150.800 37.700 ;
        RECT 159.600 37.600 160.400 37.700 ;
        RECT 180.400 38.300 181.200 38.400 ;
        RECT 198.000 38.300 198.800 38.400 ;
        RECT 180.400 37.700 198.800 38.300 ;
        RECT 180.400 37.600 181.200 37.700 ;
        RECT 198.000 37.600 198.800 37.700 ;
        RECT 158.000 32.300 158.800 32.400 ;
        RECT 164.400 32.300 165.200 32.400 ;
        RECT 158.000 31.700 165.200 32.300 ;
        RECT 158.000 31.600 158.800 31.700 ;
        RECT 164.400 31.600 165.200 31.700 ;
        RECT 41.200 30.300 42.000 30.400 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 55.600 30.300 56.400 30.400 ;
        RECT 41.200 29.700 56.400 30.300 ;
        RECT 41.200 29.600 42.000 29.700 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 55.600 29.600 56.400 29.700 ;
        RECT 84.400 30.300 85.200 30.400 ;
        RECT 89.200 30.300 90.000 30.400 ;
        RECT 84.400 29.700 90.000 30.300 ;
        RECT 84.400 29.600 85.200 29.700 ;
        RECT 89.200 29.600 90.000 29.700 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 95.600 30.300 96.400 30.400 ;
        RECT 105.200 30.300 106.000 30.400 ;
        RECT 90.800 29.700 106.000 30.300 ;
        RECT 90.800 29.600 91.600 29.700 ;
        RECT 95.600 29.600 96.400 29.700 ;
        RECT 105.200 29.600 106.000 29.700 ;
        RECT 159.600 30.300 160.400 30.400 ;
        RECT 207.600 30.300 208.400 30.400 ;
        RECT 210.800 30.300 211.600 30.400 ;
        RECT 159.600 29.700 211.600 30.300 ;
        RECT 159.600 29.600 160.400 29.700 ;
        RECT 207.600 29.600 208.400 29.700 ;
        RECT 210.800 29.600 211.600 29.700 ;
        RECT 22.000 28.300 22.800 28.400 ;
        RECT 36.400 28.300 37.200 28.400 ;
        RECT 22.000 27.700 37.200 28.300 ;
        RECT 22.000 27.600 22.800 27.700 ;
        RECT 36.400 27.600 37.200 27.700 ;
        RECT 42.800 28.300 43.600 28.400 ;
        RECT 49.200 28.300 50.000 28.400 ;
        RECT 42.800 27.700 50.000 28.300 ;
        RECT 42.800 27.600 43.600 27.700 ;
        RECT 49.200 27.600 50.000 27.700 ;
        RECT 52.400 28.300 53.200 28.400 ;
        RECT 74.800 28.300 75.600 28.400 ;
        RECT 52.400 27.700 75.600 28.300 ;
        RECT 52.400 27.600 53.200 27.700 ;
        RECT 74.800 27.600 75.600 27.700 ;
        RECT 100.400 28.300 101.200 28.400 ;
        RECT 114.800 28.300 115.600 28.400 ;
        RECT 100.400 27.700 115.600 28.300 ;
        RECT 100.400 27.600 101.200 27.700 ;
        RECT 114.800 27.600 115.600 27.700 ;
        RECT 124.400 28.300 125.200 28.400 ;
        RECT 151.600 28.300 152.400 28.400 ;
        RECT 124.400 27.700 152.400 28.300 ;
        RECT 124.400 27.600 125.200 27.700 ;
        RECT 151.600 27.600 152.400 27.700 ;
        RECT 167.600 28.300 168.400 28.400 ;
        RECT 182.000 28.300 182.800 28.400 ;
        RECT 167.600 27.700 182.800 28.300 ;
        RECT 167.600 27.600 168.400 27.700 ;
        RECT 182.000 27.600 182.800 27.700 ;
        RECT 206.000 28.300 206.800 28.400 ;
        RECT 209.200 28.300 210.000 28.400 ;
        RECT 206.000 27.700 210.000 28.300 ;
        RECT 206.000 27.600 206.800 27.700 ;
        RECT 209.200 27.600 210.000 27.700 ;
        RECT 18.800 26.300 19.600 26.400 ;
        RECT 63.600 26.300 64.400 26.400 ;
        RECT 71.600 26.300 72.400 26.400 ;
        RECT 82.800 26.300 83.600 26.400 ;
        RECT 18.800 25.700 83.600 26.300 ;
        RECT 18.800 25.600 19.600 25.700 ;
        RECT 63.600 25.600 64.400 25.700 ;
        RECT 71.600 25.600 72.400 25.700 ;
        RECT 82.800 25.600 83.600 25.700 ;
        RECT 113.200 26.300 114.000 26.400 ;
        RECT 116.400 26.300 117.200 26.400 ;
        RECT 127.600 26.300 128.400 26.400 ;
        RECT 145.200 26.300 146.000 26.400 ;
        RECT 178.800 26.300 179.600 26.400 ;
        RECT 199.600 26.300 200.400 26.400 ;
        RECT 113.200 25.700 200.400 26.300 ;
        RECT 113.200 25.600 114.000 25.700 ;
        RECT 116.400 25.600 117.200 25.700 ;
        RECT 127.600 25.600 128.400 25.700 ;
        RECT 145.200 25.600 146.000 25.700 ;
        RECT 178.800 25.600 179.600 25.700 ;
        RECT 199.600 25.600 200.400 25.700 ;
        RECT 158.000 24.300 158.800 24.400 ;
        RECT 162.800 24.300 163.600 24.400 ;
        RECT 158.000 23.700 163.600 24.300 ;
        RECT 158.000 23.600 158.800 23.700 ;
        RECT 162.800 23.600 163.600 23.700 ;
        RECT 178.800 24.300 179.600 24.400 ;
        RECT 202.800 24.300 203.600 24.400 ;
        RECT 178.800 23.700 203.600 24.300 ;
        RECT 178.800 23.600 179.600 23.700 ;
        RECT 202.800 23.600 203.600 23.700 ;
        RECT 206.000 20.300 206.800 20.400 ;
        RECT 215.600 20.300 216.400 20.400 ;
        RECT 190.100 19.700 216.400 20.300 ;
        RECT 180.400 18.300 181.200 18.400 ;
        RECT 190.100 18.300 190.700 19.700 ;
        RECT 206.000 19.600 206.800 19.700 ;
        RECT 215.600 19.600 216.400 19.700 ;
        RECT 180.400 17.700 190.700 18.300 ;
        RECT 180.400 17.600 181.200 17.700 ;
        RECT 2.800 16.300 3.600 16.400 ;
        RECT 36.400 16.300 37.200 16.400 ;
        RECT 2.800 15.700 37.200 16.300 ;
        RECT 2.800 15.600 3.600 15.700 ;
        RECT 36.400 15.600 37.200 15.700 ;
        RECT 169.200 16.300 170.000 16.400 ;
        RECT 175.600 16.300 176.400 16.400 ;
        RECT 169.200 15.700 176.400 16.300 ;
        RECT 169.200 15.600 170.000 15.700 ;
        RECT 175.600 15.600 176.400 15.700 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 44.400 14.300 45.200 14.400 ;
        RECT 22.000 13.700 45.200 14.300 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 44.400 13.600 45.200 13.700 ;
        RECT 110.000 14.300 110.800 14.400 ;
        RECT 142.000 14.300 142.800 14.400 ;
        RECT 110.000 13.700 142.800 14.300 ;
        RECT 110.000 13.600 110.800 13.700 ;
        RECT 142.000 13.600 142.800 13.700 ;
        RECT 148.400 14.300 149.200 14.400 ;
        RECT 151.600 14.300 152.400 14.400 ;
        RECT 166.000 14.300 166.800 14.400 ;
        RECT 148.400 13.700 152.400 14.300 ;
        RECT 148.400 13.600 149.200 13.700 ;
        RECT 151.600 13.600 152.400 13.700 ;
        RECT 156.500 13.700 166.800 14.300 ;
        RECT 156.500 12.400 157.100 13.700 ;
        RECT 166.000 13.600 166.800 13.700 ;
        RECT 170.800 14.300 171.600 14.400 ;
        RECT 175.600 14.300 176.400 14.400 ;
        RECT 170.800 13.700 176.400 14.300 ;
        RECT 170.800 13.600 171.600 13.700 ;
        RECT 175.600 13.600 176.400 13.700 ;
        RECT 31.600 12.300 32.400 12.400 ;
        RECT 55.600 12.300 56.400 12.400 ;
        RECT 31.600 11.700 56.400 12.300 ;
        RECT 31.600 11.600 32.400 11.700 ;
        RECT 55.600 11.600 56.400 11.700 ;
        RECT 76.400 12.300 77.200 12.400 ;
        RECT 84.400 12.300 85.200 12.400 ;
        RECT 76.400 11.700 85.200 12.300 ;
        RECT 76.400 11.600 77.200 11.700 ;
        RECT 84.400 11.600 85.200 11.700 ;
        RECT 132.400 12.300 133.200 12.400 ;
        RECT 138.800 12.300 139.600 12.400 ;
        RECT 132.400 11.700 139.600 12.300 ;
        RECT 132.400 11.600 133.200 11.700 ;
        RECT 138.800 11.600 139.600 11.700 ;
        RECT 148.400 12.300 149.200 12.400 ;
        RECT 156.400 12.300 157.200 12.400 ;
        RECT 148.400 11.700 157.200 12.300 ;
        RECT 148.400 11.600 149.200 11.700 ;
        RECT 156.400 11.600 157.200 11.700 ;
        RECT 164.400 12.300 165.200 12.400 ;
        RECT 178.800 12.300 179.600 12.400 ;
        RECT 164.400 11.700 179.600 12.300 ;
        RECT 164.400 11.600 165.200 11.700 ;
        RECT 178.800 11.600 179.600 11.700 ;
      LAYER metal4 ;
        RECT 7.400 133.400 8.600 150.600 ;
        RECT 20.200 95.400 21.400 188.600 ;
        RECT 36.200 109.400 37.400 150.600 ;
        RECT 71.400 95.400 72.600 146.600 ;
        RECT 90.600 135.400 91.800 146.600 ;
        RECT 77.800 81.400 79.000 98.600 ;
        RECT 90.600 29.400 91.800 110.600 ;
        RECT 122.600 67.400 123.800 104.600 ;
        RECT 154.600 91.400 155.800 144.600 ;
        RECT 161.000 141.400 162.200 176.600 ;
        RECT 167.400 137.400 168.600 158.600 ;
        RECT 157.800 95.400 159.000 132.600 ;
        RECT 138.600 51.400 139.800 84.600 ;
        RECT 170.600 13.400 171.800 100.600 ;
        RECT 177.000 63.400 178.200 84.600 ;
  END
END map9v3
END LIBRARY


magic
tech scmos
magscale 1 2
timestamp 1743498307
<< metal1 >>
rect 1496 5606 1502 5614
rect 1510 5606 1516 5614
rect 1524 5606 1530 5614
rect 1538 5606 1544 5614
rect 4568 5606 4574 5614
rect 4582 5606 4588 5614
rect 4596 5606 4602 5614
rect 4610 5606 4616 5614
rect 636 5537 675 5543
rect 1898 5536 1900 5544
rect 476 5532 484 5536
rect 612 5516 620 5524
rect 1940 5517 1955 5523
rect 2461 5517 2499 5523
rect 429 5497 444 5503
rect 532 5497 547 5503
rect 1821 5497 1836 5503
rect 1853 5497 1868 5503
rect 2397 5497 2435 5503
rect 2894 5497 2931 5503
rect 3453 5503 3459 5523
rect 3652 5516 3660 5524
rect 3677 5517 3715 5523
rect 3453 5497 3491 5503
rect 3597 5497 3628 5503
rect 4429 5503 4435 5523
rect 4429 5497 4467 5503
rect 4861 5503 4867 5523
rect 5316 5516 5324 5524
rect 4861 5497 4899 5503
rect 13 5477 28 5483
rect 493 5477 531 5483
rect 1917 5477 1932 5483
rect 3389 5477 3411 5483
rect 3549 5477 3571 5483
rect 4541 5477 4572 5483
rect 5261 5477 5276 5483
rect 365 5457 380 5463
rect 2349 5457 2380 5463
rect 3012 5457 3043 5463
rect 468 5436 470 5444
rect 4596 5437 4627 5443
rect 3032 5406 3038 5414
rect 3046 5406 3052 5414
rect 3060 5406 3066 5414
rect 3074 5406 3080 5414
rect 436 5356 444 5364
rect 2077 5357 2115 5363
rect 5421 5357 5436 5363
rect 493 5337 515 5343
rect 1229 5337 1244 5343
rect 1341 5337 1426 5343
rect 2237 5337 2252 5343
rect 3549 5337 3571 5343
rect 3588 5337 3603 5343
rect 3645 5337 3660 5343
rect 3741 5337 3763 5343
rect 3805 5337 3820 5343
rect 6045 5337 6067 5343
rect 1060 5317 1075 5323
rect 1149 5317 1187 5323
rect 1213 5317 1228 5323
rect 356 5297 371 5303
rect 596 5296 604 5304
rect 621 5297 659 5303
rect 1181 5297 1187 5317
rect 1309 5317 1404 5323
rect 2125 5317 2163 5323
rect 2189 5317 2227 5323
rect 2189 5297 2195 5317
rect 2973 5317 3011 5323
rect 3629 5317 3644 5323
rect 3652 5317 3683 5323
rect 3693 5317 3724 5323
rect 4557 5317 4643 5323
rect 3037 5297 3123 5303
rect 4557 5297 4563 5317
rect 4676 5317 4691 5323
rect 4740 5317 4771 5323
rect 4797 5317 4835 5323
rect 4797 5297 4803 5317
rect 4925 5317 4963 5323
rect 4925 5297 4931 5317
rect 5236 5317 5251 5323
rect 5988 5317 6019 5323
rect 5421 5297 5436 5303
rect 4532 5276 4534 5284
rect 1496 5206 1502 5214
rect 1510 5206 1516 5214
rect 1524 5206 1530 5214
rect 1538 5206 1544 5214
rect 4568 5206 4574 5214
rect 4582 5206 4588 5214
rect 4596 5206 4602 5214
rect 4610 5206 4616 5214
rect 1332 5176 1334 5184
rect 4522 5176 4524 5184
rect 4890 5176 4892 5184
rect 2340 5137 2356 5143
rect 3188 5137 3252 5143
rect 3244 5132 3252 5137
rect 3292 5132 3300 5136
rect 3718 5136 3724 5144
rect 3564 5132 3572 5136
rect 3932 5132 3940 5136
rect 4828 5132 4836 5136
rect 5460 5136 5462 5144
rect 5484 5137 5507 5143
rect 5036 5132 5044 5136
rect 548 5097 579 5103
rect 589 5097 604 5103
rect 685 5103 691 5123
rect 708 5116 716 5124
rect 612 5097 643 5103
rect 653 5097 691 5103
rect 1284 5097 1299 5103
rect 1357 5097 1372 5103
rect 3684 5097 3699 5103
rect 3853 5097 3891 5103
rect 605 5077 620 5083
rect 3853 5083 3859 5097
rect 3972 5097 4003 5103
rect 4013 5097 4028 5103
rect 4484 5097 4499 5103
rect 4925 5097 4940 5103
rect 5108 5097 5139 5103
rect 5300 5097 5331 5103
rect 5405 5097 5436 5103
rect 3837 5077 3859 5083
rect 4029 5077 4067 5083
rect 4125 5077 4140 5083
rect 4372 5077 4387 5083
rect 5300 5077 5315 5083
rect 500 5056 502 5064
rect 1428 5057 1443 5063
rect 1453 5037 1500 5043
rect 1780 5036 1784 5044
rect 3204 5037 3251 5043
rect 3306 5036 3308 5044
rect 3556 5036 3558 5044
rect 4580 5037 4627 5043
rect 4820 5036 4822 5044
rect 5706 5036 5708 5044
rect 3032 5006 3038 5014
rect 3046 5006 3052 5014
rect 3060 5006 3066 5014
rect 3074 5006 3080 5014
rect 1277 4957 1315 4963
rect 1725 4957 1740 4963
rect 77 4937 99 4943
rect 77 4923 83 4937
rect 500 4937 515 4943
rect 1261 4937 1276 4943
rect 3389 4937 3404 4943
rect 5037 4937 5059 4943
rect 45 4917 83 4923
rect 500 4917 515 4923
rect 596 4917 611 4923
rect 765 4917 796 4923
rect 909 4917 947 4923
rect 973 4917 988 4923
rect 941 4897 947 4917
rect 1229 4917 1244 4923
rect 1229 4897 1235 4917
rect 3165 4917 3180 4923
rect 3492 4917 3507 4923
rect 3629 4917 3667 4923
rect 3629 4897 3635 4917
rect 3716 4917 3731 4923
rect 4045 4917 4083 4923
rect 4045 4897 4051 4917
rect 4189 4917 4204 4923
rect 4445 4917 4483 4923
rect 4509 4917 4524 4923
rect 4477 4897 4483 4917
rect 4548 4917 4563 4923
rect 4685 4917 4723 4923
rect 4589 4897 4636 4903
rect 4717 4897 4723 4917
rect 5053 4923 5059 4937
rect 5053 4917 5091 4923
rect 5117 4917 5155 4923
rect 5117 4897 5123 4917
rect 5300 4917 5315 4923
rect 5228 4904 5236 4914
rect 5476 4896 5484 4904
rect 5516 4903 5524 4908
rect 5501 4897 5524 4903
rect 374 4876 380 4884
rect 2100 4877 2115 4883
rect 3450 4876 3452 4884
rect 1034 4856 1036 4864
rect 1162 4836 1164 4844
rect 1706 4836 1708 4844
rect 2996 4836 2998 4844
rect 3604 4836 3606 4844
rect 4564 4836 4566 4844
rect 1496 4806 1502 4814
rect 1510 4806 1516 4814
rect 1524 4806 1530 4814
rect 1538 4806 1544 4814
rect 4568 4806 4574 4814
rect 4582 4806 4588 4814
rect 4596 4806 4602 4814
rect 4610 4806 4616 4814
rect 2148 4776 2150 4784
rect 3380 4776 3382 4784
rect 4484 4776 4486 4784
rect 4900 4776 4902 4784
rect 5114 4776 5116 4784
rect 5172 4776 5174 4784
rect 1242 4756 1244 4764
rect 3546 4756 3548 4764
rect 1364 4736 1366 4744
rect 748 4732 756 4736
rect 253 4703 259 4723
rect 253 4697 291 4703
rect 589 4703 595 4723
rect 1300 4716 1308 4724
rect 557 4697 595 4703
rect 660 4697 675 4703
rect 964 4697 979 4703
rect 1101 4697 1116 4703
rect 1245 4697 1276 4703
rect 1556 4697 1571 4703
rect 1732 4697 1747 4703
rect 2077 4703 2083 4723
rect 2077 4697 2115 4703
rect 2173 4703 2179 4723
rect 3405 4717 3427 4723
rect 2173 4697 2211 4703
rect 2404 4697 2412 4703
rect 2420 4697 2435 4703
rect 3348 4697 3379 4703
rect 3517 4703 3523 4723
rect 4253 4717 4268 4723
rect 3485 4697 3523 4703
rect 3572 4697 3603 4703
rect 4365 4703 4371 4723
rect 4365 4697 4403 4703
rect 4509 4697 4604 4703
rect 4925 4697 4956 4703
rect 5085 4703 5091 4716
rect 5085 4697 5107 4703
rect 5741 4697 5788 4703
rect 804 4677 819 4683
rect 1597 4677 1628 4683
rect 2244 4677 2259 4683
rect 2436 4677 2451 4683
rect 3341 4677 3347 4696
rect 3437 4677 3452 4683
rect 1501 4657 1532 4663
rect 3437 4657 3443 4677
rect 3565 4677 3580 4683
rect 4260 4677 4275 4683
rect 4532 4677 4611 4683
rect 5341 4677 5379 4683
rect 5469 4677 5507 4683
rect 5780 4677 5810 4683
rect 5133 4657 5148 4663
rect 5325 4657 5347 4663
rect 5517 4657 5539 4663
rect 2068 4636 2070 4644
rect 4244 4636 4246 4644
rect 4708 4636 4710 4644
rect 5432 4636 5436 4644
rect 5624 4636 5628 4644
rect 3032 4606 3038 4614
rect 3046 4606 3052 4614
rect 3060 4606 3066 4614
rect 3074 4606 3080 4614
rect 1485 4577 1500 4583
rect 2074 4576 2076 4584
rect 3700 4556 3702 4564
rect 4868 4556 4870 4564
rect 2220 4552 2228 4556
rect 276 4537 291 4543
rect 781 4537 796 4543
rect 925 4537 963 4543
rect 1373 4537 1395 4543
rect 2813 4537 2851 4543
rect 3565 4537 3580 4543
rect 3588 4537 3603 4543
rect 3844 4537 3859 4543
rect 4573 4537 4643 4543
rect 5037 4537 5052 4543
rect 5213 4537 5251 4543
rect 781 4517 796 4523
rect 861 4517 899 4523
rect 836 4496 844 4504
rect 861 4497 867 4517
rect 1012 4517 1027 4523
rect 1373 4517 1388 4523
rect 1373 4497 1379 4517
rect 3821 4517 3852 4523
rect 3981 4517 3996 4523
rect 4644 4517 4659 4523
rect 4733 4517 4771 4523
rect 2045 4497 2067 4503
rect 2893 4497 2979 4503
rect 4429 4497 4444 4503
rect 4765 4497 4771 4517
rect 1117 4477 1148 4483
rect 1412 4436 1414 4444
rect 4202 4436 4204 4444
rect 4266 4436 4268 4444
rect 4324 4436 4326 4444
rect 4660 4436 4662 4444
rect 5290 4436 5292 4444
rect 1496 4406 1502 4414
rect 1510 4406 1516 4414
rect 1524 4406 1530 4414
rect 1538 4406 1544 4414
rect 4568 4406 4574 4414
rect 4582 4406 4588 4414
rect 4596 4406 4602 4414
rect 4610 4406 4616 4414
rect 282 4376 284 4384
rect 1802 4376 1804 4384
rect 3828 4376 3830 4384
rect 662 4336 668 4344
rect 1674 4336 1676 4344
rect 4708 4337 4771 4343
rect 589 4297 604 4303
rect 797 4297 835 4303
rect 29 4277 51 4283
rect 301 4277 323 4283
rect 317 4264 323 4277
rect 797 4283 803 4297
rect 861 4303 867 4323
rect 861 4297 899 4303
rect 1053 4297 1068 4303
rect 1133 4303 1139 4323
rect 1133 4297 1171 4303
rect 1645 4303 1651 4323
rect 1572 4297 1603 4303
rect 1613 4297 1651 4303
rect 1773 4303 1779 4323
rect 2365 4317 2403 4323
rect 1741 4297 1779 4303
rect 2196 4297 2227 4303
rect 2253 4297 2275 4303
rect 781 4277 803 4283
rect 1053 4277 1068 4283
rect 1229 4277 1251 4283
rect 2077 4277 2099 4283
rect 2253 4277 2259 4297
rect 2436 4297 2451 4303
rect 2653 4297 2668 4303
rect 3565 4297 3603 4303
rect 2477 4277 2499 4283
rect 3565 4283 3571 4297
rect 3629 4303 3635 4323
rect 4733 4317 4748 4323
rect 3629 4297 3667 4303
rect 3860 4297 3891 4303
rect 3949 4297 3964 4303
rect 4125 4297 4140 4303
rect 4260 4297 4275 4303
rect 4381 4297 4396 4303
rect 4509 4297 4540 4303
rect 3549 4277 3571 4283
rect 4365 4277 4387 4283
rect 5517 4277 5532 4283
rect 2509 4257 2531 4263
rect 964 4236 966 4244
rect 2356 4236 2358 4244
rect 2794 4236 2796 4244
rect 3032 4206 3038 4214
rect 3046 4206 3052 4214
rect 3060 4206 3066 4214
rect 3074 4206 3080 4214
rect 2728 4176 2732 4184
rect 4516 4176 4518 4184
rect 4808 4176 4812 4184
rect 5416 4176 5420 4184
rect 5656 4176 5660 4184
rect 2141 4157 2172 4163
rect 2189 4157 2211 4163
rect 5229 4157 5251 4163
rect 413 4137 428 4143
rect 1012 4137 1027 4143
rect 1069 4137 1084 4143
rect 1460 4137 1475 4143
rect 2285 4137 2328 4143
rect 2484 4137 2499 4143
rect 2893 4137 2915 4143
rect 2925 4137 2988 4143
rect 3853 4137 3875 4143
rect 4141 4137 4163 4143
rect 4532 4137 4547 4143
rect 4557 4137 4604 4143
rect 4989 4143 4995 4156
rect 461 4117 476 4123
rect 893 4117 931 4123
rect 333 4097 364 4103
rect 893 4097 899 4117
rect 1028 4117 1043 4123
rect 1204 4117 1219 4123
rect 1437 4117 1468 4123
rect 1748 4117 1779 4123
rect 2429 4117 2451 4123
rect 3581 4117 3619 4123
rect 3613 4097 3619 4117
rect 3741 4117 3779 4123
rect 3773 4097 3779 4117
rect 4045 4117 4060 4123
rect 4189 4117 4243 4123
rect 4525 4117 4563 4123
rect 4381 4097 4403 4103
rect 4525 4097 4531 4117
rect 4909 4123 4915 4143
rect 4973 4137 4995 4143
rect 5341 4143 5347 4163
rect 5341 4137 5356 4143
rect 5581 4137 5603 4143
rect 4909 4117 4931 4123
rect 5037 4117 5075 4123
rect 5277 4117 5299 4123
rect 5460 4117 5491 4123
rect 4580 4097 4627 4103
rect 5085 4097 5123 4103
rect 5220 4097 5235 4103
rect 2892 4077 2908 4083
rect 3494 4076 3500 4084
rect 4650 4056 4652 4064
rect 868 4036 870 4044
rect 1332 4036 1334 4044
rect 1780 4036 1782 4044
rect 2228 4036 2230 4044
rect 3802 4036 3804 4044
rect 4244 4036 4246 4044
rect 4308 4036 4310 4044
rect 4452 4036 4454 4044
rect 4714 4036 4716 4044
rect 4890 4036 4892 4044
rect 5492 4036 5494 4044
rect 1496 4006 1502 4014
rect 1510 4006 1516 4014
rect 1524 4006 1530 4014
rect 1538 4006 1544 4014
rect 4568 4006 4574 4014
rect 4582 4006 4588 4014
rect 4596 4006 4602 4014
rect 4610 4006 4616 4014
rect 5098 3976 5100 3984
rect 4468 3937 4484 3943
rect 5610 3936 5612 3944
rect 364 3932 372 3936
rect 580 3897 595 3903
rect 765 3897 796 3903
rect 877 3897 892 3903
rect 1101 3897 1116 3903
rect 1389 3903 1395 3923
rect 1357 3897 1395 3903
rect 1501 3897 1564 3903
rect 1645 3897 1682 3903
rect 2532 3897 2563 3903
rect 5524 3897 5539 3903
rect 5549 3897 5580 3903
rect 1444 3877 1475 3883
rect 2589 3877 2611 3883
rect 4436 3877 4451 3883
rect 4461 3877 4483 3883
rect 5629 3877 5651 3883
rect 333 3857 348 3863
rect 1524 3857 1571 3863
rect 378 3836 380 3844
rect 3032 3806 3038 3814
rect 3046 3806 3052 3814
rect 3060 3806 3066 3814
rect 3074 3806 3080 3814
rect 253 3737 268 3743
rect 637 3737 659 3743
rect 29 3717 44 3723
rect 189 3717 227 3723
rect 237 3717 284 3723
rect 189 3697 195 3717
rect 541 3717 556 3723
rect 653 3723 659 3737
rect 788 3737 803 3743
rect 2253 3737 2268 3743
rect 3261 3737 3283 3743
rect 3373 3737 3388 3743
rect 4196 3737 4227 3743
rect 4237 3737 4259 3743
rect 4301 3737 4316 3743
rect 4365 3737 4387 3743
rect 4397 3737 4476 3743
rect 5012 3737 5027 3743
rect 653 3717 691 3723
rect 717 3717 755 3723
rect 765 3717 812 3723
rect 477 3697 515 3703
rect 717 3697 723 3717
rect 829 3717 867 3723
rect 861 3697 867 3717
rect 1028 3717 1043 3723
rect 1341 3717 1372 3723
rect 1469 3717 1532 3723
rect 2173 3717 2188 3723
rect 2237 3717 2284 3723
rect 3149 3717 3187 3723
rect 3245 3717 3260 3723
rect 3373 3717 3411 3723
rect 4285 3717 4332 3723
rect 5181 3717 5218 3723
rect 884 3696 892 3704
rect 1133 3697 1155 3703
rect 2132 3697 2147 3703
rect 2317 3697 2355 3703
rect 4244 3697 4259 3703
rect 4365 3697 4380 3703
rect 4413 3697 4444 3703
rect 5709 3697 5747 3703
rect 6109 3677 6124 3683
rect 164 3636 166 3644
rect 292 3636 294 3644
rect 692 3636 694 3644
rect 1236 3636 1238 3644
rect 1496 3606 1502 3614
rect 1510 3606 1516 3614
rect 1524 3606 1530 3614
rect 1538 3606 1544 3614
rect 4568 3606 4574 3614
rect 4582 3606 4588 3614
rect 4596 3606 4602 3614
rect 4610 3606 4616 3614
rect 4516 3576 4518 3584
rect 541 3537 556 3543
rect 970 3536 972 3544
rect 516 3517 531 3523
rect 820 3517 835 3523
rect 845 3517 883 3523
rect 900 3516 908 3524
rect 669 3497 684 3503
rect 932 3497 963 3503
rect 973 3497 1011 3503
rect 1101 3497 1132 3503
rect 1181 3503 1187 3523
rect 4061 3517 4076 3523
rect 5620 3516 5628 3524
rect 1181 3497 1219 3503
rect 1389 3497 1420 3503
rect 1629 3497 1667 3503
rect 2765 3497 2803 3503
rect 3220 3497 3244 3503
rect 3252 3497 3267 3503
rect 3325 3497 3363 3503
rect 3828 3497 3843 3503
rect 4525 3497 4610 3503
rect 5604 3497 5619 3503
rect 6052 3497 6067 3503
rect 29 3477 51 3483
rect 1101 3477 1116 3483
rect 2132 3477 2163 3483
rect 2317 3477 2332 3483
rect 3757 3477 3779 3483
rect 3812 3477 3843 3483
rect 5460 3477 5475 3483
rect 6004 3477 6019 3483
rect 6093 3477 6124 3483
rect 452 3457 467 3463
rect 1572 3457 1619 3463
rect 2740 3456 2742 3464
rect 3300 3456 3302 3464
rect 1364 3436 1366 3444
rect 1690 3436 1692 3444
rect 4026 3436 4028 3444
rect 4116 3436 4118 3444
rect 5316 3436 5318 3444
rect 6036 3436 6038 3444
rect 3032 3406 3038 3414
rect 3046 3406 3052 3414
rect 3060 3406 3066 3414
rect 3074 3406 3080 3414
rect 333 3357 348 3363
rect 1469 3357 1555 3363
rect 980 3337 995 3343
rect 2829 3337 2851 3343
rect 2893 3337 2915 3343
rect 2957 3337 2979 3343
rect 3021 3337 3043 3343
rect 429 3317 483 3323
rect 957 3317 995 3323
rect 1133 3317 1164 3323
rect 2829 3317 2835 3337
rect 2893 3317 2899 3337
rect 2957 3317 2963 3337
rect 3021 3317 3027 3337
rect 3060 3337 3123 3343
rect 3901 3343 3907 3363
rect 4765 3357 4787 3363
rect 5037 3357 5052 3363
rect 3885 3337 3907 3343
rect 4564 3337 4643 3343
rect 4701 3337 4739 3343
rect 3181 3317 3235 3323
rect 3821 3317 3875 3323
rect 3949 3317 3986 3323
rect 4381 3317 4419 3323
rect 4541 3317 4604 3323
rect 4733 3317 4739 3337
rect 5940 3337 5955 3343
rect 5837 3317 5875 3323
rect 5981 3317 6019 3323
rect 3037 3297 3052 3303
rect 4420 3296 4428 3304
rect 5725 3297 5763 3303
rect 5773 3297 5811 3303
rect 3738 3276 3740 3284
rect 4964 3277 4979 3283
rect 4746 3236 4748 3244
rect 5018 3236 5020 3244
rect 1496 3206 1502 3214
rect 1510 3206 1516 3214
rect 1524 3206 1530 3214
rect 1538 3206 1544 3214
rect 4568 3206 4574 3214
rect 4582 3206 4588 3214
rect 4596 3206 4602 3214
rect 4610 3206 4616 3214
rect 2692 3176 2694 3184
rect 5258 3176 5260 3184
rect 3588 3137 3619 3143
rect 5028 3136 5030 3144
rect 5092 3136 5094 3144
rect 5220 3137 5236 3143
rect 1980 3124 1988 3128
rect 3357 3117 3372 3123
rect 941 3097 956 3103
rect 1021 3097 1059 3103
rect 2637 3097 2652 3103
rect 2717 3097 2748 3103
rect 2804 3097 2819 3103
rect 868 3077 883 3083
rect 1021 3077 1036 3083
rect 2388 3077 2403 3083
rect 2413 3077 2451 3083
rect 2525 3077 2540 3083
rect 2740 3077 2755 3083
rect 2813 3077 2819 3097
rect 2852 3097 2867 3103
rect 2893 3097 2924 3103
rect 3405 3103 3411 3123
rect 4701 3117 4716 3123
rect 5940 3117 5955 3123
rect 3405 3097 3443 3103
rect 3453 3097 3507 3103
rect 2909 3077 2940 3083
rect 3341 3077 3379 3083
rect 3533 3077 3555 3083
rect 3581 3077 3587 3108
rect 3652 3097 3667 3103
rect 3693 3083 3699 3108
rect 3997 3097 4028 3103
rect 4061 3097 4076 3103
rect 4221 3097 4236 3103
rect 4685 3097 4716 3103
rect 4909 3097 4947 3103
rect 4989 3097 5004 3103
rect 5124 3097 5155 3103
rect 5885 3097 5923 3103
rect 5981 3097 6019 3103
rect 3677 3077 3699 3083
rect 4733 3077 4755 3083
rect 6077 3077 6124 3083
rect 1069 3057 1107 3063
rect 1453 3057 1539 3063
rect 1972 3037 1987 3043
rect 3396 3036 3398 3044
rect 3604 3037 3619 3043
rect 3930 3036 3932 3044
rect 3032 3006 3038 3014
rect 3046 3006 3052 3014
rect 3060 3006 3066 3014
rect 3074 3006 3080 3014
rect 3364 2976 3366 2984
rect 3876 2976 3878 2984
rect 4356 2976 4358 2984
rect 4436 2976 4438 2984
rect 4980 2976 4982 2984
rect 477 2957 515 2963
rect 525 2957 563 2963
rect 941 2957 979 2963
rect 989 2957 1027 2963
rect 2509 2957 2547 2963
rect 3453 2957 3475 2963
rect 4541 2957 4588 2963
rect 1629 2937 1651 2943
rect 2030 2937 2060 2943
rect 2109 2937 2147 2943
rect 2580 2937 2595 2943
rect 2990 2937 3027 2943
rect 3037 2937 3123 2943
rect 3181 2937 3219 2943
rect 2132 2917 2163 2923
rect 2557 2917 2595 2923
rect 3060 2917 3139 2923
rect 3373 2917 3411 2923
rect 3421 2917 3443 2923
rect 2125 2897 2140 2903
rect 3236 2896 3244 2904
rect 3373 2897 3379 2917
rect 3533 2912 3539 2943
rect 3741 2937 3763 2943
rect 3757 2917 3763 2937
rect 4461 2937 4476 2943
rect 4516 2937 4531 2943
rect 4804 2937 4819 2943
rect 4893 2943 4899 2956
rect 4893 2937 4908 2943
rect 5053 2937 5068 2943
rect 5268 2937 5283 2943
rect 4484 2917 4499 2923
rect 4996 2917 5027 2923
rect 5037 2917 5084 2923
rect 3965 2897 3980 2903
rect 5117 2897 5155 2903
rect 3437 2877 3507 2883
rect 3732 2877 3763 2883
rect 3757 2857 3763 2877
rect 4676 2877 4707 2883
rect 4941 2877 4956 2883
rect 1156 2836 1158 2844
rect 3636 2836 3638 2844
rect 5194 2836 5196 2844
rect 1496 2806 1502 2814
rect 1510 2806 1516 2814
rect 1524 2806 1530 2814
rect 1538 2806 1544 2814
rect 4568 2806 4574 2814
rect 4582 2806 4588 2814
rect 4596 2806 4602 2814
rect 4610 2806 4616 2814
rect 4922 2776 4924 2784
rect 5252 2776 5254 2784
rect 5316 2776 5318 2784
rect 3444 2737 3459 2743
rect 4541 2737 4556 2743
rect 4653 2743 4659 2763
rect 4573 2737 4659 2743
rect 2884 2716 2892 2724
rect 3476 2717 3491 2723
rect 3572 2716 3580 2724
rect 4573 2717 4579 2737
rect 4708 2737 4739 2743
rect 5098 2736 5100 2744
rect 5708 2737 5724 2743
rect 4701 2717 4716 2723
rect 5597 2717 5612 2723
rect 1540 2697 1587 2703
rect 2109 2697 2124 2703
rect 2733 2697 2771 2703
rect 2788 2697 2819 2703
rect 2829 2697 2860 2703
rect 3492 2697 3507 2703
rect 3540 2697 3571 2703
rect 3604 2697 3619 2703
rect 756 2677 787 2683
rect 1373 2677 1388 2683
rect 1613 2677 1628 2683
rect 2132 2677 2147 2683
rect 2157 2677 2195 2683
rect 3021 2677 3084 2683
rect 3709 2683 3715 2703
rect 3693 2677 3715 2683
rect 3885 2677 3891 2708
rect 4020 2697 4035 2703
rect 4148 2697 4163 2703
rect 4228 2697 4243 2703
rect 5101 2697 5116 2703
rect 3997 2677 4012 2683
rect 4125 2677 4156 2683
rect 5181 2683 5187 2703
rect 5197 2697 5251 2703
rect 5149 2677 5187 2683
rect 5533 2677 5548 2683
rect 5597 2677 5619 2683
rect 5652 2677 5667 2683
rect 5709 2677 5731 2683
rect 5741 2677 5772 2683
rect 733 2657 771 2663
rect 2708 2656 2710 2664
rect 3658 2636 3660 2644
rect 5386 2636 5388 2644
rect 5514 2636 5516 2644
rect 3032 2606 3038 2614
rect 3046 2606 3052 2614
rect 3060 2606 3066 2614
rect 3074 2606 3080 2614
rect 1732 2577 1747 2583
rect 3012 2576 3014 2584
rect 3988 2576 3990 2584
rect 4330 2576 4332 2584
rect 4776 2576 4780 2584
rect 765 2557 803 2563
rect 877 2557 892 2563
rect 925 2557 963 2563
rect 2269 2557 2307 2563
rect 4244 2556 4252 2564
rect 1316 2537 1347 2543
rect 1828 2537 1843 2543
rect 1892 2537 1923 2543
rect 2340 2537 2355 2543
rect 3156 2537 3171 2543
rect 884 2517 899 2523
rect 1805 2517 1843 2523
rect 1837 2497 1843 2517
rect 2317 2517 2355 2523
rect 2413 2517 2428 2523
rect 2893 2517 2947 2523
rect 3325 2517 3379 2523
rect 3405 2512 3411 2543
rect 3901 2512 3907 2543
rect 4020 2537 4044 2543
rect 4381 2537 4396 2543
rect 4504 2537 4524 2543
rect 4660 2537 4675 2543
rect 4989 2537 5020 2543
rect 5245 2537 5260 2543
rect 5325 2537 5379 2543
rect 4221 2517 4236 2523
rect 5316 2517 5340 2523
rect 5469 2517 5507 2523
rect 4429 2497 4467 2503
rect 5396 2496 5406 2504
rect 356 2477 371 2483
rect 3242 2476 3244 2484
rect 3300 2436 3302 2444
rect 4820 2436 4822 2444
rect 5508 2436 5510 2444
rect 1496 2406 1502 2414
rect 1510 2406 1516 2414
rect 1524 2406 1530 2414
rect 1538 2406 1544 2414
rect 4568 2406 4574 2414
rect 4582 2406 4588 2414
rect 4596 2406 4602 2414
rect 4610 2406 4616 2414
rect 228 2376 230 2384
rect 164 2336 166 2344
rect 788 2337 804 2343
rect 813 2337 828 2343
rect 300 2332 308 2336
rect 796 2332 804 2337
rect 3524 2337 3555 2343
rect 4628 2337 4668 2343
rect 5053 2337 5084 2343
rect 5316 2337 5331 2343
rect 340 2316 348 2324
rect 1268 2316 1276 2324
rect 1405 2317 1427 2323
rect 2980 2316 2988 2324
rect 3140 2316 3148 2324
rect 3453 2317 3468 2323
rect 4788 2317 4803 2323
rect 5165 2317 5180 2323
rect 5549 2317 5571 2323
rect 6052 2316 6060 2324
rect 5164 2304 5172 2308
rect 109 2297 140 2303
rect 1117 2297 1148 2303
rect 1277 2297 1292 2303
rect 1348 2297 1379 2303
rect 2660 2297 2691 2303
rect 2772 2297 2787 2303
rect 2884 2297 2915 2303
rect 2925 2297 2956 2303
rect 3124 2297 3139 2303
rect 4020 2297 4035 2303
rect 4685 2297 4700 2303
rect 5636 2297 5651 2303
rect 1309 2283 1315 2296
rect 1293 2277 1315 2283
rect 1341 2277 1356 2283
rect 1341 2257 1347 2277
rect 2701 2277 2739 2283
rect 2756 2277 2771 2283
rect 3645 2277 3660 2283
rect 4141 2277 4156 2283
rect 4308 2277 4323 2283
rect 4820 2277 4851 2283
rect 2252 2264 2260 2268
rect 292 2236 294 2244
rect 3032 2206 3038 2214
rect 3046 2206 3052 2214
rect 3060 2206 3066 2214
rect 3074 2206 3080 2214
rect 1720 2176 1724 2184
rect 5338 2176 5340 2184
rect 746 2156 748 2164
rect 1588 2157 1619 2163
rect 2468 2157 2483 2163
rect 2852 2157 2867 2163
rect 29 2137 51 2143
rect 157 2143 163 2156
rect 157 2137 179 2143
rect 541 2137 556 2143
rect 1229 2137 1244 2143
rect 1629 2137 1644 2143
rect 3485 2137 3500 2143
rect 4013 2137 4051 2143
rect 4093 2137 4108 2143
rect 4221 2137 4252 2143
rect 5924 2137 5939 2143
rect 100 2117 115 2123
rect 317 2117 348 2123
rect 1037 2117 1075 2123
rect 196 2096 204 2104
rect 1037 2097 1043 2117
rect 1165 2117 1203 2123
rect 1165 2097 1171 2117
rect 1220 2117 1260 2123
rect 1277 2117 1315 2123
rect 1309 2097 1315 2117
rect 4036 2117 4067 2123
rect 5245 2117 5276 2123
rect 5293 2117 5331 2123
rect 1332 2096 1340 2104
rect 3485 2097 3523 2103
rect 4093 2097 4108 2103
rect 5325 2097 5331 2117
rect 68 2036 70 2044
rect 378 2036 380 2044
rect 1496 2006 1502 2014
rect 1510 2006 1516 2014
rect 1524 2006 1530 2014
rect 1538 2006 1544 2014
rect 4568 2006 4574 2014
rect 4582 2006 4588 2014
rect 4596 2006 4602 2014
rect 4610 2006 4616 2014
rect 1172 1976 1174 1984
rect 1332 1976 1334 1984
rect 2428 1937 2444 1943
rect 3212 1937 3251 1943
rect 4886 1936 4892 1944
rect 5021 1937 5036 1943
rect 676 1916 684 1924
rect 1092 1916 1100 1924
rect 2900 1917 2915 1923
rect 5100 1912 5108 1916
rect 461 1897 476 1903
rect 596 1897 611 1903
rect 1220 1897 1251 1903
rect 1677 1897 1724 1903
rect 2964 1897 2979 1903
rect 5213 1897 5251 1903
rect 6036 1897 6051 1903
rect 724 1877 739 1883
rect 1716 1877 1746 1883
rect 2221 1877 2236 1883
rect 2429 1877 2451 1883
rect 2461 1877 2476 1883
rect 2500 1877 2515 1883
rect 3629 1877 3644 1883
rect 6077 1877 6124 1883
rect 1476 1857 1491 1863
rect 1572 1837 1587 1843
rect 3032 1806 3038 1814
rect 3046 1806 3052 1814
rect 3060 1806 3066 1814
rect 3074 1806 3080 1814
rect 1018 1776 1020 1784
rect 1930 1776 1932 1784
rect 5556 1776 5558 1784
rect 762 1756 764 1764
rect 1277 1757 1292 1763
rect 1437 1757 1452 1763
rect 3837 1757 3860 1763
rect 1261 1743 1267 1756
rect 3852 1754 3860 1757
rect 5220 1756 5222 1764
rect 6077 1757 6124 1763
rect 1245 1737 1267 1743
rect 1860 1737 1875 1743
rect 1997 1737 2019 1743
rect 2772 1737 2803 1743
rect 2957 1737 2972 1743
rect 3588 1737 3603 1743
rect 4180 1737 4195 1743
rect 4580 1737 4643 1743
rect 4749 1737 4764 1743
rect 5524 1737 5539 1743
rect 6045 1737 6067 1743
rect 77 1717 92 1723
rect 212 1717 227 1723
rect 461 1717 499 1723
rect 861 1717 899 1723
rect 836 1696 844 1704
rect 861 1697 867 1717
rect 957 1717 972 1723
rect 1981 1717 2012 1723
rect 3645 1717 3660 1723
rect 4077 1717 4115 1723
rect 4109 1697 4115 1717
rect 4180 1717 4195 1723
rect 4509 1717 4547 1723
rect 4557 1717 4636 1723
rect 4509 1697 4515 1717
rect 4644 1717 4659 1723
rect 4756 1717 4787 1723
rect 5101 1717 5139 1723
rect 4660 1696 4668 1704
rect 5101 1697 5107 1717
rect 5613 1717 5644 1723
rect 5460 1696 5468 1704
rect 5636 1697 5667 1703
rect 1085 1677 1100 1683
rect 3821 1677 3836 1683
rect 4900 1676 4906 1684
rect 458 1636 460 1644
rect 1496 1606 1502 1614
rect 1510 1606 1516 1614
rect 1524 1606 1530 1614
rect 1538 1606 1544 1614
rect 4568 1606 4574 1614
rect 4582 1606 4588 1614
rect 4596 1606 4602 1614
rect 4610 1606 4616 1614
rect 234 1576 236 1584
rect 1380 1576 1382 1584
rect 1512 1576 1516 1584
rect 3738 1576 3740 1584
rect 3802 1576 3804 1584
rect 1124 1536 1126 1544
rect 1933 1537 1972 1543
rect 2973 1537 2988 1543
rect 3588 1537 3604 1543
rect 5204 1536 5210 1544
rect 5460 1536 5466 1544
rect 5661 1537 5676 1543
rect 6093 1537 6124 1543
rect 237 1497 284 1503
rect 333 1503 339 1523
rect 301 1497 339 1503
rect 404 1497 419 1503
rect 653 1503 659 1523
rect 892 1517 915 1523
rect 892 1512 900 1517
rect 1316 1516 1324 1524
rect 3133 1517 3148 1523
rect 3860 1516 3868 1524
rect 621 1497 659 1503
rect 1284 1497 1299 1503
rect 253 1477 268 1483
rect 404 1477 419 1483
rect 1293 1477 1299 1497
rect 1997 1497 2012 1503
rect 2109 1497 2140 1503
rect 4157 1503 4163 1523
rect 4125 1497 4163 1503
rect 4189 1497 4227 1503
rect 1437 1477 1459 1483
rect 2013 1477 2051 1483
rect 2996 1477 3011 1483
rect 3021 1477 3084 1483
rect 538 1456 540 1464
rect 3021 1457 3027 1477
rect 3133 1477 3155 1483
rect 3556 1477 3571 1483
rect 3581 1477 3603 1483
rect 4221 1483 4227 1497
rect 4500 1497 4531 1503
rect 4973 1503 4979 1523
rect 4941 1497 4979 1503
rect 5085 1503 5091 1523
rect 5085 1497 5123 1503
rect 5389 1497 5404 1503
rect 5508 1497 5539 1503
rect 4221 1477 4243 1483
rect 4365 1477 4387 1483
rect 2154 1436 2156 1444
rect 2618 1436 2620 1444
rect 3032 1406 3038 1414
rect 3046 1406 3052 1414
rect 3060 1406 3066 1414
rect 3074 1406 3080 1414
rect 1236 1376 1238 1384
rect 4564 1376 4568 1384
rect 3533 1357 3548 1363
rect 900 1337 915 1343
rect 2036 1337 2051 1343
rect 2452 1337 2467 1343
rect 3725 1337 3747 1343
rect 3757 1337 3772 1343
rect 4717 1343 4723 1363
rect 4493 1337 4531 1343
rect 4621 1337 4723 1343
rect 4836 1337 4851 1343
rect 4957 1337 4979 1343
rect 381 1317 419 1323
rect 413 1297 419 1317
rect 605 1317 643 1323
rect 637 1297 643 1317
rect 1460 1317 1491 1323
rect 4340 1317 4355 1323
rect 4797 1317 4828 1323
rect 4957 1323 4963 1337
rect 5501 1337 5516 1343
rect 5757 1337 5779 1343
rect 4925 1317 4963 1323
rect 5661 1317 5676 1323
rect 5773 1323 5779 1337
rect 5773 1317 5811 1323
rect 5821 1317 5852 1323
rect 2100 1297 2115 1303
rect 2653 1297 2691 1303
rect 4452 1297 4467 1303
rect 4916 1296 4924 1304
rect 5421 1297 5443 1303
rect 5852 1284 5860 1288
rect 1485 1277 1532 1283
rect 3724 1277 3740 1283
rect 1428 1236 1430 1244
rect 2516 1236 2518 1244
rect 4314 1236 4316 1244
rect 1496 1206 1502 1214
rect 1510 1206 1516 1214
rect 1524 1206 1530 1214
rect 1538 1206 1544 1214
rect 4568 1206 4574 1214
rect 4582 1206 4588 1214
rect 4596 1206 4602 1214
rect 4610 1206 4616 1214
rect 1044 1176 1046 1184
rect 1562 1176 1564 1184
rect 4724 1137 4755 1143
rect 5676 1137 5715 1143
rect 5036 1132 5044 1136
rect 77 1097 92 1103
rect 404 1097 419 1103
rect 557 1103 563 1123
rect 980 1116 988 1124
rect 3117 1117 3155 1123
rect 4653 1117 4675 1123
rect 4989 1117 5027 1123
rect 5108 1116 5116 1124
rect 525 1097 563 1103
rect 589 1097 627 1103
rect 317 1077 348 1083
rect 621 1083 627 1097
rect 765 1097 780 1103
rect 1012 1097 1043 1103
rect 1117 1097 1171 1103
rect 1389 1097 1404 1103
rect 1428 1097 1443 1103
rect 1565 1097 1580 1103
rect 1901 1097 1923 1103
rect 1917 1084 1923 1097
rect 2317 1097 2332 1103
rect 3533 1097 3548 1103
rect 3613 1097 3667 1103
rect 4317 1097 4355 1103
rect 621 1077 643 1083
rect 1309 1077 1324 1083
rect 1924 1077 1939 1083
rect 2093 1077 2108 1083
rect 1325 1057 1331 1076
rect 1876 1056 1878 1064
rect 2093 1057 2099 1077
rect 2260 1077 2291 1083
rect 2852 1077 2883 1083
rect 4349 1083 4355 1097
rect 4429 1097 4444 1103
rect 4477 1097 4508 1103
rect 4692 1097 4707 1103
rect 4900 1097 4915 1103
rect 4932 1097 4963 1103
rect 5076 1097 5107 1103
rect 5156 1097 5171 1103
rect 5293 1103 5299 1123
rect 5293 1097 5331 1103
rect 5661 1097 5692 1103
rect 4349 1077 4371 1083
rect 4493 1077 4515 1083
rect 4724 1077 4739 1083
rect 5597 1077 5628 1083
rect 4076 1072 4084 1076
rect 2349 1057 2364 1063
rect 1290 1036 1292 1044
rect 3108 1036 3110 1044
rect 4644 1036 4646 1044
rect 4756 1036 4758 1044
rect 3032 1006 3038 1014
rect 3046 1006 3052 1014
rect 3060 1006 3066 1014
rect 3074 1006 3080 1014
rect 1434 976 1436 984
rect 4218 976 4220 984
rect 5428 976 5430 984
rect 5668 976 5670 984
rect 2445 957 2467 963
rect 2333 937 2348 943
rect 4061 937 4076 943
rect 4093 937 4115 943
rect 4541 937 4556 943
rect 4740 937 4755 943
rect 5124 937 5139 943
rect 5245 937 5267 943
rect 557 917 588 923
rect 813 917 867 923
rect 1268 917 1283 923
rect 1341 917 1356 923
rect 2205 917 2243 923
rect 292 896 300 904
rect 957 897 979 903
rect 1580 903 1588 908
rect 1517 897 1588 903
rect 2148 896 2156 904
rect 2237 897 2243 917
rect 2276 917 2291 923
rect 2365 917 2396 923
rect 3293 917 3330 923
rect 4461 917 4492 923
rect 4829 917 4844 923
rect 4916 917 4931 923
rect 5261 923 5267 937
rect 5261 917 5299 923
rect 5325 917 5363 923
rect 5325 897 5331 917
rect 5164 884 5172 888
rect 5436 884 5444 888
rect 234 836 236 844
rect 874 836 876 844
rect 1306 836 1308 844
rect 4404 836 4406 844
rect 4932 836 4934 844
rect 5716 836 5718 844
rect 1496 806 1502 814
rect 1510 806 1516 814
rect 1524 806 1530 814
rect 1538 806 1544 814
rect 4568 806 4574 814
rect 4582 806 4588 814
rect 4596 806 4602 814
rect 4610 806 4616 814
rect 660 776 662 784
rect 1866 776 1868 784
rect 3988 776 3992 784
rect 4420 776 4422 784
rect 4554 756 4556 764
rect 189 737 204 743
rect 794 736 796 744
rect 2365 737 2404 743
rect 2508 737 2524 743
rect 3908 736 3910 744
rect 4116 736 4118 744
rect 4260 737 4307 743
rect 5364 736 5366 744
rect 5588 736 5590 744
rect 5754 736 5756 744
rect 4300 724 4308 728
rect 93 703 99 723
rect 93 697 131 703
rect 365 703 371 723
rect 365 697 403 703
rect 765 703 771 723
rect 733 697 771 703
rect 893 697 924 703
rect 973 697 988 703
rect 1469 703 1475 723
rect 1389 697 1427 703
rect 1437 697 1475 703
rect 29 677 51 683
rect 205 677 220 683
rect 916 677 947 683
rect 1389 683 1395 697
rect 1837 703 1843 723
rect 2957 717 3043 723
rect 4180 716 4188 724
rect 1805 697 1843 703
rect 2388 697 2419 703
rect 2429 697 2476 703
rect 4045 697 4083 703
rect 1373 677 1395 683
rect 1517 677 1564 683
rect 2445 677 2460 683
rect 2509 677 2531 683
rect 2541 677 2572 683
rect 3421 677 3443 683
rect 3821 677 3843 683
rect 4045 677 4051 697
rect 4452 697 4483 703
rect 4557 697 4572 703
rect 4877 703 4883 723
rect 4877 697 4915 703
rect 5021 703 5027 723
rect 5044 716 5052 724
rect 5389 717 5427 723
rect 5444 717 5459 723
rect 4932 697 4979 703
rect 4989 697 5027 703
rect 5092 697 5107 703
rect 5492 697 5507 703
rect 5556 697 5587 703
rect 5620 697 5635 703
rect 4573 677 4588 683
rect 4948 677 4963 683
rect 5693 677 5708 683
rect 868 656 870 664
rect 1940 656 1942 664
rect 5460 656 5468 664
rect 2948 636 2950 644
rect 3476 636 3480 644
rect 3860 636 3862 644
rect 4234 636 4236 644
rect 3032 606 3038 614
rect 3046 606 3052 614
rect 3060 606 3066 614
rect 3074 606 3080 614
rect 442 576 444 584
rect 730 576 732 584
rect 4596 577 4643 583
rect 1434 556 1436 564
rect 3556 537 3571 543
rect 4285 537 4307 543
rect 4685 537 4707 543
rect 356 517 387 523
rect 701 517 716 523
rect 829 517 860 523
rect 1140 517 1155 523
rect 1220 517 1235 523
rect 1373 517 1388 523
rect 1581 517 1619 523
rect 1581 497 1587 517
rect 2301 517 2339 523
rect 2365 517 2403 523
rect 2333 497 2339 517
rect 2877 517 2892 523
rect 3316 517 3331 523
rect 3421 517 3459 523
rect 3469 517 3507 523
rect 2356 496 2364 504
rect 3453 497 3459 517
rect 4484 517 4515 523
rect 4573 517 4636 523
rect 5124 517 5148 523
rect 5197 517 5212 523
rect 5341 517 5379 523
rect 4388 496 4396 504
rect 5373 497 5379 517
rect 5524 517 5555 523
rect 428 484 436 488
rect 2244 477 2259 483
rect 5402 476 5404 484
rect 388 436 390 444
rect 804 436 806 444
rect 906 436 908 444
rect 1178 436 1180 444
rect 1268 436 1270 444
rect 2804 436 2806 444
rect 2874 436 2876 444
rect 1496 406 1502 414
rect 1510 406 1516 414
rect 1524 406 1530 414
rect 1538 406 1544 414
rect 4568 406 4574 414
rect 4582 406 4588 414
rect 4596 406 4602 414
rect 4610 406 4616 414
rect 3396 376 3400 384
rect 5434 336 5436 344
rect 6109 337 6124 343
rect 573 303 579 323
rect 852 316 860 324
rect 541 297 579 303
rect 877 303 883 323
rect 1172 316 1180 324
rect 877 297 915 303
rect 1197 303 1203 323
rect 1197 297 1235 303
rect 1325 303 1331 323
rect 1268 297 1299 303
rect 1325 297 1363 303
rect 1725 303 1731 323
rect 4333 317 4348 323
rect 4461 317 4476 323
rect 1661 297 1699 303
rect 1725 297 1763 303
rect 2141 297 2172 303
rect 2269 297 2307 303
rect 3156 297 3187 303
rect 3245 297 3260 303
rect 404 277 419 283
rect 461 277 483 283
rect 1580 277 1612 283
rect 1773 277 1810 283
rect 3245 277 3251 297
rect 3325 297 3363 303
rect 3357 284 3363 297
rect 4788 297 4803 303
rect 4829 303 4835 323
rect 4829 297 4867 303
rect 4877 297 4892 303
rect 5108 297 5123 303
rect 5149 303 5155 323
rect 5396 317 5411 323
rect 5149 297 5187 303
rect 5437 297 5484 303
rect 6068 297 6083 303
rect 4061 277 4076 283
rect 5460 277 5475 283
rect 5645 277 5667 283
rect 1636 257 1651 263
rect 2653 257 2691 263
rect 3108 257 3123 263
rect 3032 206 3038 214
rect 3046 206 3052 214
rect 3060 206 3066 214
rect 3074 206 3080 214
rect 4276 176 4278 184
rect 3469 157 3507 163
rect 3549 157 3564 163
rect 3604 157 3619 163
rect 4676 156 4678 164
rect 4778 156 4780 164
rect 6093 157 6108 163
rect 477 137 499 143
rect 1276 137 1292 143
rect 3492 137 3523 143
rect 3581 137 3596 143
rect 5357 137 5395 143
rect 397 117 435 123
rect 429 97 435 117
rect 765 117 780 123
rect 829 117 867 123
rect 829 97 835 117
rect 1389 117 1474 123
rect 2126 117 2156 123
rect 2526 117 2563 123
rect 3022 117 3100 123
rect 3549 117 3571 123
rect 4701 117 4732 123
rect 4877 117 4915 123
rect 4877 97 4883 117
rect 5156 117 5171 123
rect 5293 117 5331 123
rect 5293 97 5299 117
rect 1496 6 1502 14
rect 1510 6 1516 14
rect 1524 6 1530 14
rect 1538 6 1544 14
rect 4568 6 4574 14
rect 4582 6 4588 14
rect 4596 6 4602 14
rect 4610 6 4616 14
<< m2contact >>
rect 1502 5606 1510 5614
rect 1516 5606 1524 5614
rect 1530 5606 1538 5614
rect 4574 5606 4582 5614
rect 4588 5606 4596 5614
rect 4602 5606 4610 5614
rect 76 5576 84 5584
rect 396 5576 404 5584
rect 956 5576 964 5584
rect 1468 5576 1476 5584
rect 1788 5576 1796 5584
rect 1980 5576 1988 5584
rect 2060 5576 2068 5584
rect 2524 5576 2532 5584
rect 2604 5576 2612 5584
rect 2956 5576 2964 5584
rect 3324 5576 3332 5584
rect 3964 5558 3972 5566
rect 5852 5558 5860 5566
rect 6076 5556 6084 5564
rect 476 5536 484 5544
rect 1900 5536 1908 5544
rect 4060 5536 4068 5544
rect 4940 5536 4948 5544
rect 76 5516 84 5524
rect 572 5516 580 5524
rect 604 5516 612 5524
rect 636 5516 644 5524
rect 956 5516 964 5524
rect 1468 5516 1476 5524
rect 1868 5516 1876 5524
rect 1932 5516 1940 5524
rect 1964 5516 1972 5524
rect 2060 5516 2068 5524
rect 2508 5516 2516 5524
rect 2604 5516 2612 5524
rect 3324 5516 3332 5524
rect 60 5496 68 5504
rect 284 5496 292 5504
rect 444 5496 452 5504
rect 524 5496 532 5504
rect 604 5496 612 5504
rect 748 5496 756 5504
rect 956 5496 964 5504
rect 1052 5494 1060 5502
rect 1244 5494 1252 5502
rect 1452 5496 1460 5504
rect 1676 5496 1684 5504
rect 1836 5496 1844 5504
rect 1868 5496 1876 5504
rect 1900 5496 1908 5504
rect 2012 5496 2020 5504
rect 2044 5496 2052 5504
rect 2268 5496 2276 5504
rect 2444 5496 2452 5504
rect 2556 5496 2564 5504
rect 2620 5496 2628 5504
rect 3324 5496 3332 5504
rect 3420 5496 3428 5504
rect 3468 5516 3476 5524
rect 3612 5516 3620 5524
rect 3644 5516 3652 5524
rect 3964 5512 3972 5520
rect 3500 5496 3508 5504
rect 3580 5496 3588 5504
rect 3628 5496 3636 5504
rect 3644 5496 3652 5504
rect 3996 5496 4004 5504
rect 4252 5496 4260 5504
rect 4316 5494 4324 5502
rect 4396 5496 4404 5504
rect 4412 5496 4420 5504
rect 4444 5516 4452 5524
rect 4476 5496 4484 5504
rect 4684 5496 4692 5504
rect 4748 5494 4756 5502
rect 4828 5496 4836 5504
rect 4876 5516 4884 5524
rect 5180 5516 5188 5524
rect 5292 5516 5300 5524
rect 5324 5516 5332 5524
rect 5852 5512 5860 5520
rect 4908 5496 4916 5504
rect 5052 5496 5060 5504
rect 5148 5496 5156 5504
rect 5196 5496 5204 5504
rect 5212 5496 5220 5504
rect 5260 5496 5268 5504
rect 5324 5496 5332 5504
rect 5500 5496 5508 5504
rect 5884 5496 5892 5504
rect 28 5476 36 5484
rect 172 5476 180 5484
rect 444 5476 452 5484
rect 572 5476 580 5484
rect 588 5476 596 5484
rect 860 5476 868 5484
rect 1020 5476 1028 5484
rect 1116 5476 1124 5484
rect 1212 5476 1220 5484
rect 1564 5476 1572 5484
rect 1758 5476 1766 5484
rect 1932 5476 1940 5484
rect 2156 5476 2164 5484
rect 2412 5476 2420 5484
rect 2476 5476 2484 5484
rect 2700 5476 2708 5484
rect 3228 5476 3236 5484
rect 3436 5476 3444 5484
rect 3516 5476 3524 5484
rect 3628 5476 3636 5484
rect 3900 5476 3908 5484
rect 4172 5476 4180 5484
rect 4348 5476 4356 5484
rect 4380 5476 4388 5484
rect 4492 5476 4500 5484
rect 4572 5476 4580 5484
rect 4812 5476 4820 5484
rect 4860 5476 4868 5484
rect 4924 5476 4932 5484
rect 5100 5476 5108 5484
rect 5132 5476 5140 5484
rect 5180 5476 5188 5484
rect 5276 5476 5284 5484
rect 5340 5476 5348 5484
rect 5452 5476 5460 5484
rect 5548 5476 5556 5484
rect 5788 5476 5796 5484
rect 5932 5476 5940 5484
rect 5964 5476 5972 5484
rect 28 5456 36 5464
rect 204 5456 212 5464
rect 380 5456 388 5464
rect 508 5456 516 5464
rect 828 5456 836 5464
rect 1596 5456 1604 5464
rect 1836 5456 1844 5464
rect 2188 5456 2196 5464
rect 2380 5456 2388 5464
rect 2732 5456 2740 5464
rect 3004 5456 3012 5464
rect 3196 5456 3204 5464
rect 3372 5456 3380 5464
rect 3532 5456 3540 5464
rect 3868 5456 3876 5464
rect 4556 5456 4564 5464
rect 5356 5456 5364 5464
rect 5756 5456 5764 5464
rect 5948 5456 5956 5464
rect 460 5436 468 5444
rect 1180 5436 1188 5444
rect 1372 5436 1380 5444
rect 2892 5436 2900 5444
rect 3708 5436 3716 5444
rect 4188 5436 4196 5444
rect 4508 5436 4516 5444
rect 4588 5436 4596 5444
rect 5372 5436 5380 5444
rect 5388 5436 5396 5444
rect 5596 5436 5604 5444
rect 3038 5406 3046 5414
rect 3052 5406 3060 5414
rect 3066 5406 3074 5414
rect 332 5376 340 5384
rect 1036 5376 1044 5384
rect 1180 5376 1188 5384
rect 2076 5376 2084 5384
rect 2268 5376 2276 5384
rect 2924 5376 2932 5384
rect 5276 5376 5284 5384
rect 5340 5376 5348 5384
rect 5868 5376 5876 5384
rect 172 5356 180 5364
rect 428 5356 436 5364
rect 476 5356 484 5364
rect 812 5356 820 5364
rect 1580 5356 1588 5364
rect 1916 5356 1924 5364
rect 2428 5356 2436 5364
rect 2764 5356 2772 5364
rect 2956 5356 2964 5364
rect 3324 5356 3332 5364
rect 3500 5356 3508 5364
rect 3580 5356 3588 5364
rect 3724 5356 3732 5364
rect 3996 5356 4004 5364
rect 5436 5356 5444 5364
rect 5612 5356 5620 5364
rect 6076 5356 6084 5364
rect 140 5336 148 5344
rect 364 5336 372 5344
rect 412 5336 420 5344
rect 460 5336 468 5344
rect 556 5336 564 5344
rect 572 5336 580 5344
rect 844 5336 852 5344
rect 988 5336 996 5344
rect 1052 5336 1060 5344
rect 1084 5336 1092 5344
rect 1116 5336 1124 5344
rect 1244 5336 1252 5344
rect 1612 5336 1620 5344
rect 1884 5336 1892 5344
rect 2140 5336 2148 5344
rect 2172 5336 2180 5344
rect 2252 5336 2260 5344
rect 2460 5336 2468 5344
rect 2732 5336 2740 5344
rect 2988 5336 2996 5344
rect 3020 5336 3028 5344
rect 3100 5336 3108 5344
rect 3356 5336 3364 5344
rect 3580 5336 3588 5344
rect 3660 5336 3668 5344
rect 3820 5336 3828 5344
rect 4028 5336 4036 5344
rect 4172 5336 4180 5344
rect 4300 5336 4308 5344
rect 4508 5336 4516 5344
rect 4668 5336 4676 5344
rect 4716 5336 4724 5344
rect 4748 5336 4756 5344
rect 4780 5336 4788 5344
rect 4860 5336 4868 5344
rect 4876 5336 4884 5344
rect 4924 5336 4932 5344
rect 4988 5336 4996 5344
rect 5020 5336 5028 5344
rect 5228 5336 5236 5344
rect 5372 5336 5380 5344
rect 5644 5336 5652 5344
rect 5788 5336 5796 5344
rect 5980 5336 5988 5344
rect 60 5316 68 5324
rect 396 5316 404 5324
rect 524 5316 532 5324
rect 588 5316 596 5324
rect 940 5316 948 5324
rect 1004 5316 1012 5324
rect 1052 5316 1060 5324
rect 1132 5316 1140 5324
rect 76 5300 84 5308
rect 348 5296 356 5304
rect 428 5296 436 5304
rect 556 5296 564 5304
rect 588 5296 596 5304
rect 940 5296 948 5304
rect 1036 5296 1044 5304
rect 1100 5296 1108 5304
rect 1164 5296 1172 5304
rect 1228 5316 1236 5324
rect 1404 5316 1412 5324
rect 1676 5316 1684 5324
rect 1772 5316 1780 5324
rect 1996 5316 2004 5324
rect 1708 5296 1716 5304
rect 1820 5300 1828 5308
rect 2524 5316 2532 5324
rect 2636 5316 2644 5324
rect 3452 5316 3460 5324
rect 3532 5316 3540 5324
rect 3644 5316 3652 5324
rect 3724 5316 3732 5324
rect 3772 5316 3780 5324
rect 3916 5316 3924 5324
rect 4124 5316 4132 5324
rect 4380 5316 4388 5324
rect 4444 5318 4452 5326
rect 4524 5316 4532 5324
rect 2204 5296 2212 5304
rect 2556 5296 2564 5304
rect 2636 5296 2644 5304
rect 3132 5296 3140 5304
rect 3420 5300 3428 5308
rect 3500 5296 3508 5304
rect 3596 5296 3604 5304
rect 3708 5296 3716 5304
rect 3804 5296 3812 5304
rect 4092 5300 4100 5308
rect 4652 5316 4660 5324
rect 4668 5316 4676 5324
rect 4732 5316 4740 5324
rect 4620 5296 4628 5304
rect 4844 5316 4852 5324
rect 4892 5316 4900 5324
rect 4812 5296 4820 5304
rect 4972 5316 4980 5324
rect 5052 5318 5060 5326
rect 5228 5316 5236 5324
rect 5308 5316 5316 5324
rect 5388 5316 5396 5324
rect 5724 5316 5732 5324
rect 5804 5316 5812 5324
rect 5820 5316 5828 5324
rect 5980 5316 5988 5324
rect 6028 5316 6036 5324
rect 4940 5296 4948 5304
rect 5196 5296 5204 5304
rect 5436 5296 5444 5304
rect 5740 5296 5748 5304
rect 5996 5296 6004 5304
rect 3836 5276 3844 5284
rect 4524 5276 4532 5284
rect 5180 5276 5188 5284
rect 5836 5276 5844 5284
rect 3420 5254 3428 5262
rect 76 5236 84 5244
rect 652 5236 660 5244
rect 940 5236 948 5244
rect 1420 5236 1428 5244
rect 1708 5236 1716 5244
rect 1820 5236 1828 5244
rect 2268 5236 2276 5244
rect 2556 5236 2564 5244
rect 2636 5236 2644 5244
rect 3164 5236 3172 5244
rect 4092 5236 4100 5244
rect 4316 5236 4324 5244
rect 5212 5236 5220 5244
rect 5452 5236 5460 5244
rect 5740 5236 5748 5244
rect 1502 5206 1510 5214
rect 1516 5206 1524 5214
rect 1530 5206 1538 5214
rect 4574 5206 4582 5214
rect 4588 5206 4596 5214
rect 4602 5206 4610 5214
rect 1228 5176 1236 5184
rect 1324 5176 1332 5184
rect 2028 5176 2036 5184
rect 2428 5176 2436 5184
rect 2812 5176 2820 5184
rect 2876 5176 2884 5184
rect 4060 5176 4068 5184
rect 4172 5176 4180 5184
rect 4524 5176 4532 5184
rect 4748 5176 4756 5184
rect 4892 5176 4900 5184
rect 5756 5176 5764 5184
rect 2556 5158 2564 5166
rect 6012 5158 6020 5166
rect 1532 5136 1540 5144
rect 2332 5136 2340 5144
rect 3180 5136 3188 5144
rect 3292 5136 3300 5144
rect 3564 5136 3572 5144
rect 3724 5136 3732 5144
rect 3756 5136 3764 5144
rect 3932 5136 3940 5144
rect 4828 5136 4836 5144
rect 5036 5136 5044 5144
rect 5452 5136 5460 5144
rect 444 5116 452 5124
rect 556 5116 564 5124
rect 668 5116 676 5124
rect 60 5094 68 5102
rect 124 5096 132 5104
rect 268 5096 276 5104
rect 412 5096 420 5104
rect 428 5096 436 5104
rect 460 5096 468 5104
rect 476 5096 484 5104
rect 524 5096 532 5104
rect 540 5096 548 5104
rect 604 5096 612 5104
rect 716 5116 724 5124
rect 2028 5116 2036 5124
rect 2444 5116 2452 5124
rect 2556 5112 2564 5120
rect 2876 5116 2884 5124
rect 3916 5116 3924 5124
rect 3980 5116 3988 5124
rect 4284 5116 4292 5124
rect 4364 5116 4372 5124
rect 4652 5116 4660 5124
rect 5164 5116 5172 5124
rect 5180 5116 5188 5124
rect 5260 5116 5268 5124
rect 5356 5116 5364 5124
rect 5420 5116 5428 5124
rect 5484 5116 5492 5124
rect 5692 5116 5700 5124
rect 6012 5112 6020 5120
rect 716 5096 724 5104
rect 796 5094 804 5102
rect 860 5096 868 5104
rect 1004 5096 1012 5104
rect 1052 5096 1060 5104
rect 1212 5096 1220 5104
rect 1260 5096 1268 5104
rect 1276 5096 1284 5104
rect 1308 5096 1316 5104
rect 1372 5096 1380 5104
rect 1420 5096 1428 5104
rect 1708 5096 1716 5104
rect 1724 5096 1732 5104
rect 2044 5096 2052 5104
rect 2236 5096 2244 5104
rect 2364 5096 2372 5104
rect 2380 5096 2388 5104
rect 2540 5096 2548 5104
rect 2620 5096 2628 5104
rect 2876 5096 2884 5104
rect 3166 5096 3174 5104
rect 3388 5094 3396 5102
rect 3644 5096 3652 5104
rect 3676 5096 3684 5104
rect 3772 5096 3780 5104
rect 3788 5096 3796 5104
rect 3836 5096 3844 5104
rect 220 5076 228 5084
rect 396 5076 404 5084
rect 620 5076 628 5084
rect 732 5076 740 5084
rect 1644 5076 1652 5084
rect 1740 5076 1748 5084
rect 1836 5076 1844 5084
rect 1852 5076 1860 5084
rect 2124 5076 2132 5084
rect 2396 5076 2404 5084
rect 2412 5076 2420 5084
rect 2476 5076 2484 5084
rect 2620 5076 2628 5084
rect 2972 5076 2980 5084
rect 3276 5076 3284 5084
rect 3324 5076 3332 5084
rect 3356 5076 3364 5084
rect 3532 5076 3540 5084
rect 3900 5096 3908 5104
rect 3964 5096 3972 5104
rect 4028 5096 4036 5104
rect 4092 5096 4100 5104
rect 4156 5096 4164 5104
rect 4204 5096 4212 5104
rect 4220 5096 4228 5104
rect 4252 5096 4260 5104
rect 4348 5096 4356 5104
rect 4412 5096 4420 5104
rect 4476 5096 4484 5104
rect 4540 5096 4548 5104
rect 4556 5096 4564 5104
rect 4700 5096 4708 5104
rect 4716 5096 4724 5104
rect 4764 5096 4772 5104
rect 4860 5096 4868 5104
rect 4908 5096 4916 5104
rect 4940 5096 4948 5104
rect 4988 5096 4996 5104
rect 5052 5096 5060 5104
rect 5100 5096 5108 5104
rect 5212 5096 5220 5104
rect 5228 5096 5236 5104
rect 5276 5096 5284 5104
rect 5292 5096 5300 5104
rect 5388 5096 5396 5104
rect 5436 5096 5444 5104
rect 5452 5096 5460 5104
rect 5612 5096 5620 5104
rect 5836 5096 5844 5104
rect 6044 5096 6052 5104
rect 3868 5076 3876 5084
rect 3964 5076 3972 5084
rect 4140 5076 4148 5084
rect 4236 5076 4244 5084
rect 4364 5076 4372 5084
rect 4396 5076 4404 5084
rect 4684 5076 4692 5084
rect 4796 5076 4804 5084
rect 5004 5076 5012 5084
rect 5116 5076 5124 5084
rect 5292 5076 5300 5084
rect 5372 5076 5380 5084
rect 5436 5076 5444 5084
rect 5660 5076 5668 5084
rect 5724 5076 5732 5084
rect 5948 5076 5956 5084
rect 252 5056 260 5064
rect 492 5056 500 5064
rect 1148 5056 1156 5064
rect 1164 5056 1172 5064
rect 1388 5056 1396 5064
rect 1420 5056 1428 5064
rect 1660 5056 1668 5064
rect 1676 5056 1684 5064
rect 1692 5056 1700 5064
rect 2156 5056 2164 5064
rect 2460 5056 2468 5064
rect 2652 5056 2660 5064
rect 3004 5056 3012 5064
rect 4108 5056 4116 5064
rect 4636 5056 4644 5064
rect 5196 5056 5204 5064
rect 5356 5056 5364 5064
rect 5916 5056 5924 5064
rect 188 5036 196 5044
rect 380 5036 388 5044
rect 924 5036 932 5044
rect 1116 5036 1124 5044
rect 1132 5036 1140 5044
rect 1180 5036 1188 5044
rect 1404 5036 1412 5044
rect 1500 5036 1508 5044
rect 1772 5036 1780 5044
rect 1964 5036 1972 5044
rect 2316 5036 2324 5044
rect 2812 5036 2820 5044
rect 3196 5036 3204 5044
rect 3308 5036 3316 5044
rect 3516 5036 3524 5044
rect 3548 5036 3556 5044
rect 3932 5036 3940 5044
rect 4284 5036 4292 5044
rect 4316 5036 4324 5044
rect 4444 5036 4452 5044
rect 4572 5036 4580 5044
rect 4652 5036 4660 5044
rect 4812 5036 4820 5044
rect 4956 5036 4964 5044
rect 5036 5036 5044 5044
rect 5084 5036 5092 5044
rect 5164 5036 5172 5044
rect 5708 5036 5716 5044
rect 3038 5006 3046 5014
rect 3052 5006 3060 5014
rect 3066 5006 3074 5014
rect 12 4976 20 4984
rect 412 4976 420 4984
rect 940 4976 948 4984
rect 1308 4976 1316 4984
rect 2476 4976 2484 4984
rect 2892 4976 2900 4984
rect 3292 4976 3300 4984
rect 4044 4976 4052 4984
rect 4348 4976 4356 4984
rect 5788 4976 5796 4984
rect 844 4956 852 4964
rect 1468 4956 1476 4964
rect 1740 4956 1748 4964
rect 1916 4956 1924 4964
rect 2268 4956 2276 4964
rect 2956 4956 2964 4964
rect 3196 4956 3204 4964
rect 3308 4956 3316 4964
rect 3932 4956 3940 4964
rect 4476 4956 4484 4964
rect 4716 4956 4724 4964
rect 4908 4956 4916 4964
rect 5116 4956 5124 4964
rect 5324 4956 5332 4964
rect 5436 4956 5444 4964
rect 5948 4956 5956 4964
rect 60 4936 68 4944
rect 172 4936 180 4944
rect 220 4936 228 4944
rect 252 4936 260 4944
rect 428 4936 436 4944
rect 492 4936 500 4944
rect 636 4936 644 4944
rect 716 4936 724 4944
rect 748 4936 756 4944
rect 796 4936 804 4944
rect 876 4936 884 4944
rect 988 4936 996 4944
rect 1052 4936 1060 4944
rect 1180 4936 1188 4944
rect 1196 4936 1204 4944
rect 1276 4936 1284 4944
rect 1500 4936 1508 4944
rect 1948 4936 1956 4944
rect 2300 4936 2308 4944
rect 2508 4936 2516 4944
rect 2636 4936 2644 4944
rect 2652 4936 2660 4944
rect 2780 4936 2788 4944
rect 2812 4936 2820 4944
rect 2844 4936 2852 4944
rect 2860 4936 2868 4944
rect 2908 4936 2916 4944
rect 2972 4936 2980 4944
rect 3244 4936 3252 4944
rect 3404 4936 3412 4944
rect 3468 4936 3476 4944
rect 3580 4936 3588 4944
rect 3692 4936 3700 4944
rect 3996 4936 4004 4944
rect 4108 4936 4116 4944
rect 4188 4936 4196 4944
rect 4412 4936 4420 4944
rect 4524 4936 4532 4944
rect 4540 4936 4548 4944
rect 4652 4936 4660 4944
rect 4764 4936 4772 4944
rect 92 4916 100 4924
rect 140 4916 148 4924
rect 156 4916 164 4924
rect 204 4916 212 4924
rect 300 4916 308 4924
rect 444 4916 452 4924
rect 460 4916 468 4924
rect 492 4916 500 4924
rect 556 4916 564 4924
rect 572 4916 580 4924
rect 588 4916 596 4924
rect 620 4916 628 4924
rect 652 4916 660 4924
rect 668 4916 676 4924
rect 716 4916 724 4924
rect 796 4916 804 4924
rect 892 4916 900 4924
rect 12 4896 20 4904
rect 172 4896 180 4904
rect 476 4896 484 4904
rect 588 4896 596 4904
rect 780 4896 788 4904
rect 828 4896 836 4904
rect 924 4896 932 4904
rect 988 4916 996 4924
rect 1036 4916 1044 4924
rect 1084 4916 1092 4924
rect 1164 4916 1172 4924
rect 1004 4896 1012 4904
rect 1068 4896 1076 4904
rect 1132 4896 1140 4904
rect 1244 4916 1252 4924
rect 1596 4916 1604 4924
rect 1692 4916 1700 4924
rect 1836 4916 1844 4924
rect 2044 4916 2052 4924
rect 2380 4916 2388 4924
rect 2444 4916 2452 4924
rect 2828 4916 2836 4924
rect 2924 4916 2932 4924
rect 2988 4916 2996 4924
rect 3100 4916 3108 4924
rect 3116 4916 3124 4924
rect 3148 4916 3156 4924
rect 3180 4916 3188 4924
rect 3228 4916 3236 4924
rect 3260 4916 3268 4924
rect 3324 4916 3332 4924
rect 3340 4916 3348 4924
rect 3356 4916 3364 4924
rect 3452 4916 3460 4924
rect 3484 4916 3492 4924
rect 3516 4916 3524 4924
rect 3548 4916 3556 4924
rect 3564 4916 3572 4924
rect 3596 4916 3604 4924
rect 1596 4896 1604 4904
rect 2044 4896 2052 4904
rect 2396 4896 2404 4904
rect 2796 4896 2804 4904
rect 2892 4896 2900 4904
rect 2956 4896 2964 4904
rect 3020 4896 3028 4904
rect 3292 4896 3300 4904
rect 3420 4896 3428 4904
rect 3676 4916 3684 4924
rect 3708 4916 3716 4924
rect 3740 4916 3748 4924
rect 3772 4916 3780 4924
rect 3788 4916 3796 4924
rect 3916 4916 3924 4924
rect 4012 4916 4020 4924
rect 3644 4896 3652 4904
rect 4092 4916 4100 4924
rect 4204 4916 4212 4924
rect 4332 4916 4340 4924
rect 4380 4916 4388 4924
rect 4396 4916 4404 4924
rect 4428 4916 4436 4924
rect 4060 4896 4068 4904
rect 4460 4896 4468 4904
rect 4524 4916 4532 4924
rect 4540 4916 4548 4924
rect 4668 4916 4676 4924
rect 4636 4896 4644 4904
rect 4700 4896 4708 4904
rect 4748 4916 4756 4924
rect 4892 4916 4900 4924
rect 4972 4916 4980 4924
rect 4988 4916 4996 4924
rect 5036 4916 5044 4924
rect 5068 4936 5076 4944
rect 5180 4936 5188 4944
rect 5388 4936 5396 4944
rect 5452 4936 5460 4944
rect 5676 4936 5684 4944
rect 5756 4936 5764 4944
rect 5980 4936 5988 4944
rect 5164 4916 5172 4924
rect 5292 4916 5300 4924
rect 5404 4916 5412 4924
rect 5468 4916 5476 4924
rect 5628 4916 5636 4924
rect 5724 4916 5732 4924
rect 5740 4916 5748 4924
rect 6060 4916 6068 4924
rect 5132 4896 5140 4904
rect 5228 4896 5236 4904
rect 5436 4896 5444 4904
rect 5468 4896 5476 4904
rect 5708 4896 5716 4904
rect 6044 4900 6052 4908
rect 380 4876 388 4884
rect 812 4876 820 4884
rect 1100 4876 1108 4884
rect 2092 4876 2100 4884
rect 3452 4876 3460 4884
rect 3804 4876 3812 4884
rect 4300 4876 4308 4884
rect 5196 4876 5204 4884
rect 1036 4856 1044 4864
rect 6044 4854 6052 4862
rect 860 4836 868 4844
rect 1116 4836 1124 4844
rect 1164 4836 1172 4844
rect 1212 4836 1220 4844
rect 1596 4836 1604 4844
rect 1708 4836 1716 4844
rect 1756 4836 1764 4844
rect 2044 4836 2052 4844
rect 2396 4836 2404 4844
rect 2524 4836 2532 4844
rect 2988 4836 2996 4844
rect 3596 4836 3604 4844
rect 4556 4836 4564 4844
rect 4780 4836 4788 4844
rect 5516 4836 5524 4844
rect 5788 4836 5796 4844
rect 1502 4806 1510 4814
rect 1516 4806 1524 4814
rect 1530 4806 1538 4814
rect 4574 4806 4582 4814
rect 4588 4806 4596 4814
rect 4602 4806 4610 4814
rect 908 4776 916 4784
rect 988 4776 996 4784
rect 2140 4776 2148 4784
rect 2300 4776 2308 4784
rect 3004 4776 3012 4784
rect 3372 4776 3380 4784
rect 4476 4776 4484 4784
rect 4892 4776 4900 4784
rect 5068 4776 5076 4784
rect 5116 4776 5124 4784
rect 5164 4776 5172 4784
rect 5244 4776 5252 4784
rect 6092 4776 6100 4784
rect 508 4756 516 4764
rect 1244 4756 1252 4764
rect 2668 4756 2676 4764
rect 3548 4756 3556 4764
rect 3852 4756 3860 4764
rect 188 4736 196 4744
rect 748 4736 756 4744
rect 1180 4736 1188 4744
rect 1196 4736 1204 4744
rect 1356 4736 1364 4744
rect 1852 4736 1860 4744
rect 2364 4736 2372 4744
rect 3276 4736 3284 4744
rect 3612 4736 3620 4744
rect 76 4696 84 4704
rect 124 4696 132 4704
rect 220 4696 228 4704
rect 236 4696 244 4704
rect 268 4716 276 4724
rect 572 4716 580 4724
rect 300 4696 308 4704
rect 396 4696 404 4704
rect 540 4696 548 4704
rect 1148 4716 1156 4724
rect 1212 4716 1220 4724
rect 1276 4716 1284 4724
rect 1308 4716 1316 4724
rect 1388 4716 1396 4724
rect 1500 4716 1508 4724
rect 1772 4716 1780 4724
rect 1836 4716 1844 4724
rect 620 4696 628 4704
rect 652 4696 660 4704
rect 716 4696 724 4704
rect 732 4696 740 4704
rect 812 4696 820 4704
rect 860 4696 868 4704
rect 876 4696 884 4704
rect 940 4696 948 4704
rect 956 4696 964 4704
rect 1020 4696 1028 4704
rect 1036 4696 1044 4704
rect 1116 4696 1124 4704
rect 1132 4696 1140 4704
rect 1164 4696 1172 4704
rect 1276 4696 1284 4704
rect 1308 4696 1316 4704
rect 1356 4696 1364 4704
rect 1436 4696 1444 4704
rect 1468 4696 1476 4704
rect 1548 4696 1556 4704
rect 1644 4696 1652 4704
rect 1660 4696 1668 4704
rect 1692 4696 1700 4704
rect 1708 4696 1716 4704
rect 1724 4696 1732 4704
rect 1804 4696 1812 4704
rect 1820 4696 1828 4704
rect 1964 4696 1972 4704
rect 2108 4716 2116 4724
rect 2140 4696 2148 4704
rect 2188 4716 2196 4724
rect 2508 4716 2516 4724
rect 2572 4716 2580 4724
rect 2924 4716 2932 4724
rect 3292 4716 3300 4724
rect 3500 4716 3508 4724
rect 2220 4696 2228 4704
rect 2396 4696 2404 4704
rect 2412 4696 2420 4704
rect 2476 4696 2484 4704
rect 2668 4696 2676 4704
rect 2940 4696 2948 4704
rect 3036 4696 3044 4704
rect 3164 4696 3172 4704
rect 3308 4696 3316 4704
rect 3324 4696 3332 4704
rect 3340 4696 3348 4704
rect 3468 4696 3476 4704
rect 3932 4716 3940 4724
rect 4268 4716 4276 4724
rect 4300 4716 4308 4724
rect 3548 4696 3556 4704
rect 3564 4696 3572 4704
rect 3644 4696 3652 4704
rect 3660 4696 3668 4704
rect 3740 4696 3748 4704
rect 3916 4696 3924 4704
rect 3964 4696 3972 4704
rect 4092 4696 4100 4704
rect 4332 4696 4340 4704
rect 4348 4696 4356 4704
rect 4380 4716 4388 4724
rect 4716 4716 4724 4724
rect 4780 4716 4788 4724
rect 4812 4716 4820 4724
rect 5036 4716 5044 4724
rect 5084 4716 5092 4724
rect 5532 4716 5540 4724
rect 6092 4716 6100 4724
rect 4412 4696 4420 4704
rect 4444 4696 4452 4704
rect 4460 4696 4468 4704
rect 4604 4696 4612 4704
rect 4652 4696 4660 4704
rect 4668 4696 4676 4704
rect 4748 4696 4756 4704
rect 4844 4696 4852 4704
rect 4860 4696 4868 4704
rect 4876 4696 4884 4704
rect 4956 4696 4964 4704
rect 5004 4696 5012 4704
rect 5020 4696 5028 4704
rect 5180 4696 5188 4704
rect 5196 4696 5204 4704
rect 5212 4696 5220 4704
rect 5260 4696 5268 4704
rect 5292 4696 5300 4704
rect 5308 4696 5316 4704
rect 5484 4696 5492 4704
rect 5788 4696 5796 4704
rect 5884 4696 5892 4704
rect 204 4676 212 4684
rect 316 4676 324 4684
rect 380 4676 388 4684
rect 524 4676 532 4684
rect 588 4676 596 4684
rect 636 4676 644 4684
rect 780 4676 788 4684
rect 796 4676 804 4684
rect 1260 4676 1268 4684
rect 1324 4676 1332 4684
rect 1340 4676 1348 4684
rect 1452 4676 1460 4684
rect 1628 4676 1636 4684
rect 1724 4676 1732 4684
rect 1772 4676 1780 4684
rect 1788 4676 1796 4684
rect 2012 4676 2020 4684
rect 2044 4676 2052 4684
rect 2092 4676 2100 4684
rect 2124 4676 2132 4684
rect 2236 4676 2244 4684
rect 2348 4676 2356 4684
rect 2412 4676 2420 4684
rect 2428 4676 2436 4684
rect 2668 4676 2676 4684
rect 2892 4676 2900 4684
rect 3356 4676 3364 4684
rect 1116 4656 1124 4664
rect 1404 4656 1412 4664
rect 1532 4656 1540 4664
rect 2460 4656 2468 4664
rect 2700 4656 2708 4664
rect 2972 4656 2980 4664
rect 3148 4656 3156 4664
rect 3452 4676 3460 4684
rect 3580 4676 3588 4684
rect 3724 4676 3732 4684
rect 3980 4676 3988 4684
rect 4044 4676 4052 4684
rect 4220 4676 4228 4684
rect 4252 4676 4260 4684
rect 4316 4676 4324 4684
rect 4428 4676 4436 4684
rect 4524 4676 4532 4684
rect 4684 4676 4692 4684
rect 4732 4676 4740 4684
rect 4988 4676 4996 4684
rect 5052 4676 5060 4684
rect 5564 4676 5572 4684
rect 5660 4676 5668 4684
rect 5676 4676 5684 4684
rect 5772 4676 5780 4684
rect 5996 4676 6004 4684
rect 3996 4656 4004 4664
rect 4956 4656 4964 4664
rect 5148 4656 5156 4664
rect 5356 4656 5364 4664
rect 5548 4656 5556 4664
rect 5964 4656 5972 4664
rect 684 4636 692 4644
rect 748 4636 756 4644
rect 1068 4636 1076 4644
rect 1420 4636 1428 4644
rect 2060 4636 2068 4644
rect 2364 4636 2372 4644
rect 2860 4636 2868 4644
rect 2924 4636 2932 4644
rect 2956 4636 2964 4644
rect 3404 4636 3412 4644
rect 3884 4636 3892 4644
rect 3932 4636 3940 4644
rect 4012 4636 4020 4644
rect 4204 4636 4212 4644
rect 4236 4636 4244 4644
rect 4300 4636 4308 4644
rect 4700 4636 4708 4644
rect 4780 4636 4788 4644
rect 4972 4636 4980 4644
rect 5436 4636 5444 4644
rect 5628 4636 5636 4644
rect 3038 4606 3046 4614
rect 3052 4606 3060 4614
rect 3066 4606 3074 4614
rect 380 4576 388 4584
rect 412 4576 420 4584
rect 956 4576 964 4584
rect 1308 4576 1316 4584
rect 1500 4576 1508 4584
rect 1772 4576 1780 4584
rect 2076 4576 2084 4584
rect 2252 4576 2260 4584
rect 2892 4576 2900 4584
rect 5068 4576 5076 4584
rect 5404 4576 5412 4584
rect 364 4556 372 4564
rect 1052 4556 1060 4564
rect 1292 4556 1300 4564
rect 2028 4556 2036 4564
rect 2220 4556 2228 4564
rect 2540 4556 2548 4564
rect 2764 4556 2772 4564
rect 2812 4556 2820 4564
rect 3132 4556 3140 4564
rect 3436 4556 3444 4564
rect 3500 4556 3508 4564
rect 3692 4556 3700 4564
rect 4108 4556 4116 4564
rect 4556 4556 4564 4564
rect 4860 4556 4868 4564
rect 5084 4556 5092 4564
rect 5228 4556 5236 4564
rect 5564 4556 5572 4564
rect 5916 4556 5924 4564
rect 172 4536 180 4544
rect 204 4536 212 4544
rect 268 4536 276 4544
rect 476 4536 484 4544
rect 508 4536 516 4544
rect 540 4536 548 4544
rect 796 4536 804 4544
rect 812 4536 820 4544
rect 1004 4536 1012 4544
rect 1324 4536 1332 4544
rect 1452 4536 1460 4544
rect 1708 4536 1716 4544
rect 1740 4536 1748 4544
rect 1932 4536 1940 4544
rect 2092 4536 2100 4544
rect 2108 4536 2116 4544
rect 2284 4536 2292 4544
rect 2572 4536 2580 4544
rect 2748 4536 2756 4544
rect 3164 4536 3172 4544
rect 3580 4536 3588 4544
rect 3820 4536 3828 4544
rect 3836 4536 3844 4544
rect 3900 4536 3908 4544
rect 3980 4536 3988 4544
rect 4156 4536 4164 4544
rect 4220 4536 4228 4544
rect 4284 4536 4292 4544
rect 4300 4536 4308 4544
rect 4364 4536 4372 4544
rect 4396 4536 4404 4544
rect 4700 4536 4708 4544
rect 4764 4536 4772 4544
rect 4812 4536 4820 4544
rect 4940 4536 4948 4544
rect 4972 4536 4980 4544
rect 4988 4536 4996 4544
rect 5052 4536 5060 4544
rect 5308 4536 5316 4544
rect 5596 4536 5604 4544
rect 5948 4536 5956 4544
rect 140 4518 148 4526
rect 220 4516 228 4524
rect 236 4516 244 4524
rect 284 4516 292 4524
rect 332 4516 340 4524
rect 348 4516 356 4524
rect 444 4516 452 4524
rect 492 4516 500 4524
rect 588 4516 596 4524
rect 716 4516 724 4524
rect 732 4516 740 4524
rect 796 4516 804 4524
rect 828 4516 836 4524
rect 252 4496 260 4504
rect 460 4496 468 4504
rect 828 4496 836 4504
rect 908 4516 916 4524
rect 988 4516 996 4524
rect 1004 4516 1012 4524
rect 1084 4516 1092 4524
rect 1148 4516 1156 4524
rect 1212 4516 1220 4524
rect 1260 4516 1268 4524
rect 1276 4516 1284 4524
rect 1340 4516 1348 4524
rect 876 4496 884 4504
rect 1052 4496 1060 4504
rect 1068 4496 1076 4504
rect 1132 4496 1140 4504
rect 1388 4516 1396 4524
rect 1404 4516 1412 4524
rect 1564 4516 1572 4524
rect 1612 4516 1620 4524
rect 1628 4516 1636 4524
rect 1676 4516 1684 4524
rect 1724 4516 1732 4524
rect 1884 4516 1892 4524
rect 1980 4516 1988 4524
rect 2300 4516 2308 4524
rect 2460 4516 2468 4524
rect 2780 4516 2788 4524
rect 2860 4516 2868 4524
rect 3052 4516 3060 4524
rect 3436 4518 3444 4526
rect 3532 4516 3540 4524
rect 3612 4516 3620 4524
rect 3628 4516 3636 4524
rect 3660 4516 3668 4524
rect 3676 4516 3684 4524
rect 3724 4516 3732 4524
rect 3756 4516 3764 4524
rect 3772 4516 3780 4524
rect 3852 4516 3860 4524
rect 3868 4516 3876 4524
rect 3996 4516 4004 4524
rect 4140 4516 4148 4524
rect 4204 4516 4212 4524
rect 4268 4516 4276 4524
rect 4316 4516 4324 4524
rect 4380 4516 4388 4524
rect 4444 4516 4452 4524
rect 4508 4516 4516 4524
rect 4636 4516 4644 4524
rect 4716 4516 4724 4524
rect 1436 4496 1444 4504
rect 1484 4496 1492 4504
rect 1692 4496 1700 4504
rect 1756 4496 1764 4504
rect 1964 4496 1972 4504
rect 2252 4496 2260 4504
rect 2668 4496 2676 4504
rect 3260 4496 3268 4504
rect 3644 4496 3652 4504
rect 3900 4496 3908 4504
rect 4108 4496 4116 4504
rect 4172 4496 4180 4504
rect 4236 4496 4244 4504
rect 4348 4496 4356 4504
rect 4412 4496 4420 4504
rect 4444 4496 4452 4504
rect 4492 4496 4500 4504
rect 4684 4496 4692 4504
rect 4748 4496 4756 4504
rect 4796 4516 4804 4524
rect 4828 4516 4836 4524
rect 4844 4516 4852 4524
rect 4892 4516 4900 4524
rect 4956 4516 4964 4524
rect 5004 4516 5012 4524
rect 5052 4516 5060 4524
rect 5132 4516 5140 4524
rect 5180 4516 5188 4524
rect 5196 4516 5204 4524
rect 5292 4516 5300 4524
rect 5324 4516 5332 4524
rect 5596 4516 5604 4524
rect 5836 4516 5844 4524
rect 4924 4496 4932 4504
rect 5036 4496 5044 4504
rect 5148 4496 5156 4504
rect 5164 4496 5172 4504
rect 5260 4496 5268 4504
rect 5692 4496 5700 4504
rect 6012 4500 6020 4508
rect 700 4476 708 4484
rect 1100 4476 1108 4484
rect 1148 4476 1156 4484
rect 1164 4476 1172 4484
rect 1660 4476 1668 4484
rect 1996 4476 2004 4484
rect 3308 4476 3316 4484
rect 3516 4476 3524 4484
rect 4460 4476 4468 4484
rect 4524 4476 4532 4484
rect 5116 4476 5124 4484
rect 5132 4456 5140 4464
rect 6012 4454 6020 4462
rect 12 4436 20 4444
rect 1180 4436 1188 4444
rect 1228 4436 1236 4444
rect 1404 4436 1412 4444
rect 1580 4436 1588 4444
rect 1676 4436 1684 4444
rect 1772 4436 1780 4444
rect 2012 4436 2020 4444
rect 2332 4436 2340 4444
rect 2380 4436 2388 4444
rect 2668 4436 2676 4444
rect 2716 4436 2724 4444
rect 2812 4436 2820 4444
rect 2972 4436 2980 4444
rect 3260 4436 3268 4444
rect 4092 4436 4100 4444
rect 4204 4436 4212 4444
rect 4268 4436 4276 4444
rect 4316 4436 4324 4444
rect 4444 4436 4452 4444
rect 4508 4436 4516 4444
rect 4652 4436 4660 4444
rect 5292 4436 5300 4444
rect 5356 4436 5364 4444
rect 5692 4436 5700 4444
rect 5756 4436 5764 4444
rect 1502 4406 1510 4414
rect 1516 4406 1524 4414
rect 1530 4406 1538 4414
rect 4574 4406 4582 4414
rect 4588 4406 4596 4414
rect 4602 4406 4610 4414
rect 220 4376 228 4384
rect 284 4376 292 4384
rect 1324 4376 1332 4384
rect 1804 4376 1812 4384
rect 1836 4376 1844 4384
rect 2732 4376 2740 4384
rect 2844 4376 2852 4384
rect 3164 4376 3172 4384
rect 3276 4376 3284 4384
rect 3820 4376 3828 4384
rect 4716 4376 4724 4384
rect 5116 4376 5124 4384
rect 5404 4376 5412 4384
rect 5596 4376 5604 4384
rect 5948 4376 5956 4384
rect 5020 4358 5028 4366
rect 668 4336 676 4344
rect 700 4336 708 4344
rect 1340 4336 1348 4344
rect 1676 4336 1684 4344
rect 2876 4336 2884 4344
rect 3468 4336 3476 4344
rect 4156 4336 4164 4344
rect 4620 4336 4628 4344
rect 4700 4336 4708 4344
rect 92 4316 100 4324
rect 252 4316 260 4324
rect 60 4296 68 4304
rect 284 4296 292 4304
rect 364 4296 372 4304
rect 604 4296 612 4304
rect 716 4296 724 4304
rect 732 4296 740 4304
rect 780 4296 788 4304
rect 76 4276 84 4284
rect 108 4276 116 4284
rect 332 4276 340 4284
rect 380 4276 388 4284
rect 508 4276 516 4284
rect 540 4276 548 4284
rect 844 4296 852 4304
rect 876 4316 884 4324
rect 972 4316 980 4324
rect 908 4296 916 4304
rect 988 4296 996 4304
rect 1004 4296 1012 4304
rect 1068 4296 1076 4304
rect 1100 4296 1108 4304
rect 1148 4316 1156 4324
rect 1292 4316 1300 4324
rect 1628 4316 1636 4324
rect 1180 4296 1188 4304
rect 1260 4296 1268 4304
rect 1452 4296 1460 4304
rect 1564 4296 1572 4304
rect 1756 4316 1764 4324
rect 1676 4296 1684 4304
rect 1724 4296 1732 4304
rect 2076 4316 2084 4324
rect 2140 4316 2148 4324
rect 2156 4316 2164 4324
rect 2204 4316 2212 4324
rect 2412 4316 2420 4324
rect 2428 4316 2436 4324
rect 2524 4316 2532 4324
rect 2780 4316 2788 4324
rect 3164 4316 3172 4324
rect 1804 4296 1812 4304
rect 1948 4296 1956 4304
rect 2044 4296 2052 4304
rect 2108 4296 2116 4304
rect 2188 4296 2196 4304
rect 2236 4296 2244 4304
rect 812 4276 820 4284
rect 924 4276 932 4284
rect 940 4276 948 4284
rect 1068 4276 1076 4284
rect 1084 4276 1092 4284
rect 1132 4276 1140 4284
rect 1196 4276 1204 4284
rect 1500 4276 1508 4284
rect 1580 4276 1588 4284
rect 1692 4276 1700 4284
rect 1708 4276 1716 4284
rect 1820 4276 1828 4284
rect 1932 4276 1940 4284
rect 2028 4276 2036 4284
rect 2188 4276 2196 4284
rect 2300 4296 2308 4304
rect 2428 4296 2436 4304
rect 2460 4296 2468 4304
rect 2556 4296 2564 4304
rect 2588 4296 2596 4304
rect 2604 4296 2612 4304
rect 2668 4296 2676 4304
rect 2684 4296 2692 4304
rect 2700 4296 2708 4304
rect 2748 4296 2756 4304
rect 2956 4296 2964 4304
rect 3356 4296 3364 4304
rect 3484 4296 3492 4304
rect 3500 4296 3508 4304
rect 3548 4296 3556 4304
rect 2316 4276 2324 4284
rect 2332 4276 2340 4284
rect 2380 4276 2388 4284
rect 2572 4276 2580 4284
rect 2652 4276 2660 4284
rect 2812 4276 2820 4284
rect 3068 4276 3076 4284
rect 3372 4276 3380 4284
rect 3612 4296 3620 4304
rect 3644 4316 3652 4324
rect 3852 4316 3860 4324
rect 3980 4316 3988 4324
rect 4140 4316 4148 4324
rect 4428 4316 4436 4324
rect 4748 4316 4756 4324
rect 5020 4312 5028 4320
rect 5404 4316 5412 4324
rect 5948 4316 5956 4324
rect 3676 4296 3684 4304
rect 3724 4296 3732 4304
rect 3772 4296 3780 4304
rect 3788 4296 3796 4304
rect 3820 4296 3828 4304
rect 3852 4296 3860 4304
rect 3932 4296 3940 4304
rect 3964 4296 3972 4304
rect 4012 4296 4020 4304
rect 4028 4296 4036 4304
rect 4060 4296 4068 4304
rect 4076 4296 4084 4304
rect 4108 4296 4116 4304
rect 4140 4296 4148 4304
rect 4252 4296 4260 4304
rect 4396 4296 4404 4304
rect 4540 4296 4548 4304
rect 4716 4296 4724 4304
rect 5052 4296 5060 4304
rect 5196 4296 5204 4304
rect 5420 4296 5428 4304
rect 5452 4296 5460 4304
rect 5468 4296 5476 4304
rect 5516 4296 5524 4304
rect 5548 4296 5556 4304
rect 5564 4296 5572 4304
rect 5612 4296 5620 4304
rect 5740 4296 5748 4304
rect 5852 4296 5860 4304
rect 3580 4276 3588 4284
rect 3692 4276 3700 4284
rect 3804 4276 3812 4284
rect 4092 4276 4100 4284
rect 4252 4276 4260 4284
rect 4460 4276 4468 4284
rect 4956 4276 4964 4284
rect 5308 4276 5316 4284
rect 5532 4276 5540 4284
rect 5852 4276 5860 4284
rect 6124 4276 6132 4284
rect 12 4256 20 4264
rect 316 4256 324 4264
rect 572 4256 580 4264
rect 1212 4256 1220 4264
rect 1308 4256 1316 4264
rect 2828 4256 2836 4264
rect 3036 4256 3044 4264
rect 3260 4256 3268 4264
rect 3964 4256 3972 4264
rect 4348 4256 4356 4264
rect 4924 4256 4932 4264
rect 5276 4256 5284 4264
rect 5820 4256 5828 4264
rect 956 4236 964 4244
rect 1292 4236 1300 4244
rect 2140 4236 2148 4244
rect 2156 4236 2164 4244
rect 2348 4236 2356 4244
rect 2796 4236 2804 4244
rect 3740 4236 3748 4244
rect 3900 4236 3908 4244
rect 4428 4236 4436 4244
rect 5660 4236 5668 4244
rect 6012 4236 6020 4244
rect 3038 4206 3046 4214
rect 3052 4206 3060 4214
rect 3066 4206 3074 4214
rect 364 4176 372 4184
rect 1004 4176 1012 4184
rect 1164 4176 1172 4184
rect 1244 4176 1252 4184
rect 1724 4176 1732 4184
rect 2268 4176 2276 4184
rect 2460 4176 2468 4184
rect 2540 4176 2548 4184
rect 2732 4176 2740 4184
rect 3532 4176 3540 4184
rect 4108 4176 4116 4184
rect 4508 4176 4516 4184
rect 4812 4176 4820 4184
rect 5260 4176 5268 4184
rect 5420 4176 5428 4184
rect 5660 4176 5668 4184
rect 172 4156 180 4164
rect 1276 4156 1284 4164
rect 1292 4156 1300 4164
rect 1612 4156 1620 4164
rect 1980 4156 1988 4164
rect 2172 4156 2180 4164
rect 2252 4156 2260 4164
rect 2380 4156 2388 4164
rect 2476 4156 2484 4164
rect 3164 4156 3172 4164
rect 3612 4156 3620 4164
rect 3676 4156 3684 4164
rect 3692 4156 3700 4164
rect 3836 4156 3844 4164
rect 3916 4156 3924 4164
rect 4124 4156 4132 4164
rect 4364 4156 4372 4164
rect 4412 4156 4420 4164
rect 4988 4156 4996 4164
rect 5212 4156 5220 4164
rect 140 4136 148 4144
rect 428 4136 436 4144
rect 556 4136 564 4144
rect 636 4136 644 4144
rect 668 4136 676 4144
rect 844 4136 852 4144
rect 956 4136 964 4144
rect 972 4136 980 4144
rect 1004 4136 1012 4144
rect 1084 4136 1092 4144
rect 1100 4136 1108 4144
rect 1308 4136 1316 4144
rect 1452 4136 1460 4144
rect 1564 4136 1572 4144
rect 1628 4136 1636 4144
rect 1676 4136 1684 4144
rect 1756 4136 1764 4144
rect 1948 4136 1956 4144
rect 2396 4136 2404 4144
rect 2476 4136 2484 4144
rect 2588 4136 2596 4144
rect 2620 4136 2628 4144
rect 2652 4136 2660 4144
rect 2668 4136 2676 4144
rect 2764 4136 2772 4144
rect 2780 4136 2788 4144
rect 2812 4136 2820 4144
rect 2844 4136 2852 4144
rect 2988 4136 2996 4144
rect 3132 4136 3140 4144
rect 3372 4136 3380 4144
rect 3548 4136 3556 4144
rect 3660 4136 3668 4144
rect 3708 4136 3716 4144
rect 3820 4136 3828 4144
rect 4060 4136 4068 4144
rect 4220 4136 4228 4144
rect 4284 4136 4292 4144
rect 4348 4136 4356 4144
rect 4428 4136 4436 4144
rect 4492 4136 4500 4144
rect 4524 4136 4532 4144
rect 4604 4136 4612 4144
rect 4668 4136 4676 4144
rect 4732 4136 4740 4144
rect 4748 4136 4756 4144
rect 4844 4136 4852 4144
rect 252 4116 260 4124
rect 396 4116 404 4124
rect 444 4116 452 4124
rect 476 4116 484 4124
rect 492 4116 500 4124
rect 508 4116 516 4124
rect 556 4116 564 4124
rect 604 4116 612 4124
rect 620 4116 628 4124
rect 700 4118 708 4126
rect 860 4116 868 4124
rect 44 4096 52 4104
rect 364 4096 372 4104
rect 476 4096 484 4104
rect 588 4096 596 4104
rect 940 4116 948 4124
rect 1020 4116 1028 4124
rect 1132 4116 1140 4124
rect 1196 4116 1204 4124
rect 1324 4116 1332 4124
rect 1372 4116 1380 4124
rect 1388 4116 1396 4124
rect 1468 4116 1476 4124
rect 1580 4116 1588 4124
rect 1644 4116 1652 4124
rect 1692 4116 1700 4124
rect 1740 4116 1748 4124
rect 1948 4116 1956 4124
rect 2236 4116 2244 4124
rect 2300 4116 2308 4124
rect 2348 4116 2356 4124
rect 2636 4116 2644 4124
rect 2796 4116 2804 4124
rect 2860 4116 2868 4124
rect 3036 4116 3044 4124
rect 3420 4116 3428 4124
rect 3564 4116 3572 4124
rect 908 4096 916 4104
rect 1004 4096 1012 4104
rect 1068 4096 1076 4104
rect 1356 4096 1364 4104
rect 1484 4096 1492 4104
rect 1500 4096 1508 4104
rect 1612 4096 1620 4104
rect 1676 4096 1684 4104
rect 1804 4096 1812 4104
rect 1884 4100 1892 4108
rect 2364 4096 2372 4104
rect 2428 4096 2436 4104
rect 2604 4096 2612 4104
rect 2940 4096 2948 4104
rect 3068 4100 3076 4108
rect 3596 4096 3604 4104
rect 3644 4116 3652 4124
rect 3724 4116 3732 4124
rect 3756 4096 3764 4104
rect 3804 4116 3812 4124
rect 3884 4116 3892 4124
rect 3948 4116 3956 4124
rect 4012 4116 4020 4124
rect 4060 4116 4068 4124
rect 4076 4116 4084 4124
rect 4172 4116 4180 4124
rect 4300 4116 4308 4124
rect 4444 4116 4452 4124
rect 3916 4096 3924 4104
rect 3932 4096 3940 4104
rect 3996 4096 4004 4104
rect 4108 4096 4116 4104
rect 4204 4096 4212 4104
rect 4268 4096 4276 4104
rect 4332 4096 4340 4104
rect 4476 4096 4484 4104
rect 4652 4116 4660 4124
rect 4716 4116 4724 4124
rect 4892 4116 4900 4124
rect 4956 4132 4964 4140
rect 5020 4136 5028 4144
rect 5052 4136 5060 4144
rect 5100 4136 5108 4144
rect 5324 4136 5332 4144
rect 5916 4156 5924 4164
rect 5356 4136 5364 4144
rect 5452 4136 5460 4144
rect 5468 4136 5476 4144
rect 5532 4136 5540 4144
rect 5692 4136 5700 4144
rect 5708 4136 5716 4144
rect 5884 4136 5892 4144
rect 4988 4116 4996 4124
rect 5164 4116 5172 4124
rect 5452 4116 5460 4124
rect 5548 4116 5556 4124
rect 5788 4116 5796 4124
rect 5996 4116 6004 4124
rect 4572 4096 4580 4104
rect 4684 4096 4692 4104
rect 4860 4096 4868 4104
rect 5132 4096 5140 4104
rect 5148 4096 5156 4104
rect 5212 4096 5220 4104
rect 5516 4096 5524 4104
rect 5580 4096 5588 4104
rect 5740 4096 5748 4104
rect 5820 4100 5828 4108
rect 828 4076 836 4084
rect 2188 4076 2196 4084
rect 2332 4076 2340 4084
rect 2828 4076 2836 4084
rect 2908 4076 2916 4084
rect 3324 4076 3332 4084
rect 3500 4076 3508 4084
rect 3964 4076 3972 4084
rect 4028 4076 4036 4084
rect 5180 4076 5188 4084
rect 1884 4054 1892 4062
rect 3948 4056 3956 4064
rect 4652 4056 4660 4064
rect 5164 4056 5172 4064
rect 5820 4054 5828 4062
rect 44 4036 52 4044
rect 860 4036 868 4044
rect 1324 4036 1332 4044
rect 1420 4036 1428 4044
rect 1772 4036 1780 4044
rect 2220 4036 2228 4044
rect 3068 4036 3076 4044
rect 3804 4036 3812 4044
rect 4236 4036 4244 4044
rect 4300 4036 4308 4044
rect 4444 4036 4452 4044
rect 4716 4036 4724 4044
rect 4892 4036 4900 4044
rect 5292 4036 5300 4044
rect 5484 4036 5492 4044
rect 5724 4036 5732 4044
rect 6076 4036 6084 4044
rect 1502 4006 1510 4014
rect 1516 4006 1524 4014
rect 1530 4006 1538 4014
rect 4574 4006 4582 4014
rect 4588 4006 4596 4014
rect 4602 4006 4610 4014
rect 44 3976 52 3984
rect 428 3976 436 3984
rect 652 3976 660 3984
rect 924 3976 932 3984
rect 988 3976 996 3984
rect 1580 3976 1588 3984
rect 1612 3976 1620 3984
rect 1676 3976 1684 3984
rect 1964 3976 1972 3984
rect 2028 3976 2036 3984
rect 2684 3976 2692 3984
rect 2972 3976 2980 3984
rect 3084 3976 3092 3984
rect 3372 3976 3380 3984
rect 3420 3976 3428 3984
rect 3708 3976 3716 3984
rect 3932 3976 3940 3984
rect 3964 3976 3972 3984
rect 3996 3976 4004 3984
rect 4380 3976 4388 3984
rect 4620 3976 4628 3984
rect 4908 3976 4916 3984
rect 5100 3976 5108 3984
rect 5212 3976 5220 3984
rect 5676 3976 5684 3984
rect 5772 3976 5780 3984
rect 6060 3976 6068 3984
rect 2204 3958 2212 3966
rect 364 3936 372 3944
rect 1308 3936 1316 3944
rect 2460 3936 2468 3944
rect 2540 3936 2548 3944
rect 4092 3936 4100 3944
rect 4460 3936 4468 3944
rect 5612 3936 5620 3944
rect 44 3916 52 3924
rect 732 3916 740 3924
rect 1372 3916 1380 3924
rect 252 3896 260 3904
rect 460 3896 468 3904
rect 540 3896 548 3904
rect 572 3896 580 3904
rect 668 3896 676 3904
rect 748 3896 756 3904
rect 796 3896 804 3904
rect 812 3896 820 3904
rect 860 3896 868 3904
rect 892 3896 900 3904
rect 908 3896 916 3904
rect 956 3896 964 3904
rect 972 3896 980 3904
rect 1068 3896 1076 3904
rect 1084 3896 1092 3904
rect 1116 3896 1124 3904
rect 1196 3896 1204 3904
rect 1340 3896 1348 3904
rect 1964 3916 1972 3924
rect 2044 3916 2052 3924
rect 2092 3916 2100 3924
rect 2204 3912 2212 3920
rect 2524 3916 2532 3924
rect 2684 3916 2692 3924
rect 3084 3916 3092 3924
rect 3708 3916 3716 3924
rect 4380 3916 4388 3924
rect 4428 3916 4436 3924
rect 4620 3916 4628 3924
rect 5132 3916 5140 3924
rect 5212 3916 5220 3924
rect 5580 3916 5588 3924
rect 5772 3916 5780 3924
rect 1420 3896 1428 3904
rect 1564 3896 1572 3904
rect 1948 3896 1956 3904
rect 1964 3896 1972 3904
rect 2172 3896 2180 3904
rect 2524 3896 2532 3904
rect 2572 3896 2580 3904
rect 2636 3896 2644 3904
rect 2668 3896 2676 3904
rect 2892 3896 2900 3904
rect 3116 3896 3124 3904
rect 3676 3896 3684 3904
rect 3804 3894 3812 3902
rect 3868 3896 3876 3904
rect 4012 3896 4020 3904
rect 4380 3896 4388 3904
rect 4508 3896 4516 3904
rect 4828 3896 4836 3904
rect 5084 3896 5092 3904
rect 5196 3896 5204 3904
rect 5212 3896 5220 3904
rect 5420 3896 5428 3904
rect 5502 3896 5510 3904
rect 5516 3896 5524 3904
rect 5580 3896 5588 3904
rect 5612 3896 5620 3904
rect 5756 3896 5764 3904
rect 5772 3896 5780 3904
rect 140 3876 148 3884
rect 396 3876 404 3884
rect 780 3876 788 3884
rect 1212 3876 1220 3884
rect 1324 3876 1332 3884
rect 1388 3876 1396 3884
rect 1436 3876 1444 3884
rect 1868 3876 1876 3884
rect 2076 3876 2084 3884
rect 2108 3876 2116 3884
rect 2124 3876 2132 3884
rect 2268 3876 2276 3884
rect 2492 3876 2500 3884
rect 2780 3876 2788 3884
rect 3180 3876 3188 3884
rect 3612 3876 3620 3884
rect 4284 3876 4292 3884
rect 4428 3876 4436 3884
rect 4524 3876 4532 3884
rect 4716 3876 4724 3884
rect 4940 3876 4948 3884
rect 5068 3876 5076 3884
rect 5148 3876 5156 3884
rect 5164 3876 5172 3884
rect 5308 3876 5316 3884
rect 5708 3876 5716 3884
rect 5868 3876 5876 3884
rect 172 3856 180 3864
rect 348 3856 356 3864
rect 1004 3856 1012 3864
rect 1116 3856 1124 3864
rect 1516 3856 1524 3864
rect 1836 3856 1844 3864
rect 2012 3856 2020 3864
rect 2300 3856 2308 3864
rect 2812 3856 2820 3864
rect 3212 3856 3220 3864
rect 3580 3856 3588 3864
rect 3948 3856 3956 3864
rect 3980 3856 3988 3864
rect 4252 3856 4260 3864
rect 4748 3856 4756 3864
rect 5116 3856 5124 3864
rect 5340 3856 5348 3864
rect 5564 3856 5572 3864
rect 5660 3856 5668 3864
rect 5724 3856 5732 3864
rect 5900 3856 5908 3864
rect 380 3836 388 3844
rect 428 3836 436 3844
rect 700 3836 708 3844
rect 828 3836 836 3844
rect 1036 3836 1044 3844
rect 1612 3836 1620 3844
rect 2044 3836 2052 3844
rect 2524 3836 2532 3844
rect 2604 3836 2612 3844
rect 3372 3836 3380 3844
rect 4044 3836 4052 3844
rect 4092 3836 4100 3844
rect 5548 3836 5556 3844
rect 3038 3806 3046 3814
rect 3052 3806 3060 3814
rect 3066 3806 3074 3814
rect 124 3776 132 3784
rect 396 3776 404 3784
rect 924 3776 932 3784
rect 1148 3776 1156 3784
rect 1420 3776 1428 3784
rect 1724 3776 1732 3784
rect 2140 3776 2148 3784
rect 2316 3776 2324 3784
rect 2860 3776 2868 3784
rect 3004 3776 3012 3784
rect 3132 3776 3140 3784
rect 3212 3776 3220 3784
rect 3756 3776 3764 3784
rect 5084 3776 5092 3784
rect 5148 3776 5156 3784
rect 12 3756 20 3764
rect 44 3756 52 3764
rect 332 3756 340 3764
rect 1116 3756 1124 3764
rect 1900 3756 1908 3764
rect 2508 3756 2516 3764
rect 3196 3756 3204 3764
rect 3292 3756 3300 3764
rect 3420 3756 3428 3764
rect 3596 3756 3604 3764
rect 3964 3756 3972 3764
rect 4172 3756 4180 3764
rect 4652 3756 4660 3764
rect 4844 3756 4852 3764
rect 5372 3756 5380 3764
rect 5628 3756 5636 3764
rect 5900 3756 5908 3764
rect 60 3736 68 3744
rect 76 3736 84 3744
rect 140 3736 148 3744
rect 268 3736 276 3744
rect 380 3736 388 3744
rect 444 3736 452 3744
rect 492 3736 500 3744
rect 524 3736 532 3744
rect 556 3736 564 3744
rect 44 3716 52 3724
rect 92 3716 100 3724
rect 156 3716 164 3724
rect 124 3696 132 3704
rect 284 3716 292 3724
rect 364 3716 372 3724
rect 428 3716 436 3724
rect 556 3716 564 3724
rect 572 3716 580 3724
rect 588 3716 596 3724
rect 636 3716 644 3724
rect 668 3736 676 3744
rect 780 3736 788 3744
rect 908 3736 916 3744
rect 1084 3736 1092 3744
rect 1196 3736 1204 3744
rect 1212 3736 1220 3744
rect 1372 3736 1380 3744
rect 1436 3736 1444 3744
rect 1564 3736 1572 3744
rect 1660 3736 1668 3744
rect 1868 3736 1876 3744
rect 2124 3736 2132 3744
rect 2188 3736 2196 3744
rect 2204 3736 2212 3744
rect 2268 3736 2276 3744
rect 2540 3736 2548 3744
rect 2700 3736 2708 3744
rect 2748 3736 2756 3744
rect 2892 3736 2900 3744
rect 3388 3736 3396 3744
rect 3564 3736 3572 3744
rect 3996 3736 4004 3744
rect 4188 3736 4196 3744
rect 4316 3736 4324 3744
rect 4476 3736 4484 3744
rect 4684 3736 4692 3744
rect 4988 3736 4996 3744
rect 5004 3736 5012 3744
rect 5404 3736 5412 3744
rect 5580 3736 5588 3744
rect 5644 3736 5652 3744
rect 5660 3736 5668 3744
rect 5692 3736 5700 3744
rect 5932 3736 5940 3744
rect 204 3696 212 3704
rect 316 3696 324 3704
rect 332 3696 340 3704
rect 396 3696 404 3704
rect 460 3696 468 3704
rect 812 3716 820 3724
rect 732 3696 740 3704
rect 844 3696 852 3704
rect 892 3716 900 3724
rect 1020 3716 1028 3724
rect 1180 3716 1188 3724
rect 1228 3716 1236 3724
rect 1276 3716 1284 3724
rect 1292 3716 1300 3724
rect 1372 3716 1380 3724
rect 1388 3716 1396 3724
rect 1452 3716 1460 3724
rect 1532 3716 1540 3724
rect 1596 3718 1604 3726
rect 1980 3716 1988 3724
rect 2188 3716 2196 3724
rect 2284 3716 2292 3724
rect 2636 3716 2644 3724
rect 2732 3716 2740 3724
rect 3084 3716 3092 3724
rect 3100 3716 3108 3724
rect 3260 3716 3268 3724
rect 3308 3716 3316 3724
rect 3324 3716 3332 3724
rect 3468 3716 3476 3724
rect 3676 3716 3684 3724
rect 4076 3716 4084 3724
rect 4140 3716 4148 3724
rect 4332 3716 4340 3724
rect 4572 3716 4580 3724
rect 4780 3716 4788 3724
rect 4860 3716 4868 3724
rect 5052 3716 5060 3724
rect 5116 3716 5124 3724
rect 5292 3716 5300 3724
rect 5548 3716 5556 3724
rect 5676 3716 5684 3724
rect 5820 3716 5828 3724
rect 6076 3716 6084 3724
rect 892 3696 900 3704
rect 1260 3696 1268 3704
rect 1420 3696 1428 3704
rect 1484 3696 1492 3704
rect 1804 3700 1812 3708
rect 2060 3696 2068 3704
rect 2092 3696 2100 3704
rect 2124 3696 2132 3704
rect 2636 3696 2644 3704
rect 3212 3696 3220 3704
rect 3500 3700 3508 3708
rect 3804 3696 3812 3704
rect 4060 3700 4068 3708
rect 4204 3696 4212 3704
rect 4236 3696 4244 3704
rect 4380 3696 4388 3704
rect 4444 3696 4452 3704
rect 4492 3696 4500 3704
rect 4748 3700 4756 3708
rect 5468 3700 5476 3708
rect 5612 3696 5620 3704
rect 6028 3696 6036 3704
rect 1324 3676 1332 3684
rect 2204 3676 2212 3684
rect 2316 3676 2324 3684
rect 5708 3676 5716 3684
rect 6124 3676 6132 3684
rect 1804 3654 1812 3662
rect 3500 3654 3508 3662
rect 4060 3654 4068 3662
rect 5292 3654 5300 3662
rect 156 3636 164 3644
rect 284 3636 292 3644
rect 684 3636 692 3644
rect 1228 3636 1236 3644
rect 2108 3636 2116 3644
rect 2636 3636 2644 3644
rect 2860 3636 2868 3644
rect 4748 3636 4756 3644
rect 4828 3636 4836 3644
rect 5212 3636 5220 3644
rect 6028 3636 6036 3644
rect 1502 3606 1510 3614
rect 1516 3606 1524 3614
rect 1530 3606 1538 3614
rect 4574 3606 4582 3614
rect 4588 3606 4596 3614
rect 4602 3606 4610 3614
rect 140 3576 148 3584
rect 476 3576 484 3584
rect 492 3576 500 3584
rect 572 3576 580 3584
rect 780 3576 788 3584
rect 796 3576 804 3584
rect 1532 3576 1540 3584
rect 1820 3576 1828 3584
rect 2108 3576 2116 3584
rect 2220 3576 2228 3584
rect 2380 3576 2388 3584
rect 2668 3576 2676 3584
rect 2844 3576 2852 3584
rect 3420 3576 3428 3584
rect 4444 3576 4452 3584
rect 4508 3576 4516 3584
rect 5516 3576 5524 3584
rect 5692 3576 5700 3584
rect 2924 3558 2932 3566
rect 4860 3558 4868 3566
rect 5004 3558 5012 3566
rect 428 3536 436 3544
rect 556 3536 564 3544
rect 972 3536 980 3544
rect 92 3516 100 3524
rect 140 3516 148 3524
rect 508 3516 516 3524
rect 812 3516 820 3524
rect 908 3516 916 3524
rect 940 3516 948 3524
rect 60 3496 68 3504
rect 124 3496 132 3504
rect 236 3496 244 3504
rect 684 3496 692 3504
rect 908 3496 916 3504
rect 924 3496 932 3504
rect 1036 3496 1044 3504
rect 1052 3496 1060 3504
rect 1132 3496 1140 3504
rect 1148 3496 1156 3504
rect 1196 3516 1204 3524
rect 1260 3516 1268 3524
rect 1820 3516 1828 3524
rect 2380 3516 2388 3524
rect 2924 3512 2932 3520
rect 3420 3516 3428 3524
rect 3804 3516 3812 3524
rect 3948 3516 3956 3524
rect 4012 3516 4020 3524
rect 4076 3516 4084 3524
rect 4124 3516 4132 3524
rect 4444 3516 4452 3524
rect 4860 3512 4868 3520
rect 5004 3512 5012 3520
rect 5324 3516 5332 3524
rect 5548 3516 5556 3524
rect 5612 3516 5620 3524
rect 5644 3516 5652 3524
rect 5692 3516 5700 3524
rect 6044 3516 6052 3524
rect 1228 3496 1236 3504
rect 1292 3496 1300 3504
rect 1324 3496 1332 3504
rect 1340 3496 1348 3504
rect 1420 3496 1428 3504
rect 1708 3496 1716 3504
rect 1724 3496 1732 3504
rect 1740 3496 1748 3504
rect 2028 3496 2036 3504
rect 2188 3496 2196 3504
rect 2284 3496 2292 3504
rect 2380 3496 2388 3504
rect 2588 3496 2596 3504
rect 2700 3496 2708 3504
rect 2716 3496 2724 3504
rect 2892 3496 2900 3504
rect 3100 3496 3108 3504
rect 3182 3496 3190 3504
rect 3212 3496 3220 3504
rect 3244 3496 3252 3504
rect 3276 3496 3284 3504
rect 3436 3496 3444 3504
rect 3628 3496 3636 3504
rect 3820 3496 3828 3504
rect 3884 3496 3892 3504
rect 3900 3496 3908 3504
rect 3932 3496 3940 3504
rect 3980 3496 3988 3504
rect 3996 3496 4004 3504
rect 4236 3496 4244 3504
rect 4428 3496 4436 3504
rect 4892 3496 4900 3504
rect 4956 3496 4964 3504
rect 5180 3496 5188 3504
rect 5388 3496 5396 3504
rect 5404 3496 5412 3504
rect 5596 3496 5604 3504
rect 5676 3496 5684 3504
rect 5788 3496 5796 3504
rect 5900 3496 5908 3504
rect 5982 3496 5990 3504
rect 6044 3496 6052 3504
rect 236 3476 244 3484
rect 556 3476 564 3484
rect 684 3476 692 3484
rect 860 3476 868 3484
rect 924 3476 932 3484
rect 988 3476 996 3484
rect 1116 3476 1124 3484
rect 1132 3476 1140 3484
rect 1164 3476 1172 3484
rect 1244 3476 1252 3484
rect 1276 3476 1284 3484
rect 1308 3476 1316 3484
rect 1420 3476 1428 3484
rect 1916 3476 1924 3484
rect 2124 3476 2132 3484
rect 2268 3476 2276 3484
rect 2332 3476 2340 3484
rect 2476 3476 2484 3484
rect 2988 3476 2996 3484
rect 3516 3476 3524 3484
rect 3804 3476 3812 3484
rect 4044 3476 4052 3484
rect 4092 3476 4100 3484
rect 4348 3476 4356 3484
rect 4602 3476 4610 3484
rect 4796 3476 4804 3484
rect 5068 3476 5076 3484
rect 5292 3476 5300 3484
rect 5436 3476 5444 3484
rect 5452 3476 5460 3484
rect 5580 3476 5588 3484
rect 5596 3476 5604 3484
rect 5788 3476 5796 3484
rect 5996 3476 6004 3484
rect 6124 3476 6132 3484
rect 12 3456 20 3464
rect 268 3456 276 3464
rect 444 3456 452 3464
rect 508 3456 516 3464
rect 588 3456 596 3464
rect 812 3456 820 3464
rect 1020 3456 1028 3464
rect 1564 3456 1572 3464
rect 1948 3456 1956 3464
rect 2508 3456 2516 3464
rect 2732 3456 2740 3464
rect 2812 3456 2820 3464
rect 2828 3456 2836 3464
rect 3020 3456 3028 3464
rect 3292 3456 3300 3464
rect 3372 3456 3380 3464
rect 3548 3456 3556 3464
rect 3740 3456 3748 3464
rect 4076 3456 4084 3464
rect 4156 3456 4164 3464
rect 4316 3456 4324 3464
rect 4492 3456 4500 3464
rect 4764 3456 4772 3464
rect 5100 3456 5108 3464
rect 5820 3456 5828 3464
rect 92 3436 100 3444
rect 1356 3436 1364 3444
rect 1532 3436 1540 3444
rect 1692 3436 1700 3444
rect 3708 3436 3716 3444
rect 3804 3436 3812 3444
rect 4028 3436 4036 3444
rect 4108 3436 4116 3444
rect 5260 3436 5268 3444
rect 5308 3436 5316 3444
rect 5356 3436 5364 3444
rect 5548 3436 5556 3444
rect 6028 3436 6036 3444
rect 3196 3416 3204 3424
rect 3038 3406 3046 3414
rect 3052 3406 3060 3414
rect 3066 3406 3074 3414
rect 604 3376 612 3384
rect 1244 3376 1252 3384
rect 1436 3376 1444 3384
rect 1452 3376 1460 3384
rect 1548 3376 1556 3384
rect 2268 3376 2276 3384
rect 2348 3376 2356 3384
rect 3788 3376 3796 3384
rect 5724 3376 5732 3384
rect 5804 3376 5812 3384
rect 6060 3376 6068 3384
rect 172 3356 180 3364
rect 348 3356 356 3364
rect 444 3356 452 3364
rect 556 3356 564 3364
rect 764 3356 772 3364
rect 940 3356 948 3364
rect 1708 3356 1716 3364
rect 2108 3356 2116 3364
rect 2380 3356 2388 3364
rect 2572 3356 2580 3364
rect 2732 3356 2740 3364
rect 2780 3356 2788 3364
rect 3260 3356 3268 3364
rect 3532 3356 3540 3364
rect 140 3336 148 3344
rect 796 3336 804 3344
rect 972 3336 980 3344
rect 1084 3336 1092 3344
rect 1340 3336 1348 3344
rect 1740 3336 1748 3344
rect 1916 3336 1924 3344
rect 2076 3336 2084 3344
rect 2300 3336 2308 3344
rect 2540 3336 2548 3344
rect 76 3316 84 3324
rect 412 3316 420 3324
rect 524 3316 532 3324
rect 540 3316 548 3324
rect 796 3316 804 3324
rect 1036 3316 1044 3324
rect 1052 3316 1060 3324
rect 1164 3316 1172 3324
rect 1308 3318 1316 3326
rect 1804 3316 1812 3324
rect 1836 3316 1844 3324
rect 1884 3316 1892 3324
rect 2188 3316 2196 3324
rect 2540 3316 2548 3324
rect 3052 3336 3060 3344
rect 3164 3336 3172 3344
rect 3212 3336 3220 3344
rect 3276 3336 3284 3344
rect 3292 3336 3300 3344
rect 3340 3336 3348 3344
rect 3564 3336 3572 3344
rect 3756 3336 3764 3344
rect 3772 3336 3780 3344
rect 3836 3336 3844 3344
rect 4140 3356 4148 3364
rect 4364 3356 4372 3364
rect 4668 3356 4676 3364
rect 4684 3356 4692 3364
rect 4908 3356 4916 3364
rect 5052 3356 5060 3364
rect 5228 3356 5236 3364
rect 5564 3356 5572 3364
rect 5884 3356 5892 3364
rect 6028 3356 6036 3364
rect 3916 3336 3924 3344
rect 4172 3336 4180 3344
rect 4348 3336 4356 3344
rect 4396 3336 4404 3344
rect 4460 3336 4468 3344
rect 4508 3336 4516 3344
rect 4524 3336 4532 3344
rect 4556 3336 4564 3344
rect 3148 3316 3156 3324
rect 3260 3316 3268 3324
rect 3324 3316 3332 3324
rect 3628 3316 3636 3324
rect 3740 3316 3748 3324
rect 3788 3316 3796 3324
rect 4236 3316 4244 3324
rect 4476 3316 4484 3324
rect 4604 3316 4612 3324
rect 4620 3316 4628 3324
rect 4716 3316 4724 3324
rect 4828 3336 4836 3344
rect 4844 3336 4852 3344
rect 4892 3336 4900 3344
rect 5260 3336 5268 3344
rect 5532 3336 5540 3344
rect 5788 3336 5796 3344
rect 5852 3336 5860 3344
rect 5900 3336 5908 3344
rect 5932 3336 5940 3344
rect 5996 3336 6004 3344
rect 6108 3336 6116 3344
rect 4812 3316 4820 3324
rect 4956 3316 4964 3324
rect 5004 3316 5012 3324
rect 5356 3316 5364 3324
rect 5436 3316 5444 3324
rect 44 3296 52 3304
rect 892 3296 900 3304
rect 1836 3296 1844 3304
rect 2012 3300 2020 3308
rect 2476 3300 2484 3308
rect 2844 3296 2852 3304
rect 2908 3296 2916 3304
rect 2972 3296 2980 3304
rect 3052 3296 3060 3304
rect 3196 3296 3204 3304
rect 3292 3296 3300 3304
rect 3372 3296 3380 3304
rect 3660 3296 3668 3304
rect 3708 3296 3716 3304
rect 3852 3296 3860 3304
rect 4268 3296 4276 3304
rect 4316 3296 4324 3304
rect 4412 3296 4420 3304
rect 4444 3296 4452 3304
rect 4508 3296 4516 3304
rect 4556 3296 4564 3304
rect 4780 3296 4788 3304
rect 4876 3296 4884 3304
rect 4940 3296 4948 3304
rect 5324 3300 5332 3308
rect 5436 3296 5444 3304
rect 5932 3296 5940 3304
rect 5948 3296 5956 3304
rect 2812 3276 2820 3284
rect 2876 3276 2884 3284
rect 2940 3276 2948 3284
rect 3004 3276 3012 3284
rect 3740 3276 3748 3284
rect 4668 3276 4676 3284
rect 4956 3276 4964 3284
rect 2476 3254 2484 3262
rect 5324 3254 5332 3262
rect 44 3236 52 3244
rect 380 3236 388 3244
rect 492 3236 500 3244
rect 572 3236 580 3244
rect 892 3236 900 3244
rect 1836 3236 1844 3244
rect 2012 3236 2020 3244
rect 2396 3236 2404 3244
rect 2764 3236 2772 3244
rect 2796 3236 2804 3244
rect 2892 3236 2900 3244
rect 2956 3236 2964 3244
rect 3020 3236 3028 3244
rect 3660 3236 3668 3244
rect 3980 3236 3988 3244
rect 4268 3236 4276 3244
rect 4332 3236 4340 3244
rect 4748 3236 4756 3244
rect 4860 3236 4868 3244
rect 4908 3236 4916 3244
rect 4988 3236 4996 3244
rect 5020 3236 5028 3244
rect 5068 3236 5076 3244
rect 5436 3236 5444 3244
rect 5916 3236 5924 3244
rect 1502 3206 1510 3214
rect 1516 3206 1524 3214
rect 1530 3206 1538 3214
rect 4574 3206 4582 3214
rect 4588 3206 4596 3214
rect 4602 3206 4610 3214
rect 124 3176 132 3184
rect 188 3176 196 3184
rect 476 3176 484 3184
rect 524 3176 532 3184
rect 812 3176 820 3184
rect 1100 3176 1108 3184
rect 1388 3176 1396 3184
rect 1612 3176 1620 3184
rect 1964 3176 1972 3184
rect 2364 3176 2372 3184
rect 2588 3176 2596 3184
rect 2684 3176 2692 3184
rect 4284 3176 4292 3184
rect 5260 3176 5268 3184
rect 5468 3176 5476 3184
rect 5532 3176 5540 3184
rect 1868 3158 1876 3166
rect 2076 3158 2084 3166
rect 3244 3158 3252 3166
rect 3708 3156 3716 3164
rect 4572 3156 4580 3164
rect 3580 3136 3588 3144
rect 3724 3136 3732 3144
rect 5020 3136 5028 3144
rect 5084 3136 5092 3144
rect 5212 3136 5220 3144
rect 5324 3136 5332 3144
rect 188 3116 196 3124
rect 812 3116 820 3124
rect 1388 3116 1396 3124
rect 1868 3112 1876 3120
rect 1948 3116 1956 3124
rect 1980 3116 1988 3124
rect 2076 3112 2084 3120
rect 2428 3116 2436 3124
rect 2476 3116 2484 3124
rect 2748 3116 2756 3124
rect 2844 3116 2852 3124
rect 3244 3112 3252 3120
rect 3372 3116 3380 3124
rect 188 3096 196 3104
rect 796 3096 804 3104
rect 876 3096 884 3104
rect 924 3096 932 3104
rect 956 3096 964 3104
rect 972 3096 980 3104
rect 1180 3096 1188 3104
rect 1372 3096 1380 3104
rect 1468 3096 1476 3104
rect 1580 3096 1588 3104
rect 1692 3096 1700 3104
rect 1804 3096 1812 3104
rect 1916 3096 1924 3104
rect 1964 3096 1972 3104
rect 2044 3096 2052 3104
rect 2334 3096 2342 3104
rect 2492 3096 2500 3104
rect 2572 3096 2580 3104
rect 2620 3096 2628 3104
rect 2652 3096 2660 3104
rect 2668 3096 2676 3104
rect 2748 3096 2756 3104
rect 2780 3096 2788 3104
rect 2796 3096 2804 3104
rect 12 3076 20 3084
rect 284 3076 292 3084
rect 716 3076 724 3084
rect 860 3076 868 3084
rect 1036 3076 1044 3084
rect 1292 3076 1300 3084
rect 1564 3076 1572 3084
rect 1804 3076 1812 3084
rect 2140 3076 2148 3084
rect 2380 3076 2388 3084
rect 2540 3076 2548 3084
rect 2732 3076 2740 3084
rect 2796 3076 2804 3084
rect 2844 3096 2852 3104
rect 2924 3096 2932 3104
rect 3068 3096 3076 3104
rect 3420 3116 3428 3124
rect 3484 3116 3492 3124
rect 3852 3116 3860 3124
rect 3868 3116 3876 3124
rect 4012 3116 4020 3124
rect 4076 3116 4084 3124
rect 4124 3116 4132 3124
rect 4236 3116 4244 3124
rect 4284 3116 4292 3124
rect 4716 3116 4724 3124
rect 4796 3116 4804 3124
rect 4812 3116 4820 3124
rect 4876 3116 4884 3124
rect 5052 3116 5060 3124
rect 5116 3116 5124 3124
rect 5132 3116 5140 3124
rect 5180 3116 5188 3124
rect 5372 3116 5380 3124
rect 5532 3116 5540 3124
rect 5852 3116 5860 3124
rect 5932 3116 5940 3124
rect 3516 3096 3524 3104
rect 2828 3076 2836 3084
rect 2876 3076 2884 3084
rect 2940 3076 2948 3084
rect 2986 3076 2994 3084
rect 3180 3076 3188 3084
rect 3324 3076 3332 3084
rect 3468 3076 3476 3084
rect 3596 3096 3604 3104
rect 3644 3096 3652 3104
rect 3708 3096 3716 3104
rect 3756 3096 3764 3104
rect 3788 3096 3796 3104
rect 3820 3096 3828 3104
rect 3884 3096 3892 3104
rect 3948 3096 3956 3104
rect 3980 3096 3988 3104
rect 4028 3096 4036 3104
rect 4044 3096 4052 3104
rect 4076 3096 4084 3104
rect 4156 3096 4164 3104
rect 4204 3096 4212 3104
rect 4236 3096 4244 3104
rect 4284 3096 4292 3104
rect 4492 3096 4500 3104
rect 4668 3096 4676 3104
rect 4716 3096 4724 3104
rect 4764 3096 4772 3104
rect 4844 3096 4852 3104
rect 5004 3096 5012 3104
rect 5020 3096 5028 3104
rect 5084 3096 5092 3104
rect 5116 3096 5124 3104
rect 5260 3096 5268 3104
rect 5292 3096 5300 3104
rect 5388 3096 5396 3104
rect 5740 3096 5748 3104
rect 6044 3096 6052 3104
rect 3772 3076 3780 3084
rect 3804 3076 3812 3084
rect 3836 3076 3844 3084
rect 3900 3076 3908 3084
rect 3932 3076 3940 3084
rect 3964 3076 3972 3084
rect 4028 3076 4036 3084
rect 4092 3076 4100 3084
rect 4172 3076 4180 3084
rect 4188 3076 4196 3084
rect 4380 3076 4388 3084
rect 4652 3076 4660 3084
rect 4860 3076 4868 3084
rect 4924 3076 4932 3084
rect 4972 3076 4980 3084
rect 5004 3076 5012 3084
rect 5068 3076 5076 3084
rect 5164 3076 5172 3084
rect 5212 3076 5220 3084
rect 5276 3076 5284 3084
rect 5340 3076 5348 3084
rect 5452 3076 5460 3084
rect 5628 3076 5636 3084
rect 5852 3076 5860 3084
rect 5900 3076 5908 3084
rect 5996 3076 6004 3084
rect 6124 3076 6132 3084
rect 316 3056 324 3064
rect 684 3056 692 3064
rect 1260 3056 1268 3064
rect 1436 3056 1444 3064
rect 1772 3056 1780 3064
rect 2172 3056 2180 3064
rect 2460 3056 2468 3064
rect 3148 3056 3156 3064
rect 3564 3056 3572 3064
rect 4108 3056 4116 3064
rect 4412 3056 4420 3064
rect 4716 3056 4724 3064
rect 4796 3056 4804 3064
rect 4940 3056 4948 3064
rect 5660 3056 5668 3064
rect 5820 3056 5828 3064
rect 5932 3056 5940 3064
rect 6028 3056 6036 3064
rect 1548 3036 1556 3044
rect 1612 3036 1620 3044
rect 1964 3036 1972 3044
rect 2892 3036 2900 3044
rect 3388 3036 3396 3044
rect 3596 3036 3604 3044
rect 3932 3036 3940 3044
rect 4124 3036 4132 3044
rect 4572 3036 4580 3044
rect 4812 3036 4820 3044
rect 4876 3036 4884 3044
rect 5180 3036 5188 3044
rect 5372 3036 5380 3044
rect 5420 3036 5428 3044
rect 5468 3036 5476 3044
rect 5948 3036 5956 3044
rect 3038 3006 3046 3014
rect 3052 3006 3060 3014
rect 3066 3006 3074 3014
rect 1980 2996 1988 3004
rect 1228 2976 1236 2984
rect 1692 2976 1700 2984
rect 2076 2976 2084 2984
rect 2988 2976 2996 2984
rect 3356 2976 3364 2984
rect 3692 2976 3700 2984
rect 3868 2976 3876 2984
rect 3964 2976 3972 2984
rect 3996 2976 4004 2984
rect 4348 2976 4356 2984
rect 4428 2976 4436 2984
rect 4764 2976 4772 2984
rect 4972 2976 4980 2984
rect 5116 2976 5124 2984
rect 5292 2976 5300 2984
rect 5756 2976 5764 2984
rect 316 2956 324 2964
rect 572 2956 580 2964
rect 780 2956 788 2964
rect 1084 2956 1092 2964
rect 1388 2956 1396 2964
rect 1612 2956 1620 2964
rect 1868 2956 1876 2964
rect 2348 2956 2356 2964
rect 2828 2956 2836 2964
rect 3388 2956 3396 2964
rect 4156 2956 4164 2964
rect 4508 2956 4516 2964
rect 4588 2956 4596 2964
rect 4780 2956 4788 2964
rect 4892 2956 4900 2964
rect 4908 2956 4916 2964
rect 5212 2956 5220 2964
rect 5228 2956 5236 2964
rect 5548 2956 5556 2964
rect 5932 2956 5940 2964
rect 12 2936 20 2944
rect 140 2936 148 2944
rect 284 2936 292 2944
rect 588 2936 596 2944
rect 748 2936 756 2944
rect 1052 2936 1060 2944
rect 1420 2936 1428 2944
rect 1836 2936 1844 2944
rect 2060 2936 2068 2944
rect 2092 2936 2100 2944
rect 2316 2936 2324 2944
rect 2572 2936 2580 2944
rect 2796 2936 2804 2944
rect 3164 2936 3172 2944
rect 3276 2936 3284 2944
rect 3340 2936 3348 2944
rect 188 2916 196 2924
rect 284 2916 292 2924
rect 540 2916 548 2924
rect 604 2916 612 2924
rect 684 2916 692 2924
rect 1004 2916 1012 2924
rect 1020 2916 1028 2924
rect 1068 2916 1076 2924
rect 1100 2916 1108 2924
rect 1116 2916 1124 2924
rect 1132 2916 1140 2924
rect 1180 2916 1188 2924
rect 1516 2916 1524 2924
rect 1660 2916 1668 2924
rect 1756 2916 1764 2924
rect 2124 2916 2132 2924
rect 2220 2916 2228 2924
rect 2636 2916 2644 2924
rect 2652 2916 2660 2924
rect 2700 2916 2708 2924
rect 2908 2916 2916 2924
rect 3052 2916 3060 2924
rect 3228 2916 3236 2924
rect 3292 2916 3300 2924
rect 3308 2916 3316 2924
rect 188 2896 196 2904
rect 652 2896 660 2904
rect 1484 2900 1492 2908
rect 1692 2896 1700 2904
rect 1772 2900 1780 2908
rect 2140 2896 2148 2904
rect 2172 2896 2180 2904
rect 2220 2896 2228 2904
rect 2700 2896 2708 2904
rect 3052 2896 3060 2904
rect 3148 2896 3156 2904
rect 3196 2896 3204 2904
rect 3228 2896 3236 2904
rect 3260 2896 3268 2904
rect 3324 2896 3332 2904
rect 3484 2916 3492 2924
rect 3724 2936 3732 2944
rect 3548 2916 3556 2924
rect 3596 2916 3604 2924
rect 3612 2916 3620 2924
rect 3660 2916 3668 2924
rect 3804 2936 3812 2944
rect 3868 2936 3876 2944
rect 3900 2936 3908 2944
rect 3932 2936 3940 2944
rect 4188 2936 4196 2944
rect 4348 2936 4356 2944
rect 4380 2936 4388 2944
rect 4428 2936 4436 2944
rect 4476 2936 4484 2944
rect 4508 2936 4516 2944
rect 4636 2936 4644 2944
rect 4748 2936 4756 2944
rect 4796 2936 4804 2944
rect 4828 2936 4836 2944
rect 4860 2936 4868 2944
rect 4908 2936 4916 2944
rect 4956 2936 4964 2944
rect 5068 2936 5076 2944
rect 5132 2936 5140 2944
rect 5260 2936 5268 2944
rect 5324 2936 5332 2944
rect 5356 2936 5364 2944
rect 5580 2936 5588 2944
rect 5724 2936 5732 2944
rect 5900 2936 5908 2944
rect 3852 2916 3860 2924
rect 3916 2916 3924 2924
rect 4284 2916 4292 2924
rect 4332 2916 4340 2924
rect 4396 2916 4404 2924
rect 4412 2916 4420 2924
rect 4476 2916 4484 2924
rect 4620 2916 4628 2924
rect 4684 2916 4692 2924
rect 4732 2916 4740 2924
rect 4844 2916 4852 2924
rect 4892 2916 4900 2924
rect 4940 2916 4948 2924
rect 4988 2916 4996 2924
rect 5084 2916 5092 2924
rect 5180 2916 5188 2924
rect 5260 2916 5268 2924
rect 5340 2916 5348 2924
rect 5580 2916 5588 2924
rect 5692 2916 5700 2924
rect 5788 2916 5796 2924
rect 6012 2916 6020 2924
rect 3468 2896 3476 2904
rect 3516 2896 3524 2904
rect 3692 2896 3700 2904
rect 3740 2896 3748 2904
rect 3980 2896 3988 2904
rect 4284 2896 4292 2904
rect 4604 2896 4612 2904
rect 4668 2896 4676 2904
rect 4796 2896 4804 2904
rect 4988 2896 4996 2904
rect 5004 2896 5012 2904
rect 5164 2896 5172 2904
rect 5308 2896 5316 2904
rect 5388 2896 5396 2904
rect 5644 2900 5652 2908
rect 5756 2896 5764 2904
rect 5804 2896 5812 2904
rect 3564 2876 3572 2884
rect 3724 2876 3732 2884
rect 3548 2856 3556 2864
rect 3772 2876 3780 2884
rect 4636 2876 4644 2884
rect 4668 2876 4676 2884
rect 4956 2876 4964 2884
rect 5644 2854 5652 2862
rect 188 2836 196 2844
rect 476 2836 484 2844
rect 652 2836 660 2844
rect 940 2836 948 2844
rect 1148 2836 1156 2844
rect 1228 2836 1236 2844
rect 1484 2836 1492 2844
rect 1772 2836 1780 2844
rect 2076 2836 2084 2844
rect 2220 2836 2228 2844
rect 2508 2836 2516 2844
rect 2700 2836 2708 2844
rect 3628 2836 3636 2844
rect 3820 2836 3828 2844
rect 3996 2836 4004 2844
rect 4284 2836 4292 2844
rect 4716 2836 4724 2844
rect 5196 2836 5204 2844
rect 5260 2836 5268 2844
rect 5292 2836 5300 2844
rect 5804 2836 5812 2844
rect 6092 2836 6100 2844
rect 1502 2806 1510 2814
rect 1516 2806 1524 2814
rect 1530 2806 1538 2814
rect 4574 2806 4582 2814
rect 4588 2806 4596 2814
rect 4602 2806 4610 2814
rect 44 2776 52 2784
rect 668 2776 676 2784
rect 844 2776 852 2784
rect 1132 2776 1140 2784
rect 1260 2776 1268 2784
rect 1644 2776 1652 2784
rect 1788 2776 1796 2784
rect 2284 2776 2292 2784
rect 2348 2776 2356 2784
rect 2940 2776 2948 2784
rect 3804 2776 3812 2784
rect 3836 2776 3844 2784
rect 3900 2776 3908 2784
rect 4332 2776 4340 2784
rect 4412 2776 4420 2784
rect 4524 2776 4532 2784
rect 4748 2776 4756 2784
rect 4924 2776 4932 2784
rect 5052 2776 5060 2784
rect 5244 2776 5252 2784
rect 5308 2776 5316 2784
rect 3164 2758 3172 2766
rect 3996 2756 4004 2764
rect 3436 2736 3444 2744
rect 3724 2736 3732 2744
rect 3788 2736 3796 2744
rect 3852 2736 3860 2744
rect 3916 2736 3924 2744
rect 4076 2736 4084 2744
rect 4172 2736 4180 2744
rect 4348 2736 4356 2744
rect 4396 2736 4404 2744
rect 4556 2736 4564 2744
rect 4780 2756 4788 2764
rect 5004 2756 5012 2764
rect 5788 2756 5796 2764
rect 6044 2758 6052 2766
rect 44 2716 52 2724
rect 668 2716 676 2724
rect 1132 2716 1140 2724
rect 1692 2716 1700 2724
rect 1788 2716 1796 2724
rect 2172 2716 2180 2724
rect 2220 2716 2228 2724
rect 2348 2716 2356 2724
rect 2796 2716 2804 2724
rect 2876 2716 2884 2724
rect 2908 2716 2916 2724
rect 3164 2712 3172 2720
rect 3468 2716 3476 2724
rect 3564 2716 3572 2724
rect 3596 2716 3604 2724
rect 3644 2716 3652 2724
rect 3692 2716 3700 2724
rect 3756 2716 3764 2724
rect 3820 2716 3828 2724
rect 4140 2716 4148 2724
rect 4316 2716 4324 2724
rect 4428 2716 4436 2724
rect 4460 2716 4468 2724
rect 4668 2736 4676 2744
rect 4700 2736 4708 2744
rect 4796 2736 4804 2744
rect 4828 2736 4836 2744
rect 5100 2736 5108 2744
rect 5724 2736 5732 2744
rect 4636 2716 4644 2724
rect 4716 2716 4724 2724
rect 4764 2716 4772 2724
rect 5068 2716 5076 2724
rect 5276 2716 5284 2724
rect 5372 2716 5380 2724
rect 5452 2716 5460 2724
rect 5500 2716 5508 2724
rect 5612 2716 5620 2724
rect 5644 2716 5652 2724
rect 5756 2716 5764 2724
rect 6044 2712 6052 2720
rect 252 2696 260 2704
rect 460 2696 468 2704
rect 652 2696 660 2704
rect 748 2696 756 2704
rect 812 2696 820 2704
rect 924 2696 932 2704
rect 1132 2696 1140 2704
rect 1228 2696 1236 2704
rect 1532 2696 1540 2704
rect 1644 2696 1652 2704
rect 1788 2696 1796 2704
rect 1996 2696 2004 2704
rect 2124 2696 2132 2704
rect 2556 2696 2564 2704
rect 2668 2696 2676 2704
rect 2684 2696 2692 2704
rect 2780 2696 2788 2704
rect 2860 2696 2868 2704
rect 2876 2696 2884 2704
rect 2956 2696 2964 2704
rect 2972 2696 2980 2704
rect 3020 2696 3028 2704
rect 3228 2696 3236 2704
rect 3484 2696 3492 2704
rect 3516 2696 3524 2704
rect 3532 2696 3540 2704
rect 3596 2696 3604 2704
rect 140 2676 148 2684
rect 572 2676 580 2684
rect 748 2676 756 2684
rect 796 2676 804 2684
rect 1036 2676 1044 2684
rect 1212 2676 1220 2684
rect 1388 2676 1396 2684
rect 1628 2676 1636 2684
rect 1724 2676 1732 2684
rect 1884 2676 1892 2684
rect 2078 2676 2086 2684
rect 2124 2676 2132 2684
rect 2300 2676 2308 2684
rect 2444 2676 2452 2684
rect 2844 2676 2852 2684
rect 2860 2676 2868 2684
rect 3084 2676 3092 2684
rect 3228 2676 3236 2684
rect 3532 2676 3540 2684
rect 3548 2676 3556 2684
rect 3676 2676 3684 2684
rect 3772 2696 3780 2704
rect 3836 2696 3844 2704
rect 3724 2676 3732 2684
rect 3900 2696 3908 2704
rect 3948 2696 3956 2704
rect 4012 2696 4020 2704
rect 4092 2696 4100 2704
rect 4140 2696 4148 2704
rect 4220 2696 4228 2704
rect 4268 2696 4276 2704
rect 4300 2696 4308 2704
rect 4332 2696 4340 2704
rect 4412 2696 4420 2704
rect 4444 2696 4452 2704
rect 4508 2696 4516 2704
rect 4540 2696 4548 2704
rect 4652 2696 4660 2704
rect 4716 2696 4724 2704
rect 4780 2696 4788 2704
rect 4828 2696 4836 2704
rect 4892 2696 4900 2704
rect 4924 2696 4932 2704
rect 4956 2696 4964 2704
rect 5052 2696 5060 2704
rect 5116 2696 5124 2704
rect 5164 2696 5172 2704
rect 3964 2676 3972 2684
rect 4012 2676 4020 2684
rect 4044 2676 4052 2684
rect 4076 2676 4084 2684
rect 4108 2676 4116 2684
rect 4156 2676 4164 2684
rect 4172 2676 4180 2684
rect 4204 2676 4212 2684
rect 4252 2676 4260 2684
rect 4284 2676 4292 2684
rect 4460 2676 4468 2684
rect 4492 2676 4500 2684
rect 4876 2676 4884 2684
rect 4940 2676 4948 2684
rect 4972 2676 4980 2684
rect 5116 2676 5124 2684
rect 5308 2696 5316 2704
rect 5340 2696 5348 2704
rect 5564 2696 5572 2704
rect 5676 2696 5684 2704
rect 5868 2696 5876 2704
rect 5228 2676 5236 2684
rect 5292 2676 5300 2684
rect 5356 2676 5364 2684
rect 5404 2676 5412 2684
rect 5484 2676 5492 2684
rect 5548 2676 5556 2684
rect 5644 2676 5652 2684
rect 5772 2676 5780 2684
rect 5980 2676 5988 2684
rect 172 2656 180 2664
rect 540 2656 548 2664
rect 716 2656 724 2664
rect 1004 2656 1012 2664
rect 1180 2656 1188 2664
rect 1676 2656 1684 2664
rect 1740 2656 1748 2664
rect 1916 2656 1924 2664
rect 2204 2656 2212 2664
rect 2476 2656 2484 2664
rect 2636 2656 2644 2664
rect 2700 2656 2708 2664
rect 2780 2656 2788 2664
rect 2924 2656 2932 2664
rect 3260 2656 3268 2664
rect 3468 2656 3476 2664
rect 3628 2656 3636 2664
rect 4860 2656 4868 2664
rect 5004 2656 5012 2664
rect 5020 2656 5028 2664
rect 5132 2656 5140 2664
rect 5148 2656 5156 2664
rect 5212 2656 5220 2664
rect 5436 2656 5444 2664
rect 5948 2656 5956 2664
rect 332 2636 340 2644
rect 380 2636 388 2644
rect 1196 2636 1204 2644
rect 1260 2636 1268 2644
rect 1500 2636 1508 2644
rect 2252 2636 2260 2644
rect 3420 2636 3428 2644
rect 3660 2636 3668 2644
rect 4844 2636 4852 2644
rect 5388 2636 5396 2644
rect 5420 2636 5428 2644
rect 5452 2636 5460 2644
rect 5516 2636 5524 2644
rect 5644 2636 5652 2644
rect 3260 2616 3268 2624
rect 3038 2606 3046 2614
rect 3052 2606 3060 2614
rect 3066 2606 3074 2614
rect 812 2576 820 2584
rect 908 2576 916 2584
rect 1724 2576 1732 2584
rect 2860 2576 2868 2584
rect 2956 2576 2964 2584
rect 3004 2576 3012 2584
rect 3116 2576 3124 2584
rect 3868 2576 3876 2584
rect 3980 2576 3988 2584
rect 4332 2576 4340 2584
rect 4556 2576 4564 2584
rect 4684 2576 4692 2584
rect 4780 2576 4788 2584
rect 4812 2576 4820 2584
rect 4924 2576 4932 2584
rect 5148 2576 5156 2584
rect 5196 2576 5204 2584
rect 5276 2576 5284 2584
rect 5468 2576 5476 2584
rect 5708 2576 5716 2584
rect 6076 2576 6084 2584
rect 172 2556 180 2564
rect 380 2556 388 2564
rect 556 2556 564 2564
rect 748 2556 756 2564
rect 892 2556 900 2564
rect 1116 2556 1124 2564
rect 1308 2556 1316 2564
rect 1612 2556 1620 2564
rect 2108 2556 2116 2564
rect 2668 2556 2676 2564
rect 3084 2556 3092 2564
rect 3132 2556 3140 2564
rect 3500 2556 3508 2564
rect 3676 2556 3684 2564
rect 3884 2556 3892 2564
rect 4236 2556 4244 2564
rect 4796 2556 4804 2564
rect 4876 2556 4884 2564
rect 4892 2556 4900 2564
rect 4908 2556 4916 2564
rect 4940 2556 4948 2564
rect 5004 2556 5012 2564
rect 5164 2556 5172 2564
rect 5340 2556 5348 2564
rect 5868 2556 5876 2564
rect 140 2536 148 2544
rect 524 2536 532 2544
rect 828 2536 836 2544
rect 1148 2536 1156 2544
rect 1308 2536 1316 2544
rect 1644 2536 1652 2544
rect 1788 2536 1796 2544
rect 1820 2536 1828 2544
rect 1884 2536 1892 2544
rect 1932 2536 1940 2544
rect 2076 2536 2084 2544
rect 2332 2536 2340 2544
rect 2700 2536 2708 2544
rect 2844 2536 2852 2544
rect 2908 2536 2916 2544
rect 2972 2536 2980 2544
rect 2988 2536 2996 2544
rect 3100 2536 3108 2544
rect 3148 2536 3156 2544
rect 3260 2536 3268 2544
rect 3276 2536 3284 2544
rect 3340 2536 3348 2544
rect 3388 2536 3396 2544
rect 252 2516 260 2524
rect 412 2516 420 2524
rect 636 2516 644 2524
rect 780 2516 788 2524
rect 844 2516 852 2524
rect 876 2516 884 2524
rect 1244 2516 1252 2524
rect 1372 2516 1380 2524
rect 1740 2516 1748 2524
rect 44 2496 52 2504
rect 460 2500 468 2508
rect 1212 2500 1220 2508
rect 1708 2500 1716 2508
rect 1820 2496 1828 2504
rect 1868 2516 1876 2524
rect 1996 2516 2004 2524
rect 2396 2516 2404 2524
rect 2428 2516 2436 2524
rect 2476 2516 2484 2524
rect 2588 2516 2596 2524
rect 2860 2516 2868 2524
rect 2956 2516 2964 2524
rect 3196 2516 3204 2524
rect 3244 2516 3252 2524
rect 3292 2516 3300 2524
rect 3644 2536 3652 2544
rect 3420 2516 3428 2524
rect 3468 2516 3476 2524
rect 3564 2516 3572 2524
rect 3980 2536 3988 2544
rect 4012 2536 4020 2544
rect 4044 2536 4052 2544
rect 4060 2536 4068 2544
rect 4092 2536 4100 2544
rect 4124 2536 4132 2544
rect 4268 2536 4276 2544
rect 4300 2536 4308 2544
rect 4332 2536 4340 2544
rect 4364 2536 4372 2544
rect 4396 2536 4404 2544
rect 4444 2536 4452 2544
rect 4524 2536 4532 2544
rect 4540 2536 4548 2544
rect 4572 2536 4580 2544
rect 4652 2536 4660 2544
rect 4700 2536 4708 2544
rect 4972 2536 4980 2544
rect 5020 2536 5028 2544
rect 5052 2536 5060 2544
rect 5180 2536 5188 2544
rect 5260 2536 5268 2544
rect 5436 2536 5444 2544
rect 5452 2536 5460 2544
rect 5484 2536 5492 2544
rect 5548 2536 5556 2544
rect 5900 2536 5908 2544
rect 3916 2516 3924 2524
rect 3964 2516 3972 2524
rect 4028 2516 4036 2524
rect 4044 2516 4052 2524
rect 4076 2516 4084 2524
rect 4108 2516 4116 2524
rect 4188 2516 4196 2524
rect 4236 2516 4244 2524
rect 4284 2516 4292 2524
rect 4348 2516 4356 2524
rect 4476 2516 4484 2524
rect 4524 2516 4532 2524
rect 4588 2516 4596 2524
rect 4652 2516 4660 2524
rect 4716 2516 4724 2524
rect 4748 2516 4756 2524
rect 4828 2516 4836 2524
rect 4844 2516 4852 2524
rect 4956 2516 4964 2524
rect 5100 2516 5108 2524
rect 5132 2516 5140 2524
rect 5196 2516 5204 2524
rect 5228 2516 5236 2524
rect 5276 2516 5284 2524
rect 5308 2516 5316 2524
rect 5340 2516 5348 2524
rect 5388 2516 5396 2524
rect 5420 2516 5428 2524
rect 5788 2516 5796 2524
rect 6044 2516 6052 2524
rect 2012 2500 2020 2508
rect 2796 2496 2804 2504
rect 2924 2496 2932 2504
rect 3020 2496 3028 2504
rect 3212 2496 3220 2504
rect 3356 2496 3364 2504
rect 3580 2500 3588 2508
rect 4140 2496 4148 2504
rect 4156 2496 4164 2504
rect 4172 2496 4180 2504
rect 4236 2496 4244 2504
rect 4396 2496 4404 2504
rect 4412 2496 4420 2504
rect 4732 2496 4740 2504
rect 5020 2496 5028 2504
rect 5116 2496 5124 2504
rect 5388 2496 5396 2504
rect 5532 2496 5540 2504
rect 5964 2500 5972 2508
rect 348 2476 356 2484
rect 3244 2476 3252 2484
rect 3436 2476 3444 2484
rect 3932 2476 3940 2484
rect 4204 2476 4212 2484
rect 4492 2476 4500 2484
rect 4764 2476 4772 2484
rect 5084 2476 5092 2484
rect 460 2454 468 2462
rect 1212 2454 1220 2462
rect 1708 2454 1716 2462
rect 3580 2454 3588 2462
rect 3916 2456 3924 2464
rect 5964 2454 5972 2462
rect 44 2436 52 2444
rect 332 2436 340 2444
rect 716 2436 724 2444
rect 860 2436 868 2444
rect 956 2436 964 2444
rect 1292 2436 1300 2444
rect 1452 2436 1460 2444
rect 2012 2436 2020 2444
rect 2268 2436 2276 2444
rect 2444 2436 2452 2444
rect 2508 2436 2516 2444
rect 2796 2436 2804 2444
rect 3132 2436 3140 2444
rect 3164 2436 3172 2444
rect 3292 2436 3300 2444
rect 3420 2436 3428 2444
rect 3836 2436 3844 2444
rect 4812 2436 4820 2444
rect 4844 2436 4852 2444
rect 5036 2436 5044 2444
rect 5068 2436 5076 2444
rect 5500 2436 5508 2444
rect 5660 2436 5668 2444
rect 1502 2406 1510 2414
rect 1516 2406 1524 2414
rect 1530 2406 1538 2414
rect 4574 2406 4582 2414
rect 4588 2406 4596 2414
rect 4602 2406 4610 2414
rect 220 2376 228 2384
rect 476 2376 484 2384
rect 1820 2376 1828 2384
rect 1868 2376 1876 2384
rect 1916 2376 1924 2384
rect 2204 2376 2212 2384
rect 2348 2376 2356 2384
rect 2860 2376 2868 2384
rect 3196 2376 3204 2384
rect 3260 2376 3268 2384
rect 3404 2376 3412 2384
rect 4188 2376 4196 2384
rect 4732 2376 4740 2384
rect 4908 2376 4916 2384
rect 5132 2376 5140 2384
rect 5244 2376 5252 2384
rect 5356 2376 5364 2384
rect 5548 2376 5556 2384
rect 5580 2376 5588 2384
rect 5980 2376 5988 2384
rect 1564 2358 1572 2366
rect 3532 2356 3540 2364
rect 3740 2358 3748 2366
rect 5068 2356 5076 2364
rect 5308 2356 5316 2364
rect 156 2336 164 2344
rect 300 2336 308 2344
rect 780 2336 788 2344
rect 828 2336 836 2344
rect 3212 2336 3220 2344
rect 3420 2336 3428 2344
rect 3484 2336 3492 2344
rect 3516 2336 3524 2344
rect 3996 2336 4004 2344
rect 4620 2336 4628 2344
rect 4668 2336 4676 2344
rect 4748 2336 4756 2344
rect 4876 2336 4884 2344
rect 4924 2336 4932 2344
rect 5084 2336 5092 2344
rect 5116 2336 5124 2344
rect 5196 2336 5204 2344
rect 5260 2336 5268 2344
rect 5308 2336 5316 2344
rect 5372 2336 5380 2344
rect 5436 2336 5444 2344
rect 5596 2336 5604 2344
rect 124 2316 132 2324
rect 188 2316 196 2324
rect 252 2316 260 2324
rect 332 2316 340 2324
rect 364 2316 372 2324
rect 476 2316 484 2324
rect 1244 2316 1252 2324
rect 1276 2316 1284 2324
rect 1564 2312 1572 2320
rect 1916 2316 1924 2324
rect 2348 2316 2356 2324
rect 2668 2316 2676 2324
rect 2716 2316 2724 2324
rect 2796 2316 2804 2324
rect 2892 2316 2900 2324
rect 2972 2316 2980 2324
rect 3004 2316 3012 2324
rect 3052 2316 3060 2324
rect 3132 2316 3140 2324
rect 3164 2316 3172 2324
rect 3180 2316 3188 2324
rect 3388 2316 3396 2324
rect 3468 2316 3476 2324
rect 3516 2316 3524 2324
rect 3740 2312 3748 2320
rect 4060 2316 4068 2324
rect 4076 2316 4084 2324
rect 4700 2316 4708 2324
rect 4716 2316 4724 2324
rect 4780 2316 4788 2324
rect 4812 2316 4820 2324
rect 4956 2316 4964 2324
rect 5084 2316 5092 2324
rect 5148 2316 5156 2324
rect 5180 2316 5188 2324
rect 5228 2316 5236 2324
rect 5292 2316 5300 2324
rect 5404 2316 5412 2324
rect 5468 2316 5476 2324
rect 5484 2316 5492 2324
rect 5628 2316 5636 2324
rect 5980 2316 5988 2324
rect 6044 2316 6052 2324
rect 6076 2316 6084 2324
rect 92 2296 100 2304
rect 140 2296 148 2304
rect 156 2296 164 2304
rect 220 2296 228 2304
rect 332 2296 340 2304
rect 476 2296 484 2304
rect 684 2296 692 2304
rect 766 2296 774 2304
rect 988 2296 996 2304
rect 1148 2296 1156 2304
rect 1292 2296 1300 2304
rect 1308 2296 1316 2304
rect 1340 2296 1348 2304
rect 1740 2296 1748 2304
rect 2124 2296 2132 2304
rect 2444 2296 2452 2304
rect 2556 2296 2564 2304
rect 2652 2296 2660 2304
rect 2764 2296 2772 2304
rect 2828 2296 2836 2304
rect 2876 2296 2884 2304
rect 2956 2296 2964 2304
rect 2972 2296 2980 2304
rect 3116 2296 3124 2304
rect 3196 2296 3204 2304
rect 3404 2296 3412 2304
rect 3468 2296 3476 2304
rect 3532 2296 3540 2304
rect 3580 2296 3588 2304
rect 3596 2296 3604 2304
rect 3644 2296 3652 2304
rect 3708 2296 3716 2304
rect 4012 2296 4020 2304
rect 4108 2296 4116 2304
rect 4460 2296 4468 2304
rect 4492 2296 4500 2304
rect 4524 2296 4532 2304
rect 4540 2296 4548 2304
rect 4572 2296 4580 2304
rect 4604 2296 4612 2304
rect 4700 2296 4708 2304
rect 4732 2296 4740 2304
rect 4828 2296 4836 2304
rect 4892 2296 4900 2304
rect 4940 2296 4948 2304
rect 4972 2296 4980 2304
rect 5020 2296 5028 2304
rect 5068 2296 5076 2304
rect 5132 2296 5140 2304
rect 5164 2296 5172 2304
rect 5180 2296 5188 2304
rect 5244 2296 5252 2304
rect 5308 2296 5316 2304
rect 5388 2296 5396 2304
rect 5420 2296 5428 2304
rect 5452 2296 5460 2304
rect 5580 2296 5588 2304
rect 5628 2296 5636 2304
rect 5772 2296 5780 2304
rect 6044 2296 6052 2304
rect 28 2276 36 2284
rect 76 2276 84 2284
rect 140 2276 148 2284
rect 204 2276 212 2284
rect 268 2276 276 2284
rect 316 2276 324 2284
rect 428 2276 436 2284
rect 572 2276 580 2284
rect 828 2276 836 2284
rect 844 2276 852 2284
rect 1020 2276 1028 2284
rect 1068 2276 1076 2284
rect 12 2256 20 2264
rect 44 2256 52 2264
rect 60 2256 68 2264
rect 396 2256 404 2264
rect 412 2256 420 2264
rect 604 2256 612 2264
rect 1356 2276 1364 2284
rect 1388 2276 1396 2284
rect 1628 2276 1636 2284
rect 2012 2276 2020 2284
rect 2300 2276 2308 2284
rect 2444 2276 2452 2284
rect 2638 2276 2646 2284
rect 2748 2276 2756 2284
rect 2844 2276 2852 2284
rect 2940 2276 2948 2284
rect 2956 2276 2964 2284
rect 3020 2276 3028 2284
rect 3036 2276 3044 2284
rect 3116 2276 3124 2284
rect 3372 2276 3380 2284
rect 3484 2276 3492 2284
rect 3660 2276 3668 2284
rect 3804 2276 3812 2284
rect 4092 2276 4100 2284
rect 4156 2276 4164 2284
rect 4300 2276 4308 2284
rect 4476 2276 4484 2284
rect 4508 2276 4516 2284
rect 4556 2276 4564 2284
rect 4588 2276 4596 2284
rect 4668 2276 4676 2284
rect 4780 2276 4788 2284
rect 4812 2276 4820 2284
rect 4876 2276 4884 2284
rect 5004 2276 5012 2284
rect 5196 2276 5204 2284
rect 5516 2276 5524 2284
rect 5532 2276 5540 2284
rect 5660 2276 5668 2284
rect 5884 2276 5892 2284
rect 6028 2276 6036 2284
rect 1436 2256 1444 2264
rect 1660 2256 1668 2264
rect 1852 2256 1860 2264
rect 2044 2256 2052 2264
rect 2252 2256 2260 2264
rect 2476 2256 2484 2264
rect 2876 2256 2884 2264
rect 3836 2256 3844 2264
rect 4044 2256 4052 2264
rect 4972 2256 4980 2264
rect 5852 2256 5860 2264
rect 284 2236 292 2244
rect 380 2236 388 2244
rect 956 2236 964 2244
rect 1228 2236 1236 2244
rect 1324 2236 1332 2244
rect 2204 2236 2212 2244
rect 2796 2236 2804 2244
rect 3260 2236 3268 2244
rect 4428 2236 4436 2244
rect 5484 2236 5492 2244
rect 5692 2236 5700 2244
rect 3038 2206 3046 2214
rect 3052 2206 3060 2214
rect 3066 2206 3074 2214
rect 668 2176 676 2184
rect 1164 2176 1172 2184
rect 1724 2176 1732 2184
rect 2444 2176 2452 2184
rect 2492 2176 2500 2184
rect 3100 2176 3108 2184
rect 3516 2176 3524 2184
rect 4012 2176 4020 2184
rect 4812 2176 4820 2184
rect 5196 2176 5204 2184
rect 5340 2176 5348 2184
rect 5388 2176 5396 2184
rect 6044 2176 6052 2184
rect 12 2156 20 2164
rect 156 2156 164 2164
rect 748 2156 756 2164
rect 924 2156 932 2164
rect 1500 2156 1508 2164
rect 1580 2156 1588 2164
rect 1948 2156 1956 2164
rect 2284 2156 2292 2164
rect 2460 2156 2468 2164
rect 2668 2156 2676 2164
rect 2844 2156 2852 2164
rect 2876 2156 2884 2164
rect 3260 2156 3268 2164
rect 3676 2156 3684 2164
rect 3868 2156 3876 2164
rect 4108 2156 4116 2164
rect 4428 2156 4436 2164
rect 4652 2156 4660 2164
rect 4684 2156 4692 2164
rect 4716 2156 4724 2164
rect 4748 2156 4756 2164
rect 4780 2156 4788 2164
rect 5036 2156 5044 2164
rect 5228 2156 5236 2164
rect 5548 2156 5556 2164
rect 140 2136 148 2144
rect 236 2136 244 2144
rect 332 2136 340 2144
rect 396 2136 404 2144
rect 556 2136 564 2144
rect 988 2136 996 2144
rect 1020 2136 1028 2144
rect 1100 2136 1108 2144
rect 1116 2136 1124 2144
rect 1244 2136 1252 2144
rect 1356 2136 1364 2144
rect 1644 2136 1652 2144
rect 1660 2136 1668 2144
rect 1756 2136 1764 2144
rect 1980 2136 1988 2144
rect 2252 2136 2260 2144
rect 2636 2136 2644 2144
rect 3020 2136 3028 2144
rect 3292 2136 3300 2144
rect 3436 2136 3444 2144
rect 3500 2136 3508 2144
rect 3708 2136 3716 2144
rect 3852 2136 3860 2144
rect 3900 2136 3908 2144
rect 4108 2136 4116 2144
rect 4204 2136 4212 2144
rect 4252 2136 4260 2144
rect 4460 2136 4468 2144
rect 4860 2136 4868 2144
rect 5004 2136 5012 2144
rect 5260 2136 5268 2144
rect 5356 2136 5364 2144
rect 5580 2136 5588 2144
rect 5724 2136 5732 2144
rect 5788 2136 5796 2144
rect 5916 2136 5924 2144
rect 60 2116 68 2124
rect 92 2116 100 2124
rect 188 2116 196 2124
rect 300 2116 308 2124
rect 348 2116 356 2124
rect 380 2116 388 2124
rect 412 2116 420 2124
rect 684 2116 692 2124
rect 716 2116 724 2124
rect 764 2116 772 2124
rect 780 2116 788 2124
rect 924 2118 932 2126
rect 1004 2116 1012 2124
rect 92 2096 100 2104
rect 188 2096 196 2104
rect 220 2096 228 2104
rect 268 2096 276 2104
rect 284 2096 292 2104
rect 348 2096 356 2104
rect 1084 2116 1092 2124
rect 1132 2116 1140 2124
rect 1052 2096 1060 2104
rect 1212 2116 1220 2124
rect 1260 2116 1268 2124
rect 1180 2096 1188 2104
rect 1292 2096 1300 2104
rect 1340 2116 1348 2124
rect 1484 2116 1492 2124
rect 1644 2116 1652 2124
rect 2044 2116 2052 2124
rect 2156 2116 2164 2124
rect 2556 2116 2564 2124
rect 2748 2116 2756 2124
rect 3180 2116 3188 2124
rect 3404 2116 3412 2124
rect 3452 2116 3460 2124
rect 3788 2116 3796 2124
rect 3980 2116 3988 2124
rect 4028 2116 4036 2124
rect 4140 2116 4148 2124
rect 4348 2116 4356 2124
rect 4844 2116 4852 2124
rect 5116 2116 5124 2124
rect 5276 2116 5284 2124
rect 1340 2096 1348 2104
rect 2076 2096 2084 2104
rect 2156 2096 2164 2104
rect 2572 2100 2580 2108
rect 3388 2096 3396 2104
rect 3772 2100 3780 2108
rect 3884 2096 3892 2104
rect 4108 2096 4116 2104
rect 4236 2096 4244 2104
rect 4268 2096 4276 2104
rect 4524 2100 4532 2108
rect 4940 2100 4948 2108
rect 5308 2096 5316 2104
rect 5676 2116 5684 2124
rect 5740 2116 5748 2124
rect 5756 2116 5764 2124
rect 5644 2100 5652 2108
rect 5772 2096 5780 2104
rect 252 2076 260 2084
rect 796 2076 804 2084
rect 1372 2076 1380 2084
rect 2828 2056 2836 2064
rect 4524 2054 4532 2062
rect 4940 2054 4948 2062
rect 5644 2054 5652 2062
rect 60 2036 68 2044
rect 380 2036 388 2044
rect 1788 2036 1796 2044
rect 2076 2036 2084 2044
rect 2156 2036 2164 2044
rect 2444 2036 2452 2044
rect 2572 2036 2580 2044
rect 2908 2036 2916 2044
rect 3100 2036 3108 2044
rect 3388 2036 3396 2044
rect 3772 2036 3780 2044
rect 3916 2036 3924 2044
rect 4124 2036 4132 2044
rect 4172 2036 4180 2044
rect 4668 2036 4676 2044
rect 4700 2036 4708 2044
rect 4732 2036 4740 2044
rect 4764 2036 4772 2044
rect 4796 2036 4804 2044
rect 1502 2006 1510 2014
rect 1516 2006 1524 2014
rect 1530 2006 1538 2014
rect 4574 2006 4582 2014
rect 4588 2006 4596 2014
rect 4602 2006 4610 2014
rect 44 1976 52 1984
rect 332 1976 340 1984
rect 828 1976 836 1984
rect 1164 1976 1172 1984
rect 1324 1976 1332 1984
rect 1420 1976 1428 1984
rect 1452 1976 1460 1984
rect 1580 1976 1588 1984
rect 2028 1976 2036 1984
rect 2092 1976 2100 1984
rect 2588 1976 2596 1984
rect 3004 1976 3012 1984
rect 3100 1976 3108 1984
rect 3244 1976 3252 1984
rect 3948 1976 3956 1984
rect 4380 1976 4388 1984
rect 5580 1976 5588 1984
rect 572 1956 580 1964
rect 3500 1958 3508 1966
rect 4060 1958 4068 1966
rect 5692 1958 5700 1966
rect 2172 1936 2180 1944
rect 2364 1936 2372 1944
rect 2444 1936 2452 1944
rect 2876 1936 2884 1944
rect 3580 1936 3588 1944
rect 3660 1936 3668 1944
rect 4892 1936 4900 1944
rect 5036 1936 5044 1944
rect 44 1916 52 1924
rect 588 1916 596 1924
rect 668 1916 676 1924
rect 700 1916 708 1924
rect 1084 1916 1092 1924
rect 1116 1916 1124 1924
rect 1228 1916 1236 1924
rect 2028 1916 2036 1924
rect 2076 1916 2084 1924
rect 2476 1916 2484 1924
rect 2588 1916 2596 1924
rect 2892 1916 2900 1924
rect 3500 1912 3508 1920
rect 3948 1916 3956 1924
rect 4060 1912 4068 1920
rect 4380 1916 4388 1924
rect 4988 1916 4996 1924
rect 5004 1916 5012 1924
rect 5100 1916 5108 1924
rect 5180 1916 5188 1924
rect 5580 1916 5588 1924
rect 5692 1912 5700 1920
rect 5980 1916 5988 1924
rect 252 1896 260 1904
rect 476 1896 484 1904
rect 588 1896 596 1904
rect 620 1896 628 1904
rect 668 1896 676 1904
rect 732 1896 740 1904
rect 780 1896 788 1904
rect 796 1896 804 1904
rect 860 1896 868 1904
rect 940 1896 948 1904
rect 1084 1896 1092 1904
rect 1132 1896 1140 1904
rect 1148 1896 1156 1904
rect 1196 1896 1204 1904
rect 1212 1896 1220 1904
rect 1260 1896 1268 1904
rect 1292 1896 1300 1904
rect 1308 1896 1316 1904
rect 1356 1896 1364 1904
rect 1388 1896 1396 1904
rect 1516 1896 1524 1904
rect 1724 1896 1732 1904
rect 1820 1896 1828 1904
rect 2044 1896 2052 1904
rect 2140 1896 2148 1904
rect 2188 1896 2196 1904
rect 2332 1896 2340 1904
rect 2348 1896 2356 1904
rect 2396 1896 2404 1904
rect 2540 1896 2548 1904
rect 2588 1896 2596 1904
rect 2940 1896 2948 1904
rect 2956 1896 2964 1904
rect 3132 1896 3140 1904
rect 3148 1896 3156 1904
rect 3180 1896 3188 1904
rect 3324 1896 3332 1904
rect 3612 1896 3620 1904
rect 3740 1896 3748 1904
rect 3964 1896 3972 1904
rect 4044 1896 4052 1904
rect 4380 1896 4388 1904
rect 4796 1894 4804 1902
rect 4956 1896 4964 1904
rect 5132 1896 5140 1904
rect 5372 1896 5380 1904
rect 5596 1896 5604 1904
rect 5660 1896 5668 1904
rect 5950 1896 5958 1904
rect 6012 1896 6020 1904
rect 6028 1896 6036 1904
rect 140 1876 148 1884
rect 412 1876 420 1884
rect 636 1876 644 1884
rect 652 1876 660 1884
rect 716 1876 724 1884
rect 892 1876 900 1884
rect 1068 1876 1076 1884
rect 1276 1876 1284 1884
rect 1612 1876 1620 1884
rect 1708 1876 1716 1884
rect 1932 1876 1940 1884
rect 2108 1876 2116 1884
rect 2124 1876 2132 1884
rect 2156 1876 2164 1884
rect 2236 1876 2244 1884
rect 2300 1876 2308 1884
rect 2316 1876 2324 1884
rect 2380 1876 2388 1884
rect 2476 1876 2484 1884
rect 2492 1876 2500 1884
rect 2684 1876 2692 1884
rect 2956 1876 2964 1884
rect 3004 1876 3012 1884
rect 3164 1876 3172 1884
rect 3436 1876 3444 1884
rect 3644 1876 3652 1884
rect 3852 1876 3860 1884
rect 4124 1876 4132 1884
rect 4476 1876 4484 1884
rect 4812 1876 4820 1884
rect 4940 1876 4948 1884
rect 5036 1876 5044 1884
rect 5116 1876 5124 1884
rect 5196 1876 5204 1884
rect 5228 1876 5236 1884
rect 5484 1876 5492 1884
rect 5756 1876 5764 1884
rect 6028 1876 6036 1884
rect 6124 1876 6132 1884
rect 172 1856 180 1864
rect 380 1856 388 1864
rect 1468 1856 1476 1864
rect 1500 1856 1508 1864
rect 1596 1856 1604 1864
rect 1900 1856 1908 1864
rect 2716 1856 2724 1864
rect 3084 1856 3092 1864
rect 3116 1856 3124 1864
rect 3404 1856 3412 1864
rect 3820 1856 3828 1864
rect 4156 1856 4164 1864
rect 4508 1856 4516 1864
rect 5164 1856 5172 1864
rect 5260 1856 5268 1864
rect 5452 1856 5460 1864
rect 5788 1856 5796 1864
rect 364 1836 372 1844
rect 828 1836 836 1844
rect 1052 1836 1060 1844
rect 1452 1836 1460 1844
rect 1564 1836 1572 1844
rect 2252 1836 2260 1844
rect 2908 1836 2916 1844
rect 3212 1836 3220 1844
rect 3580 1836 3588 1844
rect 4316 1836 4324 1844
rect 4668 1836 4676 1844
rect 4924 1836 4932 1844
rect 4988 1836 4996 1844
rect 5148 1836 5156 1844
rect 5292 1836 5300 1844
rect 5980 1836 5988 1844
rect 3038 1806 3046 1814
rect 3052 1806 3060 1814
rect 3066 1806 3074 1814
rect 380 1776 388 1784
rect 524 1776 532 1784
rect 1020 1776 1028 1784
rect 1212 1776 1220 1784
rect 1324 1776 1332 1784
rect 1932 1776 1940 1784
rect 2748 1776 2756 1784
rect 3404 1776 3412 1784
rect 3628 1776 3636 1784
rect 3740 1776 3748 1784
rect 3804 1776 3812 1784
rect 3852 1776 3860 1784
rect 5100 1776 5108 1784
rect 5500 1776 5508 1784
rect 5548 1776 5556 1784
rect 60 1756 68 1764
rect 508 1756 516 1764
rect 764 1756 772 1764
rect 940 1756 948 1764
rect 1068 1756 1076 1764
rect 1148 1756 1156 1764
rect 1180 1756 1188 1764
rect 1260 1756 1268 1764
rect 1292 1756 1300 1764
rect 1372 1756 1380 1764
rect 1452 1756 1460 1764
rect 1676 1756 1684 1764
rect 2252 1756 2260 1764
rect 2588 1756 2596 1764
rect 3180 1756 3188 1764
rect 3500 1756 3508 1764
rect 252 1736 260 1744
rect 476 1736 484 1744
rect 684 1736 692 1744
rect 812 1736 820 1744
rect 924 1736 932 1744
rect 1100 1736 1108 1744
rect 4108 1756 4116 1764
rect 5212 1756 5220 1764
rect 5516 1756 5524 1764
rect 5820 1756 5828 1764
rect 6124 1756 6132 1764
rect 1708 1736 1716 1744
rect 1852 1736 1860 1744
rect 1948 1736 1956 1744
rect 2060 1736 2068 1744
rect 2284 1736 2292 1744
rect 2556 1736 2564 1744
rect 2764 1736 2772 1744
rect 2812 1736 2820 1744
rect 2972 1736 2980 1744
rect 3148 1736 3156 1744
rect 3372 1736 3380 1744
rect 3436 1736 3444 1744
rect 3468 1736 3476 1744
rect 3484 1736 3492 1744
rect 3564 1736 3572 1744
rect 3580 1736 3588 1744
rect 3644 1736 3652 1744
rect 3692 1736 3700 1744
rect 3772 1736 3780 1744
rect 4012 1736 4020 1744
rect 4044 1736 4052 1744
rect 4156 1736 4164 1744
rect 4172 1736 4180 1744
rect 4332 1736 4340 1744
rect 4460 1736 4468 1744
rect 4572 1736 4580 1744
rect 4700 1736 4708 1744
rect 4764 1736 4772 1744
rect 4780 1736 4788 1744
rect 5020 1736 5028 1744
rect 5052 1736 5060 1744
rect 5164 1736 5172 1744
rect 5372 1736 5380 1744
rect 5436 1736 5444 1744
rect 5516 1736 5524 1744
rect 5580 1736 5588 1744
rect 5852 1736 5860 1744
rect 5996 1736 6004 1744
rect 92 1716 100 1724
rect 204 1716 212 1724
rect 236 1716 244 1724
rect 268 1716 276 1724
rect 284 1716 292 1724
rect 316 1716 324 1724
rect 332 1716 340 1724
rect 412 1716 420 1724
rect 652 1718 660 1726
rect 732 1716 740 1724
rect 780 1716 788 1724
rect 796 1716 804 1724
rect 828 1716 836 1724
rect 204 1696 212 1704
rect 428 1696 436 1704
rect 828 1696 836 1704
rect 908 1716 916 1724
rect 972 1716 980 1724
rect 988 1716 996 1724
rect 1036 1716 1044 1724
rect 1052 1716 1060 1724
rect 1292 1716 1300 1724
rect 1356 1716 1364 1724
rect 1404 1716 1412 1724
rect 1804 1716 1812 1724
rect 1900 1716 1908 1724
rect 2012 1716 2020 1724
rect 2044 1716 2052 1724
rect 2380 1716 2388 1724
rect 2492 1716 2500 1724
rect 3260 1716 3268 1724
rect 3452 1716 3460 1724
rect 3532 1716 3540 1724
rect 3660 1716 3668 1724
rect 3708 1716 3716 1724
rect 3980 1718 3988 1726
rect 4060 1716 4068 1724
rect 876 1696 884 1704
rect 1132 1696 1140 1704
rect 1212 1696 1220 1704
rect 1804 1696 1812 1704
rect 1916 1696 1924 1704
rect 1964 1696 1972 1704
rect 2012 1696 2020 1704
rect 2092 1696 2100 1704
rect 2348 1700 2356 1708
rect 2460 1696 2468 1704
rect 2780 1696 2788 1704
rect 3084 1700 3092 1708
rect 3340 1696 3348 1704
rect 3404 1696 3412 1704
rect 3420 1696 3428 1704
rect 3516 1696 3524 1704
rect 3628 1696 3636 1704
rect 3692 1696 3700 1704
rect 3804 1696 3812 1704
rect 4092 1696 4100 1704
rect 4140 1716 4148 1724
rect 4172 1716 4180 1724
rect 4236 1716 4244 1724
rect 4252 1716 4260 1724
rect 4332 1716 4340 1724
rect 4476 1716 4484 1724
rect 4492 1716 4500 1724
rect 4636 1716 4644 1724
rect 4716 1716 4724 1724
rect 4748 1716 4756 1724
rect 4828 1716 4836 1724
rect 4844 1716 4852 1724
rect 4972 1716 4980 1724
rect 5068 1716 5076 1724
rect 4524 1696 4532 1704
rect 4652 1696 4660 1704
rect 4684 1696 4692 1704
rect 4748 1696 4756 1704
rect 5148 1716 5156 1724
rect 5180 1716 5188 1724
rect 5196 1716 5204 1724
rect 5244 1716 5252 1724
rect 5276 1716 5284 1724
rect 5292 1716 5300 1724
rect 5340 1716 5348 1724
rect 5388 1716 5396 1724
rect 5404 1716 5412 1724
rect 5452 1716 5460 1724
rect 5596 1716 5604 1724
rect 5644 1716 5652 1724
rect 5740 1716 5748 1724
rect 5948 1716 5956 1724
rect 6028 1716 6036 1724
rect 5116 1696 5124 1704
rect 5420 1696 5428 1704
rect 5452 1696 5460 1704
rect 5484 1696 5492 1704
rect 5564 1696 5572 1704
rect 5628 1696 5636 1704
rect 5916 1700 5924 1708
rect 5996 1696 6004 1704
rect 188 1676 196 1684
rect 1100 1676 1108 1684
rect 3836 1676 3844 1684
rect 4860 1676 4868 1684
rect 4892 1676 4900 1684
rect 1516 1656 1524 1664
rect 2348 1654 2356 1662
rect 3084 1654 3092 1662
rect 380 1636 388 1644
rect 460 1636 468 1644
rect 1116 1636 1124 1644
rect 1164 1636 1172 1644
rect 1196 1636 1204 1644
rect 1388 1636 1396 1644
rect 1404 1636 1412 1644
rect 1804 1636 1812 1644
rect 2460 1636 2468 1644
rect 2844 1636 2852 1644
rect 4444 1636 4452 1644
rect 5324 1636 5332 1644
rect 5916 1636 5924 1644
rect 1502 1606 1510 1614
rect 1516 1606 1524 1614
rect 1530 1606 1538 1614
rect 4574 1606 4582 1614
rect 4588 1606 4596 1614
rect 4602 1606 4610 1614
rect 236 1576 244 1584
rect 1372 1576 1380 1584
rect 1516 1576 1524 1584
rect 1932 1576 1940 1584
rect 2684 1576 2692 1584
rect 3740 1576 3748 1584
rect 3804 1576 3812 1584
rect 4460 1576 4468 1584
rect 4796 1576 4804 1584
rect 5420 1576 5428 1584
rect 5980 1576 5988 1584
rect 1676 1558 1684 1566
rect 2316 1558 2324 1566
rect 2572 1556 2580 1564
rect 3260 1558 3268 1566
rect 4028 1556 4036 1564
rect 4604 1556 4612 1564
rect 892 1536 900 1544
rect 940 1536 948 1544
rect 1068 1536 1076 1544
rect 1116 1536 1124 1544
rect 2236 1536 2244 1544
rect 2988 1536 2996 1544
rect 3516 1536 3524 1544
rect 3580 1536 3588 1544
rect 3980 1536 3988 1544
rect 4044 1536 4052 1544
rect 4876 1536 4884 1544
rect 5164 1536 5172 1544
rect 5196 1536 5204 1544
rect 5452 1536 5460 1544
rect 5676 1536 5684 1544
rect 6124 1536 6132 1544
rect 204 1516 212 1524
rect 316 1516 324 1524
rect 76 1496 84 1504
rect 284 1496 292 1504
rect 636 1516 644 1524
rect 364 1496 372 1504
rect 396 1496 404 1504
rect 460 1496 468 1504
rect 476 1496 484 1504
rect 508 1496 516 1504
rect 556 1496 564 1504
rect 572 1496 580 1504
rect 604 1496 612 1504
rect 956 1516 964 1524
rect 1020 1516 1028 1524
rect 1036 1516 1044 1524
rect 1084 1516 1092 1524
rect 1148 1516 1156 1524
rect 1164 1516 1172 1524
rect 1276 1516 1284 1524
rect 1308 1516 1316 1524
rect 1340 1516 1348 1524
rect 1404 1516 1412 1524
rect 1676 1512 1684 1520
rect 2140 1516 2148 1524
rect 2316 1512 2324 1520
rect 2604 1516 2612 1524
rect 2684 1516 2692 1524
rect 3148 1516 3156 1524
rect 3180 1516 3188 1524
rect 3260 1512 3268 1520
rect 3548 1516 3556 1524
rect 3692 1516 3700 1524
rect 3708 1516 3716 1524
rect 3772 1516 3780 1524
rect 3852 1516 3860 1524
rect 3884 1516 3892 1524
rect 3900 1516 3908 1524
rect 3964 1516 3972 1524
rect 4012 1516 4020 1524
rect 4076 1516 4084 1524
rect 4140 1516 4148 1524
rect 668 1496 676 1504
rect 684 1496 692 1504
rect 764 1494 772 1502
rect 924 1496 932 1504
rect 988 1496 996 1504
rect 1052 1496 1060 1504
rect 1116 1496 1124 1504
rect 1180 1496 1188 1504
rect 1196 1496 1204 1504
rect 1244 1496 1252 1504
rect 1276 1496 1284 1504
rect 60 1476 68 1484
rect 268 1476 276 1484
rect 332 1476 340 1484
rect 380 1476 388 1484
rect 396 1476 404 1484
rect 588 1476 596 1484
rect 700 1476 708 1484
rect 732 1476 740 1484
rect 972 1476 980 1484
rect 1100 1476 1108 1484
rect 1212 1476 1220 1484
rect 1228 1476 1236 1484
rect 1276 1476 1284 1484
rect 1308 1496 1316 1504
rect 1372 1496 1380 1504
rect 1852 1496 1860 1504
rect 2012 1496 2020 1504
rect 2076 1496 2084 1504
rect 2092 1496 2100 1504
rect 2140 1496 2148 1504
rect 2204 1496 2212 1504
rect 2380 1496 2388 1504
rect 2492 1496 2500 1504
rect 2668 1496 2676 1504
rect 2892 1496 2900 1504
rect 3100 1496 3108 1504
rect 3324 1496 3332 1504
rect 3436 1496 3444 1504
rect 3628 1496 3636 1504
rect 3740 1496 3748 1504
rect 3804 1496 3812 1504
rect 3852 1496 3860 1504
rect 3932 1496 3940 1504
rect 3996 1496 4004 1504
rect 4060 1496 4068 1504
rect 4108 1496 4116 1504
rect 4316 1516 4324 1524
rect 4508 1516 4516 1524
rect 4956 1516 4964 1524
rect 1356 1476 1364 1484
rect 1420 1476 1428 1484
rect 1548 1476 1556 1484
rect 1740 1476 1748 1484
rect 2172 1476 2180 1484
rect 2188 1476 2196 1484
rect 2220 1476 2228 1484
rect 2380 1476 2388 1484
rect 2636 1476 2644 1484
rect 2780 1476 2788 1484
rect 2988 1476 2996 1484
rect 540 1456 548 1464
rect 764 1456 772 1464
rect 1772 1456 1780 1464
rect 2044 1456 2052 1464
rect 2124 1456 2132 1464
rect 2412 1456 2420 1464
rect 2812 1456 2820 1464
rect 3084 1476 3092 1484
rect 3324 1476 3332 1484
rect 3548 1476 3556 1484
rect 3644 1476 3652 1484
rect 3660 1476 3668 1484
rect 3756 1476 3764 1484
rect 3820 1476 3828 1484
rect 3836 1476 3844 1484
rect 3900 1476 3908 1484
rect 3948 1476 3956 1484
rect 4092 1476 4100 1484
rect 4172 1476 4180 1484
rect 4204 1476 4212 1484
rect 4236 1496 4244 1504
rect 4284 1496 4292 1504
rect 4300 1496 4308 1504
rect 4348 1496 4356 1504
rect 4412 1496 4420 1504
rect 4428 1496 4436 1504
rect 4476 1496 4484 1504
rect 4492 1496 4500 1504
rect 4716 1496 4724 1504
rect 4828 1496 4836 1504
rect 4844 1496 4852 1504
rect 4892 1496 4900 1504
rect 5004 1496 5012 1504
rect 5052 1496 5060 1504
rect 5100 1516 5108 1524
rect 5404 1516 5412 1524
rect 5980 1516 5988 1524
rect 5132 1496 5140 1504
rect 5276 1496 5284 1504
rect 5372 1496 5380 1504
rect 5404 1496 5412 1504
rect 5500 1496 5508 1504
rect 5948 1496 5956 1504
rect 5980 1496 5988 1504
rect 6060 1496 6068 1504
rect 4540 1476 4548 1484
rect 4764 1476 4772 1484
rect 4924 1476 4932 1484
rect 5020 1476 5028 1484
rect 5036 1476 5044 1484
rect 5084 1476 5092 1484
rect 5148 1476 5156 1484
rect 5324 1476 5332 1484
rect 5356 1476 5364 1484
rect 5532 1476 5540 1484
rect 5628 1476 5636 1484
rect 5884 1476 5892 1484
rect 3356 1456 3364 1464
rect 4396 1456 4404 1464
rect 4812 1456 4820 1464
rect 5292 1456 5300 1464
rect 5612 1456 5620 1464
rect 5852 1456 5860 1464
rect 6044 1456 6052 1464
rect 188 1436 196 1444
rect 1020 1436 1028 1444
rect 1436 1436 1444 1444
rect 1964 1436 1972 1444
rect 2108 1436 2116 1444
rect 2156 1436 2164 1444
rect 2620 1436 2628 1444
rect 2972 1436 2980 1444
rect 3180 1436 3188 1444
rect 3692 1436 3700 1444
rect 4316 1436 4324 1444
rect 4972 1436 4980 1444
rect 5692 1436 5700 1444
rect 6028 1436 6036 1444
rect 3038 1406 3046 1414
rect 3052 1406 3060 1414
rect 3066 1406 3074 1414
rect 956 1376 964 1384
rect 1228 1376 1236 1384
rect 1612 1376 1620 1384
rect 1980 1376 1988 1384
rect 4556 1376 4564 1384
rect 5068 1376 5076 1384
rect 5180 1376 5188 1384
rect 5596 1376 5604 1384
rect 5852 1376 5860 1384
rect 6076 1376 6084 1384
rect 188 1356 196 1364
rect 412 1356 420 1364
rect 1260 1356 1268 1364
rect 1388 1356 1396 1364
rect 1804 1356 1812 1364
rect 2268 1356 2276 1364
rect 2476 1356 2484 1364
rect 2492 1356 2500 1364
rect 2844 1356 2852 1364
rect 3372 1356 3380 1364
rect 3548 1356 3556 1364
rect 3596 1356 3604 1364
rect 3948 1356 3956 1364
rect 4476 1356 4484 1364
rect 4700 1356 4708 1364
rect 220 1336 228 1344
rect 364 1336 372 1344
rect 460 1336 468 1344
rect 572 1336 580 1344
rect 684 1336 692 1344
rect 764 1336 772 1344
rect 892 1336 900 1344
rect 1004 1336 1012 1344
rect 1036 1336 1044 1344
rect 1212 1336 1220 1344
rect 1276 1336 1284 1344
rect 1292 1336 1300 1344
rect 1340 1336 1348 1344
rect 1404 1336 1412 1344
rect 1500 1336 1508 1344
rect 1564 1336 1572 1344
rect 1836 1336 1844 1344
rect 2012 1336 2020 1344
rect 2028 1336 2036 1344
rect 2300 1336 2308 1344
rect 2444 1336 2452 1344
rect 2604 1336 2612 1344
rect 2636 1336 2644 1344
rect 2876 1336 2884 1344
rect 3196 1336 3204 1344
rect 3340 1336 3348 1344
rect 3628 1336 3636 1344
rect 3676 1336 3684 1344
rect 3772 1336 3780 1344
rect 3916 1336 3924 1344
rect 4140 1336 4148 1344
rect 4268 1336 4276 1344
rect 4332 1336 4340 1344
rect 4380 1336 4388 1344
rect 4732 1356 4740 1364
rect 5452 1356 5460 1364
rect 5564 1356 5572 1364
rect 5612 1356 5620 1364
rect 4764 1336 4772 1344
rect 4828 1336 4836 1344
rect 4940 1336 4948 1344
rect 108 1316 116 1324
rect 300 1316 308 1324
rect 316 1296 324 1304
rect 396 1296 404 1304
rect 444 1316 452 1324
rect 492 1316 500 1324
rect 540 1316 548 1324
rect 556 1316 564 1324
rect 588 1316 596 1324
rect 620 1296 628 1304
rect 652 1316 660 1324
rect 668 1316 676 1324
rect 748 1318 756 1326
rect 940 1316 948 1324
rect 988 1316 996 1324
rect 1068 1318 1076 1326
rect 1356 1316 1364 1324
rect 1420 1316 1428 1324
rect 1452 1316 1460 1324
rect 1580 1316 1588 1324
rect 1836 1316 1844 1324
rect 1932 1316 1940 1324
rect 2076 1316 2084 1324
rect 2188 1316 2196 1324
rect 2444 1316 2452 1324
rect 2524 1316 2532 1324
rect 2540 1316 2548 1324
rect 2620 1316 2628 1324
rect 2764 1316 2772 1324
rect 2876 1316 2884 1324
rect 3068 1316 3076 1324
rect 3228 1316 3236 1324
rect 3452 1316 3460 1324
rect 3564 1316 3572 1324
rect 3660 1316 3668 1324
rect 3692 1316 3700 1324
rect 3820 1316 3828 1324
rect 4316 1316 4324 1324
rect 4332 1316 4340 1324
rect 4444 1316 4452 1324
rect 4508 1316 4516 1324
rect 4748 1316 4756 1324
rect 4780 1316 4788 1324
rect 4828 1316 4836 1324
rect 4876 1316 4884 1324
rect 5116 1336 5124 1344
rect 5292 1336 5300 1344
rect 5372 1336 5380 1344
rect 5516 1336 5524 1344
rect 5628 1336 5636 1344
rect 4972 1316 4980 1324
rect 5020 1316 5028 1324
rect 5036 1316 5044 1324
rect 5100 1316 5108 1324
rect 5132 1316 5140 1324
rect 5148 1316 5156 1324
rect 5292 1316 5300 1324
rect 5388 1316 5396 1324
rect 5404 1316 5412 1324
rect 5468 1316 5476 1324
rect 5532 1316 5540 1324
rect 5644 1316 5652 1324
rect 5676 1316 5684 1324
rect 5692 1316 5700 1324
rect 5708 1316 5716 1324
rect 5756 1316 5764 1324
rect 5788 1336 5796 1344
rect 5884 1336 5892 1344
rect 5916 1336 5924 1344
rect 5852 1316 5860 1324
rect 5948 1318 5956 1326
rect 956 1296 964 1304
rect 1244 1296 1252 1304
rect 1324 1296 1332 1304
rect 1388 1296 1396 1304
rect 1452 1296 1460 1304
rect 1468 1296 1476 1304
rect 1612 1296 1620 1304
rect 1900 1300 1908 1308
rect 1980 1296 1988 1304
rect 2092 1296 2100 1304
rect 2396 1296 2404 1304
rect 2940 1300 2948 1308
rect 3244 1296 3252 1304
rect 3772 1296 3780 1304
rect 3852 1300 3860 1308
rect 4284 1296 4292 1304
rect 4444 1296 4452 1304
rect 4812 1296 4820 1304
rect 4892 1296 4900 1304
rect 4924 1296 4932 1304
rect 5164 1296 5172 1304
rect 5676 1296 5684 1304
rect 5836 1296 5844 1304
rect 1308 1276 1316 1284
rect 1532 1276 1540 1284
rect 2652 1276 2660 1284
rect 3740 1276 3748 1284
rect 4108 1276 4116 1284
rect 4428 1276 4436 1284
rect 5852 1276 5860 1284
rect 1900 1254 1908 1262
rect 2940 1254 2948 1262
rect 28 1236 36 1244
rect 316 1236 324 1244
rect 508 1236 516 1244
rect 876 1236 884 1244
rect 1196 1236 1204 1244
rect 1420 1236 1428 1244
rect 1644 1236 1652 1244
rect 2396 1236 2404 1244
rect 2508 1236 2516 1244
rect 2572 1236 2580 1244
rect 3244 1236 3252 1244
rect 3532 1236 3540 1244
rect 3852 1236 3860 1244
rect 4156 1236 4164 1244
rect 4316 1236 4324 1244
rect 4444 1236 4452 1244
rect 5500 1236 5508 1244
rect 1502 1206 1510 1214
rect 1516 1206 1524 1214
rect 1530 1206 1538 1214
rect 4574 1206 4582 1214
rect 4588 1206 4596 1214
rect 4602 1206 4610 1214
rect 348 1176 356 1184
rect 428 1176 436 1184
rect 940 1176 948 1184
rect 1036 1176 1044 1184
rect 1340 1176 1348 1184
rect 1564 1176 1572 1184
rect 1708 1176 1716 1184
rect 3148 1176 3156 1184
rect 3740 1176 3748 1184
rect 4060 1176 4068 1184
rect 4268 1176 4276 1184
rect 4812 1176 4820 1184
rect 5052 1176 5060 1184
rect 2188 1156 2196 1164
rect 2684 1158 2692 1166
rect 3404 1158 3412 1166
rect 5964 1158 5972 1166
rect 188 1136 196 1144
rect 860 1136 868 1144
rect 924 1136 932 1144
rect 2204 1136 2212 1144
rect 2236 1136 2244 1144
rect 2764 1136 2772 1144
rect 4716 1136 4724 1144
rect 5036 1136 5044 1144
rect 5372 1136 5380 1144
rect 204 1116 212 1124
rect 268 1116 276 1124
rect 540 1116 548 1124
rect 92 1096 100 1104
rect 220 1096 228 1104
rect 236 1096 244 1104
rect 300 1096 308 1104
rect 380 1096 388 1104
rect 396 1096 404 1104
rect 460 1096 468 1104
rect 476 1096 484 1104
rect 508 1096 516 1104
rect 732 1116 740 1124
rect 876 1116 884 1124
rect 892 1116 900 1124
rect 956 1116 964 1124
rect 988 1116 996 1124
rect 1068 1116 1076 1124
rect 1132 1116 1140 1124
rect 1196 1116 1204 1124
rect 1276 1116 1284 1124
rect 1356 1116 1364 1124
rect 1420 1116 1428 1124
rect 1532 1116 1540 1124
rect 2172 1116 2180 1124
rect 2380 1116 2388 1124
rect 2508 1112 2516 1120
rect 2796 1116 2804 1124
rect 3404 1112 3412 1120
rect 3692 1116 3700 1124
rect 3740 1116 3748 1124
rect 4284 1116 4292 1124
rect 4444 1116 4452 1124
rect 4508 1116 4516 1124
rect 4764 1116 4772 1124
rect 4828 1116 4836 1124
rect 4892 1116 4900 1124
rect 5100 1116 5108 1124
rect 5132 1116 5140 1124
rect 572 1096 580 1104
rect 60 1076 68 1084
rect 252 1076 260 1084
rect 268 1076 276 1084
rect 348 1076 356 1084
rect 492 1076 500 1084
rect 604 1076 612 1084
rect 636 1096 644 1104
rect 684 1096 692 1104
rect 700 1096 708 1104
rect 780 1096 788 1104
rect 828 1096 836 1104
rect 908 1096 916 1104
rect 988 1096 996 1104
rect 1004 1096 1012 1104
rect 1100 1096 1108 1104
rect 1180 1096 1188 1104
rect 1212 1096 1220 1104
rect 1404 1096 1412 1104
rect 1420 1096 1428 1104
rect 1452 1096 1460 1104
rect 1580 1096 1588 1104
rect 1740 1096 1748 1104
rect 1756 1096 1764 1104
rect 1804 1096 1812 1104
rect 1836 1096 1844 1104
rect 1852 1096 1860 1104
rect 1980 1096 1988 1104
rect 2156 1096 2164 1104
rect 2188 1096 2196 1104
rect 2332 1096 2340 1104
rect 2364 1096 2372 1104
rect 2412 1096 2420 1104
rect 2684 1096 2692 1104
rect 2828 1096 2836 1104
rect 2908 1096 2916 1104
rect 3228 1096 3236 1104
rect 3436 1096 3444 1104
rect 3548 1096 3556 1104
rect 3948 1096 3956 1104
rect 4188 1094 4196 1102
rect 844 1076 852 1084
rect 1004 1076 1012 1084
rect 1020 1076 1028 1084
rect 1084 1076 1092 1084
rect 1148 1076 1156 1084
rect 1324 1076 1332 1084
rect 1372 1076 1380 1084
rect 1404 1076 1412 1084
rect 1468 1076 1476 1084
rect 1580 1076 1588 1084
rect 1596 1076 1604 1084
rect 1916 1076 1924 1084
rect 2028 1076 2036 1084
rect 2076 1076 2084 1084
rect 1244 1056 1252 1064
rect 1868 1056 1876 1064
rect 2108 1076 2116 1084
rect 2140 1076 2148 1084
rect 2252 1076 2260 1084
rect 2428 1076 2436 1084
rect 2572 1076 2580 1084
rect 2812 1076 2820 1084
rect 2844 1076 2852 1084
rect 2924 1076 2932 1084
rect 3020 1076 3028 1084
rect 3084 1076 3092 1084
rect 3340 1076 3348 1084
rect 3500 1076 3508 1084
rect 3644 1076 3652 1084
rect 3692 1076 3700 1084
rect 3836 1076 3844 1084
rect 4076 1076 4084 1084
rect 4156 1076 4164 1084
rect 4284 1076 4292 1084
rect 4332 1076 4340 1084
rect 4364 1096 4372 1104
rect 4412 1096 4420 1104
rect 4444 1096 4452 1104
rect 4508 1096 4516 1104
rect 4540 1096 4548 1104
rect 4684 1096 4692 1104
rect 4812 1096 4820 1104
rect 4860 1096 4868 1104
rect 4892 1096 4900 1104
rect 4924 1096 4932 1104
rect 5068 1096 5076 1104
rect 5148 1096 5156 1104
rect 5180 1096 5188 1104
rect 5212 1096 5220 1104
rect 5228 1096 5236 1104
rect 5260 1096 5268 1104
rect 5308 1116 5316 1124
rect 5676 1116 5684 1124
rect 5964 1112 5972 1120
rect 6044 1116 6052 1124
rect 5340 1096 5348 1104
rect 5484 1096 5492 1104
rect 5564 1096 5572 1104
rect 5644 1096 5652 1104
rect 5692 1096 5700 1104
rect 5788 1096 5796 1104
rect 5980 1096 5988 1104
rect 6076 1096 6084 1104
rect 4556 1076 4564 1084
rect 4620 1076 4628 1084
rect 4716 1076 4724 1084
rect 4876 1076 4884 1084
rect 4924 1076 4932 1084
rect 4940 1076 4948 1084
rect 5004 1076 5012 1084
rect 5084 1076 5092 1084
rect 5244 1076 5252 1084
rect 5292 1076 5300 1084
rect 5356 1076 5364 1084
rect 5532 1076 5540 1084
rect 5628 1076 5636 1084
rect 5900 1076 5908 1084
rect 6044 1076 6052 1084
rect 6092 1076 6100 1084
rect 2108 1056 2116 1064
rect 2252 1056 2260 1064
rect 2268 1056 2276 1064
rect 2332 1056 2340 1064
rect 2364 1056 2372 1064
rect 2604 1056 2612 1064
rect 3308 1056 3316 1064
rect 3628 1056 3636 1064
rect 3868 1056 3876 1064
rect 4252 1056 4260 1064
rect 4444 1056 4452 1064
rect 4684 1056 4692 1064
rect 4716 1056 4724 1064
rect 4780 1056 4788 1064
rect 5068 1056 5076 1064
rect 5868 1056 5876 1064
rect 796 1036 804 1044
rect 1292 1036 1300 1044
rect 1788 1036 1796 1044
rect 2044 1036 2052 1044
rect 2124 1036 2132 1044
rect 2380 1036 2388 1044
rect 2972 1036 2980 1044
rect 3100 1036 3108 1044
rect 3580 1036 3588 1044
rect 4028 1036 4036 1044
rect 4636 1036 4644 1044
rect 4748 1036 4756 1044
rect 4828 1036 4836 1044
rect 4988 1036 4996 1044
rect 5132 1036 5140 1044
rect 3038 1006 3046 1014
rect 3052 1006 3060 1014
rect 3066 1006 3074 1014
rect 204 976 212 984
rect 428 976 436 984
rect 972 976 980 984
rect 1148 976 1156 984
rect 1212 976 1220 984
rect 1404 976 1412 984
rect 1436 976 1444 984
rect 2092 976 2100 984
rect 2236 976 2244 984
rect 2476 976 2484 984
rect 3324 976 3332 984
rect 4012 976 4020 984
rect 4220 976 4228 984
rect 4284 976 4292 984
rect 4332 976 4340 984
rect 4492 976 4500 984
rect 5164 976 5172 984
rect 5420 976 5428 984
rect 5660 976 5668 984
rect 6076 976 6084 984
rect 684 956 692 964
rect 796 956 804 964
rect 1132 956 1140 964
rect 1932 956 1940 964
rect 2508 956 2516 964
rect 2668 956 2676 964
rect 3004 956 3012 964
rect 3484 956 3492 964
rect 3820 956 3828 964
rect 4076 956 4084 964
rect 4300 956 4308 964
rect 4476 956 4484 964
rect 4764 956 4772 964
rect 5100 956 5108 964
rect 5916 956 5924 964
rect 124 936 132 944
rect 252 936 260 944
rect 268 936 276 944
rect 476 936 484 944
rect 556 936 564 944
rect 732 936 740 944
rect 892 936 900 944
rect 1020 936 1028 944
rect 1196 936 1204 944
rect 1244 936 1252 944
rect 1356 936 1364 944
rect 1452 936 1460 944
rect 1692 936 1700 944
rect 1900 936 1908 944
rect 2172 936 2180 944
rect 2188 936 2196 944
rect 2268 936 2276 944
rect 2316 932 2324 940
rect 2348 936 2356 944
rect 2380 936 2388 944
rect 2396 936 2404 944
rect 2700 936 2708 944
rect 2972 936 2980 944
rect 3166 936 3174 944
rect 3516 936 3524 944
rect 3788 936 3796 944
rect 4076 936 4084 944
rect 4140 936 4148 944
rect 4380 936 4388 944
rect 4556 936 4564 944
rect 4588 936 4596 944
rect 4732 936 4740 944
rect 4908 936 4916 944
rect 5116 936 5124 944
rect 140 918 148 926
rect 236 916 244 924
rect 284 916 292 924
rect 348 916 356 924
rect 364 916 372 924
rect 396 916 404 924
rect 412 916 420 924
rect 460 916 468 924
rect 588 916 596 924
rect 716 916 724 924
rect 748 916 756 924
rect 764 916 772 924
rect 876 916 884 924
rect 924 916 932 924
rect 1004 916 1012 924
rect 1052 916 1060 924
rect 1100 916 1108 924
rect 1180 916 1188 924
rect 1260 916 1268 924
rect 1324 916 1332 924
rect 1356 916 1364 924
rect 1372 916 1380 924
rect 1500 916 1508 924
rect 1708 918 1716 926
rect 1820 916 1828 924
rect 2012 916 2020 924
rect 2156 916 2164 924
rect 204 896 212 904
rect 284 896 292 904
rect 316 896 324 904
rect 428 896 436 904
rect 684 896 692 904
rect 844 896 852 904
rect 908 896 916 904
rect 1036 896 1044 904
rect 1116 896 1124 904
rect 1148 896 1156 904
rect 1212 896 1220 904
rect 1404 896 1412 904
rect 1420 896 1428 904
rect 1836 900 1844 908
rect 2124 896 2132 904
rect 2156 896 2164 904
rect 2220 896 2228 904
rect 2268 916 2276 924
rect 2396 916 2404 924
rect 2412 916 2420 924
rect 2796 916 2804 924
rect 2860 916 2868 924
rect 2876 916 2884 924
rect 3404 916 3412 924
rect 3692 916 3700 924
rect 4044 916 4052 924
rect 4124 916 4132 924
rect 4188 916 4196 924
rect 4236 916 4244 924
rect 4252 916 4260 924
rect 4268 916 4276 924
rect 4364 916 4372 924
rect 4396 916 4404 924
rect 4444 916 4452 924
rect 4492 916 4500 924
rect 4524 916 4532 924
rect 4652 916 4660 924
rect 4668 916 4676 924
rect 4716 916 4724 924
rect 4844 916 4852 924
rect 4908 916 4916 924
rect 4972 916 4980 924
rect 4988 916 4996 924
rect 5036 916 5044 924
rect 5068 916 5076 924
rect 5180 916 5188 924
rect 5196 916 5204 924
rect 5244 916 5252 924
rect 5276 936 5284 944
rect 5324 936 5332 944
rect 5388 936 5396 944
rect 5404 936 5412 944
rect 5612 936 5620 944
rect 5644 936 5652 944
rect 5692 936 5700 944
rect 5884 936 5892 944
rect 2348 896 2356 904
rect 2444 896 2452 904
rect 2764 900 2772 908
rect 2876 896 2884 904
rect 3580 900 3588 908
rect 3724 900 3732 908
rect 4012 896 4020 904
rect 4156 896 4164 904
rect 4428 896 4436 904
rect 4492 896 4500 904
rect 4556 896 4564 904
rect 4572 896 4580 904
rect 4956 896 4964 904
rect 5372 916 5380 924
rect 5564 916 5572 924
rect 5708 916 5716 924
rect 5788 916 5796 924
rect 5884 916 5892 924
rect 5340 896 5348 904
rect 5676 896 5684 904
rect 5740 896 5748 904
rect 5820 900 5828 908
rect 12 876 20 884
rect 668 876 676 884
rect 940 876 948 884
rect 1068 876 1076 884
rect 1084 876 1092 884
rect 1468 876 1476 884
rect 1484 876 1492 884
rect 5164 876 5172 884
rect 5436 876 5444 884
rect 5452 876 5460 884
rect 1836 854 1844 862
rect 3404 854 3412 862
rect 3724 854 3732 862
rect 5820 854 5828 862
rect 236 836 244 844
rect 876 836 884 844
rect 1308 836 1316 844
rect 1580 836 1588 844
rect 2764 836 2772 844
rect 2876 836 2884 844
rect 3260 836 3268 844
rect 3980 836 3988 844
rect 4396 836 4404 844
rect 4700 836 4708 844
rect 4796 836 4804 844
rect 4876 836 4884 844
rect 4924 836 4932 844
rect 5020 836 5028 844
rect 5708 836 5716 844
rect 1502 806 1510 814
rect 1516 806 1524 814
rect 1530 806 1538 814
rect 4574 806 4582 814
rect 4588 806 4596 814
rect 4602 806 4610 814
rect 652 776 660 784
rect 1004 776 1012 784
rect 1036 776 1044 784
rect 1068 776 1076 784
rect 1276 776 1284 784
rect 1324 776 1332 784
rect 1756 776 1764 784
rect 1868 776 1876 784
rect 2076 776 2084 784
rect 3324 776 3332 784
rect 3980 776 3988 784
rect 4284 776 4292 784
rect 4412 776 4420 784
rect 5996 776 6004 784
rect 2844 758 2852 766
rect 4556 756 4564 764
rect 5148 756 5156 764
rect 204 736 212 744
rect 620 736 628 744
rect 796 736 804 744
rect 2524 736 2532 744
rect 2588 736 2596 744
rect 3036 736 3044 744
rect 3548 736 3556 744
rect 3900 736 3908 744
rect 4108 736 4116 744
rect 4252 736 4260 744
rect 4636 736 4644 744
rect 5356 736 5364 744
rect 5580 736 5588 744
rect 5756 736 5764 744
rect 5964 736 5972 744
rect 60 696 68 704
rect 108 716 116 724
rect 172 716 180 724
rect 140 696 148 704
rect 236 696 244 704
rect 252 696 260 704
rect 284 696 292 704
rect 300 696 308 704
rect 332 696 340 704
rect 380 716 388 724
rect 684 716 692 724
rect 748 716 756 724
rect 412 696 420 704
rect 492 694 500 702
rect 556 696 564 704
rect 652 696 660 704
rect 716 696 724 704
rect 1452 716 1460 724
rect 796 696 804 704
rect 828 696 836 704
rect 844 696 852 704
rect 924 696 932 704
rect 988 696 996 704
rect 1196 696 1204 704
rect 1340 696 1348 704
rect 1820 716 1828 724
rect 156 676 164 684
rect 220 676 228 684
rect 316 676 324 684
rect 364 676 372 684
rect 428 676 436 684
rect 636 676 644 684
rect 700 676 708 684
rect 812 676 820 684
rect 908 676 916 684
rect 1180 676 1188 684
rect 1500 696 1508 704
rect 1628 694 1636 702
rect 1788 696 1796 704
rect 1996 716 2004 724
rect 2076 716 2084 724
rect 2556 716 2564 724
rect 2844 712 2852 720
rect 3324 716 3332 724
rect 3420 716 3428 724
rect 3644 716 3652 724
rect 3740 716 3748 724
rect 3820 716 3828 724
rect 3868 716 3876 724
rect 3932 716 3940 724
rect 4140 716 4148 724
rect 4172 716 4180 724
rect 4204 716 4212 724
rect 4220 716 4228 724
rect 4268 716 4276 724
rect 4300 716 4308 724
rect 4444 716 4452 724
rect 4460 716 4468 724
rect 4524 716 4532 724
rect 1868 696 1876 704
rect 1900 696 1908 704
rect 1916 696 1924 704
rect 1964 696 1972 704
rect 2076 696 2084 704
rect 2380 696 2388 704
rect 2476 696 2484 704
rect 2860 696 2868 704
rect 3116 696 3124 704
rect 3228 696 3236 704
rect 3388 696 3396 704
rect 3580 696 3588 704
rect 3756 696 3764 704
rect 3788 696 3796 704
rect 3900 696 3908 704
rect 1404 676 1412 684
rect 1468 676 1476 684
rect 1564 676 1572 684
rect 1772 676 1780 684
rect 1884 676 1892 684
rect 2012 676 2020 684
rect 2028 676 2036 684
rect 2172 676 2180 684
rect 2460 676 2468 684
rect 2572 676 2580 684
rect 2780 676 2788 684
rect 2924 676 2932 684
rect 3228 676 3236 684
rect 3372 676 3380 684
rect 3532 676 3540 684
rect 3564 676 3572 684
rect 3596 676 3604 684
rect 3612 676 3620 684
rect 3676 676 3684 684
rect 3772 676 3780 684
rect 3884 676 3892 684
rect 3948 676 3956 684
rect 4108 696 4116 704
rect 4172 696 4180 704
rect 4284 696 4292 704
rect 4380 696 4388 704
rect 4412 696 4420 704
rect 4444 696 4452 704
rect 4492 696 4500 704
rect 4572 696 4580 704
rect 4748 696 4756 704
rect 4844 696 4852 704
rect 4892 716 4900 724
rect 5004 716 5012 724
rect 4924 696 4932 704
rect 5052 716 5060 724
rect 5132 716 5140 724
rect 5436 716 5444 724
rect 5612 716 5620 724
rect 5724 716 5732 724
rect 6012 716 6020 724
rect 6028 716 6036 724
rect 5052 696 5060 704
rect 5084 696 5092 704
rect 5260 696 5268 704
rect 5356 696 5364 704
rect 5484 696 5492 704
rect 5548 696 5556 704
rect 5612 696 5620 704
rect 5644 696 5652 704
rect 5692 696 5700 704
rect 5756 696 5764 704
rect 5836 694 5844 702
rect 6060 696 6068 704
rect 4060 676 4068 684
rect 4076 676 4084 684
rect 4092 676 4100 684
rect 4156 676 4164 684
rect 4252 676 4260 684
rect 4396 676 4404 684
rect 4508 676 4516 684
rect 4588 676 4596 684
rect 4732 676 4740 684
rect 4828 676 4836 684
rect 4940 676 4948 684
rect 5068 676 5076 684
rect 5084 676 5092 684
rect 5260 676 5268 684
rect 5340 676 5348 684
rect 5404 676 5412 684
rect 5484 676 5492 684
rect 5564 676 5572 684
rect 5708 676 5716 684
rect 5772 676 5780 684
rect 5804 676 5812 684
rect 5980 676 5988 684
rect 6076 676 6084 684
rect 12 656 20 664
rect 492 656 500 664
rect 860 656 868 664
rect 988 656 996 664
rect 1020 656 1028 664
rect 1052 656 1060 664
rect 1292 656 1300 664
rect 1308 656 1316 664
rect 1628 656 1636 664
rect 1932 656 1940 664
rect 2204 656 2212 664
rect 2748 656 2756 664
rect 3196 656 3204 664
rect 3628 656 3636 664
rect 3660 656 3668 664
rect 3724 656 3732 664
rect 5452 656 5460 664
rect 92 636 100 644
rect 1084 636 1092 644
rect 1372 636 1380 644
rect 2364 636 2372 644
rect 2940 636 2948 644
rect 3468 636 3476 644
rect 3708 636 3716 644
rect 3852 636 3860 644
rect 4236 636 4244 644
rect 4348 636 4356 644
rect 4876 636 4884 644
rect 5132 636 5140 644
rect 5532 636 5540 644
rect 6028 636 6036 644
rect 3038 606 3046 614
rect 3052 606 3060 614
rect 3066 606 3074 614
rect 332 576 340 584
rect 444 576 452 584
rect 492 576 500 584
rect 732 576 740 584
rect 972 576 980 584
rect 1004 576 1012 584
rect 2124 576 2132 584
rect 3532 576 3540 584
rect 3676 576 3684 584
rect 3708 576 3716 584
rect 4044 576 4052 584
rect 4252 576 4260 584
rect 4348 576 4356 584
rect 4588 576 4596 584
rect 5004 576 5012 584
rect 5036 576 5044 584
rect 5436 576 5444 584
rect 5788 576 5796 584
rect 172 556 180 564
rect 956 556 964 564
rect 1436 556 1444 564
rect 1964 556 1972 564
rect 2204 556 2212 564
rect 2220 556 2228 564
rect 2412 556 2420 564
rect 2588 556 2596 564
rect 2748 556 2756 564
rect 3116 556 3124 564
rect 3548 556 3556 564
rect 3612 556 3620 564
rect 3692 556 3700 564
rect 3884 556 3892 564
rect 4268 556 4276 564
rect 4428 556 4436 564
rect 4524 556 4532 564
rect 4716 556 4724 564
rect 5020 556 5028 564
rect 5948 556 5956 564
rect 140 536 148 544
rect 364 536 372 544
rect 460 536 468 544
rect 604 536 612 544
rect 748 536 756 544
rect 1116 536 1124 544
rect 1532 536 1540 544
rect 1644 536 1652 544
rect 1660 536 1668 544
rect 1788 536 1796 544
rect 1932 536 1940 544
rect 2156 536 2164 544
rect 2236 536 2244 544
rect 2284 536 2292 544
rect 2380 536 2388 544
rect 2556 536 2564 544
rect 2780 536 2788 544
rect 2892 536 2900 544
rect 3084 536 3092 544
rect 3404 536 3412 544
rect 3484 536 3492 544
rect 3516 536 3524 544
rect 3548 536 3556 544
rect 3628 536 3636 544
rect 3852 536 3860 544
rect 4092 536 4100 544
rect 4412 536 4420 544
rect 4476 536 4484 544
rect 4844 536 4852 544
rect 5164 536 5172 544
rect 5308 536 5316 544
rect 5420 536 5428 544
rect 5596 536 5604 544
rect 5756 536 5764 544
rect 5980 536 5988 544
rect 76 516 84 524
rect 348 516 356 524
rect 636 516 644 524
rect 684 516 692 524
rect 716 516 724 524
rect 764 516 772 524
rect 780 516 788 524
rect 860 516 868 524
rect 876 516 884 524
rect 924 516 932 524
rect 940 516 948 524
rect 1132 516 1140 524
rect 1196 516 1204 524
rect 1212 516 1220 524
rect 1244 516 1252 524
rect 1292 516 1300 524
rect 1388 516 1396 524
rect 1404 516 1412 524
rect 1452 516 1460 524
rect 1468 516 1476 524
rect 1548 516 1556 524
rect 1564 516 1572 524
rect 44 496 52 504
rect 412 496 420 504
rect 716 496 724 504
rect 1628 516 1636 524
rect 1852 516 1860 524
rect 2044 516 2052 524
rect 1596 496 1604 504
rect 1836 496 1844 504
rect 2188 496 2196 504
rect 2268 496 2276 504
rect 2316 496 2324 504
rect 2460 516 2468 524
rect 2796 516 2804 524
rect 2892 516 2900 524
rect 2972 516 2980 524
rect 3196 516 3204 524
rect 3308 516 3316 524
rect 3372 516 3380 524
rect 3388 516 3396 524
rect 2364 496 2372 504
rect 2460 496 2468 504
rect 2828 496 2836 504
rect 2844 496 2852 504
rect 3020 500 3028 508
rect 3276 496 3284 504
rect 3436 496 3444 504
rect 3580 516 3588 524
rect 3644 516 3652 524
rect 3756 516 3764 524
rect 3852 516 3860 524
rect 4140 516 4148 524
rect 4188 516 4196 524
rect 4316 516 4324 524
rect 4396 516 4404 524
rect 4460 516 4468 524
rect 4476 516 4484 524
rect 4556 516 4564 524
rect 4636 516 4644 524
rect 4668 516 4676 524
rect 4732 516 4740 524
rect 4748 516 4756 524
rect 4796 516 4804 524
rect 4876 518 4884 526
rect 5052 516 5060 524
rect 5068 516 5076 524
rect 5116 516 5124 524
rect 5148 516 5156 524
rect 5212 516 5220 524
rect 5228 516 5236 524
rect 5276 516 5284 524
rect 5292 516 5300 524
rect 5324 516 5332 524
rect 3612 496 3620 504
rect 3788 500 3796 508
rect 4348 496 4356 504
rect 4364 496 4372 504
rect 4396 496 4404 504
rect 4428 496 4436 504
rect 4636 496 4644 504
rect 5244 496 5252 504
rect 5356 496 5364 504
rect 5404 516 5412 524
rect 5500 516 5508 524
rect 5516 516 5524 524
rect 5868 516 5876 524
rect 5980 516 5988 524
rect 6044 500 6052 508
rect 428 476 436 484
rect 2236 476 2244 484
rect 5404 476 5412 484
rect 3020 454 3028 462
rect 6044 454 6052 462
rect 44 436 52 444
rect 380 436 388 444
rect 652 436 660 444
rect 796 436 804 444
rect 908 436 916 444
rect 1004 436 1012 444
rect 1180 436 1188 444
rect 1260 436 1268 444
rect 1340 436 1348 444
rect 1836 436 1844 444
rect 2172 436 2180 444
rect 2460 436 2468 444
rect 2748 436 2756 444
rect 2796 436 2804 444
rect 2876 436 2884 444
rect 3340 436 3348 444
rect 3788 436 3796 444
rect 4780 436 4788 444
rect 5100 436 5108 444
rect 5644 436 5652 444
rect 1502 406 1510 414
rect 1516 406 1524 414
rect 1530 406 1538 414
rect 4574 406 4582 414
rect 4588 406 4596 414
rect 4602 406 4610 414
rect 92 376 100 384
rect 380 376 388 384
rect 1132 376 1140 384
rect 1404 376 1412 384
rect 2700 376 2708 384
rect 3132 376 3140 384
rect 3308 376 3316 384
rect 3388 376 3396 384
rect 3516 376 3524 384
rect 3564 376 3572 384
rect 3884 376 3892 384
rect 4188 376 4196 384
rect 4316 376 4324 384
rect 4444 376 4452 384
rect 4764 376 4772 384
rect 5084 376 5092 384
rect 5372 376 5380 384
rect 6044 376 6052 384
rect 636 356 644 364
rect 2060 358 2068 366
rect 2396 358 2404 366
rect 2780 358 2788 366
rect 5708 356 5716 364
rect 5964 358 5972 366
rect 3500 336 3508 344
rect 4300 336 4308 344
rect 4428 336 4436 344
rect 5436 336 5444 344
rect 6124 336 6132 344
rect 92 316 100 324
rect 412 316 420 324
rect 556 316 564 324
rect 44 296 52 304
rect 92 296 100 304
rect 300 296 308 304
rect 444 296 452 304
rect 524 296 532 304
rect 844 316 852 324
rect 604 296 612 304
rect 764 294 772 302
rect 844 296 852 304
rect 892 316 900 324
rect 1164 316 1172 324
rect 924 296 932 304
rect 1020 296 1028 304
rect 1164 296 1172 304
rect 1212 316 1220 324
rect 1244 296 1252 304
rect 1260 296 1268 304
rect 1340 316 1348 324
rect 1372 296 1380 304
rect 1468 296 1476 304
rect 1740 316 1748 324
rect 2060 312 2068 320
rect 2172 316 2180 324
rect 2236 316 2244 324
rect 2396 312 2404 320
rect 2780 312 2788 320
rect 3468 316 3476 324
rect 3884 316 3892 324
rect 4268 316 4276 324
rect 4348 316 4356 324
rect 4476 316 4484 324
rect 1532 294 1540 302
rect 1802 296 1810 304
rect 1884 296 1892 304
rect 2172 296 2180 304
rect 2204 296 2212 304
rect 2572 296 2580 304
rect 2956 296 2964 304
rect 3148 296 3156 304
rect 12 276 20 284
rect 188 276 196 284
rect 396 276 404 284
rect 508 276 516 284
rect 620 276 628 284
rect 828 276 836 284
rect 940 276 948 284
rect 1004 276 1012 284
rect 1148 276 1156 284
rect 1260 276 1268 284
rect 1276 276 1284 284
rect 1388 276 1396 284
rect 1612 276 1620 284
rect 1676 276 1684 284
rect 1996 276 2004 284
rect 2220 276 2228 284
rect 2284 276 2292 284
rect 2460 276 2468 284
rect 2844 276 2852 284
rect 3038 276 3046 284
rect 3148 276 3156 284
rect 3260 296 3268 304
rect 3276 296 3284 304
rect 3484 296 3492 304
rect 3564 296 3572 304
rect 3676 296 3684 304
rect 3852 296 3860 304
rect 4236 296 4244 304
rect 4316 296 4324 304
rect 4364 296 4372 304
rect 4380 296 4388 304
rect 4444 296 4452 304
rect 4508 296 4516 304
rect 4652 296 4660 304
rect 4700 296 4708 304
rect 4780 296 4788 304
rect 4812 296 4820 304
rect 4844 316 4852 324
rect 4892 296 4900 304
rect 4972 296 4980 304
rect 5020 296 5028 304
rect 5100 296 5108 304
rect 5132 296 5140 304
rect 5164 316 5172 324
rect 5388 316 5396 324
rect 5516 316 5524 324
rect 5532 316 5540 324
rect 5596 316 5604 324
rect 5964 312 5972 320
rect 5196 296 5204 304
rect 5484 296 5492 304
rect 5564 296 5572 304
rect 5628 296 5636 304
rect 5980 296 5988 304
rect 6012 296 6020 304
rect 6060 296 6068 304
rect 3356 276 3364 284
rect 3452 276 3460 284
rect 3788 276 3796 284
rect 4076 276 4084 284
rect 4220 276 4228 284
rect 4252 276 4260 284
rect 4396 276 4404 284
rect 4492 276 4500 284
rect 4524 276 4532 284
rect 4780 276 4788 284
rect 4892 276 4900 284
rect 5100 276 5108 284
rect 5212 276 5220 284
rect 5228 276 5236 284
rect 5356 276 5364 284
rect 5452 276 5460 284
rect 5516 276 5524 284
rect 5580 276 5588 284
rect 5612 276 5620 284
rect 5900 276 5908 284
rect 220 256 228 264
rect 492 256 500 264
rect 764 256 772 264
rect 1628 256 1636 264
rect 1964 256 1972 264
rect 2156 256 2164 264
rect 2316 256 2324 264
rect 2492 256 2500 264
rect 2876 256 2884 264
rect 3100 256 3108 264
rect 3532 256 3540 264
rect 3596 256 3604 264
rect 3756 256 3764 264
rect 5388 256 5396 264
rect 5676 256 5684 264
rect 5868 256 5876 264
rect 6060 256 6068 264
rect 572 236 580 244
rect 1324 236 1332 244
rect 1724 236 1732 244
rect 2172 236 2180 244
rect 2236 236 2244 244
rect 2652 236 2660 244
rect 3948 236 3956 244
rect 5532 236 5540 244
rect 3038 206 3046 214
rect 3052 206 3060 214
rect 3066 206 3074 214
rect 700 176 708 184
rect 732 176 740 184
rect 908 176 916 184
rect 1100 176 1108 184
rect 1308 176 1316 184
rect 1468 176 1476 184
rect 2524 176 2532 184
rect 3468 176 3476 184
rect 3964 176 3972 184
rect 4268 176 4276 184
rect 4332 176 4340 184
rect 5388 176 5396 184
rect 5436 176 5444 184
rect 5628 176 5636 184
rect 5708 176 5716 184
rect 5740 176 5748 184
rect 6076 176 6084 184
rect 172 156 180 164
rect 332 156 340 164
rect 508 156 516 164
rect 1628 156 1636 164
rect 1964 156 1972 164
rect 2364 156 2372 164
rect 2860 156 2868 164
rect 3308 156 3316 164
rect 3564 156 3572 164
rect 3596 156 3604 164
rect 3628 156 3636 164
rect 3804 156 3812 164
rect 4092 156 4100 164
rect 4460 156 4468 164
rect 4668 156 4676 164
rect 4780 156 4788 164
rect 5644 156 5652 164
rect 5900 156 5908 164
rect 6108 156 6116 164
rect 140 136 148 144
rect 364 136 372 144
rect 428 136 436 144
rect 540 136 548 144
rect 780 136 788 144
rect 828 136 836 144
rect 892 136 900 144
rect 1004 136 1012 144
rect 1292 136 1300 144
rect 1660 136 1668 144
rect 1932 136 1940 144
rect 2332 136 2340 144
rect 2828 136 2836 144
rect 3276 136 3284 144
rect 3484 136 3492 144
rect 3596 136 3604 144
rect 3772 136 3780 144
rect 4524 136 4532 144
rect 4572 136 4580 144
rect 4828 136 4836 144
rect 4876 136 4884 144
rect 4940 136 4948 144
rect 5020 136 5028 144
rect 5244 136 5252 144
rect 5292 136 5300 144
rect 5596 136 5604 144
rect 5660 136 5668 144
rect 5932 136 5940 144
rect 76 116 84 124
rect 380 116 388 124
rect 44 96 52 104
rect 412 96 420 104
rect 460 116 468 124
rect 572 118 580 126
rect 780 116 788 124
rect 796 116 804 124
rect 876 116 884 124
rect 1020 116 1028 124
rect 1164 116 1172 124
rect 1228 118 1236 126
rect 1340 116 1348 124
rect 1548 116 1556 124
rect 1772 116 1780 124
rect 1836 116 1844 124
rect 2044 116 2052 124
rect 2156 116 2164 124
rect 2236 116 2244 124
rect 2604 116 2612 124
rect 2652 116 2660 124
rect 2732 116 2740 124
rect 3100 116 3108 124
rect 3180 116 3188 124
rect 3676 116 3684 124
rect 3996 116 4004 124
rect 4108 116 4116 124
rect 4236 116 4244 124
rect 4252 116 4260 124
rect 4300 116 4308 124
rect 4460 118 4468 126
rect 4556 116 4564 124
rect 4636 116 4644 124
rect 4652 116 4660 124
rect 4732 116 4740 124
rect 4748 116 4756 124
rect 4796 116 4804 124
rect 4812 116 4820 124
rect 4844 116 4852 124
rect 844 96 852 104
rect 1756 96 1764 104
rect 1868 100 1876 108
rect 2236 96 2244 104
rect 2764 100 2772 108
rect 3212 100 3220 108
rect 3676 96 3684 104
rect 4524 96 4532 104
rect 4924 116 4932 124
rect 5004 118 5012 126
rect 5148 116 5156 124
rect 5212 116 5220 124
rect 5228 116 5236 124
rect 5260 116 5268 124
rect 4892 96 4900 104
rect 5180 96 5188 104
rect 5340 116 5348 124
rect 5420 116 5428 124
rect 5548 116 5556 124
rect 5676 116 5684 124
rect 6012 116 6020 124
rect 5308 96 5316 104
rect 5708 96 5716 104
rect 5996 100 6004 108
rect 4220 76 4228 84
rect 5132 76 5140 84
rect 2764 54 2772 62
rect 44 36 52 44
rect 1356 36 1364 44
rect 1756 36 1764 44
rect 1868 36 1876 44
rect 2188 36 2196 44
rect 2236 36 2244 44
rect 2588 36 2596 44
rect 2636 36 2644 44
rect 2684 36 2692 44
rect 3132 36 3140 44
rect 3212 36 3220 44
rect 3676 36 3684 44
rect 4028 36 4036 44
rect 5996 36 6004 44
rect 1502 6 1510 14
rect 1516 6 1524 14
rect 1530 6 1538 14
rect 4574 6 4582 14
rect 4588 6 4596 14
rect 4602 6 4610 14
<< metal2 >>
rect 397 5637 419 5643
rect 461 5637 483 5643
rect 397 5584 403 5637
rect 77 5524 83 5576
rect 461 5523 467 5637
rect 461 5517 483 5523
rect 29 5284 35 5456
rect 61 5324 67 5496
rect 285 5464 291 5496
rect 173 5364 179 5456
rect 333 5384 339 5496
rect 13 4984 19 5036
rect 13 4904 19 4916
rect 13 4324 19 4436
rect 29 4304 35 5276
rect 77 5244 83 5300
rect 61 5044 67 5094
rect 125 5084 131 5096
rect 173 5084 179 5356
rect 333 5304 339 5376
rect 349 5304 355 5356
rect 381 5323 387 5456
rect 381 5317 396 5323
rect 413 5224 419 5336
rect 445 5324 451 5476
rect 461 5364 467 5436
rect 477 5364 483 5517
rect 509 5464 515 5643
rect 1789 5637 1811 5643
rect 1981 5637 2003 5643
rect 2525 5637 2547 5643
rect 2941 5637 2963 5643
rect 1496 5606 1502 5614
rect 1510 5606 1516 5614
rect 1524 5606 1530 5614
rect 1538 5606 1544 5614
rect 1789 5584 1795 5637
rect 1981 5584 1987 5637
rect 2525 5584 2531 5637
rect 2957 5584 2963 5637
rect 637 5524 643 5536
rect 957 5524 963 5576
rect 1469 5524 1475 5576
rect 525 5324 531 5496
rect 589 5463 595 5476
rect 573 5457 595 5463
rect 573 5344 579 5457
rect 525 5284 531 5316
rect 573 5224 579 5336
rect 605 5323 611 5496
rect 749 5464 755 5496
rect 957 5464 963 5496
rect 941 5457 956 5463
rect 829 5423 835 5456
rect 813 5417 835 5423
rect 813 5364 819 5417
rect 596 5317 611 5323
rect 61 4864 67 4936
rect 93 4484 99 4916
rect 125 4704 131 5076
rect 189 5024 195 5036
rect 157 4924 163 4996
rect 173 4924 179 4936
rect 141 4904 147 4916
rect 157 4844 163 4916
rect 189 4903 195 5016
rect 253 4944 259 5056
rect 205 4904 211 4916
rect 180 4897 195 4903
rect 125 4404 131 4696
rect 205 4684 211 4856
rect 221 4804 227 4936
rect 269 4724 275 4736
rect 301 4704 307 4896
rect 317 4804 323 5216
rect 813 5144 819 5356
rect 941 5324 947 5457
rect 989 5304 995 5336
rect 941 5244 947 5296
rect 452 5117 460 5123
rect 541 5104 547 5116
rect 381 5044 387 5076
rect 173 4544 179 4556
rect 205 4544 211 4676
rect 221 4644 227 4696
rect 13 4264 19 4296
rect 45 4044 51 4096
rect 45 3924 51 3976
rect 61 3764 67 4296
rect 77 4144 83 4276
rect 93 4244 99 4316
rect 173 4164 179 4536
rect 221 4524 227 4536
rect 221 4384 227 4396
rect 141 3823 147 3876
rect 173 3864 179 4156
rect 253 3904 259 4116
rect 125 3817 147 3823
rect 125 3784 131 3817
rect 13 3744 19 3756
rect 45 3743 51 3756
rect 29 3737 51 3743
rect 29 3704 35 3737
rect 77 3724 83 3736
rect 93 3724 99 3756
rect 93 3604 99 3716
rect 125 3704 131 3756
rect 61 3504 67 3596
rect 93 3524 99 3576
rect 141 3524 147 3576
rect 13 3464 19 3496
rect 93 3424 99 3436
rect 125 3404 131 3496
rect 157 3484 163 3636
rect 205 3624 211 3696
rect 253 3583 259 3896
rect 269 3824 275 4476
rect 285 4384 291 4496
rect 301 4303 307 4696
rect 317 4684 323 4796
rect 333 4524 339 4536
rect 349 4524 355 4956
rect 381 4684 387 4876
rect 397 4864 403 5076
rect 413 5064 419 5096
rect 461 5004 467 5096
rect 477 5084 483 5096
rect 413 4904 419 4976
rect 429 4864 435 4936
rect 445 4924 451 4936
rect 477 4904 483 4916
rect 493 4883 499 4916
rect 525 4884 531 5096
rect 557 5084 563 5116
rect 557 4924 563 4976
rect 605 4923 611 5096
rect 621 4943 627 5076
rect 669 5004 675 5116
rect 797 5102 803 5116
rect 861 5104 867 5136
rect 621 4937 636 4943
rect 653 4924 659 4956
rect 669 4924 675 4996
rect 717 4944 723 5096
rect 733 5044 739 5076
rect 605 4917 620 4923
rect 557 4904 563 4916
rect 477 4877 499 4883
rect 477 4844 483 4877
rect 397 4704 403 4716
rect 381 4584 387 4596
rect 413 4584 419 4676
rect 365 4544 371 4556
rect 333 4324 339 4516
rect 445 4444 451 4516
rect 461 4504 467 4576
rect 477 4544 483 4836
rect 573 4824 579 4916
rect 573 4724 579 4756
rect 573 4684 579 4716
rect 589 4684 595 4716
rect 653 4704 659 4876
rect 717 4844 723 4916
rect 733 4864 739 5036
rect 749 4944 755 5016
rect 797 4944 803 5076
rect 845 4964 851 4996
rect 804 4917 851 4923
rect 845 4904 851 4917
rect 877 4903 883 4936
rect 893 4924 899 5216
rect 877 4897 899 4903
rect 717 4804 723 4836
rect 717 4704 723 4736
rect 733 4704 739 4816
rect 749 4744 755 4896
rect 829 4784 835 4896
rect 861 4824 867 4836
rect 861 4704 867 4796
rect 877 4704 883 4836
rect 621 4664 627 4696
rect 637 4624 643 4676
rect 653 4603 659 4696
rect 637 4597 659 4603
rect 541 4544 547 4556
rect 493 4484 499 4516
rect 445 4304 451 4436
rect 292 4297 307 4303
rect 285 4164 291 4296
rect 381 4264 387 4276
rect 317 4224 323 4256
rect 365 4184 371 4236
rect 397 4124 403 4276
rect 429 4144 435 4216
rect 365 3944 371 4096
rect 397 3904 403 4116
rect 429 3984 435 4136
rect 445 4124 451 4156
rect 461 3984 467 4476
rect 493 4124 499 4356
rect 541 4284 547 4536
rect 589 4504 595 4516
rect 637 4284 643 4597
rect 733 4543 739 4696
rect 813 4684 819 4696
rect 717 4537 739 4543
rect 717 4524 723 4537
rect 733 4484 739 4516
rect 509 4104 515 4116
rect 349 3704 355 3856
rect 365 3724 371 3896
rect 381 3763 387 3836
rect 397 3784 403 3816
rect 381 3757 403 3763
rect 397 3704 403 3757
rect 429 3744 435 3836
rect 317 3684 323 3696
rect 285 3584 291 3636
rect 237 3577 259 3583
rect 237 3504 243 3577
rect 349 3484 355 3676
rect 77 3324 83 3396
rect 141 3344 147 3416
rect 173 3364 179 3456
rect 349 3364 355 3476
rect 45 3244 51 3296
rect 173 3244 179 3356
rect 413 3324 419 3556
rect 429 3544 435 3616
rect 477 3584 483 3836
rect 525 3744 531 4236
rect 557 4024 563 4116
rect 541 3904 547 3916
rect 573 3904 579 4256
rect 637 4244 643 4276
rect 669 4144 675 4336
rect 717 4304 723 4356
rect 733 4324 739 4336
rect 733 4304 739 4316
rect 621 4124 627 4136
rect 717 4124 723 4156
rect 589 4104 595 4116
rect 749 4043 755 4636
rect 781 4544 787 4676
rect 797 4664 803 4676
rect 813 4544 819 4616
rect 861 4544 867 4696
rect 781 4304 787 4456
rect 733 4037 755 4043
rect 765 4297 780 4303
rect 653 3984 659 4036
rect 669 3904 675 3976
rect 733 3924 739 4037
rect 749 3904 755 4016
rect 557 3744 563 3876
rect 701 3764 707 3836
rect 573 3724 579 3736
rect 493 3584 499 3716
rect 557 3703 563 3716
rect 589 3704 595 3716
rect 557 3697 579 3703
rect 573 3584 579 3697
rect 637 3644 643 3716
rect 669 3664 675 3736
rect 765 3644 771 4297
rect 797 4024 803 4516
rect 813 4344 819 4536
rect 829 4524 835 4536
rect 877 4523 883 4696
rect 893 4584 899 4897
rect 909 4784 915 5036
rect 925 5004 931 5036
rect 941 4984 947 5036
rect 989 4944 995 5296
rect 1005 5284 1011 5316
rect 1021 5144 1027 5476
rect 1053 5423 1059 5494
rect 1453 5464 1459 5496
rect 1565 5484 1571 5536
rect 2061 5524 2067 5576
rect 2605 5524 2611 5576
rect 3325 5524 3331 5576
rect 1037 5417 1059 5423
rect 1037 5384 1043 5417
rect 1037 5304 1043 5356
rect 1085 5344 1091 5356
rect 1053 5224 1059 5316
rect 1101 5304 1107 5436
rect 1165 5304 1171 5396
rect 1181 5384 1187 5416
rect 1373 5404 1379 5436
rect 1597 5423 1603 5456
rect 1581 5417 1603 5423
rect 1581 5364 1587 5417
rect 1581 5344 1587 5356
rect 1053 5104 1059 5136
rect 1101 5124 1107 5296
rect 1005 5044 1011 5096
rect 1149 5064 1155 5116
rect 1165 5084 1171 5296
rect 1229 5184 1235 5316
rect 1245 5304 1251 5336
rect 1325 5184 1331 5276
rect 1309 5104 1315 5116
rect 1421 5104 1427 5236
rect 1261 5084 1267 5096
rect 1165 5064 1171 5076
rect 1053 4944 1059 4996
rect 925 4824 931 4896
rect 989 4784 995 4916
rect 1021 4824 1027 4936
rect 1069 4904 1075 4976
rect 1117 4944 1123 5036
rect 1133 5004 1139 5036
rect 1181 4944 1187 5036
rect 1197 4944 1203 5056
rect 1245 4924 1251 5036
rect 1277 4964 1283 5096
rect 1277 4944 1283 4956
rect 941 4684 947 4696
rect 957 4663 963 4696
rect 941 4657 963 4663
rect 877 4517 899 4523
rect 877 4484 883 4496
rect 813 4284 819 4336
rect 893 4304 899 4517
rect 909 4304 915 4516
rect 941 4464 947 4657
rect 973 4324 979 4776
rect 1021 4704 1027 4816
rect 1005 4544 1011 4596
rect 989 4444 995 4516
rect 1005 4323 1011 4516
rect 1021 4504 1027 4696
rect 1037 4684 1043 4696
rect 1069 4624 1075 4636
rect 1085 4524 1091 4916
rect 1133 4884 1139 4896
rect 1005 4317 1027 4323
rect 813 4144 819 4276
rect 829 4084 835 4096
rect 861 4064 867 4116
rect 861 3924 867 4036
rect 893 3904 899 4296
rect 909 4224 915 4296
rect 941 4284 947 4316
rect 925 4244 931 4276
rect 925 4164 931 4236
rect 957 4204 963 4236
rect 973 4184 979 4316
rect 1005 4284 1011 4296
rect 1005 4184 1011 4256
rect 957 4144 963 4156
rect 989 4137 1004 4143
rect 957 4103 963 4136
rect 973 4104 979 4136
rect 941 4097 963 4103
rect 909 4044 915 4096
rect 925 3984 931 4056
rect 781 3764 787 3796
rect 781 3744 787 3756
rect 781 3684 787 3696
rect 429 3524 435 3536
rect 509 3484 515 3516
rect 685 3504 691 3636
rect 781 3584 787 3676
rect 797 3584 803 3896
rect 813 3784 819 3896
rect 893 3844 899 3896
rect 829 3764 835 3836
rect 845 3704 851 3776
rect 909 3763 915 3896
rect 941 3804 947 4097
rect 957 3904 963 4036
rect 989 3984 995 4137
rect 1021 4124 1027 4317
rect 1053 4264 1059 4496
rect 1069 4484 1075 4496
rect 1101 4484 1107 4876
rect 1117 4764 1123 4836
rect 1165 4804 1171 4836
rect 1149 4724 1155 4736
rect 1117 4704 1123 4716
rect 1165 4624 1171 4696
rect 1181 4644 1187 4736
rect 1213 4724 1219 4756
rect 1277 4724 1283 4736
rect 1261 4684 1267 4696
rect 1277 4664 1283 4696
rect 1149 4617 1164 4623
rect 1149 4524 1155 4617
rect 1149 4484 1155 4496
rect 1181 4483 1187 4636
rect 1293 4583 1299 4996
rect 1309 4984 1315 5056
rect 1316 4717 1347 4723
rect 1341 4684 1347 4717
rect 1309 4677 1324 4683
rect 1309 4584 1315 4677
rect 1277 4577 1299 4583
rect 1213 4524 1219 4536
rect 1261 4524 1267 4536
rect 1277 4524 1283 4577
rect 1172 4477 1187 4483
rect 1085 4284 1091 4336
rect 1101 4284 1107 4296
rect 1133 4284 1139 4316
rect 1149 4304 1155 4316
rect 1037 4104 1043 4176
rect 1069 4104 1075 4196
rect 1165 4184 1171 4416
rect 1181 4344 1187 4436
rect 1181 4224 1187 4296
rect 1197 4244 1203 4276
rect 1229 4264 1235 4436
rect 1277 4364 1283 4516
rect 1293 4404 1299 4556
rect 1325 4384 1331 4536
rect 1341 4524 1347 4656
rect 1341 4424 1347 4516
rect 1341 4344 1347 4396
rect 1293 4324 1299 4336
rect 1341 4304 1347 4336
rect 1213 4164 1219 4256
rect 1245 4224 1251 4276
rect 1261 4244 1267 4296
rect 1245 4184 1251 4216
rect 1293 4183 1299 4236
rect 1309 4224 1315 4256
rect 1293 4177 1315 4183
rect 1101 4124 1107 4136
rect 1117 4117 1132 4123
rect 1117 3924 1123 4117
rect 1277 4044 1283 4156
rect 1309 4144 1315 4177
rect 1325 4124 1331 4136
rect 1357 4104 1363 4596
rect 1373 4464 1379 5096
rect 1421 5064 1427 5096
rect 1405 5004 1411 5036
rect 1469 4964 1475 5336
rect 1613 5324 1619 5336
rect 1773 5324 1779 5496
rect 1837 5484 1843 5496
rect 1837 5464 1843 5476
rect 1933 5424 1939 5476
rect 1965 5404 1971 5516
rect 2013 5384 2019 5496
rect 1885 5344 1891 5356
rect 1917 5344 1923 5356
rect 1677 5244 1683 5316
rect 1709 5244 1715 5296
rect 1496 5206 1502 5214
rect 1510 5206 1516 5214
rect 1524 5206 1530 5214
rect 1538 5206 1544 5214
rect 1597 4924 1603 5236
rect 1725 5104 1731 5296
rect 1821 5244 1827 5300
rect 1693 5044 1699 5056
rect 1693 4924 1699 5036
rect 1725 5024 1731 5096
rect 1837 5084 1843 5096
rect 1741 5064 1747 5076
rect 1741 4964 1747 5056
rect 1773 4944 1779 5036
rect 1917 5004 1923 5336
rect 2045 5324 2051 5496
rect 2157 5484 2163 5496
rect 2269 5484 2275 5496
rect 2189 5364 2195 5456
rect 2413 5424 2419 5476
rect 2477 5424 2483 5476
rect 2509 5444 2515 5516
rect 2557 5464 2563 5496
rect 2621 5484 2627 5496
rect 2173 5344 2179 5356
rect 2205 5344 2211 5416
rect 2269 5384 2275 5396
rect 2205 5304 2211 5336
rect 2029 5124 2035 5176
rect 1965 5004 1971 5036
rect 1389 4604 1395 4716
rect 1405 4624 1411 4656
rect 1437 4644 1443 4696
rect 1453 4684 1459 4776
rect 1469 4704 1475 4916
rect 1597 4844 1603 4896
rect 1496 4806 1502 4814
rect 1510 4806 1516 4814
rect 1524 4806 1530 4814
rect 1538 4806 1544 4814
rect 1405 4524 1411 4556
rect 1389 4504 1395 4516
rect 1421 4504 1427 4636
rect 1437 4504 1443 4596
rect 1469 4584 1475 4696
rect 1485 4524 1491 4676
rect 1501 4584 1507 4716
rect 1549 4704 1555 4716
rect 1693 4704 1699 4716
rect 1709 4704 1715 4836
rect 1405 4364 1411 4436
rect 1373 4124 1379 4356
rect 1421 4184 1427 4496
rect 1549 4444 1555 4696
rect 1496 4406 1502 4414
rect 1510 4406 1516 4414
rect 1524 4406 1530 4414
rect 1538 4406 1544 4414
rect 1565 4324 1571 4516
rect 1581 4324 1587 4436
rect 1453 4304 1459 4316
rect 1389 4124 1395 4136
rect 1469 4124 1475 4316
rect 1565 4284 1571 4296
rect 1501 4204 1507 4276
rect 1325 3944 1331 4036
rect 1309 3924 1315 3936
rect 1389 3923 1395 4116
rect 1380 3917 1395 3923
rect 973 3904 979 3916
rect 1069 3904 1075 3916
rect 1117 3904 1123 3916
rect 1421 3904 1427 4036
rect 909 3757 931 3763
rect 893 3724 899 3756
rect 909 3664 915 3736
rect 909 3524 915 3636
rect 925 3504 931 3757
rect 941 3524 947 3536
rect 445 3364 451 3456
rect 509 3364 515 3456
rect 13 3084 19 3196
rect 125 3184 131 3236
rect 189 3124 195 3176
rect 13 2944 19 3076
rect 45 2724 51 2776
rect 173 2664 179 2936
rect 189 2924 195 3096
rect 317 3064 323 3236
rect 381 3204 387 3236
rect 445 3184 451 3356
rect 493 3084 499 3236
rect 509 3183 515 3356
rect 525 3324 531 3456
rect 525 3224 531 3316
rect 509 3177 524 3183
rect 573 3104 579 3236
rect 589 2964 595 3456
rect 605 3384 611 3416
rect 685 3364 691 3476
rect 813 3424 819 3456
rect 909 3404 915 3496
rect 989 3484 995 3876
rect 1005 3684 1011 3856
rect 1037 3724 1043 3836
rect 1085 3744 1091 3816
rect 1117 3764 1123 3796
rect 1149 3784 1155 3876
rect 1181 3724 1187 3896
rect 1213 3864 1219 3876
rect 1197 3744 1203 3856
rect 1213 3824 1219 3856
rect 1021 3704 1027 3716
rect 1197 3584 1203 3736
rect 1053 3504 1059 3516
rect 1133 3504 1139 3516
rect 1117 3463 1123 3476
rect 1149 3463 1155 3496
rect 1117 3457 1155 3463
rect 941 3364 947 3416
rect 285 2944 291 2956
rect 317 2944 323 2956
rect 189 2844 195 2896
rect 285 2704 291 2916
rect 541 2904 547 2916
rect 589 2904 595 2936
rect 605 2924 611 3216
rect 685 3064 691 3356
rect 797 3124 803 3316
rect 893 3244 899 3296
rect 813 3124 819 3176
rect 797 3104 803 3116
rect 957 3104 963 3316
rect 1021 3184 1027 3456
rect 1085 3344 1091 3356
rect 1165 3324 1171 3476
rect 1197 3424 1203 3516
rect 1213 3503 1219 3716
rect 1229 3524 1235 3636
rect 1213 3497 1228 3503
rect 1245 3484 1251 3736
rect 1277 3724 1283 3836
rect 1325 3804 1331 3876
rect 1341 3844 1347 3896
rect 1389 3884 1395 3896
rect 1293 3724 1299 3756
rect 1389 3724 1395 3836
rect 1421 3724 1427 3756
rect 1437 3744 1443 3876
rect 1261 3644 1267 3696
rect 1277 3504 1283 3716
rect 1389 3704 1395 3716
rect 1421 3704 1427 3716
rect 1437 3664 1443 3736
rect 1453 3684 1459 3716
rect 1245 3384 1251 3416
rect 1277 3324 1283 3476
rect 1293 3444 1299 3496
rect 1309 3484 1315 3656
rect 1341 3504 1347 3536
rect 1421 3504 1427 3636
rect 1469 3544 1475 4116
rect 1501 4104 1507 4176
rect 1565 4144 1571 4156
rect 1597 4123 1603 4576
rect 1613 4504 1619 4516
rect 1629 4324 1635 4496
rect 1645 4464 1651 4696
rect 1661 4484 1667 4636
rect 1677 4564 1683 4616
rect 1709 4563 1715 4696
rect 1693 4557 1715 4563
rect 1677 4524 1683 4556
rect 1693 4524 1699 4557
rect 1741 4544 1747 4696
rect 1757 4564 1763 4836
rect 1773 4704 1779 4716
rect 1789 4684 1795 4756
rect 1821 4704 1827 4976
rect 1917 4964 1923 4996
rect 1853 4724 1859 4736
rect 1805 4664 1811 4696
rect 1837 4664 1843 4716
rect 1837 4604 1843 4656
rect 1853 4604 1859 4716
rect 1965 4684 1971 4696
rect 2013 4684 2019 4956
rect 2045 4924 2051 5096
rect 2045 4844 2051 4896
rect 2045 4684 2051 4696
rect 2093 4684 2099 4876
rect 2125 4844 2131 5076
rect 2157 5004 2163 5056
rect 2237 5024 2243 5096
rect 2253 5044 2259 5336
rect 2333 5144 2339 5236
rect 2429 5184 2435 5336
rect 2621 5323 2627 5476
rect 2701 5404 2707 5476
rect 3373 5464 3379 5643
rect 2733 5364 2739 5456
rect 2893 5364 2899 5436
rect 2925 5384 2931 5416
rect 2989 5364 2995 5416
rect 2621 5317 2636 5323
rect 2381 5064 2387 5096
rect 2413 5084 2419 5096
rect 2141 4784 2147 4936
rect 2189 4704 2195 4716
rect 1773 4544 1779 4576
rect 1853 4544 1859 4596
rect 1677 4384 1683 4436
rect 1677 4304 1683 4316
rect 1709 4284 1715 4536
rect 1725 4304 1731 4516
rect 1757 4504 1763 4516
rect 1773 4323 1779 4436
rect 1805 4384 1811 4516
rect 1837 4384 1843 4496
rect 1764 4317 1779 4323
rect 1693 4264 1699 4276
rect 1588 4117 1603 4123
rect 1496 4006 1502 4014
rect 1510 4006 1516 4014
rect 1524 4006 1530 4014
rect 1538 4006 1544 4014
rect 1565 3904 1571 4116
rect 1581 3984 1587 4056
rect 1613 3984 1619 4076
rect 1629 4064 1635 4136
rect 1645 4124 1651 4216
rect 1709 4084 1715 4276
rect 1725 4184 1731 4256
rect 1805 4244 1811 4296
rect 1933 4284 1939 4536
rect 1965 4504 1971 4596
rect 2045 4563 2051 4676
rect 2036 4557 2051 4563
rect 1981 4524 1987 4556
rect 2029 4524 2035 4556
rect 2013 4344 2019 4436
rect 1949 4304 1955 4336
rect 2061 4303 2067 4636
rect 2077 4584 2083 4636
rect 2093 4544 2099 4676
rect 2093 4484 2099 4536
rect 2109 4504 2115 4536
rect 2125 4344 2131 4676
rect 2141 4644 2147 4696
rect 2221 4684 2227 4696
rect 2237 4684 2243 4716
rect 2253 4584 2259 4836
rect 2301 4784 2307 4936
rect 2365 4744 2371 5036
rect 2381 4724 2387 4916
rect 2397 4844 2403 4896
rect 2413 4704 2419 5056
rect 2445 4984 2451 5116
rect 2461 5064 2467 5076
rect 2525 5064 2531 5316
rect 2557 5244 2563 5296
rect 2557 5120 2563 5158
rect 2621 5104 2627 5317
rect 2637 5244 2643 5296
rect 2284 4664 2292 4670
rect 2221 4544 2227 4556
rect 2301 4524 2307 4636
rect 2365 4544 2371 4636
rect 2397 4544 2403 4696
rect 2413 4664 2419 4676
rect 2077 4324 2083 4336
rect 2141 4324 2147 4376
rect 2253 4364 2259 4496
rect 2205 4324 2211 4336
rect 2301 4324 2307 4516
rect 2189 4304 2195 4316
rect 2052 4297 2067 4303
rect 1821 4264 1827 4276
rect 1933 4204 1939 4276
rect 2045 4224 2051 4296
rect 2141 4204 2147 4236
rect 1981 4164 1987 4196
rect 1741 4124 1747 4156
rect 2157 4144 2163 4236
rect 2173 4164 2179 4236
rect 2253 4164 2259 4256
rect 2269 4184 2275 4296
rect 2301 4244 2307 4296
rect 2381 4284 2387 4436
rect 2429 4384 2435 4676
rect 2445 4644 2451 4916
rect 2461 4884 2467 5056
rect 2477 5024 2483 5056
rect 2477 4984 2483 5016
rect 2509 4944 2515 4956
rect 2461 4664 2467 4876
rect 2477 4644 2483 4696
rect 2509 4604 2515 4716
rect 2525 4664 2531 4836
rect 2541 4704 2547 5096
rect 2653 5064 2659 5356
rect 2989 5344 2995 5356
rect 2733 5224 2739 5336
rect 3005 5224 3011 5456
rect 3032 5406 3038 5414
rect 3046 5406 3052 5414
rect 3060 5406 3066 5414
rect 3074 5406 3080 5414
rect 3021 5344 3027 5376
rect 3197 5364 3203 5456
rect 3421 5404 3427 5496
rect 3101 5344 3107 5356
rect 2813 5184 2819 5216
rect 2877 5124 2883 5176
rect 3133 5104 3139 5296
rect 3181 5243 3187 5296
rect 3172 5237 3187 5243
rect 3181 5144 3187 5237
rect 3197 5124 3203 5356
rect 3357 5344 3363 5356
rect 3453 5324 3459 5496
rect 3421 5262 3427 5300
rect 3469 5224 3475 5516
rect 3501 5484 3507 5496
rect 3517 5464 3523 5476
rect 3533 5464 3539 5643
rect 3501 5304 3507 5336
rect 3533 5324 3539 5396
rect 3565 5383 3571 5643
rect 3581 5404 3587 5496
rect 3645 5484 3651 5496
rect 3629 5464 3635 5476
rect 3565 5377 3587 5383
rect 3581 5364 3587 5377
rect 3645 5324 3651 5476
rect 3661 5344 3667 5456
rect 3709 5384 3715 5436
rect 3725 5364 3731 5643
rect 4568 5606 4574 5614
rect 4582 5606 4588 5614
rect 4596 5606 4602 5614
rect 4610 5606 4616 5614
rect 3965 5520 3971 5558
rect 3901 5484 3907 5496
rect 3293 5144 3299 5216
rect 3565 5144 3571 5276
rect 3661 5224 3667 5336
rect 2653 4944 2659 5056
rect 2797 4904 2803 5096
rect 2813 4984 2819 5036
rect 2669 4704 2675 4756
rect 2525 4603 2531 4656
rect 2669 4623 2675 4676
rect 2653 4617 2675 4623
rect 2525 4597 2547 4603
rect 2461 4524 2467 4596
rect 2541 4564 2547 4597
rect 2573 4524 2579 4536
rect 2653 4484 2659 4617
rect 2749 4544 2755 4556
rect 2765 4544 2771 4556
rect 2781 4524 2787 4636
rect 2829 4544 2835 4916
rect 2845 4884 2851 4936
rect 2429 4324 2435 4376
rect 2317 4264 2323 4276
rect 2333 4244 2339 4276
rect 2349 4144 2355 4236
rect 2381 4164 2387 4276
rect 2381 4144 2387 4156
rect 2301 4124 2307 4136
rect 1805 4104 1811 4116
rect 1885 4062 1891 4100
rect 1773 4004 1779 4036
rect 1565 3884 1571 3896
rect 1869 3884 1875 3996
rect 1949 3904 1955 4116
rect 2237 4104 2243 4116
rect 2381 4103 2387 4136
rect 2397 4124 2403 4136
rect 2413 4123 2419 4316
rect 2461 4304 2467 4476
rect 2669 4444 2675 4496
rect 2461 4184 2467 4296
rect 2477 4164 2483 4236
rect 2404 4117 2419 4123
rect 2372 4097 2387 4103
rect 2029 3984 2035 4016
rect 2221 4004 2227 4036
rect 1965 3924 1971 3976
rect 2045 3924 2051 3976
rect 2093 3924 2099 3936
rect 2205 3920 2211 3958
rect 2493 3944 2499 4416
rect 2717 4344 2723 4436
rect 2733 4384 2739 4516
rect 2781 4384 2787 4516
rect 2525 4244 2531 4316
rect 2557 4304 2563 4316
rect 2685 4304 2691 4336
rect 2781 4324 2787 4356
rect 2541 4244 2547 4296
rect 2589 4264 2595 4296
rect 2653 4284 2659 4296
rect 2669 4284 2675 4296
rect 2596 4257 2611 4263
rect 2541 4184 2547 4236
rect 2589 4124 2595 4136
rect 2605 4104 2611 4257
rect 2701 4244 2707 4296
rect 2733 4184 2739 4276
rect 2621 4144 2627 4156
rect 2669 4144 2675 4156
rect 2765 4144 2771 4316
rect 2813 4304 2819 4436
rect 2845 4384 2851 4856
rect 2877 4724 2883 5096
rect 2893 4984 2899 5076
rect 3197 5064 3203 5116
rect 3032 5006 3038 5014
rect 3046 5006 3052 5014
rect 3060 5006 3066 5014
rect 3074 5006 3080 5014
rect 2893 4744 2899 4896
rect 2925 4864 2931 4916
rect 2925 4724 2931 4736
rect 2941 4704 2947 4976
rect 3021 4904 3027 4976
rect 3149 4964 3155 5016
rect 3197 4984 3203 5036
rect 3293 4984 3299 5096
rect 3357 5084 3363 5116
rect 3677 5104 3683 5356
rect 3773 5324 3779 5396
rect 3869 5364 3875 5456
rect 4125 5324 4131 5496
rect 4173 5464 4179 5476
rect 4205 5443 4211 5516
rect 4253 5504 4259 5536
rect 4941 5524 4947 5536
rect 5220 5517 5235 5523
rect 4196 5437 4211 5443
rect 4173 5344 4179 5356
rect 3725 5304 3731 5316
rect 3709 5284 3715 5296
rect 4093 5244 4099 5300
rect 4125 5244 4131 5316
rect 3325 5043 3331 5076
rect 3325 5037 3347 5043
rect 3309 4984 3315 5036
rect 3149 4924 3155 4956
rect 3245 4944 3251 4956
rect 3101 4904 3107 4916
rect 2989 4824 2995 4836
rect 3005 4784 3011 4876
rect 3165 4704 3171 4756
rect 2893 4584 2899 4676
rect 2861 4544 2867 4556
rect 2925 4544 2931 4636
rect 2957 4564 2963 4636
rect 2861 4524 2867 4536
rect 2797 4184 2803 4236
rect 2781 4144 2787 4156
rect 2813 4144 2819 4276
rect 2829 4224 2835 4256
rect 2637 4124 2643 4136
rect 2653 4124 2659 4136
rect 2781 4124 2787 4136
rect 2637 4044 2643 4116
rect 2829 4104 2835 4176
rect 2845 4164 2851 4296
rect 2845 4144 2851 4156
rect 2861 4124 2867 4516
rect 2973 4464 2979 4656
rect 3037 4644 3043 4696
rect 3149 4623 3155 4656
rect 3133 4617 3155 4623
rect 3032 4606 3038 4614
rect 3046 4606 3052 4614
rect 3060 4606 3066 4614
rect 3074 4606 3080 4614
rect 3133 4564 3139 4617
rect 3181 4604 3187 4916
rect 3229 4864 3235 4916
rect 3293 4884 3299 4896
rect 3309 4844 3315 4956
rect 3341 4944 3347 5037
rect 3341 4924 3347 4936
rect 3357 4924 3363 5056
rect 3517 5004 3523 5036
rect 3405 4924 3411 4936
rect 3341 4704 3347 4916
rect 3421 4904 3427 4996
rect 3581 4944 3587 4956
rect 3693 4944 3699 5216
rect 4061 5184 4067 5216
rect 4173 5184 4179 5276
rect 3460 4917 3475 4923
rect 3325 4684 3331 4696
rect 3357 4684 3363 4836
rect 3373 4784 3379 4856
rect 3053 4444 3059 4516
rect 2877 4324 2883 4336
rect 2957 4304 2963 4436
rect 2973 4404 2979 4436
rect 1972 3897 1980 3903
rect 1485 3704 1491 3776
rect 1517 3644 1523 3856
rect 1613 3744 1619 3836
rect 1661 3744 1667 3856
rect 1725 3784 1731 3836
rect 1725 3764 1731 3776
rect 1496 3606 1502 3614
rect 1510 3606 1516 3614
rect 1524 3606 1530 3614
rect 1538 3606 1544 3614
rect 1565 3584 1571 3736
rect 1613 3544 1619 3736
rect 1981 3724 1987 3896
rect 2077 3864 2083 3876
rect 2013 3844 2019 3856
rect 2045 3744 2051 3836
rect 1805 3662 1811 3700
rect 1981 3624 1987 3716
rect 2093 3704 2099 3916
rect 2125 3884 2131 3916
rect 2573 3904 2579 4036
rect 2685 3924 2691 3976
rect 2141 3784 2147 3856
rect 2189 3744 2195 3776
rect 2269 3744 2275 3776
rect 2285 3724 2291 3816
rect 2301 3764 2307 3856
rect 2493 3804 2499 3876
rect 2525 3803 2531 3836
rect 2573 3824 2579 3896
rect 2525 3797 2547 3803
rect 2317 3784 2323 3796
rect 2509 3764 2515 3796
rect 1821 3524 1827 3576
rect 1428 3497 1443 3503
rect 1341 3344 1347 3356
rect 1037 3224 1043 3316
rect 1421 3204 1427 3476
rect 1437 3384 1443 3497
rect 1549 3457 1564 3463
rect 1453 3384 1459 3396
rect 1533 3364 1539 3436
rect 1549 3384 1555 3457
rect 1496 3206 1502 3214
rect 1510 3206 1516 3214
rect 1524 3206 1530 3214
rect 1538 3206 1544 3214
rect 1389 3124 1395 3176
rect 1181 3104 1187 3116
rect 1373 3104 1379 3116
rect 1581 3104 1587 3496
rect 1693 3424 1699 3436
rect 1725 3404 1731 3496
rect 1741 3444 1747 3496
rect 1917 3484 1923 3596
rect 2029 3504 2035 3616
rect 2109 3604 2115 3636
rect 2189 3504 2195 3616
rect 2205 3584 2211 3676
rect 2221 3584 2227 3616
rect 2125 3484 2131 3496
rect 1949 3424 1955 3456
rect 1741 3344 1747 3416
rect 1917 3324 1923 3336
rect 1693 3104 1699 3116
rect 1805 3104 1811 3316
rect 1885 3304 1891 3316
rect 1837 3244 1843 3296
rect 1965 3184 1971 3396
rect 2109 3364 2115 3416
rect 2013 3244 2019 3300
rect 2077 3244 2083 3336
rect 2109 3224 2115 3356
rect 2205 3324 2211 3576
rect 2269 3384 2275 3416
rect 2301 3344 2307 3476
rect 2189 3264 2195 3316
rect 2301 3284 2307 3336
rect 2317 3304 2323 3676
rect 2333 3484 2339 3496
rect 2349 3384 2355 3596
rect 2381 3524 2387 3576
rect 2509 3464 2515 3756
rect 2541 3744 2547 3797
rect 2605 3744 2611 3836
rect 2669 3724 2675 3896
rect 2781 3884 2787 4096
rect 2829 3984 2835 4076
rect 2893 3904 2899 4156
rect 2941 4104 2947 4196
rect 2957 4164 2963 4296
rect 3133 4264 3139 4556
rect 3261 4444 3267 4496
rect 3277 4384 3283 4676
rect 3357 4644 3363 4676
rect 3405 4624 3411 4636
rect 3421 4564 3427 4896
rect 3437 4564 3443 4836
rect 3469 4704 3475 4917
rect 3309 4484 3315 4496
rect 3165 4324 3171 4376
rect 3469 4364 3475 4696
rect 3485 4644 3491 4916
rect 3549 4884 3555 4916
rect 3565 4904 3571 4916
rect 3549 4704 3555 4736
rect 3565 4704 3571 4796
rect 3533 4524 3539 4616
rect 3469 4324 3475 4336
rect 3485 4304 3491 4436
rect 3565 4384 3571 4696
rect 3581 4684 3587 4936
rect 3645 4884 3651 4896
rect 3597 4704 3603 4836
rect 3645 4764 3651 4876
rect 3645 4704 3651 4716
rect 3661 4704 3667 4776
rect 3677 4744 3683 4916
rect 3709 4804 3715 4916
rect 3725 4844 3731 5136
rect 3757 5124 3763 5136
rect 3789 5104 3795 5116
rect 3917 5104 3923 5116
rect 4093 5104 4099 5136
rect 3757 5097 3772 5103
rect 3725 4724 3731 4836
rect 3757 4784 3763 5097
rect 3789 4924 3795 5036
rect 3837 5024 3843 5096
rect 3837 4984 3843 5016
rect 3869 4964 3875 5076
rect 3773 4884 3779 4916
rect 3869 4904 3875 4956
rect 3917 4924 3923 5016
rect 3933 5004 3939 5036
rect 3965 4944 3971 5076
rect 3645 4664 3651 4696
rect 3501 4304 3507 4376
rect 3549 4304 3555 4316
rect 3032 4206 3038 4214
rect 3046 4206 3052 4214
rect 3060 4206 3066 4214
rect 3074 4206 3080 4214
rect 3165 4164 3171 4256
rect 3037 4124 3043 4156
rect 3165 4124 3171 4156
rect 2813 3804 2819 3856
rect 2637 3644 2643 3696
rect 2589 3504 2595 3516
rect 2701 3504 2707 3696
rect 2733 3684 2739 3716
rect 2733 3564 2739 3676
rect 2813 3584 2819 3776
rect 2845 3584 2851 3816
rect 2861 3784 2867 3796
rect 3005 3784 3011 4116
rect 3069 4044 3075 4100
rect 3261 4004 3267 4256
rect 3373 4144 3379 4276
rect 3373 4124 3379 4136
rect 3421 4124 3427 4156
rect 3533 4104 3539 4176
rect 3549 4144 3555 4276
rect 3565 4124 3571 4356
rect 3581 4284 3587 4536
rect 3613 4524 3619 4536
rect 3645 4504 3651 4556
rect 3661 4524 3667 4696
rect 3725 4684 3731 4716
rect 3789 4704 3795 4896
rect 3917 4704 3923 4796
rect 3933 4724 3939 4756
rect 3965 4723 3971 4936
rect 3997 4904 4003 4936
rect 4029 4744 4035 5096
rect 4109 5064 4115 5116
rect 4045 4984 4051 5016
rect 4189 4964 4195 5336
rect 4205 5104 4211 5437
rect 4301 5344 4307 5456
rect 4349 5444 4355 5476
rect 4349 5344 4355 5436
rect 4381 5384 4387 5476
rect 4301 5224 4307 5336
rect 4381 5324 4387 5336
rect 4317 5204 4323 5236
rect 4260 5097 4275 5103
rect 4205 4983 4211 5096
rect 4221 5044 4227 5096
rect 4221 5024 4227 5036
rect 4205 4977 4227 4983
rect 4189 4944 4195 4956
rect 4061 4884 4067 4896
rect 4061 4844 4067 4876
rect 3965 4717 3987 4723
rect 3693 4544 3699 4556
rect 3725 4524 3731 4576
rect 3757 4524 3763 4596
rect 3773 4524 3779 4576
rect 3677 4504 3683 4516
rect 3757 4444 3763 4516
rect 3581 4184 3587 4276
rect 3645 4204 3651 4316
rect 3677 4304 3683 4356
rect 3725 4304 3731 4376
rect 3789 4304 3795 4696
rect 3885 4644 3891 4676
rect 3821 4384 3827 4496
rect 3821 4304 3827 4356
rect 3645 4124 3651 4156
rect 3661 4144 3667 4176
rect 3677 4164 3683 4196
rect 3741 4164 3747 4236
rect 3773 4204 3779 4296
rect 3700 4157 3731 4163
rect 3725 4144 3731 4157
rect 3373 3984 3379 3996
rect 3085 3924 3091 3976
rect 3032 3806 3038 3814
rect 3046 3806 3052 3814
rect 3060 3806 3066 3814
rect 3074 3806 3080 3814
rect 3117 3724 3123 3896
rect 3181 3824 3187 3876
rect 3133 3784 3139 3816
rect 3213 3784 3219 3836
rect 3293 3764 3299 3976
rect 3501 3864 3507 4076
rect 3709 4004 3715 4136
rect 3757 4104 3763 4116
rect 3773 4104 3779 4196
rect 3837 4183 3843 4536
rect 3869 4524 3875 4536
rect 3853 4444 3859 4516
rect 3853 4324 3859 4436
rect 3828 4177 3843 4183
rect 3805 4124 3811 4156
rect 3821 4144 3827 4176
rect 3853 4163 3859 4296
rect 3885 4284 3891 4636
rect 3933 4304 3939 4636
rect 3965 4624 3971 4696
rect 3981 4684 3987 4717
rect 4045 4684 4051 4716
rect 3997 4664 4003 4676
rect 4045 4664 4051 4676
rect 3965 4304 3971 4596
rect 3981 4544 3987 4656
rect 3997 4524 4003 4536
rect 4013 4504 4019 4636
rect 4061 4304 4067 4336
rect 4077 4304 4083 4776
rect 4093 4704 4099 4756
rect 4109 4724 4115 4936
rect 4205 4924 4211 4956
rect 4109 4624 4115 4716
rect 4125 4523 4131 4556
rect 4141 4524 4147 4736
rect 4221 4684 4227 4977
rect 4269 4844 4275 5097
rect 4285 5084 4291 5116
rect 4333 5043 4339 5316
rect 4381 5204 4387 5296
rect 4397 5284 4403 5496
rect 4477 5344 4483 5496
rect 4493 5464 4499 5476
rect 4509 5404 4515 5436
rect 4509 5344 4515 5376
rect 4557 5364 4563 5456
rect 4445 5284 4451 5318
rect 4349 5064 4355 5096
rect 4333 5037 4355 5043
rect 4253 4684 4259 4836
rect 4269 4724 4275 4796
rect 4205 4644 4211 4656
rect 4157 4544 4163 4616
rect 4116 4517 4131 4523
rect 4237 4523 4243 4636
rect 4285 4563 4291 5036
rect 4301 4804 4307 4856
rect 4301 4724 4307 4796
rect 4317 4744 4323 5036
rect 4349 4984 4355 5037
rect 4333 4924 4339 4976
rect 4381 4924 4387 5196
rect 4525 5184 4531 5256
rect 4541 5104 4547 5316
rect 4573 5284 4579 5476
rect 4589 5324 4595 5436
rect 4568 5206 4574 5214
rect 4582 5206 4588 5214
rect 4596 5206 4602 5214
rect 4610 5206 4616 5214
rect 4333 4704 4339 4796
rect 4381 4764 4387 4916
rect 4349 4704 4355 4756
rect 4381 4684 4387 4716
rect 4397 4704 4403 4916
rect 4413 4903 4419 4936
rect 4445 4924 4451 5036
rect 4477 4984 4483 5096
rect 4541 5084 4547 5096
rect 4436 4917 4444 4923
rect 4413 4897 4435 4903
rect 4413 4704 4419 4736
rect 4429 4724 4435 4897
rect 4461 4884 4467 4896
rect 4461 4744 4467 4876
rect 4477 4784 4483 4796
rect 4493 4784 4499 5036
rect 4557 5024 4563 5096
rect 4637 5064 4643 5516
rect 5213 5504 5219 5516
rect 4685 5444 4691 5496
rect 4669 5344 4675 5356
rect 4749 5344 4755 5376
rect 4781 5344 4787 5496
rect 4813 5384 4819 5476
rect 4653 5324 4659 5336
rect 4829 5324 4835 5496
rect 4861 5484 4867 5496
rect 4861 5344 4867 5436
rect 4877 5344 4883 5376
rect 4909 5344 4915 5496
rect 4925 5444 4931 5476
rect 4925 5364 4931 5436
rect 5101 5424 5107 5476
rect 5133 5444 5139 5476
rect 4989 5344 4995 5356
rect 5021 5344 5027 5416
rect 5149 5344 5155 5496
rect 4845 5324 4851 5336
rect 4925 5324 4931 5336
rect 4973 5324 4979 5336
rect 5197 5324 5203 5496
rect 5229 5464 5235 5517
rect 5229 5344 5235 5456
rect 5261 5364 5267 5496
rect 5277 5484 5283 5496
rect 5293 5484 5299 5516
rect 5277 5384 5283 5436
rect 4653 5124 4659 5216
rect 4669 5104 4675 5316
rect 4733 5264 4739 5316
rect 4749 5184 4755 5316
rect 4829 5144 4835 5156
rect 4685 5084 4691 5116
rect 4701 5044 4707 5096
rect 4717 5064 4723 5096
rect 4797 5064 4803 5076
rect 4525 4944 4531 4976
rect 4541 4944 4547 4956
rect 4301 4624 4307 4636
rect 4413 4624 4419 4696
rect 4429 4684 4435 4716
rect 4461 4684 4467 4696
rect 4269 4557 4291 4563
rect 4269 4524 4275 4557
rect 4221 4517 4243 4523
rect 4109 4504 4115 4516
rect 3844 4157 3859 4163
rect 3837 4124 3843 4156
rect 3885 4124 3891 4236
rect 3901 4164 3907 4236
rect 3965 4224 3971 4256
rect 3709 3924 3715 3976
rect 3805 3902 3811 4036
rect 3613 3844 3619 3876
rect 3373 3764 3379 3836
rect 3421 3764 3427 3796
rect 3597 3764 3603 3816
rect 3677 3724 3683 3896
rect 3757 3784 3763 3796
rect 3085 3704 3091 3716
rect 3101 3664 3107 3716
rect 3117 3643 3123 3716
rect 3101 3637 3123 3643
rect 1869 3120 1875 3158
rect 2077 3120 2083 3158
rect 1917 3104 1923 3116
rect 925 3064 931 3096
rect 781 2944 787 2956
rect 749 2924 755 2936
rect 173 2564 179 2656
rect 381 2564 387 2636
rect 45 2444 51 2496
rect 13 2264 19 2336
rect 125 2324 131 2336
rect 93 2304 99 2316
rect 141 2304 147 2536
rect 221 2384 227 2396
rect 333 2364 339 2436
rect 189 2324 195 2356
rect 301 2344 307 2356
rect 221 2304 227 2316
rect 45 2264 51 2296
rect 13 2104 19 2156
rect 93 2124 99 2296
rect 189 2284 195 2296
rect 141 2163 147 2276
rect 141 2157 156 2163
rect 141 2124 147 2136
rect 189 2124 195 2276
rect 205 2264 211 2276
rect 221 2264 227 2296
rect 237 2144 243 2296
rect 269 2284 275 2296
rect 333 2284 339 2296
rect 45 1924 51 1976
rect 61 1884 67 2036
rect 141 1904 147 2116
rect 285 2104 291 2236
rect 317 2164 323 2276
rect 253 1904 259 1916
rect 61 1764 67 1856
rect 253 1764 259 1896
rect 301 1784 307 2116
rect 317 1824 323 2156
rect 349 2124 355 2476
rect 365 2324 371 2416
rect 397 2264 403 2836
rect 541 2704 547 2896
rect 653 2844 659 2896
rect 669 2724 675 2776
rect 685 2724 691 2916
rect 653 2704 659 2716
rect 813 2704 819 2796
rect 861 2783 867 2956
rect 852 2777 867 2783
rect 781 2683 787 2696
rect 781 2677 796 2683
rect 573 2664 579 2676
rect 541 2603 547 2656
rect 717 2644 723 2656
rect 541 2597 563 2603
rect 557 2564 563 2597
rect 461 2462 467 2500
rect 477 2324 483 2376
rect 381 2124 387 2236
rect 333 1984 339 2096
rect 349 2084 355 2096
rect 381 1944 387 2036
rect 381 1884 387 1936
rect 413 1884 419 2116
rect 61 1484 67 1756
rect 205 1524 211 1676
rect 237 1584 243 1696
rect 61 1364 67 1476
rect 189 1444 195 1476
rect 253 1444 259 1736
rect 269 1604 275 1716
rect 285 1684 291 1716
rect 285 1584 291 1676
rect 269 1484 275 1536
rect 29 1244 35 1296
rect 13 664 19 696
rect 29 644 35 1236
rect 61 1084 67 1356
rect 221 1344 227 1356
rect 109 744 115 1316
rect 205 1084 211 1116
rect 237 1104 243 1156
rect 269 1124 275 1136
rect 285 1123 291 1496
rect 301 1324 307 1756
rect 333 1724 339 1876
rect 413 1864 419 1876
rect 381 1844 387 1856
rect 365 1524 371 1836
rect 381 1784 387 1816
rect 381 1544 387 1636
rect 317 1484 323 1516
rect 397 1504 403 1776
rect 461 1763 467 2136
rect 477 1924 483 2296
rect 461 1757 483 1763
rect 413 1684 419 1716
rect 333 1484 339 1496
rect 365 1464 371 1496
rect 381 1444 387 1476
rect 397 1464 403 1476
rect 413 1424 419 1676
rect 349 1337 364 1343
rect 317 1244 323 1296
rect 285 1117 300 1123
rect 301 1104 307 1116
rect 253 1064 259 1076
rect 205 984 211 1036
rect 45 444 51 496
rect 61 304 67 696
rect 77 524 83 736
rect 93 624 99 636
rect 125 604 131 936
rect 141 904 147 918
rect 205 744 211 896
rect 141 644 147 696
rect 157 624 163 676
rect 173 664 179 716
rect 221 684 227 936
rect 237 924 243 956
rect 269 944 275 1056
rect 237 704 243 836
rect 269 724 275 936
rect 317 904 323 976
rect 333 944 339 1316
rect 349 1184 355 1337
rect 381 1104 387 1416
rect 429 1303 435 1696
rect 461 1663 467 1757
rect 477 1744 483 1757
rect 445 1657 467 1663
rect 445 1324 451 1657
rect 461 1524 467 1636
rect 493 1523 499 1856
rect 509 1764 515 2436
rect 525 2404 531 2536
rect 781 2524 787 2677
rect 813 2584 819 2656
rect 829 2544 835 2676
rect 845 2524 851 2736
rect 877 2524 883 2676
rect 893 2564 899 2836
rect 925 2744 931 3056
rect 957 2904 963 3096
rect 973 3084 979 3096
rect 1037 3084 1043 3096
rect 1293 3084 1299 3096
rect 1565 3084 1571 3096
rect 973 2804 979 3076
rect 1229 2984 1235 3016
rect 1261 2964 1267 3056
rect 1437 3024 1443 3056
rect 1005 2924 1011 2936
rect 925 2704 931 2716
rect 1005 2684 1011 2916
rect 1069 2864 1075 2916
rect 1117 2904 1123 2916
rect 1133 2864 1139 2916
rect 1133 2724 1139 2776
rect 1149 2704 1155 2836
rect 1037 2684 1043 2696
rect 1133 2684 1139 2696
rect 1213 2684 1219 2916
rect 1229 2764 1235 2836
rect 1261 2784 1267 2956
rect 1549 2944 1555 3036
rect 1565 2924 1571 3076
rect 1581 3024 1587 3096
rect 1613 2964 1619 3036
rect 1693 2984 1699 3036
rect 1773 2964 1779 3056
rect 1805 3044 1811 3076
rect 1869 2964 1875 3036
rect 1485 2844 1491 2900
rect 1517 2884 1523 2916
rect 1229 2704 1235 2736
rect 909 2584 915 2656
rect 1005 2564 1011 2656
rect 1197 2604 1203 2636
rect 1149 2544 1155 2596
rect 1245 2524 1251 2676
rect 1261 2564 1267 2636
rect 1309 2564 1315 2756
rect 1309 2524 1315 2536
rect 685 2304 691 2516
rect 1213 2462 1219 2500
rect 717 2424 723 2436
rect 781 2344 787 2416
rect 685 2264 691 2296
rect 829 2284 835 2296
rect 557 2144 563 2216
rect 605 2204 611 2256
rect 845 2224 851 2276
rect 669 2184 675 2196
rect 637 1764 643 1876
rect 653 1824 659 1876
rect 669 1824 675 1896
rect 685 1884 691 2116
rect 701 1924 707 1956
rect 717 1944 723 2116
rect 765 2084 771 2116
rect 781 2024 787 2116
rect 829 1984 835 2116
rect 733 1904 739 1936
rect 781 1904 787 1916
rect 717 1884 723 1896
rect 685 1744 691 1876
rect 781 1804 787 1896
rect 797 1864 803 1896
rect 829 1824 835 1836
rect 653 1704 659 1718
rect 477 1517 499 1523
rect 477 1504 483 1517
rect 509 1504 515 1516
rect 557 1504 563 1536
rect 573 1504 579 1596
rect 685 1564 691 1736
rect 733 1724 739 1776
rect 829 1764 835 1816
rect 765 1744 771 1756
rect 813 1744 819 1756
rect 845 1744 851 2016
rect 861 1984 867 2436
rect 1245 2324 1251 2336
rect 989 2304 995 2316
rect 1156 2297 1171 2303
rect 877 1963 883 2236
rect 957 2184 963 2236
rect 1069 2184 1075 2276
rect 1165 2184 1171 2297
rect 925 2164 931 2176
rect 1229 2164 1235 2236
rect 925 2126 931 2136
rect 989 1984 995 2136
rect 1005 2124 1011 2156
rect 1053 2084 1059 2096
rect 861 1957 883 1963
rect 861 1904 867 1957
rect 941 1904 947 1916
rect 781 1664 787 1716
rect 637 1524 643 1536
rect 493 1497 508 1503
rect 461 1484 467 1496
rect 461 1404 467 1476
rect 477 1324 483 1496
rect 493 1324 499 1497
rect 541 1464 547 1476
rect 589 1343 595 1476
rect 580 1337 595 1343
rect 605 1323 611 1496
rect 596 1317 611 1323
rect 429 1297 451 1303
rect 349 924 355 936
rect 381 824 387 1096
rect 397 1044 403 1096
rect 397 924 403 1016
rect 413 924 419 1236
rect 429 1184 435 1276
rect 445 1044 451 1297
rect 461 1104 467 1236
rect 477 1104 483 1316
rect 541 1264 547 1316
rect 509 1164 515 1236
rect 541 1144 547 1256
rect 509 1104 515 1116
rect 541 1104 547 1116
rect 573 1104 579 1296
rect 589 1124 595 1316
rect 621 1244 627 1296
rect 637 1104 643 1496
rect 685 1484 691 1496
rect 733 1484 739 1556
rect 781 1524 787 1656
rect 701 1463 707 1476
rect 685 1457 707 1463
rect 685 1444 691 1457
rect 685 1364 691 1436
rect 685 1344 691 1356
rect 669 1284 675 1316
rect 685 1104 691 1236
rect 717 1103 723 1416
rect 765 1344 771 1456
rect 781 1104 787 1376
rect 813 1364 819 1736
rect 829 1724 835 1736
rect 845 1583 851 1736
rect 829 1577 851 1583
rect 829 1424 835 1577
rect 861 1384 867 1896
rect 877 1704 883 1776
rect 909 1724 915 1756
rect 925 1744 931 1876
rect 1021 1784 1027 1896
rect 1053 1863 1059 2076
rect 1117 1984 1123 2136
rect 1165 1984 1171 2116
rect 1181 2104 1187 2156
rect 1213 2104 1219 2116
rect 1069 1884 1075 1976
rect 1149 1904 1155 1936
rect 1053 1857 1075 1863
rect 1037 1837 1052 1843
rect 1037 1784 1043 1837
rect 941 1764 947 1776
rect 1037 1724 1043 1776
rect 1069 1764 1075 1857
rect 1133 1844 1139 1896
rect 1101 1744 1107 1796
rect 1053 1724 1059 1736
rect 1133 1724 1139 1836
rect 1149 1764 1155 1776
rect 1181 1764 1187 2096
rect 1213 1904 1219 1916
rect 1197 1763 1203 1896
rect 1213 1784 1219 1836
rect 1229 1784 1235 1916
rect 1245 1884 1251 2136
rect 1261 1904 1267 2116
rect 1277 1904 1283 2316
rect 1293 2304 1299 2436
rect 1357 2284 1363 2436
rect 1325 2117 1340 2123
rect 1293 2083 1299 2096
rect 1293 2077 1308 2083
rect 1309 1904 1315 2076
rect 1325 1984 1331 2117
rect 1357 1984 1363 2136
rect 1293 1764 1299 1896
rect 1325 1784 1331 1876
rect 1188 1757 1203 1763
rect 1293 1744 1299 1756
rect 941 1544 947 1556
rect 925 1423 931 1496
rect 909 1417 931 1423
rect 893 1344 899 1356
rect 877 1224 883 1236
rect 829 1104 835 1116
rect 708 1097 723 1103
rect 477 944 483 1076
rect 605 1064 611 1076
rect 605 984 611 1056
rect 397 904 403 916
rect 413 764 419 916
rect 285 704 291 736
rect 301 704 307 756
rect 381 724 387 736
rect 141 544 147 616
rect 237 604 243 696
rect 317 684 323 716
rect 365 684 371 716
rect 461 704 467 916
rect 493 702 499 716
rect 557 704 563 936
rect 589 924 595 956
rect 637 944 643 1096
rect 621 744 627 836
rect 637 744 643 936
rect 669 884 675 896
rect 685 884 691 896
rect 653 784 659 876
rect 669 723 675 876
rect 701 724 707 1096
rect 717 924 723 956
rect 733 944 739 976
rect 765 904 771 916
rect 669 717 684 723
rect 429 664 435 676
rect 173 564 179 596
rect 333 584 339 656
rect 77 303 83 516
rect 173 384 179 556
rect 349 524 355 636
rect 365 624 371 656
rect 365 544 371 616
rect 445 584 451 636
rect 461 544 467 676
rect 493 584 499 656
rect 493 564 499 576
rect 93 324 99 376
rect 77 297 92 303
rect 13 284 19 296
rect 45 124 51 296
rect 77 124 83 297
rect 221 264 227 376
rect 221 204 227 256
rect 301 224 307 296
rect 173 164 179 196
rect 349 124 355 516
rect 365 184 371 536
rect 397 497 412 503
rect 381 404 387 436
rect 397 383 403 497
rect 388 377 403 383
rect 413 324 419 396
rect 365 144 371 176
rect 429 163 435 476
rect 525 304 531 696
rect 637 664 643 676
rect 701 664 707 676
rect 605 544 611 556
rect 637 524 643 596
rect 685 524 691 636
rect 717 524 723 676
rect 733 584 739 856
rect 781 824 787 1096
rect 845 1084 851 1216
rect 877 1124 883 1156
rect 797 984 803 1036
rect 893 1024 899 1116
rect 909 1104 915 1417
rect 941 1343 947 1536
rect 973 1484 979 1716
rect 989 1664 995 1716
rect 1213 1704 1219 1716
rect 1037 1524 1043 1576
rect 1069 1564 1075 1656
rect 1069 1544 1075 1556
rect 989 1464 995 1496
rect 1101 1484 1107 1676
rect 1117 1564 1123 1636
rect 1117 1484 1123 1496
rect 925 1337 947 1343
rect 925 1144 931 1337
rect 989 1324 995 1456
rect 1005 1324 1011 1336
rect 941 1297 956 1303
rect 941 1184 947 1297
rect 989 1224 995 1316
rect 1069 1304 1075 1318
rect 1037 1184 1043 1216
rect 932 1137 947 1143
rect 804 977 819 983
rect 749 684 755 716
rect 749 544 755 616
rect 765 524 771 536
rect 781 524 787 736
rect 797 664 803 696
rect 813 684 819 977
rect 909 963 915 1096
rect 909 957 924 963
rect 829 724 835 936
rect 845 864 851 896
rect 829 704 835 716
rect 829 544 835 696
rect 845 604 851 696
rect 861 524 867 536
rect 877 524 883 836
rect 893 624 899 936
rect 925 924 931 956
rect 941 904 947 1137
rect 957 1124 963 1136
rect 1069 1124 1075 1136
rect 996 1117 1011 1123
rect 1005 1104 1011 1117
rect 1101 1104 1107 1316
rect 1133 1304 1139 1696
rect 1165 1564 1171 1636
rect 1149 1524 1155 1556
rect 1197 1523 1203 1636
rect 1341 1564 1347 1856
rect 1373 1764 1379 2076
rect 1389 1904 1395 2276
rect 1437 2264 1443 2836
rect 1496 2806 1502 2814
rect 1510 2806 1516 2814
rect 1524 2806 1530 2814
rect 1538 2806 1544 2814
rect 1645 2784 1651 2916
rect 1645 2704 1651 2716
rect 1533 2524 1539 2696
rect 1629 2684 1635 2696
rect 1661 2604 1667 2916
rect 1757 2884 1763 2916
rect 1693 2624 1699 2716
rect 1725 2584 1731 2676
rect 1741 2664 1747 2756
rect 1757 2704 1763 2876
rect 1773 2844 1779 2900
rect 1869 2824 1875 2956
rect 1789 2724 1795 2776
rect 1757 2523 1763 2696
rect 1917 2664 1923 2816
rect 1949 2804 1955 3116
rect 1965 2904 1971 3036
rect 1981 3004 1987 3116
rect 2045 3104 2051 3116
rect 2141 3064 2147 3076
rect 2173 3064 2179 3216
rect 2365 3184 2371 3456
rect 2381 3364 2387 3416
rect 2509 3404 2515 3456
rect 2573 3364 2579 3396
rect 2477 3262 2483 3300
rect 2541 3264 2547 3316
rect 2397 3124 2403 3236
rect 2381 3084 2387 3096
rect 2077 2984 2083 3056
rect 2173 3044 2179 3056
rect 2349 2964 2355 3036
rect 2045 2923 2051 2936
rect 2045 2917 2124 2923
rect 1997 2704 2003 2916
rect 2429 2904 2435 3116
rect 2477 3104 2483 3116
rect 2125 2704 2131 2736
rect 1885 2624 1891 2656
rect 1917 2644 1923 2656
rect 1748 2517 1763 2523
rect 1709 2462 1715 2500
rect 1496 2406 1502 2414
rect 1510 2406 1516 2414
rect 1524 2406 1530 2414
rect 1538 2406 1544 2414
rect 1565 2320 1571 2358
rect 1629 2284 1635 2416
rect 1741 2304 1747 2516
rect 1789 2444 1795 2536
rect 1821 2424 1827 2496
rect 1853 2284 1859 2596
rect 1869 2524 1875 2616
rect 1885 2544 1891 2616
rect 1933 2544 1939 2596
rect 1869 2384 1875 2416
rect 1933 2384 1939 2536
rect 1997 2524 2003 2696
rect 2109 2564 2115 2636
rect 2141 2624 2147 2896
rect 2173 2744 2179 2896
rect 2221 2844 2227 2896
rect 2285 2784 2291 2816
rect 2173 2624 2179 2716
rect 2301 2684 2307 2776
rect 2349 2724 2355 2776
rect 2253 2524 2259 2636
rect 2013 2444 2019 2500
rect 2205 2384 2211 2416
rect 2269 2384 2275 2436
rect 1917 2324 1923 2376
rect 1853 2264 1859 2276
rect 1437 2144 1443 2256
rect 1661 2184 1667 2256
rect 2013 2224 2019 2276
rect 1501 2164 1507 2176
rect 1485 2104 1491 2116
rect 1453 1984 1459 2076
rect 1496 2006 1502 2014
rect 1510 2006 1516 2014
rect 1524 2006 1530 2014
rect 1538 2006 1544 2014
rect 1581 1984 1587 2156
rect 1981 2144 1987 2176
rect 2045 2164 2051 2256
rect 1645 1984 1651 2116
rect 1661 2084 1667 2136
rect 1389 1804 1395 1896
rect 1597 1864 1603 1896
rect 1613 1884 1619 1976
rect 1709 1884 1715 1896
rect 1725 1884 1731 1896
rect 1453 1764 1459 1836
rect 1469 1764 1475 1856
rect 1565 1724 1571 1836
rect 1357 1684 1363 1716
rect 1373 1584 1379 1696
rect 1677 1684 1683 1756
rect 1197 1517 1219 1523
rect 1197 1464 1203 1496
rect 1213 1484 1219 1517
rect 1229 1484 1235 1556
rect 1261 1517 1276 1523
rect 1245 1484 1251 1496
rect 1229 1384 1235 1456
rect 1133 1164 1139 1296
rect 1213 1264 1219 1336
rect 1245 1324 1251 1476
rect 1261 1464 1267 1517
rect 1293 1503 1299 1536
rect 1293 1497 1308 1503
rect 1341 1464 1347 1516
rect 1373 1484 1379 1496
rect 1357 1444 1363 1476
rect 1261 1244 1267 1356
rect 1293 1344 1299 1396
rect 1389 1383 1395 1636
rect 1405 1604 1411 1636
rect 1405 1564 1411 1596
rect 1405 1464 1411 1516
rect 1421 1484 1427 1656
rect 1496 1606 1502 1614
rect 1510 1606 1516 1614
rect 1524 1606 1530 1614
rect 1538 1606 1544 1614
rect 1389 1377 1411 1383
rect 1405 1344 1411 1377
rect 1421 1344 1427 1476
rect 1484 1464 1492 1470
rect 1437 1404 1443 1436
rect 1437 1297 1452 1303
rect 1325 1243 1331 1296
rect 1309 1237 1331 1243
rect 1133 1084 1139 1116
rect 1181 1104 1187 1156
rect 1197 1124 1203 1136
rect 1213 1104 1219 1116
rect 1220 1097 1235 1103
rect 989 1077 1004 1083
rect 973 984 979 1076
rect 909 844 915 896
rect 941 884 947 896
rect 909 684 915 696
rect 925 684 931 696
rect 452 297 467 303
rect 420 157 435 163
rect 413 104 419 156
rect 461 124 467 297
rect 621 284 627 336
rect 653 304 659 436
rect 685 383 691 516
rect 685 377 707 383
rect 701 324 707 377
rect 45 44 51 96
rect 493 -17 499 256
rect 509 184 515 276
rect 477 -23 499 -17
rect 509 -23 515 156
rect 541 144 547 196
rect 573 126 579 236
rect 701 184 707 316
rect 765 302 771 316
rect 765 204 771 256
rect 781 144 787 156
rect 797 124 803 436
rect 829 284 835 336
rect 829 164 835 276
rect 861 244 867 516
rect 877 504 883 516
rect 909 464 915 676
rect 925 664 931 676
rect 973 584 979 936
rect 989 903 995 1077
rect 1085 1064 1091 1076
rect 1149 984 1155 1076
rect 1213 984 1219 1076
rect 989 897 1011 903
rect 989 704 995 816
rect 1005 784 1011 897
rect 1021 863 1027 936
rect 1053 924 1059 956
rect 1101 904 1107 916
rect 1037 884 1043 896
rect 1069 884 1075 896
rect 1149 884 1155 896
rect 1021 857 1043 863
rect 1037 784 1043 857
rect 1069 784 1075 856
rect 1229 824 1235 1097
rect 1277 1084 1283 1116
rect 1245 884 1251 936
rect 1261 843 1267 916
rect 1245 837 1267 843
rect 1197 704 1203 736
rect 989 644 995 656
rect 1005 584 1011 676
rect 1053 584 1059 656
rect 1085 644 1091 656
rect 925 524 931 576
rect 957 544 963 556
rect 1117 544 1123 556
rect 1197 524 1203 556
rect 1213 524 1219 716
rect 1245 524 1251 837
rect 1277 784 1283 936
rect 1293 924 1299 1036
rect 1309 904 1315 1237
rect 1341 1184 1347 1296
rect 1389 1284 1395 1296
rect 1357 1144 1363 1256
rect 1421 1143 1427 1236
rect 1405 1137 1427 1143
rect 1357 1124 1363 1136
rect 1325 1084 1331 1116
rect 1405 1104 1411 1137
rect 1325 964 1331 1076
rect 1373 1004 1379 1076
rect 1405 984 1411 1076
rect 1437 984 1443 1297
rect 1501 1244 1507 1336
rect 1549 1284 1555 1476
rect 1613 1384 1619 1616
rect 1709 1604 1715 1736
rect 1773 1684 1779 1856
rect 1789 1764 1795 2036
rect 2029 1924 2035 1976
rect 1821 1724 1827 1896
rect 1853 1724 1859 1736
rect 1901 1724 1907 1816
rect 1949 1744 1955 1756
rect 1677 1520 1683 1558
rect 1773 1464 1779 1676
rect 1805 1644 1811 1696
rect 1773 1424 1779 1456
rect 1565 1344 1571 1376
rect 1805 1364 1811 1416
rect 1853 1404 1859 1496
rect 1901 1364 1907 1716
rect 1917 1624 1923 1696
rect 1933 1584 1939 1736
rect 1997 1704 2003 1916
rect 2045 1904 2051 2116
rect 2077 2044 2083 2096
rect 2093 1984 2099 2216
rect 2125 2124 2131 2296
rect 2301 2284 2307 2676
rect 2365 2544 2371 2836
rect 2477 2664 2483 2956
rect 2493 2824 2499 3096
rect 2541 3084 2547 3256
rect 2589 3184 2595 3236
rect 2685 3184 2691 3336
rect 2701 3144 2707 3496
rect 2717 3404 2723 3496
rect 2733 3464 2739 3476
rect 2813 3464 2819 3576
rect 2861 3504 2867 3636
rect 2925 3520 2931 3558
rect 2893 3504 2899 3516
rect 3101 3504 3107 3637
rect 3213 3504 3219 3696
rect 3021 3464 3027 3496
rect 2829 3364 2835 3456
rect 3032 3406 3038 3414
rect 3046 3406 3052 3414
rect 3060 3406 3066 3414
rect 3074 3406 3080 3414
rect 2813 3284 2819 3296
rect 2877 3284 2883 3316
rect 2909 3304 2915 3316
rect 2573 3104 2579 3116
rect 2653 3104 2659 3136
rect 2724 3117 2739 3123
rect 2548 3077 2563 3083
rect 2557 2924 2563 3077
rect 2637 3024 2643 3036
rect 2637 2924 2643 3016
rect 2557 2704 2563 2916
rect 2653 2703 2659 2916
rect 2669 2864 2675 3096
rect 2733 3084 2739 3117
rect 2765 3103 2771 3236
rect 2797 3104 2803 3236
rect 2893 3144 2899 3236
rect 2925 3104 2931 3376
rect 2941 3284 2947 3396
rect 3053 3324 3059 3336
rect 3165 3324 3171 3336
rect 2973 3304 2979 3316
rect 3053 3304 3059 3316
rect 2756 3097 2771 3103
rect 2669 2824 2675 2856
rect 2685 2704 2691 3076
rect 2781 3024 2787 3096
rect 2797 2924 2803 2936
rect 2909 2924 2915 3056
rect 2941 2984 2947 3076
rect 2701 2844 2707 2896
rect 2765 2704 2771 2816
rect 2797 2724 2803 2796
rect 2861 2717 2876 2723
rect 2781 2704 2787 2716
rect 2861 2704 2867 2717
rect 2653 2697 2668 2703
rect 2397 2524 2403 2536
rect 2429 2524 2435 2576
rect 2477 2564 2483 2656
rect 2669 2644 2675 2696
rect 2701 2664 2707 2676
rect 2669 2584 2675 2636
rect 2701 2544 2707 2576
rect 2589 2484 2595 2516
rect 2445 2444 2451 2476
rect 2349 2324 2355 2376
rect 2445 2304 2451 2436
rect 2669 2304 2675 2316
rect 2765 2304 2771 2696
rect 2845 2664 2851 2676
rect 2781 2404 2787 2656
rect 2797 2444 2803 2496
rect 2813 2423 2819 2636
rect 2877 2564 2883 2696
rect 2845 2544 2851 2556
rect 2797 2417 2819 2423
rect 2845 2517 2860 2523
rect 2797 2324 2803 2417
rect 2845 2303 2851 2517
rect 2861 2384 2867 2496
rect 2893 2324 2899 2796
rect 2909 2724 2915 2876
rect 2925 2683 2931 2896
rect 2941 2784 2947 2936
rect 2957 2744 2963 3236
rect 2973 2704 2979 3096
rect 3021 3043 3027 3236
rect 3149 3224 3155 3316
rect 3197 3304 3203 3416
rect 3213 3344 3219 3436
rect 3245 3424 3251 3496
rect 3261 3444 3267 3716
rect 3309 3704 3315 3716
rect 3277 3464 3283 3496
rect 3293 3464 3299 3476
rect 3325 3384 3331 3716
rect 3421 3524 3427 3576
rect 3437 3504 3443 3716
rect 3501 3662 3507 3700
rect 3373 3464 3379 3476
rect 3517 3464 3523 3476
rect 3261 3344 3267 3356
rect 3213 3264 3219 3336
rect 3277 3284 3283 3336
rect 3293 3324 3299 3336
rect 3245 3120 3251 3158
rect 3341 3144 3347 3336
rect 3069 3064 3075 3096
rect 3149 3044 3155 3056
rect 3181 3044 3187 3076
rect 3005 3037 3027 3043
rect 2909 2677 2931 2683
rect 2909 2584 2915 2677
rect 2909 2544 2915 2576
rect 2925 2523 2931 2656
rect 2957 2644 2963 2696
rect 2957 2524 2963 2576
rect 2989 2544 2995 2736
rect 3005 2684 3011 3037
rect 3032 3006 3038 3014
rect 3046 3006 3052 3014
rect 3060 3006 3066 3014
rect 3074 3006 3080 3014
rect 3165 2944 3171 2976
rect 3021 2704 3027 2736
rect 3005 2584 3011 2656
rect 3032 2606 3038 2614
rect 3046 2606 3052 2614
rect 3060 2606 3066 2614
rect 3074 2606 3080 2614
rect 3101 2577 3116 2583
rect 3085 2544 3091 2556
rect 3101 2544 3107 2577
rect 3133 2564 3139 2856
rect 3197 2844 3203 2896
rect 3149 2683 3155 2836
rect 3245 2783 3251 3056
rect 3357 2984 3363 3416
rect 3373 3244 3379 3276
rect 3373 3124 3379 3236
rect 3405 3224 3411 3256
rect 3293 2924 3299 2936
rect 3261 2804 3267 2896
rect 3293 2864 3299 2916
rect 3325 2904 3331 2976
rect 3341 2904 3347 2936
rect 3341 2864 3347 2896
rect 3229 2777 3251 2783
rect 3165 2720 3171 2758
rect 3229 2704 3235 2777
rect 3149 2677 3171 2683
rect 2973 2524 2979 2536
rect 2909 2517 2931 2523
rect 2836 2297 2851 2303
rect 2157 2044 2163 2096
rect 2173 1944 2179 2236
rect 2445 2184 2451 2236
rect 2477 2184 2483 2256
rect 2493 2184 2499 2216
rect 2285 2164 2291 2176
rect 2077 1904 2083 1916
rect 2125 1864 2131 1876
rect 2045 1724 2051 1836
rect 2061 1744 2067 1856
rect 2141 1844 2147 1896
rect 2189 1804 2195 1896
rect 2253 1824 2259 1836
rect 2045 1504 2051 1716
rect 2077 1504 2083 1796
rect 2285 1784 2291 2156
rect 2301 1884 2307 2036
rect 2365 1944 2371 2036
rect 2333 1844 2339 1896
rect 2397 1844 2403 1896
rect 2253 1764 2259 1776
rect 1581 1324 1587 1356
rect 1533 1244 1539 1276
rect 1469 1103 1475 1236
rect 1496 1206 1502 1214
rect 1510 1206 1516 1214
rect 1524 1206 1530 1214
rect 1538 1206 1544 1214
rect 1565 1184 1571 1316
rect 1613 1284 1619 1296
rect 1469 1097 1491 1103
rect 1453 1044 1459 1096
rect 1341 937 1356 943
rect 1325 884 1331 916
rect 1341 843 1347 937
rect 1357 884 1363 916
rect 1405 884 1411 896
rect 1325 837 1347 843
rect 1309 764 1315 836
rect 1325 784 1331 837
rect 1293 524 1299 656
rect 845 237 860 243
rect 845 104 851 237
rect 877 124 883 456
rect 893 324 899 356
rect 909 304 915 436
rect 925 324 931 516
rect 1005 284 1011 436
rect 1133 384 1139 516
rect 1245 504 1251 516
rect 1133 364 1139 376
rect 1021 304 1027 316
rect 1149 284 1155 336
rect 1181 303 1187 436
rect 1213 324 1219 356
rect 1261 304 1267 436
rect 1172 297 1187 303
rect 1277 284 1283 336
rect 1293 324 1299 516
rect 1309 364 1315 656
rect 1357 524 1363 876
rect 1373 504 1379 636
rect 1389 524 1395 816
rect 1437 723 1443 856
rect 1453 744 1459 936
rect 1485 884 1491 1097
rect 1501 924 1507 1116
rect 1533 1104 1539 1116
rect 1581 1104 1587 1236
rect 1645 1124 1651 1236
rect 1805 1204 1811 1356
rect 1933 1324 1939 1396
rect 1965 1344 1971 1436
rect 1981 1384 1987 1476
rect 2029 1324 2035 1336
rect 2077 1324 2083 1356
rect 2093 1324 2099 1496
rect 2125 1464 2131 1756
rect 2253 1684 2259 1756
rect 2461 1744 2467 2156
rect 2557 2124 2563 2296
rect 2829 2264 2835 2296
rect 2909 2283 2915 2517
rect 2925 2444 2931 2496
rect 3005 2324 3011 2456
rect 3021 2364 3027 2496
rect 3037 2324 3043 2536
rect 2957 2317 2972 2323
rect 2957 2304 2963 2317
rect 3021 2284 3027 2316
rect 3053 2284 3059 2316
rect 2893 2277 2915 2283
rect 2749 2124 2755 2156
rect 2797 2144 2803 2236
rect 2845 2164 2851 2276
rect 2861 2257 2876 2263
rect 2573 2044 2579 2100
rect 2589 1924 2595 1976
rect 2493 1884 2499 1896
rect 2285 1724 2291 1736
rect 2493 1724 2499 1876
rect 2541 1824 2547 1896
rect 2717 1864 2723 1956
rect 2861 1944 2867 2257
rect 2877 2064 2883 2156
rect 2893 1924 2899 2277
rect 2957 2224 2963 2276
rect 3032 2206 3038 2214
rect 3046 2206 3052 2214
rect 3060 2206 3066 2214
rect 3074 2206 3080 2214
rect 3101 2184 3107 2436
rect 3133 2343 3139 2436
rect 3117 2337 3139 2343
rect 3117 2304 3123 2337
rect 3149 2323 3155 2496
rect 3165 2484 3171 2677
rect 3181 2504 3187 2576
rect 3261 2544 3267 2616
rect 3277 2544 3283 2556
rect 3341 2544 3347 2796
rect 3245 2504 3251 2516
rect 3165 2444 3171 2456
rect 3165 2343 3171 2436
rect 3197 2384 3203 2476
rect 3213 2444 3219 2496
rect 3293 2484 3299 2516
rect 3261 2384 3267 2436
rect 3165 2337 3187 2343
rect 3181 2324 3187 2337
rect 3149 2317 3164 2323
rect 3117 2224 3123 2276
rect 2909 1964 2915 2036
rect 2893 1784 2899 1916
rect 2349 1662 2355 1700
rect 2237 1544 2243 1556
rect 2317 1520 2323 1558
rect 2381 1504 2387 1716
rect 2461 1644 2467 1696
rect 2189 1464 2195 1476
rect 2381 1444 2387 1476
rect 2413 1464 2419 1596
rect 2493 1504 2499 1716
rect 2589 1604 2595 1756
rect 2909 1744 2915 1836
rect 2685 1524 2691 1576
rect 2781 1544 2787 1696
rect 2845 1604 2851 1636
rect 1709 1184 1715 1196
rect 1837 1143 1843 1316
rect 1901 1262 1907 1300
rect 1821 1137 1843 1143
rect 1496 806 1502 814
rect 1510 806 1516 814
rect 1524 806 1530 814
rect 1538 806 1544 814
rect 1437 717 1452 723
rect 1469 684 1475 696
rect 1444 557 1468 563
rect 1405 524 1411 556
rect 1341 444 1347 456
rect 1341 344 1347 436
rect 893 144 899 276
rect 909 184 915 236
rect 1005 204 1011 276
rect 1261 204 1267 276
rect 1005 144 1011 196
rect 1293 144 1299 256
rect 1309 184 1315 196
rect 1005 124 1011 136
rect 1021 124 1027 136
rect 1325 124 1331 236
rect 1341 184 1347 316
rect 1373 304 1379 496
rect 1453 484 1459 516
rect 1485 484 1491 736
rect 1501 704 1507 756
rect 1565 744 1571 1056
rect 1581 1044 1587 1076
rect 1581 784 1587 836
rect 1565 684 1571 736
rect 1453 384 1459 476
rect 1533 464 1539 536
rect 1549 524 1555 556
rect 1597 544 1603 1076
rect 1741 1044 1747 1096
rect 1805 1084 1811 1096
rect 1789 944 1795 1036
rect 1629 623 1635 656
rect 1613 617 1635 623
rect 1496 406 1502 414
rect 1510 406 1516 414
rect 1524 406 1530 414
rect 1538 406 1544 414
rect 1565 304 1571 516
rect 1597 484 1603 496
rect 1389 204 1395 276
rect 1469 264 1475 296
rect 1613 284 1619 617
rect 1629 524 1635 596
rect 1645 544 1651 676
rect 1693 544 1699 936
rect 1821 924 1827 1137
rect 1837 1064 1843 1096
rect 1869 1064 1875 1076
rect 1933 964 1939 1176
rect 1981 1164 1987 1296
rect 2029 1084 2035 1096
rect 2109 1084 2115 1436
rect 2493 1364 2499 1456
rect 2189 1324 2195 1336
rect 2189 1124 2195 1156
rect 2237 1144 2243 1196
rect 2269 1184 2275 1356
rect 2269 1144 2275 1176
rect 2141 1084 2147 1116
rect 1709 824 1715 918
rect 1837 862 1843 900
rect 1757 784 1763 856
rect 1869 784 1875 816
rect 1821 724 1827 776
rect 1821 704 1827 716
rect 1629 504 1635 516
rect 1629 244 1635 256
rect 1469 184 1475 236
rect 1341 124 1347 156
rect 1549 124 1555 216
rect 1645 204 1651 536
rect 1741 324 1747 616
rect 1789 604 1795 696
rect 1869 684 1875 696
rect 1885 684 1891 736
rect 1901 704 1907 796
rect 1997 724 2003 736
rect 1965 704 1971 716
rect 2013 704 2019 916
rect 2045 904 2051 1036
rect 2077 804 2083 1076
rect 2093 984 2099 1076
rect 2157 1044 2163 1096
rect 2173 1084 2179 1116
rect 2125 924 2131 1036
rect 2189 944 2195 1076
rect 2221 944 2227 1096
rect 2253 1084 2259 1096
rect 2269 1064 2275 1076
rect 2237 984 2243 1036
rect 2253 963 2259 1056
rect 2269 984 2275 1056
rect 2253 957 2268 963
rect 2269 944 2275 956
rect 2173 924 2179 936
rect 2221 904 2227 936
rect 2077 724 2083 776
rect 2029 684 2035 716
rect 1933 664 1939 676
rect 1965 564 1971 656
rect 2221 564 2227 576
rect 2285 563 2291 1216
rect 2381 1164 2387 1276
rect 2397 1244 2403 1296
rect 2381 1124 2387 1156
rect 2445 1104 2451 1316
rect 2477 1204 2483 1356
rect 2493 1344 2499 1356
rect 2525 1324 2531 1496
rect 2541 1324 2547 1356
rect 2621 1344 2627 1436
rect 2637 1344 2643 1476
rect 2573 1244 2579 1296
rect 2413 1064 2419 1096
rect 2317 943 2323 956
rect 2333 943 2339 1056
rect 2349 944 2355 1056
rect 2429 1044 2435 1076
rect 2381 944 2387 1036
rect 2477 984 2483 1036
rect 2397 944 2403 976
rect 2317 940 2339 943
rect 2324 937 2339 940
rect 2413 924 2419 936
rect 2445 904 2451 956
rect 2381 704 2387 716
rect 2461 684 2467 796
rect 2493 703 2499 1176
rect 2509 1164 2515 1236
rect 2573 1124 2579 1236
rect 2621 1184 2627 1316
rect 2653 1224 2659 1276
rect 2669 1204 2675 1496
rect 2605 1104 2611 1136
rect 2685 1104 2691 1158
rect 2573 1064 2579 1076
rect 2605 1064 2611 1096
rect 2605 1004 2611 1056
rect 2717 1024 2723 1536
rect 2813 1464 2819 1596
rect 2925 1564 2931 1856
rect 2941 1844 2947 1896
rect 2973 1744 2979 2136
rect 3005 1984 3011 2176
rect 3261 2164 3267 2236
rect 3181 2124 3187 2156
rect 3293 2144 3299 2436
rect 3341 2264 3347 2536
rect 3357 2504 3363 2816
rect 3373 2564 3379 3116
rect 3389 2764 3395 2956
rect 3405 2804 3411 3216
rect 3421 2864 3427 3116
rect 3453 2924 3459 3456
rect 3549 3423 3555 3456
rect 3533 3417 3555 3423
rect 3533 3384 3539 3417
rect 3533 3364 3539 3376
rect 3629 3324 3635 3496
rect 3485 2924 3491 2956
rect 3517 2944 3523 3096
rect 3581 3043 3587 3136
rect 3597 3104 3603 3176
rect 3645 3104 3651 3316
rect 3661 3244 3667 3296
rect 3565 3037 3587 3043
rect 3524 2937 3539 2943
rect 3469 2864 3475 2896
rect 3357 2344 3363 2496
rect 3373 2484 3379 2556
rect 3389 2544 3395 2556
rect 3389 2324 3395 2536
rect 3405 2384 3411 2676
rect 3421 2544 3427 2636
rect 3437 2523 3443 2676
rect 3428 2517 3443 2523
rect 3453 2503 3459 2736
rect 3469 2724 3475 2856
rect 3485 2704 3491 2716
rect 3517 2704 3523 2716
rect 3533 2704 3539 2937
rect 3549 2924 3555 2936
rect 3565 2884 3571 3037
rect 3597 2984 3603 3036
rect 3597 2904 3603 2916
rect 3549 2864 3555 2876
rect 3565 2744 3571 2876
rect 3597 2764 3603 2896
rect 3613 2723 3619 2776
rect 3604 2717 3619 2723
rect 3469 2544 3475 2656
rect 3501 2583 3507 2696
rect 3549 2684 3555 2696
rect 3629 2683 3635 2836
rect 3645 2824 3651 3096
rect 3677 2944 3683 3596
rect 3805 3484 3811 3516
rect 3821 3504 3827 3996
rect 3837 3984 3843 4116
rect 3949 4104 3955 4116
rect 3917 4084 3923 4096
rect 3965 4084 3971 4116
rect 3949 4064 3955 4076
rect 3981 4063 3987 4276
rect 3997 4104 4003 4196
rect 4013 4157 4051 4163
rect 4013 4144 4019 4157
rect 4045 4143 4051 4157
rect 4045 4137 4060 4143
rect 4029 4124 4035 4136
rect 4077 4124 4083 4216
rect 4093 4184 4099 4276
rect 4125 4164 4131 4336
rect 4141 4324 4147 4376
rect 4173 4343 4179 4496
rect 4205 4384 4211 4436
rect 4164 4337 4179 4343
rect 4221 4163 4227 4517
rect 4301 4504 4307 4536
rect 4205 4157 4227 4163
rect 4157 4124 4163 4156
rect 4173 4124 4179 4156
rect 4013 4104 4019 4116
rect 4029 4084 4035 4116
rect 4109 4104 4115 4116
rect 4205 4104 4211 4157
rect 4221 4124 4227 4136
rect 4237 4084 4243 4496
rect 4317 4464 4323 4516
rect 4349 4504 4355 4616
rect 4365 4484 4371 4536
rect 3965 4057 3987 4063
rect 3965 3984 3971 4057
rect 3997 3984 4003 4056
rect 3869 3824 3875 3896
rect 4253 3864 4259 4276
rect 4269 4204 4275 4436
rect 4285 4144 4291 4176
rect 4317 4123 4323 4436
rect 4349 4264 4355 4436
rect 4381 4303 4387 4516
rect 4461 4503 4467 4676
rect 4452 4497 4467 4503
rect 4477 4503 4483 4756
rect 4525 4684 4531 4916
rect 4541 4844 4547 4916
rect 4557 4904 4563 5016
rect 4573 4964 4579 5036
rect 4653 4963 4659 5036
rect 4637 4957 4659 4963
rect 4637 4904 4643 4957
rect 4765 4944 4771 4976
rect 4797 4944 4803 5056
rect 4477 4497 4492 4503
rect 4413 4444 4419 4496
rect 4509 4483 4515 4516
rect 4493 4477 4515 4483
rect 4445 4343 4451 4436
rect 4429 4337 4451 4343
rect 4429 4324 4435 4337
rect 4381 4297 4396 4303
rect 4381 4224 4387 4297
rect 4365 4124 4371 4156
rect 4308 4117 4323 4123
rect 4413 4104 4419 4156
rect 4429 4144 4435 4236
rect 4445 4124 4451 4176
rect 4493 4164 4499 4477
rect 4525 4364 4531 4476
rect 4541 4464 4547 4836
rect 4568 4806 4574 4814
rect 4582 4806 4588 4814
rect 4596 4806 4602 4814
rect 4610 4806 4616 4814
rect 4653 4724 4659 4936
rect 4669 4784 4675 4896
rect 4701 4884 4707 4896
rect 4669 4704 4675 4776
rect 4605 4644 4611 4696
rect 4653 4684 4659 4696
rect 4685 4684 4691 4736
rect 4717 4724 4723 4816
rect 4717 4664 4723 4716
rect 4733 4684 4739 4936
rect 4749 4904 4755 4916
rect 4605 4584 4611 4636
rect 4701 4563 4707 4636
rect 4685 4557 4707 4563
rect 4637 4464 4643 4516
rect 4685 4504 4691 4557
rect 4717 4524 4723 4616
rect 4749 4544 4755 4696
rect 4765 4564 4771 4936
rect 4781 4844 4787 4876
rect 4781 4824 4787 4836
rect 4813 4744 4819 5036
rect 4781 4724 4787 4736
rect 4845 4704 4851 5136
rect 4877 5104 4883 5276
rect 4893 5184 4899 5316
rect 4941 5284 4947 5296
rect 4909 5124 4915 5276
rect 4989 5184 4995 5296
rect 5197 5224 5203 5296
rect 5213 5204 5219 5236
rect 4909 5104 4915 5116
rect 4989 5104 4995 5176
rect 5037 5144 5043 5176
rect 5053 5104 5059 5136
rect 5165 5124 5171 5196
rect 5229 5144 5235 5316
rect 5309 5304 5315 5316
rect 5268 5117 5299 5123
rect 4861 4764 4867 5096
rect 4909 4964 4915 5016
rect 4893 4924 4899 4956
rect 4893 4784 4899 4896
rect 4941 4844 4947 5096
rect 5005 5064 5011 5076
rect 4957 4984 4963 5036
rect 5005 4944 5011 5056
rect 5037 4964 5043 5036
rect 5069 4984 5075 5036
rect 5085 5004 5091 5036
rect 5069 4944 5075 4976
rect 4973 4904 4979 4916
rect 4884 4757 4899 4763
rect 4861 4704 4867 4716
rect 4877 4704 4883 4756
rect 4813 4544 4819 4556
rect 4749 4504 4755 4516
rect 4568 4406 4574 4414
rect 4582 4406 4588 4414
rect 4596 4406 4602 4414
rect 4610 4406 4616 4414
rect 4509 4184 4515 4296
rect 4493 4144 4499 4156
rect 4525 4144 4531 4356
rect 4541 4304 4547 4376
rect 4573 4104 4579 4156
rect 4637 4124 4643 4456
rect 4653 4184 4659 4436
rect 4717 4384 4723 4496
rect 4701 4344 4707 4356
rect 4749 4344 4755 4496
rect 4765 4384 4771 4536
rect 4797 4524 4803 4536
rect 4829 4524 4835 4696
rect 4845 4564 4851 4696
rect 4861 4604 4867 4696
rect 4861 4544 4867 4556
rect 4893 4524 4899 4757
rect 4925 4524 4931 4836
rect 4941 4784 4947 4836
rect 4957 4704 4963 4816
rect 4973 4724 4979 4896
rect 4989 4884 4995 4916
rect 5005 4723 5011 4936
rect 5037 4884 5043 4916
rect 4989 4717 5011 4723
rect 4957 4664 4963 4696
rect 4989 4684 4995 4717
rect 5021 4704 5027 4876
rect 5069 4784 5075 4896
rect 5005 4684 5011 4696
rect 5021 4684 5027 4696
rect 4973 4544 4979 4636
rect 5053 4584 5059 4676
rect 5069 4584 5075 4656
rect 5085 4524 5091 4556
rect 4957 4444 4963 4516
rect 4749 4324 4755 4336
rect 4957 4304 4963 4436
rect 5021 4320 5027 4358
rect 4717 4164 4723 4296
rect 4813 4184 4819 4276
rect 4989 4164 4995 4196
rect 4269 4084 4275 4096
rect 4333 4084 4339 4096
rect 4653 4084 4659 4116
rect 4685 4063 4691 4096
rect 4733 4084 4739 4136
rect 4845 4104 4851 4136
rect 4660 4057 4691 4063
rect 4301 3984 4307 4036
rect 4381 3924 4387 3976
rect 4429 3924 4435 3976
rect 3949 3804 3955 3856
rect 3965 3764 3971 3816
rect 3981 3804 3987 3856
rect 4253 3844 4259 3856
rect 4045 3804 4051 3836
rect 4077 3724 4083 3776
rect 4061 3662 4067 3700
rect 3933 3504 3939 3536
rect 4093 3504 4099 3836
rect 4317 3744 4323 3816
rect 4381 3784 4387 3896
rect 4445 3864 4451 4036
rect 4568 4006 4574 4014
rect 4582 4006 4588 4014
rect 4596 4006 4602 4014
rect 4610 4006 4616 4014
rect 4621 3924 4627 3976
rect 4141 3684 4147 3716
rect 4205 3704 4211 3716
rect 4445 3704 4451 3856
rect 4509 3724 4515 3896
rect 4717 3884 4723 4036
rect 4845 4004 4851 4096
rect 4861 4084 4867 4096
rect 4893 3924 4899 4036
rect 4909 3984 4915 4156
rect 5021 4104 5027 4136
rect 5037 4004 5043 4496
rect 5053 4484 5059 4516
rect 5053 4364 5059 4476
rect 5085 4164 5091 4516
rect 5101 4464 5107 5096
rect 5117 5084 5123 5116
rect 5229 5104 5235 5116
rect 5293 5104 5299 5117
rect 5213 5084 5219 5096
rect 5165 4984 5171 5036
rect 5181 4944 5187 4996
rect 5213 4904 5219 5076
rect 5229 5064 5235 5096
rect 5277 5084 5283 5096
rect 5277 5023 5283 5076
rect 5293 5044 5299 5076
rect 5261 5017 5283 5023
rect 5117 4784 5123 4896
rect 5133 4884 5139 4896
rect 5165 4784 5171 4836
rect 5181 4704 5187 4736
rect 5149 4584 5155 4656
rect 5213 4604 5219 4696
rect 5229 4564 5235 4896
rect 5245 4784 5251 4836
rect 5261 4704 5267 5017
rect 5261 4684 5267 4696
rect 5277 4523 5283 4976
rect 5293 4924 5299 4956
rect 5309 4723 5315 5296
rect 5325 5024 5331 5416
rect 5341 5384 5347 5476
rect 5357 5464 5363 5643
rect 5853 5520 5859 5558
rect 5501 5504 5507 5516
rect 5389 5444 5395 5456
rect 5373 5344 5379 5436
rect 5453 5424 5459 5476
rect 5549 5464 5555 5476
rect 5389 5324 5395 5396
rect 5613 5364 5619 5456
rect 5869 5384 5875 5456
rect 5645 5344 5651 5356
rect 5357 5124 5363 5136
rect 5421 5124 5427 5156
rect 5437 5104 5443 5296
rect 5725 5244 5731 5316
rect 5741 5244 5747 5296
rect 5453 5164 5459 5236
rect 5460 5097 5475 5103
rect 5325 4964 5331 5016
rect 5373 5004 5379 5076
rect 5389 4944 5395 5036
rect 5437 5004 5443 5076
rect 5444 4997 5459 5003
rect 5453 4944 5459 4997
rect 5405 4844 5411 4916
rect 5453 4764 5459 4936
rect 5469 4924 5475 5097
rect 5613 5064 5619 5096
rect 5661 5003 5667 5076
rect 5661 4997 5676 5003
rect 5629 4924 5635 4956
rect 5677 4944 5683 4996
rect 5709 4904 5715 5036
rect 5757 4944 5763 5076
rect 5789 4984 5795 5116
rect 5741 4924 5747 4936
rect 5309 4717 5331 4723
rect 5293 4704 5299 4716
rect 5309 4524 5315 4536
rect 5325 4524 5331 4717
rect 5485 4684 5491 4696
rect 5357 4584 5363 4656
rect 5437 4584 5443 4636
rect 5277 4517 5292 4523
rect 5149 4504 5155 4516
rect 5165 4484 5171 4496
rect 5133 4464 5139 4476
rect 5197 4444 5203 4516
rect 5293 4384 5299 4436
rect 5357 4404 5363 4436
rect 5405 4324 5411 4376
rect 5421 4304 5427 4516
rect 5485 4404 5491 4676
rect 5517 4604 5523 4836
rect 5549 4704 5555 4736
rect 5549 4664 5555 4696
rect 5773 4684 5779 4696
rect 5789 4684 5795 4696
rect 5565 4664 5571 4676
rect 5629 4604 5635 4636
rect 5597 4544 5603 4576
rect 5453 4304 5459 4396
rect 5517 4304 5523 4396
rect 5597 4384 5603 4496
rect 5661 4424 5667 4676
rect 5693 4444 5699 4496
rect 5053 4124 5059 4136
rect 5133 4104 5139 4116
rect 5149 4104 5155 4136
rect 5165 4064 5171 4096
rect 5181 4084 5187 4096
rect 4525 3824 4531 3876
rect 4749 3864 4755 3876
rect 4749 3844 4755 3856
rect 4573 3724 4579 3776
rect 4653 3724 4659 3756
rect 4829 3744 4835 3896
rect 5069 3884 5075 3956
rect 5085 3904 5091 4016
rect 5101 3984 5107 3996
rect 5165 3884 5171 3936
rect 5197 3904 5203 4296
rect 5309 4224 5315 4276
rect 5261 4184 5267 4216
rect 5453 4204 5459 4296
rect 5469 4184 5475 4296
rect 5325 4124 5331 4136
rect 5453 4124 5459 4136
rect 5501 4103 5507 4156
rect 5517 4144 5523 4296
rect 5533 4144 5539 4236
rect 5549 4183 5555 4296
rect 5613 4284 5619 4296
rect 5549 4177 5571 4183
rect 5501 4097 5516 4103
rect 5293 3984 5299 4036
rect 5213 3924 5219 3976
rect 5485 3924 5491 4036
rect 5501 3904 5507 4097
rect 5517 3904 5523 3976
rect 4845 3824 4851 3836
rect 4845 3764 4851 3816
rect 5069 3764 5075 3876
rect 5117 3844 5123 3856
rect 5085 3784 5091 3816
rect 5149 3784 5155 3836
rect 5213 3824 5219 3896
rect 5341 3824 5347 3856
rect 5373 3764 5379 3816
rect 5421 3804 5427 3896
rect 5533 3844 5539 4136
rect 5549 4024 5555 4116
rect 5565 4084 5571 4177
rect 5581 4104 5587 4196
rect 5661 4184 5667 4216
rect 5693 4144 5699 4236
rect 5709 4144 5715 4276
rect 5693 4124 5699 4136
rect 5725 4123 5731 4536
rect 5757 4404 5763 4436
rect 5805 4424 5811 5316
rect 5741 4163 5747 4296
rect 5821 4284 5827 5316
rect 5837 5264 5843 5276
rect 5885 5244 5891 5496
rect 5837 5104 5843 5236
rect 5917 5064 5923 5556
rect 6061 5543 6067 5643
rect 6093 5604 6099 5643
rect 6061 5537 6083 5543
rect 5949 5404 5955 5456
rect 5965 5343 5971 5476
rect 5965 5337 5980 5343
rect 6029 5324 6035 5396
rect 6077 5364 6083 5537
rect 5981 5204 5987 5316
rect 5949 5084 5955 5196
rect 6013 5120 6019 5158
rect 6052 5097 6067 5103
rect 5917 5004 5923 5056
rect 5949 4964 5955 4996
rect 5949 4783 5955 4956
rect 5981 4924 5987 4936
rect 6061 4924 6067 5097
rect 6045 4862 6051 4900
rect 5949 4777 5971 4783
rect 5885 4664 5891 4696
rect 5965 4664 5971 4777
rect 5837 4524 5843 4656
rect 5965 4604 5971 4656
rect 5917 4564 5923 4596
rect 5837 4423 5843 4516
rect 5949 4504 5955 4536
rect 6013 4462 6019 4500
rect 6061 4424 6067 4916
rect 6093 4724 6099 4776
rect 5837 4417 5859 4423
rect 5853 4304 5859 4417
rect 5949 4324 5955 4376
rect 5821 4164 5827 4256
rect 5853 4224 5859 4276
rect 5741 4157 5763 4163
rect 5725 4117 5747 4123
rect 5741 4104 5747 4117
rect 5549 3884 5555 4016
rect 5581 3924 5587 3996
rect 5677 3984 5683 4076
rect 5565 3864 5571 3896
rect 4989 3744 4995 3756
rect 4781 3724 4787 3736
rect 4141 3544 4147 3676
rect 4381 3604 4387 3696
rect 4509 3584 4515 3716
rect 4749 3644 4755 3700
rect 4568 3606 4574 3614
rect 4582 3606 4588 3614
rect 4596 3606 4602 3614
rect 4610 3606 4616 3614
rect 4445 3524 4451 3576
rect 3741 3464 3747 3476
rect 3709 3304 3715 3436
rect 3789 3384 3795 3456
rect 3805 3364 3811 3436
rect 3709 3124 3715 3156
rect 3725 3144 3731 3296
rect 3757 3203 3763 3336
rect 3773 3244 3779 3336
rect 3789 3284 3795 3316
rect 3741 3197 3763 3203
rect 3693 2984 3699 3076
rect 3709 2924 3715 3096
rect 3741 2944 3747 3197
rect 3757 3144 3763 3176
rect 3821 3104 3827 3396
rect 3837 3224 3843 3336
rect 3917 3304 3923 3336
rect 3981 3324 3987 3496
rect 3997 3284 4003 3496
rect 4013 3344 4019 3456
rect 4029 3404 4035 3436
rect 3981 3204 3987 3236
rect 3629 2677 3651 2683
rect 3533 2624 3539 2676
rect 3629 2604 3635 2656
rect 3501 2577 3523 2583
rect 3444 2497 3459 2503
rect 3437 2484 3443 2496
rect 3453 2444 3459 2476
rect 3421 2363 3427 2436
rect 3405 2357 3427 2363
rect 3405 2324 3411 2357
rect 3469 2324 3475 2456
rect 3517 2384 3523 2577
rect 3645 2544 3651 2677
rect 3661 2663 3667 2916
rect 3693 2844 3699 2896
rect 3725 2884 3731 2936
rect 3741 2904 3747 2936
rect 3757 2863 3763 3096
rect 3773 2884 3779 2976
rect 3821 2884 3827 3096
rect 3837 3084 3843 3096
rect 3869 2984 3875 3116
rect 3885 3104 3891 3156
rect 3885 2984 3891 3096
rect 3901 3024 3907 3076
rect 3757 2857 3779 2863
rect 3725 2744 3731 2756
rect 3773 2724 3779 2857
rect 3789 2744 3795 2816
rect 3805 2784 3811 2876
rect 3853 2864 3859 2916
rect 3821 2744 3827 2836
rect 3837 2784 3843 2836
rect 3853 2744 3859 2816
rect 3757 2704 3763 2716
rect 3773 2704 3779 2716
rect 3821 2704 3827 2716
rect 3677 2684 3683 2696
rect 3725 2684 3731 2696
rect 3661 2657 3683 2663
rect 3661 2624 3667 2636
rect 3677 2624 3683 2657
rect 3677 2564 3683 2596
rect 3757 2564 3763 2696
rect 3773 2644 3779 2696
rect 3869 2664 3875 2936
rect 3901 2864 3907 2936
rect 3917 2924 3923 3096
rect 3949 3064 3955 3096
rect 3965 3084 3971 3116
rect 3981 3084 3987 3096
rect 3933 2944 3939 3036
rect 3965 2984 3971 3056
rect 3997 2984 4003 3176
rect 4013 3124 4019 3336
rect 4045 3184 4051 3476
rect 4109 3424 4115 3436
rect 4141 3384 4147 3416
rect 4141 3364 4147 3376
rect 4029 3104 4035 3156
rect 4045 3084 4051 3096
rect 4029 3064 4035 3076
rect 3997 2964 4003 2976
rect 3917 2763 3923 2916
rect 3901 2757 3923 2763
rect 3901 2704 3907 2757
rect 3924 2737 3939 2743
rect 3869 2584 3875 2616
rect 3373 2224 3379 2276
rect 3373 2144 3379 2216
rect 3469 2204 3475 2296
rect 3517 2184 3523 2196
rect 3405 2124 3411 2156
rect 3389 2044 3395 2096
rect 3108 2037 3123 2043
rect 3101 1984 3107 2016
rect 3117 1864 3123 2037
rect 3245 1984 3251 2036
rect 3032 1806 3038 1814
rect 3046 1806 3052 1814
rect 3060 1806 3066 1814
rect 3074 1806 3080 1814
rect 3149 1764 3155 1896
rect 3165 1824 3171 1876
rect 3213 1804 3219 1836
rect 2973 1604 2979 1736
rect 2989 1544 2995 1756
rect 3325 1724 3331 1896
rect 3405 1864 3411 1956
rect 3437 1944 3443 2136
rect 3453 2044 3459 2116
rect 3501 1920 3507 1958
rect 3533 1944 3539 2296
rect 3549 2264 3555 2316
rect 3565 2284 3571 2516
rect 3581 2462 3587 2500
rect 3837 2404 3843 2436
rect 3885 2404 3891 2556
rect 3901 2503 3907 2576
rect 3917 2524 3923 2576
rect 3901 2497 3923 2503
rect 3917 2464 3923 2497
rect 3933 2484 3939 2737
rect 3949 2523 3955 2696
rect 3965 2684 3971 2856
rect 3981 2584 3987 2896
rect 4013 2704 4019 2976
rect 3997 2697 4012 2703
rect 3981 2544 3987 2556
rect 3997 2524 4003 2697
rect 4013 2664 4019 2676
rect 4029 2604 4035 2916
rect 4061 2864 4067 3316
rect 4109 3064 4115 3076
rect 4141 3064 4147 3356
rect 4173 3324 4179 3336
rect 4237 3324 4243 3496
rect 4349 3484 4355 3516
rect 4317 3424 4323 3456
rect 4349 3384 4355 3476
rect 4317 3304 4323 3376
rect 4269 3244 4275 3296
rect 4349 3284 4355 3336
rect 4365 3304 4371 3356
rect 4333 3204 4339 3236
rect 4125 3024 4131 3036
rect 4157 3004 4163 3096
rect 4173 3084 4179 3096
rect 4189 3084 4195 3156
rect 4237 3124 4243 3196
rect 4365 3184 4371 3296
rect 4429 3244 4435 3496
rect 4461 3344 4467 3516
rect 4765 3464 4771 3716
rect 5053 3664 5059 3716
rect 5117 3664 5123 3716
rect 5293 3662 5299 3716
rect 4829 3604 4835 3636
rect 4797 3484 4803 3596
rect 4861 3520 4867 3558
rect 5005 3520 5011 3558
rect 5213 3524 5219 3636
rect 5325 3544 5331 3596
rect 5325 3524 5331 3536
rect 5293 3464 5299 3476
rect 4493 3444 4499 3456
rect 4525 3344 4531 3396
rect 4557 3344 4563 3356
rect 4477 3304 4483 3316
rect 4557 3304 4563 3336
rect 4621 3324 4627 3396
rect 5229 3364 5235 3456
rect 5261 3424 5267 3436
rect 5309 3404 5315 3436
rect 4685 3344 4691 3356
rect 4445 3204 4451 3296
rect 4285 3124 4291 3176
rect 4493 3104 4499 3236
rect 4205 3024 4211 3096
rect 4189 2944 4195 3016
rect 4285 2924 4291 3096
rect 4381 3084 4387 3096
rect 4509 3044 4515 3196
rect 4541 3164 4547 3276
rect 4605 3264 4611 3316
rect 4568 3206 4574 3214
rect 4582 3206 4588 3214
rect 4596 3206 4602 3214
rect 4610 3206 4616 3214
rect 4349 2984 4355 2996
rect 4429 2984 4435 3016
rect 4285 2844 4291 2896
rect 4333 2784 4339 2916
rect 4349 2884 4355 2936
rect 4109 2684 4115 2736
rect 4141 2724 4147 2736
rect 3949 2517 3964 2523
rect 4013 2464 4019 2536
rect 4029 2524 4035 2596
rect 4045 2544 4051 2676
rect 4077 2664 4083 2676
rect 4061 2564 4067 2636
rect 4061 2544 4067 2556
rect 4125 2544 4131 2696
rect 4141 2604 4147 2696
rect 4205 2684 4211 2776
rect 4317 2704 4323 2716
rect 4333 2704 4339 2756
rect 4397 2744 4403 2856
rect 4413 2784 4419 2916
rect 4429 2784 4435 2936
rect 4429 2704 4435 2716
rect 4445 2704 4451 2716
rect 4461 2704 4467 2716
rect 4173 2644 4179 2676
rect 4205 2604 4211 2676
rect 4141 2544 4147 2596
rect 4093 2464 4099 2536
rect 4109 2444 4115 2516
rect 3597 2304 3603 2376
rect 3741 2320 3747 2358
rect 3709 2284 3715 2296
rect 3565 2164 3571 2276
rect 3661 2263 3667 2276
rect 3725 2263 3731 2276
rect 4045 2264 4051 2336
rect 4061 2324 4067 2436
rect 4109 2424 4115 2436
rect 4093 2284 4099 2356
rect 3661 2257 3731 2263
rect 3837 2204 3843 2256
rect 3677 2164 3683 2196
rect 4013 2184 4019 2216
rect 4109 2164 4115 2256
rect 3677 1964 3683 2156
rect 3709 2144 3715 2156
rect 3901 2124 3907 2136
rect 3773 2044 3779 2100
rect 3789 2024 3795 2116
rect 3901 2044 3907 2116
rect 3741 1904 3747 2016
rect 3437 1844 3443 1876
rect 3373 1744 3379 1796
rect 3405 1784 3411 1836
rect 3469 1784 3475 1816
rect 3469 1744 3475 1776
rect 3533 1724 3539 1796
rect 3565 1744 3571 1776
rect 3581 1744 3587 1836
rect 3629 1784 3635 1876
rect 3645 1744 3651 1876
rect 3661 1724 3667 1896
rect 3741 1784 3747 1896
rect 3821 1864 3827 1956
rect 3805 1784 3811 1816
rect 3917 1784 3923 2036
rect 3949 1924 3955 1976
rect 3965 1884 3971 1896
rect 3981 1804 3987 2116
rect 4029 1904 4035 2116
rect 4125 2104 4131 2536
rect 4157 2504 4163 2596
rect 4189 2524 4195 2556
rect 4205 2484 4211 2516
rect 4221 2444 4227 2696
rect 4253 2644 4259 2676
rect 4269 2544 4275 2616
rect 4285 2604 4291 2676
rect 4301 2624 4307 2696
rect 4413 2684 4419 2696
rect 4301 2544 4307 2556
rect 4285 2504 4291 2516
rect 4317 2503 4323 2636
rect 4333 2584 4339 2676
rect 4413 2564 4419 2596
rect 4365 2544 4371 2556
rect 4333 2504 4339 2536
rect 4317 2497 4332 2503
rect 4189 2384 4195 2416
rect 4285 2324 4291 2496
rect 4141 2124 4147 2296
rect 4061 1920 4067 1958
rect 4125 1944 4131 2036
rect 4173 1984 4179 2036
rect 4045 1884 4051 1896
rect 3709 1724 3715 1776
rect 3652 1717 3660 1723
rect 3085 1662 3091 1700
rect 3181 1524 3187 1656
rect 2893 1464 2899 1496
rect 2813 1404 2819 1456
rect 3085 1444 3091 1476
rect 2845 1324 2851 1356
rect 2973 1344 2979 1436
rect 3032 1406 3038 1414
rect 3046 1406 3052 1414
rect 3060 1406 3066 1414
rect 3074 1406 3080 1414
rect 2765 1304 2771 1316
rect 2797 1084 2803 1116
rect 2829 1104 2835 1176
rect 2845 1104 2851 1316
rect 2484 697 2499 703
rect 2365 564 2371 636
rect 2461 584 2467 676
rect 2525 624 2531 736
rect 2557 724 2563 996
rect 2669 964 2675 996
rect 2669 664 2675 956
rect 2701 924 2707 936
rect 2765 844 2771 900
rect 2845 804 2851 1076
rect 2877 924 2883 1316
rect 2941 1262 2947 1300
rect 3149 1184 3155 1516
rect 2909 1104 2915 1136
rect 3181 1084 3187 1436
rect 3197 1344 3203 1596
rect 3261 1520 3267 1558
rect 3325 1504 3331 1716
rect 3405 1664 3411 1696
rect 3517 1684 3523 1696
rect 3229 1324 3235 1456
rect 3373 1364 3379 1376
rect 3245 1244 3251 1296
rect 3373 1204 3379 1356
rect 3453 1244 3459 1316
rect 3085 1064 3091 1076
rect 2845 720 2851 758
rect 2861 704 2867 916
rect 2877 844 2883 896
rect 2893 684 2899 1056
rect 2973 944 2979 1036
rect 3032 1006 3038 1014
rect 3046 1006 3052 1014
rect 3060 1006 3066 1014
rect 3074 1006 3080 1014
rect 2269 557 2291 563
rect 1933 544 1939 556
rect 1965 544 1971 556
rect 1837 444 1843 496
rect 1677 284 1683 316
rect 1803 304 1809 316
rect 1725 144 1731 236
rect 1853 204 1859 516
rect 1885 204 1891 296
rect 1965 264 1971 536
rect 2189 504 2195 536
rect 2269 504 2275 557
rect 2061 320 2067 358
rect 2173 324 2179 436
rect 2237 324 2243 476
rect 2221 284 2227 316
rect 2285 284 2291 536
rect 2317 504 2323 556
rect 2557 504 2563 536
rect 2461 444 2467 496
rect 2397 320 2403 358
rect 2461 284 2467 396
rect 1837 124 1843 196
rect 1965 164 1971 256
rect 2157 124 2163 256
rect 2173 144 2179 236
rect 2237 144 2243 236
rect 2317 224 2323 256
rect 2493 184 2499 256
rect 2525 184 2531 216
rect 2589 184 2595 556
rect 2701 384 2707 516
rect 2845 504 2851 636
rect 2893 544 2899 676
rect 3101 644 3107 1036
rect 3229 704 3235 1096
rect 3309 1064 3315 1196
rect 3405 1120 3411 1158
rect 3309 964 3315 1056
rect 3485 1004 3491 1456
rect 3533 1324 3539 1716
rect 3549 1524 3555 1696
rect 3549 1364 3555 1456
rect 3565 1324 3571 1556
rect 3597 1364 3603 1496
rect 3549 1317 3564 1323
rect 3501 1084 3507 1096
rect 3533 1084 3539 1236
rect 3549 1104 3555 1317
rect 3485 964 3491 996
rect 3581 924 3587 1036
rect 3405 862 3411 916
rect 3581 908 3587 916
rect 3261 804 3267 836
rect 3325 724 3331 776
rect 2893 444 2899 516
rect 2941 504 2947 636
rect 3032 606 3038 614
rect 3046 606 3052 614
rect 3060 606 3066 614
rect 3074 606 3080 614
rect 3117 584 3123 696
rect 3373 684 3379 796
rect 3229 664 3235 676
rect 2365 164 2371 176
rect 2605 124 2611 196
rect 2653 124 2659 236
rect 2733 124 2739 296
rect 2749 204 2755 436
rect 2797 404 2803 436
rect 2781 320 2787 358
rect 2845 284 2851 296
rect 2877 284 2883 436
rect 2973 303 2979 516
rect 3021 462 3027 500
rect 2964 297 2979 303
rect 2877 223 2883 256
rect 2861 217 2883 223
rect 2861 184 2867 217
rect 2861 164 2867 176
rect 2973 124 2979 297
rect 3032 206 3038 214
rect 3046 206 3052 214
rect 3060 206 3066 214
rect 3074 206 3080 214
rect 3101 124 3107 256
rect 3117 184 3123 556
rect 3197 524 3203 576
rect 3133 384 3139 436
rect 3261 304 3267 576
rect 3389 524 3395 636
rect 3421 584 3427 716
rect 3597 684 3603 796
rect 3613 784 3619 1676
rect 3645 1503 3651 1716
rect 3693 1704 3699 1716
rect 3709 1564 3715 1716
rect 3853 1704 3859 1776
rect 3981 1726 3987 1756
rect 4045 1744 4051 1836
rect 4125 1824 4131 1876
rect 4237 1823 4243 2096
rect 4221 1817 4243 1823
rect 3741 1584 3747 1696
rect 3805 1584 3811 1656
rect 3636 1497 3651 1503
rect 3629 1384 3635 1496
rect 3661 1484 3667 1536
rect 3645 1444 3651 1476
rect 3693 1464 3699 1516
rect 3645 1344 3651 1436
rect 3693 1404 3699 1436
rect 3693 1324 3699 1376
rect 3693 1164 3699 1316
rect 3629 1024 3635 1056
rect 3645 724 3651 776
rect 3661 704 3667 1156
rect 3693 1124 3699 1136
rect 3309 384 3315 516
rect 3373 503 3379 516
rect 3373 497 3395 503
rect 3277 304 3283 316
rect 3341 204 3347 436
rect 3389 384 3395 497
rect 3405 464 3411 536
rect 3437 504 3443 676
rect 3661 664 3667 696
rect 3677 684 3683 796
rect 3709 724 3715 1516
rect 3741 1444 3747 1496
rect 3757 1484 3763 1496
rect 3805 1424 3811 1496
rect 3837 1484 3843 1676
rect 4045 1584 4051 1736
rect 4141 1724 4147 1756
rect 4173 1744 4179 1756
rect 4061 1624 4067 1716
rect 4157 1684 4163 1736
rect 4173 1704 4179 1716
rect 3901 1524 3907 1556
rect 3933 1404 3939 1496
rect 3821 1324 3827 1356
rect 3773 1224 3779 1296
rect 3853 1244 3859 1300
rect 3741 1124 3747 1176
rect 3949 1104 3955 1236
rect 3869 1064 3875 1096
rect 3869 1004 3875 1056
rect 3821 964 3827 996
rect 4013 984 4019 1216
rect 4045 1103 4051 1536
rect 4077 1524 4083 1636
rect 4061 1324 4067 1496
rect 4093 1484 4099 1576
rect 4109 1504 4115 1616
rect 4093 1344 4099 1476
rect 4109 1384 4115 1496
rect 4125 1484 4131 1576
rect 4205 1484 4211 1676
rect 4061 1184 4067 1216
rect 4045 1097 4067 1103
rect 4029 1024 4035 1036
rect 3725 862 3731 900
rect 3789 824 3795 936
rect 4045 924 4051 1036
rect 3981 784 3987 816
rect 3869 724 3875 736
rect 4013 724 4019 896
rect 4061 844 4067 1097
rect 4077 964 4083 1076
rect 4125 924 4131 1396
rect 4141 1344 4147 1356
rect 4157 1104 4163 1236
rect 4221 1184 4227 1817
rect 4237 1724 4243 1776
rect 4237 1504 4243 1716
rect 4253 1204 4259 1716
rect 4285 1583 4291 2276
rect 4349 2244 4355 2516
rect 4365 2404 4371 2536
rect 4413 2504 4419 2556
rect 4445 2544 4451 2696
rect 4493 2684 4499 3036
rect 4509 2964 4515 2996
rect 4573 2964 4579 3036
rect 4589 2964 4595 3156
rect 4605 2904 4611 3176
rect 4653 3164 4659 3336
rect 4685 3304 4691 3336
rect 4525 2784 4531 2876
rect 4653 2844 4659 3076
rect 4701 3004 4707 3296
rect 4717 3264 4723 3316
rect 4781 3304 4787 3316
rect 4717 3124 4723 3256
rect 4749 3124 4755 3236
rect 4781 3144 4787 3296
rect 4813 3184 4819 3316
rect 4829 3304 4835 3336
rect 4845 3324 4851 3336
rect 4877 3264 4883 3296
rect 4813 3124 4819 3136
rect 4845 3104 4851 3136
rect 4861 3124 4867 3236
rect 4877 3124 4883 3156
rect 4717 3004 4723 3056
rect 4861 3024 4867 3076
rect 4669 2904 4675 2956
rect 4568 2806 4574 2814
rect 4582 2806 4588 2814
rect 4596 2806 4602 2814
rect 4610 2806 4616 2814
rect 4509 2704 4515 2736
rect 4541 2704 4547 2716
rect 4413 2204 4419 2496
rect 4445 2264 4451 2536
rect 4461 2503 4467 2676
rect 4477 2524 4483 2536
rect 4493 2503 4499 2676
rect 4509 2564 4515 2696
rect 4541 2544 4547 2596
rect 4557 2584 4563 2736
rect 4637 2724 4643 2836
rect 4653 2704 4659 2776
rect 4669 2764 4675 2876
rect 4685 2784 4691 2916
rect 4717 2864 4723 2996
rect 4765 2984 4771 3016
rect 4733 2924 4739 2936
rect 4781 2924 4787 2956
rect 4669 2744 4675 2756
rect 4685 2737 4700 2743
rect 4557 2504 4563 2536
rect 4461 2497 4483 2503
rect 4493 2497 4515 2503
rect 4477 2464 4483 2497
rect 4461 2244 4467 2296
rect 4477 2284 4483 2456
rect 4493 2304 4499 2476
rect 4509 2343 4515 2497
rect 4525 2464 4531 2496
rect 4637 2424 4643 2616
rect 4653 2544 4659 2596
rect 4685 2584 4691 2737
rect 4717 2724 4723 2836
rect 4797 2824 4803 2896
rect 4749 2784 4755 2796
rect 4749 2704 4755 2756
rect 4781 2724 4787 2756
rect 4717 2624 4723 2696
rect 4653 2504 4659 2516
rect 4669 2484 4675 2576
rect 4717 2524 4723 2576
rect 4749 2524 4755 2696
rect 4765 2684 4771 2716
rect 4797 2664 4803 2736
rect 4568 2406 4574 2414
rect 4582 2406 4588 2414
rect 4596 2406 4602 2414
rect 4610 2406 4616 2414
rect 4509 2337 4531 2343
rect 4509 2284 4515 2316
rect 4525 2304 4531 2337
rect 4541 2304 4547 2396
rect 4573 2337 4620 2343
rect 4573 2304 4579 2337
rect 4429 2164 4435 2236
rect 4557 2164 4563 2276
rect 4589 2244 4595 2276
rect 4605 2204 4611 2296
rect 4637 2204 4643 2376
rect 4653 2164 4659 2476
rect 4733 2384 4739 2496
rect 4749 2404 4755 2516
rect 4765 2484 4771 2656
rect 4781 2584 4787 2616
rect 4813 2584 4819 2836
rect 4829 2704 4835 2716
rect 4829 2564 4835 2696
rect 4845 2664 4851 2916
rect 4861 2704 4867 2936
rect 4877 2824 4883 3036
rect 4893 3004 4899 3336
rect 4941 3284 4947 3296
rect 4909 3224 4915 3236
rect 4909 3084 4915 3176
rect 4957 3104 4963 3276
rect 4989 3123 4995 3236
rect 5005 3164 5011 3316
rect 5053 3304 5059 3356
rect 5261 3344 5267 3396
rect 5021 3184 5027 3236
rect 5053 3183 5059 3296
rect 5069 3204 5075 3236
rect 5053 3177 5075 3183
rect 4973 3117 4995 3123
rect 4973 3084 4979 3117
rect 5053 3104 5059 3116
rect 4925 3064 4931 3076
rect 4941 2984 4947 3056
rect 4973 2984 4979 3016
rect 4893 2964 4899 2976
rect 4916 2957 4931 2963
rect 4893 2924 4899 2936
rect 4909 2804 4915 2936
rect 4925 2924 4931 2957
rect 4989 2924 4995 3096
rect 5021 3063 5027 3096
rect 5069 3084 5075 3177
rect 5085 3083 5091 3096
rect 5101 3083 5107 3316
rect 5133 3124 5139 3176
rect 5181 3124 5187 3216
rect 5213 3144 5219 3196
rect 5213 3084 5219 3116
rect 5085 3077 5107 3083
rect 5005 3057 5027 3063
rect 5005 2964 5011 3057
rect 4925 2784 4931 2916
rect 4957 2884 4963 2896
rect 4877 2684 4883 2756
rect 4893 2704 4899 2736
rect 4909 2697 4924 2703
rect 4861 2664 4867 2676
rect 4845 2624 4851 2636
rect 4861 2563 4867 2656
rect 4909 2564 4915 2697
rect 4973 2703 4979 2816
rect 4989 2763 4995 2896
rect 5005 2864 5011 2896
rect 5005 2784 5011 2856
rect 4989 2757 5004 2763
rect 5021 2724 5027 2996
rect 5069 2964 5075 3076
rect 5069 2824 5075 2936
rect 5053 2784 5059 2796
rect 4973 2697 4995 2703
rect 4941 2644 4947 2676
rect 4957 2664 4963 2696
rect 4941 2564 4947 2636
rect 4861 2557 4876 2563
rect 4829 2504 4835 2516
rect 4813 2424 4819 2436
rect 4829 2424 4835 2496
rect 4845 2444 4851 2456
rect 4676 2337 4723 2343
rect 4717 2324 4723 2337
rect 4749 2324 4755 2336
rect 4708 2297 4732 2303
rect 4669 2264 4675 2276
rect 4685 2164 4691 2236
rect 4717 2164 4723 2276
rect 4765 2263 4771 2336
rect 4845 2324 4851 2436
rect 4781 2284 4787 2296
rect 4829 2284 4835 2296
rect 4765 2257 4787 2263
rect 4749 2164 4755 2196
rect 4781 2164 4787 2257
rect 4813 2184 4819 2276
rect 4829 2184 4835 2276
rect 4813 2164 4819 2176
rect 4317 1724 4323 1836
rect 4333 1744 4339 1996
rect 4349 1884 4355 2116
rect 4429 2004 4435 2156
rect 4861 2144 4867 2557
rect 4877 2284 4883 2316
rect 4893 2304 4899 2536
rect 4909 2444 4915 2556
rect 4957 2524 4963 2616
rect 4957 2504 4963 2516
rect 4909 2384 4915 2396
rect 4957 2324 4963 2376
rect 4973 2204 4979 2256
rect 4989 2203 4995 2697
rect 5005 2604 5011 2656
rect 5021 2644 5027 2656
rect 5021 2624 5027 2636
rect 5037 2604 5043 2696
rect 5053 2644 5059 2696
rect 5069 2584 5075 2716
rect 5085 2704 5091 2916
rect 5101 2744 5107 3077
rect 5117 2984 5123 3056
rect 5181 2944 5187 3036
rect 5213 3024 5219 3076
rect 5213 2964 5219 2976
rect 5229 2964 5235 3176
rect 5117 2937 5132 2943
rect 5117 2704 5123 2937
rect 5213 2924 5219 2956
rect 5181 2904 5187 2916
rect 5005 2464 5011 2556
rect 5021 2544 5027 2576
rect 5053 2544 5059 2556
rect 5085 2524 5091 2636
rect 5117 2584 5123 2676
rect 5133 2664 5139 2816
rect 5165 2744 5171 2896
rect 5197 2784 5203 2836
rect 5165 2664 5171 2696
rect 5213 2664 5219 2856
rect 5229 2684 5235 2796
rect 5245 2784 5251 3216
rect 5261 3184 5267 3316
rect 5325 3262 5331 3300
rect 5261 3044 5267 3096
rect 5277 3084 5283 3136
rect 5293 3104 5299 3116
rect 5341 3104 5347 3536
rect 5357 3324 5363 3436
rect 5373 3364 5379 3756
rect 5469 3708 5475 3796
rect 5549 3744 5555 3836
rect 5581 3724 5587 3736
rect 5549 3664 5555 3716
rect 5517 3584 5523 3656
rect 5389 3504 5395 3556
rect 5405 3504 5411 3516
rect 5373 3124 5379 3336
rect 5405 3123 5411 3496
rect 5396 3117 5411 3123
rect 5389 3104 5395 3116
rect 5325 3077 5340 3083
rect 5261 2944 5267 3016
rect 5261 2723 5267 2836
rect 5277 2764 5283 3076
rect 5293 2984 5299 3076
rect 5325 2944 5331 3077
rect 5421 3064 5427 3576
rect 5517 3564 5523 3576
rect 5549 3524 5555 3596
rect 5597 3544 5603 3876
rect 5661 3864 5667 3916
rect 5725 3904 5731 4036
rect 5613 3704 5619 3856
rect 5661 3744 5667 3836
rect 5581 3484 5587 3516
rect 5597 3504 5603 3536
rect 5453 3404 5459 3476
rect 5549 3403 5555 3436
rect 5533 3397 5555 3403
rect 5437 3244 5443 3296
rect 5453 3084 5459 3396
rect 5533 3344 5539 3397
rect 5645 3384 5651 3516
rect 5661 3484 5667 3736
rect 5677 3724 5683 3876
rect 5709 3844 5715 3876
rect 5725 3864 5731 3876
rect 5693 3524 5699 3576
rect 5709 3344 5715 3676
rect 5741 3624 5747 4096
rect 5757 3904 5763 4157
rect 5773 3924 5779 3976
rect 5773 3724 5779 3896
rect 5789 3504 5795 4116
rect 5821 4062 5827 4100
rect 5917 3983 5923 4156
rect 5997 4124 6003 4416
rect 6125 4284 6131 5336
rect 6013 4164 6019 4236
rect 5901 3977 5923 3983
rect 5869 3884 5875 3896
rect 5901 3864 5907 3977
rect 5901 3764 5907 3856
rect 5933 3744 5939 3756
rect 5901 3484 5907 3496
rect 5789 3423 5795 3476
rect 5789 3417 5811 3423
rect 5805 3384 5811 3417
rect 5789 3324 5795 3336
rect 5821 3303 5827 3456
rect 5853 3344 5859 3416
rect 5933 3344 5939 3716
rect 6029 3644 6035 3696
rect 6045 3524 6051 3996
rect 6061 3984 6067 3996
rect 6077 3724 6083 4036
rect 6125 3964 6131 4276
rect 5853 3324 5859 3336
rect 5933 3304 5939 3316
rect 5949 3304 5955 3376
rect 5981 3364 5987 3496
rect 5997 3344 6003 3476
rect 5997 3324 6003 3336
rect 5805 3297 5827 3303
rect 5469 3184 5475 3236
rect 5533 3124 5539 3176
rect 5341 2924 5347 3036
rect 5373 2964 5379 3036
rect 5421 2944 5427 3036
rect 5293 2804 5299 2836
rect 5309 2784 5315 2816
rect 5261 2717 5276 2723
rect 5213 2644 5219 2656
rect 5149 2584 5155 2596
rect 5197 2584 5203 2616
rect 5101 2524 5107 2556
rect 5005 2304 5011 2416
rect 5021 2304 5027 2496
rect 5085 2484 5091 2516
rect 5117 2504 5123 2516
rect 5037 2424 5043 2436
rect 5053 2364 5059 2456
rect 5069 2384 5075 2436
rect 5005 2224 5011 2276
rect 5053 2204 5059 2356
rect 5085 2344 5091 2476
rect 5085 2284 5091 2316
rect 5101 2283 5107 2456
rect 5133 2384 5139 2516
rect 5165 2504 5171 2556
rect 5181 2544 5187 2576
rect 5229 2524 5235 2596
rect 5117 2344 5123 2356
rect 5149 2324 5155 2396
rect 5181 2324 5187 2516
rect 5229 2324 5235 2396
rect 5245 2384 5251 2656
rect 5277 2584 5283 2696
rect 5293 2584 5299 2676
rect 5309 2604 5315 2696
rect 5261 2503 5267 2536
rect 5309 2524 5315 2596
rect 5261 2497 5283 2503
rect 5261 2344 5267 2356
rect 5245 2304 5251 2316
rect 5133 2284 5139 2296
rect 5092 2277 5107 2283
rect 4989 2197 5011 2203
rect 5005 2144 5011 2197
rect 4525 2062 4531 2100
rect 5037 2104 5043 2156
rect 5117 2124 5123 2156
rect 5165 2144 5171 2296
rect 5181 2224 5187 2296
rect 5197 2184 5203 2256
rect 5197 2124 5203 2176
rect 5229 2164 5235 2216
rect 5261 2144 5267 2256
rect 5277 2124 5283 2497
rect 5293 2224 5299 2316
rect 5309 2304 5315 2316
rect 5309 2104 5315 2236
rect 5325 2184 5331 2776
rect 5341 2764 5347 2916
rect 5453 2844 5459 3076
rect 5741 3064 5747 3096
rect 5661 3044 5667 3056
rect 5341 2704 5347 2736
rect 5373 2724 5379 2796
rect 5357 2624 5363 2676
rect 5357 2523 5363 2556
rect 5373 2544 5379 2716
rect 5389 2644 5395 2696
rect 5405 2684 5411 2716
rect 5389 2524 5395 2636
rect 5421 2624 5427 2636
rect 5421 2583 5427 2616
rect 5421 2577 5443 2583
rect 5421 2524 5427 2556
rect 5437 2544 5443 2577
rect 5453 2564 5459 2636
rect 5469 2604 5475 3036
rect 5549 2964 5555 3036
rect 5581 2944 5587 2956
rect 5725 2944 5731 3016
rect 5757 2984 5763 3116
rect 5501 2543 5507 2716
rect 5549 2684 5555 2936
rect 5789 2924 5795 3056
rect 5805 3044 5811 3297
rect 5917 3123 5923 3236
rect 5917 3117 5932 3123
rect 5997 3084 6003 3316
rect 5901 3024 5907 3076
rect 5901 2944 5907 2996
rect 5933 2964 5939 3036
rect 5949 3004 5955 3036
rect 5645 2862 5651 2900
rect 5565 2704 5571 2756
rect 5645 2724 5651 2736
rect 5492 2537 5507 2543
rect 5348 2517 5363 2523
rect 5453 2464 5459 2536
rect 5501 2463 5507 2537
rect 5517 2503 5523 2636
rect 5556 2537 5571 2543
rect 5517 2497 5532 2503
rect 5501 2457 5523 2463
rect 5357 2384 5363 2436
rect 5373 2344 5379 2416
rect 5405 2324 5411 2376
rect 5501 2324 5507 2436
rect 5453 2304 5459 2316
rect 5341 2184 5347 2276
rect 5469 2224 5475 2316
rect 5517 2284 5523 2457
rect 5517 2264 5523 2276
rect 5389 2184 5395 2196
rect 5469 2144 5475 2216
rect 5533 2204 5539 2276
rect 5565 2204 5571 2537
rect 5581 2384 5587 2636
rect 5613 2584 5619 2716
rect 5677 2704 5683 2756
rect 5693 2704 5699 2916
rect 5757 2764 5763 2896
rect 5805 2844 5811 2896
rect 5933 2843 5939 2956
rect 6013 2924 6019 3476
rect 6029 3384 6035 3436
rect 6061 3384 6067 3476
rect 6077 3364 6083 3716
rect 6125 3684 6131 3696
rect 6125 3484 6131 3496
rect 6109 3344 6115 3396
rect 6045 3064 6051 3096
rect 5933 2837 5955 2843
rect 5725 2744 5731 2756
rect 5757 2724 5763 2736
rect 5613 2484 5619 2576
rect 5645 2544 5651 2636
rect 5661 2384 5667 2436
rect 5597 2284 5603 2336
rect 5661 2284 5667 2356
rect 5773 2304 5779 2596
rect 5789 2524 5795 2696
rect 5949 2664 5955 2837
rect 6029 2824 6035 3056
rect 6045 2720 6051 2758
rect 5869 2564 5875 2656
rect 5869 2443 5875 2556
rect 6045 2524 6051 2676
rect 5965 2462 5971 2500
rect 5853 2437 5875 2443
rect 5693 2224 5699 2236
rect 5549 2144 5555 2156
rect 5581 2144 5587 2176
rect 4568 2006 4574 2014
rect 4582 2006 4588 2014
rect 4596 2006 4602 2014
rect 4610 2006 4616 2014
rect 4381 1924 4387 1976
rect 4381 1884 4387 1896
rect 4509 1884 4515 1996
rect 4669 1904 4675 2036
rect 4269 1577 4291 1583
rect 4269 1344 4275 1577
rect 4285 1524 4291 1556
rect 4285 1504 4291 1516
rect 4317 1324 4323 1376
rect 4333 1304 4339 1316
rect 4269 1184 4275 1256
rect 4285 1224 4291 1296
rect 4317 1164 4323 1236
rect 4285 1124 4291 1156
rect 4157 1084 4163 1096
rect 4189 924 4195 996
rect 4221 984 4227 1116
rect 4285 1084 4291 1096
rect 4333 1084 4339 1276
rect 3677 664 3683 676
rect 3469 544 3475 636
rect 3773 624 3779 676
rect 3533 584 3539 596
rect 3709 584 3715 616
rect 3549 564 3555 576
rect 3629 544 3635 576
rect 3789 544 3795 696
rect 3853 564 3859 636
rect 3885 584 3891 676
rect 3901 604 3907 696
rect 3933 644 3939 716
rect 3949 684 3955 716
rect 4061 684 4067 836
rect 4093 644 4099 676
rect 4125 664 4131 916
rect 4157 884 4163 896
rect 4205 724 4211 956
rect 4253 943 4259 1056
rect 4333 984 4339 1076
rect 4349 1024 4355 1496
rect 4381 1464 4387 1856
rect 4477 1824 4483 1876
rect 4509 1864 4515 1876
rect 4445 1644 4451 1696
rect 4461 1684 4467 1736
rect 4477 1663 4483 1716
rect 4461 1657 4483 1663
rect 4429 1637 4444 1643
rect 4429 1504 4435 1637
rect 4461 1584 4467 1657
rect 4509 1544 4515 1816
rect 4573 1684 4579 1736
rect 4484 1517 4499 1523
rect 4493 1504 4499 1517
rect 4397 1404 4403 1456
rect 4413 1364 4419 1496
rect 4365 1104 4371 1216
rect 4413 1144 4419 1356
rect 4429 1303 4435 1496
rect 4429 1297 4444 1303
rect 4253 937 4275 943
rect 4269 924 4275 937
rect 4237 804 4243 916
rect 4253 844 4259 896
rect 4173 644 4179 696
rect 3485 524 3491 536
rect 3444 497 3452 503
rect 3389 324 3395 376
rect 3453 284 3459 496
rect 3469 324 3475 456
rect 3517 384 3523 536
rect 3549 464 3555 536
rect 3565 384 3571 536
rect 3581 504 3587 516
rect 3613 504 3619 516
rect 3629 504 3635 536
rect 3357 264 3363 276
rect 3469 264 3475 316
rect 3485 284 3491 296
rect 3277 144 3283 196
rect 3469 184 3475 256
rect 3309 164 3315 176
rect 3485 144 3491 276
rect 3501 164 3507 336
rect 3565 164 3571 296
rect 3613 264 3619 496
rect 3789 444 3795 500
rect 3853 304 3859 516
rect 3885 324 3891 376
rect 3629 164 3635 256
rect 3677 124 3683 296
rect 3757 224 3763 256
rect 3805 164 3811 216
rect 3949 184 3955 236
rect 3997 124 4003 616
rect 4045 584 4051 596
rect 4093 544 4099 556
rect 4093 164 4099 536
rect 4141 524 4147 536
rect 4189 524 4195 616
rect 4205 604 4211 716
rect 4221 684 4227 716
rect 4237 704 4243 796
rect 4253 744 4259 836
rect 4269 764 4275 916
rect 4285 784 4291 876
rect 4301 844 4307 956
rect 4333 944 4339 976
rect 4397 924 4403 1116
rect 4413 1004 4419 1096
rect 4429 1084 4435 1276
rect 4477 1264 4483 1356
rect 4525 1344 4531 1676
rect 4541 1484 4547 1656
rect 4568 1606 4574 1614
rect 4582 1606 4588 1614
rect 4596 1606 4602 1614
rect 4610 1606 4616 1614
rect 4557 1384 4563 1536
rect 4637 1444 4643 1716
rect 4669 1564 4675 1836
rect 4701 1764 4707 2036
rect 4685 1664 4691 1696
rect 4701 1604 4707 1736
rect 4637 1384 4643 1436
rect 4445 1164 4451 1236
rect 4461 1144 4467 1196
rect 4461 1103 4467 1136
rect 4452 1097 4467 1103
rect 4429 923 4435 1076
rect 4493 1064 4499 1316
rect 4509 1284 4515 1316
rect 4509 1124 4515 1156
rect 4477 964 4483 1056
rect 4493 984 4499 1036
rect 4509 1004 4515 1096
rect 4525 1044 4531 1296
rect 4568 1206 4574 1214
rect 4582 1206 4588 1214
rect 4596 1206 4602 1214
rect 4610 1206 4616 1214
rect 4429 917 4444 923
rect 4253 684 4259 716
rect 4269 704 4275 716
rect 4285 684 4291 696
rect 4237 644 4243 656
rect 4189 384 4195 516
rect 4221 504 4227 596
rect 4237 524 4243 636
rect 4253 563 4259 576
rect 4253 557 4268 563
rect 4221 284 4227 496
rect 4285 304 4291 676
rect 4301 344 4307 716
rect 4317 384 4323 496
rect 4109 124 4115 136
rect 4237 124 4243 216
rect 4253 144 4259 276
rect 4269 184 4275 296
rect 4333 224 4339 916
rect 4381 704 4387 776
rect 4397 704 4403 836
rect 4413 784 4419 916
rect 4445 904 4451 916
rect 4429 703 4435 896
rect 4461 744 4467 796
rect 4445 724 4451 736
rect 4461 724 4467 736
rect 4429 697 4444 703
rect 4349 604 4355 636
rect 4397 584 4403 676
rect 4413 644 4419 696
rect 4477 684 4483 936
rect 4525 924 4531 956
rect 4397 557 4428 563
rect 4365 504 4371 556
rect 4397 544 4403 557
rect 4381 517 4396 523
rect 4333 184 4339 196
rect 1757 44 1763 96
rect 1869 44 1875 100
rect 2237 44 2243 96
rect 2765 62 2771 100
rect 3213 44 3219 100
rect 3677 44 3683 96
rect 4253 84 4259 116
rect 4349 84 4355 316
rect 4365 304 4371 316
rect 4381 304 4387 517
rect 4413 283 4419 536
rect 4445 504 4451 556
rect 4461 524 4467 556
rect 4477 544 4483 676
rect 4493 604 4499 696
rect 4493 524 4499 596
rect 4509 544 4515 676
rect 4541 664 4547 1096
rect 4557 1084 4563 1096
rect 4637 1024 4643 1036
rect 4637 964 4643 1016
rect 4669 964 4675 1496
rect 4701 1364 4707 1556
rect 4717 1484 4723 1496
rect 4701 1083 4707 1356
rect 4717 1144 4723 1456
rect 4733 1384 4739 2036
rect 4765 1924 4771 2036
rect 4797 1964 4803 2036
rect 4893 1944 4899 2096
rect 4941 2062 4947 2100
rect 5117 2044 5123 2096
rect 4957 1904 4963 1916
rect 4749 1724 4755 1776
rect 4765 1744 4771 1896
rect 4941 1884 4947 1896
rect 5005 1844 5011 1916
rect 4925 1744 4931 1836
rect 4781 1724 4787 1736
rect 4829 1724 4835 1736
rect 4973 1724 4979 1796
rect 4989 1784 4995 1836
rect 5021 1784 5027 1916
rect 5117 1884 5123 2036
rect 5037 1864 5043 1876
rect 5165 1864 5171 2056
rect 5181 1924 5187 1936
rect 5229 1864 5235 1876
rect 5261 1864 5267 1936
rect 5373 1904 5379 1916
rect 5165 1844 5171 1856
rect 5293 1844 5299 1896
rect 5149 1824 5155 1836
rect 5101 1784 5107 1796
rect 4765 1484 4771 1696
rect 4829 1664 4835 1716
rect 4845 1684 4851 1716
rect 4893 1684 4899 1696
rect 4845 1504 4851 1556
rect 4893 1504 4899 1516
rect 4813 1464 4819 1476
rect 4829 1464 4835 1496
rect 4893 1484 4899 1496
rect 4781 1344 4787 1436
rect 4781 1324 4787 1336
rect 4749 1284 4755 1316
rect 4756 1277 4771 1283
rect 4765 1124 4771 1277
rect 4765 1104 4771 1116
rect 4701 1077 4716 1083
rect 4781 1064 4787 1076
rect 4557 904 4563 916
rect 4589 864 4595 936
rect 4669 924 4675 956
rect 4717 924 4723 1056
rect 4749 924 4755 1036
rect 4568 806 4574 814
rect 4582 806 4588 814
rect 4596 806 4602 814
rect 4610 806 4616 814
rect 4573 704 4579 756
rect 4589 584 4595 676
rect 4557 524 4563 556
rect 4653 524 4659 916
rect 4701 724 4707 836
rect 4717 744 4723 916
rect 4765 904 4771 956
rect 4781 844 4787 1056
rect 4797 924 4803 1376
rect 4813 1304 4819 1376
rect 4845 1323 4851 1336
rect 4836 1317 4851 1323
rect 4813 1184 4819 1216
rect 4829 1104 4835 1116
rect 4829 1004 4835 1036
rect 4845 924 4851 1296
rect 4861 1104 4867 1456
rect 4877 1304 4883 1316
rect 4893 1304 4899 1336
rect 4861 1024 4867 1096
rect 4877 1084 4883 1196
rect 4893 1124 4899 1176
rect 4909 1103 4915 1496
rect 4925 1484 4931 1676
rect 4941 1324 4947 1336
rect 4957 1184 4963 1516
rect 4973 1424 4979 1436
rect 4989 1323 4995 1776
rect 5213 1744 5219 1756
rect 5293 1744 5299 1836
rect 5485 1823 5491 1876
rect 5549 1864 5555 2136
rect 5677 2124 5683 2156
rect 5725 2144 5731 2276
rect 5645 2062 5651 2100
rect 5725 2044 5731 2136
rect 5773 2124 5779 2296
rect 5853 2264 5859 2437
rect 5885 2284 5891 2376
rect 5917 2144 5923 2196
rect 5741 2104 5747 2116
rect 5581 1924 5587 1976
rect 5693 1920 5699 1958
rect 5757 1924 5763 2116
rect 5773 1984 5779 2096
rect 5485 1817 5507 1823
rect 5501 1784 5507 1817
rect 5549 1803 5555 1856
rect 5533 1797 5555 1803
rect 5021 1664 5027 1736
rect 5053 1703 5059 1736
rect 5069 1724 5075 1736
rect 5133 1717 5148 1723
rect 5053 1697 5075 1703
rect 5069 1604 5075 1697
rect 5133 1604 5139 1717
rect 5165 1703 5171 1736
rect 5373 1724 5379 1736
rect 5149 1697 5171 1703
rect 5053 1504 5059 1536
rect 5005 1464 5011 1496
rect 5069 1484 5075 1596
rect 5133 1504 5139 1596
rect 5085 1484 5091 1496
rect 5149 1484 5155 1697
rect 5181 1584 5187 1716
rect 5197 1704 5203 1716
rect 5245 1704 5251 1716
rect 5197 1544 5203 1656
rect 5245 1564 5251 1696
rect 5293 1684 5299 1716
rect 5341 1704 5347 1716
rect 5293 1644 5299 1676
rect 5165 1524 5171 1536
rect 5325 1504 5331 1636
rect 5389 1604 5395 1716
rect 5405 1524 5411 1716
rect 5421 1684 5427 1696
rect 5421 1584 5427 1676
rect 5021 1404 5027 1476
rect 5069 1384 5075 1476
rect 5021 1324 5027 1376
rect 5149 1364 5155 1476
rect 5357 1464 5363 1476
rect 4980 1317 4995 1323
rect 5037 1224 5043 1316
rect 5053 1184 5059 1196
rect 5037 1144 5043 1156
rect 5069 1104 5075 1256
rect 4909 1097 4924 1103
rect 4909 944 4915 1076
rect 4925 924 4931 1076
rect 4957 904 4963 996
rect 4973 924 4979 976
rect 4989 943 4995 1036
rect 5037 944 5043 1096
rect 5085 1084 5091 1336
rect 5133 1324 5139 1356
rect 5101 1224 5107 1316
rect 5133 1083 5139 1116
rect 5149 1104 5155 1316
rect 5133 1077 5155 1083
rect 4989 937 5011 943
rect 4797 704 4803 836
rect 4845 704 4851 716
rect 4669 524 4675 656
rect 4733 624 4739 676
rect 4797 604 4803 696
rect 4877 663 4883 836
rect 4925 804 4931 836
rect 4893 724 4899 736
rect 4893 684 4899 716
rect 4877 657 4899 663
rect 4500 517 4515 523
rect 4477 504 4483 516
rect 4445 384 4451 476
rect 4404 277 4419 283
rect 4461 164 4467 276
rect 4477 204 4483 316
rect 4509 304 4515 517
rect 4644 517 4652 523
rect 4557 444 4563 516
rect 4749 504 4755 516
rect 4733 497 4748 503
rect 4637 484 4643 496
rect 4568 406 4574 414
rect 4582 406 4588 414
rect 4596 406 4602 414
rect 4610 406 4616 414
rect 4701 284 4707 296
rect 4461 126 4467 136
rect 4493 104 4499 276
rect 4525 244 4531 276
rect 4573 144 4579 256
rect 4557 124 4563 136
rect 4637 124 4643 216
rect 4653 124 4659 196
rect 4669 144 4675 156
rect 4733 124 4739 497
rect 4749 124 4755 436
rect 4765 384 4771 556
rect 4797 524 4803 556
rect 4845 544 4851 616
rect 4877 526 4883 636
rect 4765 324 4771 376
rect 4781 304 4787 436
rect 4893 304 4899 657
rect 4941 544 4947 676
rect 4973 524 4979 916
rect 4989 764 4995 916
rect 5005 824 5011 937
rect 5037 924 5043 936
rect 5069 924 5075 976
rect 4989 723 4995 756
rect 4989 717 5004 723
rect 5021 704 5027 836
rect 5069 784 5075 916
rect 5085 704 5091 1016
rect 5117 944 5123 1076
rect 5149 1044 5155 1077
rect 5133 884 5139 1036
rect 5165 984 5171 1296
rect 5229 1144 5235 1236
rect 5213 1104 5219 1116
rect 5229 1104 5235 1136
rect 5213 1064 5219 1096
rect 5005 584 5011 676
rect 5037 584 5043 676
rect 5069 663 5075 676
rect 5069 657 5091 663
rect 5021 404 5027 556
rect 5069 383 5075 516
rect 5085 404 5091 657
rect 5117 524 5123 796
rect 5133 664 5139 716
rect 5165 584 5171 876
rect 5117 504 5123 516
rect 5069 377 5084 383
rect 5085 344 5091 376
rect 5101 304 5107 436
rect 4781 264 4787 276
rect 4781 144 4787 156
rect 4829 144 4835 256
rect 4893 244 4899 276
rect 4893 144 4899 236
rect 4845 124 4851 136
rect 4797 104 4803 116
rect 4877 84 4883 136
rect 4925 124 4931 296
rect 5021 284 5027 296
rect 5021 144 5027 276
rect 5101 264 5107 276
rect 5149 124 5155 516
rect 5165 324 5171 336
rect 5181 124 5187 916
rect 5197 904 5203 916
rect 5213 524 5219 1016
rect 5229 924 5235 1096
rect 5245 1084 5251 1456
rect 5293 1344 5299 1456
rect 5357 1424 5363 1456
rect 5373 1344 5379 1436
rect 5437 1344 5443 1736
rect 5453 1724 5459 1756
rect 5453 1564 5459 1696
rect 5453 1484 5459 1536
rect 5485 1384 5491 1696
rect 5517 1344 5523 1596
rect 5533 1484 5539 1797
rect 5581 1724 5587 1736
rect 5661 1724 5667 1896
rect 5581 1364 5587 1716
rect 5597 1684 5603 1716
rect 5645 1704 5651 1716
rect 5677 1684 5683 1756
rect 5629 1484 5635 1676
rect 5677 1544 5683 1676
rect 5620 1457 5635 1463
rect 5597 1384 5603 1396
rect 5629 1364 5635 1457
rect 5693 1444 5699 1476
rect 5389 1324 5395 1336
rect 5517 1324 5523 1336
rect 5293 1304 5299 1316
rect 5469 1284 5475 1316
rect 5533 1304 5539 1316
rect 5613 1304 5619 1356
rect 5629 1344 5635 1356
rect 5501 1144 5507 1236
rect 5341 1104 5347 1136
rect 5373 1124 5379 1136
rect 5565 1104 5571 1296
rect 5693 1244 5699 1316
rect 5709 1304 5715 1316
rect 5677 1124 5683 1156
rect 5693 1104 5699 1116
rect 5293 1084 5299 1096
rect 5245 964 5251 1076
rect 5341 964 5347 1096
rect 5277 944 5283 956
rect 5245 884 5251 916
rect 5229 524 5235 816
rect 5261 704 5267 716
rect 5197 304 5203 316
rect 5213 304 5219 516
rect 5261 444 5267 676
rect 5277 604 5283 936
rect 5325 924 5331 936
rect 5373 924 5379 956
rect 5389 944 5395 1076
rect 5533 1064 5539 1076
rect 5565 1024 5571 1096
rect 5421 984 5427 996
rect 5629 984 5635 1076
rect 5661 984 5667 1036
rect 5453 884 5459 896
rect 5437 764 5443 876
rect 5437 724 5443 736
rect 5277 524 5283 556
rect 5309 544 5315 616
rect 5325 524 5331 536
rect 5213 244 5219 276
rect 5245 264 5251 396
rect 5261 284 5267 436
rect 5325 324 5331 516
rect 5341 484 5347 676
rect 5357 504 5363 556
rect 5357 364 5363 456
rect 5373 384 5379 476
rect 5389 384 5395 576
rect 5421 544 5427 596
rect 5437 584 5443 676
rect 5437 564 5443 576
rect 5405 504 5411 516
rect 5332 317 5347 323
rect 5245 144 5251 256
rect 5213 124 5219 136
rect 5293 124 5299 136
rect 5005 84 5011 118
rect 5261 104 5267 116
rect 5309 104 5315 136
rect 5341 124 5347 317
rect 5357 284 5363 356
rect 5389 324 5395 376
rect 5469 324 5475 756
rect 5485 704 5491 976
rect 5613 944 5619 956
rect 5693 944 5699 976
rect 5709 924 5715 1096
rect 5725 1044 5731 1816
rect 5789 1804 5795 1856
rect 5821 1764 5827 1796
rect 5917 1764 5923 2136
rect 5949 1904 5955 1936
rect 5821 1604 5827 1756
rect 5917 1644 5923 1700
rect 5757 1324 5763 1556
rect 5853 1464 5859 1596
rect 5949 1504 5955 1716
rect 5853 1424 5859 1456
rect 5789 1344 5795 1416
rect 5837 1304 5843 1316
rect 5853 1184 5859 1276
rect 5789 924 5795 1096
rect 5869 1064 5875 1416
rect 5917 1344 5923 1416
rect 5965 1204 5971 2336
rect 5981 2324 5987 2376
rect 6045 2344 6051 2516
rect 6045 2184 6051 2256
rect 6013 1863 6019 1896
rect 6013 1857 6035 1863
rect 5981 1604 5987 1836
rect 5981 1524 5987 1576
rect 5965 1120 5971 1158
rect 5981 1104 5987 1496
rect 5997 1104 6003 1676
rect 6013 1083 6019 1836
rect 6029 1724 6035 1857
rect 6029 1684 6035 1716
rect 6061 1504 6067 2816
rect 6077 2584 6083 3336
rect 6125 3084 6131 3096
rect 6093 2824 6099 2836
rect 6077 1844 6083 2316
rect 6125 1884 6131 1896
rect 6125 1704 6131 1756
rect 6125 1524 6131 1536
rect 6045 1464 6051 1476
rect 6029 1404 6035 1436
rect 6077 1304 6083 1376
rect 5997 1077 6019 1083
rect 5885 944 5891 976
rect 5613 724 5619 856
rect 5501 444 5507 516
rect 5517 484 5523 516
rect 5533 404 5539 636
rect 5549 544 5555 696
rect 5565 624 5571 676
rect 5597 544 5603 636
rect 5517 324 5523 356
rect 5533 324 5539 336
rect 5629 324 5635 816
rect 5645 704 5651 716
rect 5677 584 5683 896
rect 5693 704 5699 876
rect 5821 862 5827 900
rect 5709 764 5715 836
rect 5725 724 5731 736
rect 5837 702 5843 736
rect 5709 684 5715 696
rect 5773 604 5779 676
rect 5805 644 5811 676
rect 5885 603 5891 916
rect 5917 784 5923 956
rect 5997 784 6003 1077
rect 5869 597 5891 603
rect 5757 464 5763 536
rect 5869 524 5875 597
rect 5949 564 5955 776
rect 5965 724 5971 736
rect 6013 724 6019 916
rect 6061 824 6067 1096
rect 6093 1084 6099 1396
rect 6029 724 6035 756
rect 6013 684 6019 716
rect 6061 704 6067 816
rect 6029 604 6035 636
rect 5949 504 5955 556
rect 5981 544 5987 596
rect 5565 304 5571 316
rect 5389 264 5395 276
rect 5389 184 5395 236
rect 5421 124 5427 296
rect 5597 284 5603 316
rect 5629 304 5635 316
rect 5437 184 5443 276
rect 5453 244 5459 276
rect 5581 264 5587 276
rect 5437 144 5443 176
rect 5533 164 5539 236
rect 5629 184 5635 256
rect 5645 184 5651 436
rect 5597 144 5603 176
rect 5133 84 5139 96
rect 1357 -17 1363 36
rect 1496 6 1502 14
rect 1510 6 1516 14
rect 1524 6 1530 14
rect 1538 6 1544 14
rect 2189 -17 2195 36
rect 2589 -17 2595 36
rect 2637 -17 2643 36
rect 2685 -17 2691 36
rect 3133 -17 3139 36
rect 4029 -17 4035 36
rect 4568 6 4574 14
rect 4582 6 4588 14
rect 4596 6 4602 14
rect 4610 6 4616 14
rect 5645 -17 5651 156
rect 5677 144 5683 256
rect 5709 184 5715 336
rect 5741 184 5747 376
rect 5869 264 5875 496
rect 5965 320 5971 358
rect 5981 304 5987 516
rect 6045 462 6051 500
rect 6045 384 6051 416
rect 6061 304 6067 676
rect 5901 184 5907 256
rect 5901 164 5907 176
rect 5933 144 5939 156
rect 6013 124 6019 296
rect 6061 264 6067 276
rect 6077 184 6083 676
rect 6125 324 6131 336
rect 6109 104 6115 156
rect 5997 44 6003 100
rect 1357 -23 1379 -17
rect 2173 -23 2195 -17
rect 2573 -23 2595 -17
rect 2621 -23 2643 -17
rect 2669 -23 2691 -17
rect 3117 -23 3139 -17
rect 4013 -23 4035 -17
rect 5629 -23 5651 -17
rect 5661 -23 5667 16
<< m3contact >>
rect 476 5536 484 5544
rect 332 5496 340 5504
rect 444 5496 452 5504
rect 28 5476 36 5484
rect 172 5476 180 5484
rect 172 5456 180 5464
rect 204 5456 212 5464
rect 284 5456 292 5464
rect 140 5336 148 5344
rect 28 5276 36 5284
rect 12 5036 20 5044
rect 12 4916 20 4924
rect 12 4316 20 4324
rect 348 5356 356 5364
rect 364 5336 372 5344
rect 428 5356 436 5364
rect 412 5336 420 5344
rect 396 5316 404 5324
rect 332 5296 340 5304
rect 1502 5606 1510 5614
rect 1516 5606 1524 5614
rect 1530 5606 1538 5614
rect 636 5536 644 5544
rect 1564 5536 1572 5544
rect 1900 5536 1908 5544
rect 572 5516 580 5524
rect 604 5516 612 5524
rect 604 5496 612 5504
rect 1244 5502 1252 5504
rect 460 5356 468 5364
rect 460 5336 468 5344
rect 572 5476 580 5484
rect 556 5336 564 5344
rect 444 5316 452 5324
rect 428 5296 436 5304
rect 556 5296 564 5304
rect 524 5276 532 5284
rect 860 5476 868 5484
rect 1244 5496 1252 5502
rect 748 5456 756 5464
rect 588 5296 596 5304
rect 652 5236 660 5244
rect 316 5216 324 5224
rect 412 5216 420 5224
rect 572 5216 580 5224
rect 268 5096 276 5104
rect 124 5076 132 5084
rect 172 5076 180 5084
rect 220 5076 228 5084
rect 60 5036 68 5044
rect 60 4856 68 4864
rect 76 4696 84 4704
rect 188 5016 196 5024
rect 156 4996 164 5004
rect 172 4916 180 4924
rect 140 4896 148 4904
rect 172 4896 180 4904
rect 204 4896 212 4904
rect 204 4856 212 4864
rect 156 4836 164 4844
rect 188 4736 196 4744
rect 92 4476 100 4484
rect 300 4916 308 4924
rect 300 4896 308 4904
rect 220 4796 228 4804
rect 268 4736 276 4744
rect 844 5336 852 5344
rect 956 5456 964 5464
rect 988 5296 996 5304
rect 892 5216 900 5224
rect 812 5136 820 5144
rect 860 5136 868 5144
rect 460 5116 468 5124
rect 540 5116 548 5124
rect 716 5116 724 5124
rect 796 5116 804 5124
rect 428 5096 436 5104
rect 524 5096 532 5104
rect 380 5076 388 5084
rect 348 4956 356 4964
rect 316 4796 324 4804
rect 236 4696 244 4704
rect 300 4696 308 4704
rect 172 4556 180 4564
rect 220 4636 228 4644
rect 220 4536 228 4544
rect 268 4536 276 4544
rect 140 4518 148 4524
rect 140 4516 148 4518
rect 124 4396 132 4404
rect 12 4296 20 4304
rect 28 4296 36 4304
rect 60 4296 68 4304
rect 108 4276 116 4284
rect 92 4236 100 4244
rect 236 4516 244 4524
rect 284 4516 292 4524
rect 252 4496 260 4504
rect 284 4496 292 4504
rect 268 4476 276 4484
rect 220 4396 228 4404
rect 252 4316 260 4324
rect 76 4136 84 4144
rect 140 4136 148 4144
rect 252 4116 260 4124
rect 60 3756 68 3764
rect 92 3756 100 3764
rect 124 3756 132 3764
rect 12 3736 20 3744
rect 60 3736 68 3744
rect 44 3716 52 3724
rect 76 3716 84 3724
rect 92 3716 100 3724
rect 28 3696 36 3704
rect 140 3736 148 3744
rect 156 3716 164 3724
rect 60 3596 68 3604
rect 92 3596 100 3604
rect 92 3576 100 3584
rect 12 3496 20 3504
rect 92 3416 100 3424
rect 204 3616 212 3624
rect 316 4676 324 4684
rect 332 4536 340 4544
rect 412 5056 420 5064
rect 476 5076 484 5084
rect 492 5056 500 5064
rect 460 4996 468 5004
rect 444 4936 452 4944
rect 492 4936 500 4944
rect 412 4896 420 4904
rect 460 4916 468 4924
rect 476 4916 484 4924
rect 556 5076 564 5084
rect 556 4976 564 4984
rect 588 4916 596 4924
rect 668 4996 676 5004
rect 652 4956 660 4964
rect 636 4936 644 4944
rect 796 5076 804 5084
rect 732 5036 740 5044
rect 620 4916 628 4924
rect 556 4896 564 4904
rect 396 4856 404 4864
rect 428 4856 436 4864
rect 524 4876 532 4884
rect 476 4836 484 4844
rect 396 4716 404 4724
rect 412 4676 420 4684
rect 380 4596 388 4604
rect 460 4576 468 4584
rect 364 4536 372 4544
rect 588 4896 596 4904
rect 652 4876 660 4884
rect 572 4816 580 4824
rect 508 4756 516 4764
rect 572 4756 580 4764
rect 588 4716 596 4724
rect 540 4696 548 4704
rect 748 5016 756 5024
rect 844 4996 852 5004
rect 876 4936 884 4944
rect 748 4896 756 4904
rect 780 4896 788 4904
rect 828 4896 836 4904
rect 844 4896 852 4904
rect 908 5036 916 5044
rect 940 5036 948 5044
rect 892 4916 900 4924
rect 732 4856 740 4864
rect 716 4836 724 4844
rect 732 4816 740 4824
rect 716 4796 724 4804
rect 716 4736 724 4744
rect 812 4876 820 4884
rect 876 4836 884 4844
rect 860 4816 868 4824
rect 860 4796 868 4804
rect 828 4776 836 4784
rect 732 4696 740 4704
rect 524 4676 532 4684
rect 572 4676 580 4684
rect 620 4656 628 4664
rect 636 4616 644 4624
rect 684 4636 692 4644
rect 540 4556 548 4564
rect 508 4536 516 4544
rect 460 4476 468 4484
rect 492 4476 500 4484
rect 444 4436 452 4444
rect 332 4316 340 4324
rect 364 4296 372 4304
rect 444 4296 452 4304
rect 332 4276 340 4284
rect 396 4276 404 4284
rect 380 4256 388 4264
rect 364 4236 372 4244
rect 316 4216 324 4224
rect 284 4156 292 4164
rect 428 4216 436 4224
rect 444 4156 452 4164
rect 492 4356 500 4364
rect 588 4496 596 4504
rect 604 4296 612 4304
rect 812 4676 820 4684
rect 700 4476 708 4484
rect 732 4476 740 4484
rect 716 4356 724 4364
rect 700 4336 708 4344
rect 508 4276 516 4284
rect 540 4276 548 4284
rect 636 4276 644 4284
rect 524 4236 532 4244
rect 476 4116 484 4124
rect 476 4096 484 4104
rect 508 4096 516 4104
rect 460 3976 468 3984
rect 364 3896 372 3904
rect 396 3896 404 3904
rect 460 3896 468 3904
rect 268 3816 276 3824
rect 332 3756 340 3764
rect 268 3736 276 3744
rect 284 3716 292 3724
rect 396 3876 404 3884
rect 476 3836 484 3844
rect 396 3816 404 3824
rect 380 3736 388 3744
rect 364 3716 372 3724
rect 428 3736 436 3744
rect 444 3736 452 3744
rect 428 3716 436 3724
rect 332 3696 340 3704
rect 348 3696 356 3704
rect 460 3696 468 3704
rect 316 3676 324 3684
rect 348 3676 356 3684
rect 284 3576 292 3584
rect 428 3616 436 3624
rect 412 3556 420 3564
rect 156 3476 164 3484
rect 236 3476 244 3484
rect 348 3476 356 3484
rect 172 3456 180 3464
rect 268 3456 276 3464
rect 140 3416 148 3424
rect 76 3396 84 3404
rect 124 3396 132 3404
rect 556 4136 564 4144
rect 556 4016 564 4024
rect 540 3916 548 3924
rect 636 4236 644 4244
rect 732 4336 740 4344
rect 732 4316 740 4324
rect 716 4156 724 4164
rect 620 4136 628 4144
rect 636 4136 644 4144
rect 588 4116 596 4124
rect 604 4116 612 4124
rect 700 4118 708 4124
rect 700 4116 708 4118
rect 716 4116 724 4124
rect 652 4036 660 4044
rect 796 4656 804 4664
rect 812 4616 820 4624
rect 780 4536 788 4544
rect 796 4536 804 4544
rect 828 4536 836 4544
rect 860 4536 868 4544
rect 796 4516 804 4524
rect 780 4456 788 4464
rect 668 3976 676 3984
rect 748 4016 756 4024
rect 668 3896 676 3904
rect 748 3896 756 3904
rect 556 3876 564 3884
rect 700 3756 708 3764
rect 492 3736 500 3744
rect 556 3736 564 3744
rect 572 3736 580 3744
rect 492 3716 500 3724
rect 588 3696 596 3704
rect 732 3696 740 3704
rect 668 3656 676 3664
rect 924 4996 932 5004
rect 1004 5276 1012 5284
rect 1116 5476 1124 5484
rect 1212 5476 1220 5484
rect 1868 5516 1876 5524
rect 1932 5516 1940 5524
rect 1676 5496 1684 5504
rect 1772 5496 1780 5504
rect 1868 5496 1876 5504
rect 1900 5496 1908 5504
rect 1756 5476 1758 5484
rect 1758 5476 1764 5484
rect 1452 5456 1460 5464
rect 1100 5436 1108 5444
rect 1180 5436 1188 5444
rect 1036 5356 1044 5364
rect 1084 5356 1092 5364
rect 1052 5336 1060 5344
rect 1052 5316 1060 5324
rect 1180 5416 1188 5424
rect 1164 5396 1172 5404
rect 1116 5336 1124 5344
rect 1132 5316 1140 5324
rect 1372 5396 1380 5404
rect 1468 5336 1476 5344
rect 1580 5336 1588 5344
rect 1052 5216 1060 5224
rect 1020 5136 1028 5144
rect 1052 5136 1060 5144
rect 1100 5116 1108 5124
rect 1148 5116 1156 5124
rect 1404 5316 1412 5324
rect 1244 5296 1252 5304
rect 1324 5276 1332 5284
rect 1308 5116 1316 5124
rect 1212 5096 1220 5104
rect 1164 5076 1172 5084
rect 1260 5076 1268 5084
rect 1196 5056 1204 5064
rect 1004 5036 1012 5044
rect 1052 4996 1060 5004
rect 1068 4976 1076 4984
rect 1020 4936 1028 4944
rect 924 4816 932 4824
rect 1004 4896 1012 4904
rect 1036 4916 1044 4924
rect 1132 4996 1140 5004
rect 1244 5036 1252 5044
rect 1116 4936 1124 4944
rect 1308 5056 1316 5064
rect 1292 4996 1300 5004
rect 1276 4956 1284 4964
rect 1164 4916 1172 4924
rect 1036 4856 1044 4864
rect 1020 4816 1028 4824
rect 972 4776 980 4784
rect 940 4676 948 4684
rect 892 4576 900 4584
rect 828 4496 836 4504
rect 876 4476 884 4484
rect 812 4336 820 4344
rect 876 4316 884 4324
rect 956 4576 964 4584
rect 940 4456 948 4464
rect 1036 4696 1044 4704
rect 1004 4596 1012 4604
rect 1004 4516 1012 4524
rect 988 4436 996 4444
rect 940 4316 948 4324
rect 1036 4676 1044 4684
rect 1068 4616 1076 4624
rect 1052 4556 1060 4564
rect 1132 4876 1140 4884
rect 1084 4516 1092 4524
rect 1020 4496 1028 4504
rect 844 4296 852 4304
rect 892 4296 900 4304
rect 812 4136 820 4144
rect 844 4136 852 4144
rect 828 4096 836 4104
rect 860 4056 868 4064
rect 796 4016 804 4024
rect 860 3916 868 3924
rect 924 4236 932 4244
rect 908 4216 916 4224
rect 956 4196 964 4204
rect 988 4296 996 4304
rect 1004 4276 1012 4284
rect 1004 4256 1012 4264
rect 972 4176 980 4184
rect 924 4156 932 4164
rect 956 4156 964 4164
rect 940 4116 948 4124
rect 924 4056 932 4064
rect 908 4036 916 4044
rect 860 3896 868 3904
rect 780 3876 788 3884
rect 780 3796 788 3804
rect 780 3756 788 3764
rect 780 3696 788 3704
rect 780 3676 788 3684
rect 636 3636 644 3644
rect 764 3636 772 3644
rect 556 3536 564 3544
rect 428 3516 436 3524
rect 892 3836 900 3844
rect 812 3776 820 3784
rect 844 3776 852 3784
rect 828 3756 836 3764
rect 812 3716 820 3724
rect 892 3756 900 3764
rect 972 4096 980 4104
rect 956 4036 964 4044
rect 1212 4836 1220 4844
rect 1164 4796 1172 4804
rect 1116 4756 1124 4764
rect 1212 4756 1220 4764
rect 1244 4756 1252 4764
rect 1148 4736 1156 4744
rect 1196 4736 1204 4744
rect 1116 4716 1124 4724
rect 1132 4696 1140 4704
rect 1116 4656 1124 4664
rect 1276 4736 1284 4744
rect 1260 4696 1268 4704
rect 1276 4696 1284 4704
rect 1276 4656 1284 4664
rect 1180 4636 1188 4644
rect 1164 4616 1172 4624
rect 1148 4516 1156 4524
rect 1132 4496 1140 4504
rect 1148 4496 1156 4504
rect 1068 4476 1076 4484
rect 1100 4476 1108 4484
rect 1164 4476 1172 4484
rect 1356 4736 1364 4744
rect 1308 4696 1316 4704
rect 1356 4696 1364 4704
rect 1340 4656 1348 4664
rect 1212 4536 1220 4544
rect 1260 4536 1268 4544
rect 1164 4416 1172 4424
rect 1084 4336 1092 4344
rect 1068 4296 1076 4304
rect 1132 4316 1140 4324
rect 1148 4296 1156 4304
rect 1068 4276 1076 4284
rect 1100 4276 1108 4284
rect 1052 4256 1060 4264
rect 1068 4196 1076 4204
rect 1036 4176 1044 4184
rect 1180 4336 1188 4344
rect 1292 4396 1300 4404
rect 1356 4596 1364 4604
rect 1340 4416 1348 4424
rect 1340 4396 1348 4404
rect 1276 4356 1284 4364
rect 1292 4336 1300 4344
rect 1340 4296 1348 4304
rect 1244 4276 1252 4284
rect 1228 4256 1236 4264
rect 1196 4236 1204 4244
rect 1180 4216 1188 4224
rect 1260 4236 1268 4244
rect 1244 4216 1252 4224
rect 1308 4216 1316 4224
rect 1212 4156 1220 4164
rect 1292 4156 1300 4164
rect 1084 4136 1092 4144
rect 1100 4116 1108 4124
rect 1004 4096 1012 4104
rect 1036 4096 1044 4104
rect 1132 4116 1140 4124
rect 1196 4116 1204 4124
rect 1324 4136 1332 4144
rect 1388 5056 1396 5064
rect 1404 4996 1412 5004
rect 1836 5476 1844 5484
rect 1932 5416 1940 5424
rect 2156 5496 2164 5504
rect 2444 5496 2452 5504
rect 1964 5396 1972 5404
rect 2012 5376 2020 5384
rect 1884 5356 1892 5364
rect 1916 5336 1924 5344
rect 1612 5316 1620 5324
rect 1724 5296 1732 5304
rect 1596 5236 1604 5244
rect 1676 5236 1684 5244
rect 1502 5206 1510 5214
rect 1516 5206 1524 5214
rect 1530 5206 1538 5214
rect 1532 5136 1540 5144
rect 1500 5036 1508 5044
rect 1500 4936 1508 4944
rect 1708 5096 1716 5104
rect 1836 5096 1844 5104
rect 1644 5076 1652 5084
rect 1660 5056 1668 5064
rect 1676 5056 1684 5064
rect 1692 5036 1700 5044
rect 1852 5076 1860 5084
rect 1740 5056 1748 5064
rect 1724 5016 1732 5024
rect 2268 5476 2276 5484
rect 2380 5456 2388 5464
rect 2076 5376 2084 5384
rect 3324 5496 3332 5504
rect 2620 5476 2628 5484
rect 3228 5476 3236 5484
rect 2556 5456 2564 5464
rect 2508 5436 2516 5444
rect 2204 5416 2212 5424
rect 2412 5416 2420 5424
rect 2476 5416 2484 5424
rect 2172 5356 2180 5364
rect 2188 5356 2196 5364
rect 2268 5396 2276 5404
rect 2428 5356 2436 5364
rect 2140 5336 2148 5344
rect 2204 5336 2212 5344
rect 2428 5336 2436 5344
rect 2460 5336 2468 5344
rect 1996 5316 2004 5324
rect 2044 5316 2052 5324
rect 1916 4996 1924 5004
rect 1964 4996 1972 5004
rect 1820 4976 1828 4984
rect 1772 4936 1780 4944
rect 1468 4916 1476 4924
rect 1596 4916 1604 4924
rect 1452 4776 1460 4784
rect 1502 4806 1510 4814
rect 1516 4806 1524 4814
rect 1530 4806 1538 4814
rect 1548 4716 1556 4724
rect 1692 4716 1700 4724
rect 1436 4636 1444 4644
rect 1404 4616 1412 4624
rect 1388 4596 1396 4604
rect 1404 4556 1412 4564
rect 1436 4596 1444 4604
rect 1484 4676 1492 4684
rect 1468 4576 1476 4584
rect 1452 4536 1460 4544
rect 1660 4696 1668 4704
rect 1724 4696 1732 4704
rect 1740 4696 1748 4704
rect 1532 4656 1540 4664
rect 1484 4516 1492 4524
rect 1388 4496 1396 4504
rect 1420 4496 1428 4504
rect 1484 4496 1492 4504
rect 1372 4456 1380 4464
rect 1372 4356 1380 4364
rect 1404 4356 1412 4364
rect 1628 4676 1636 4684
rect 1596 4576 1604 4584
rect 1548 4436 1556 4444
rect 1502 4406 1510 4414
rect 1516 4406 1524 4414
rect 1530 4406 1538 4414
rect 1452 4316 1460 4324
rect 1468 4316 1476 4324
rect 1564 4316 1572 4324
rect 1580 4316 1588 4324
rect 1420 4176 1428 4184
rect 1388 4136 1396 4144
rect 1452 4136 1460 4144
rect 1564 4296 1572 4304
rect 1564 4276 1572 4284
rect 1580 4276 1588 4284
rect 1500 4196 1508 4204
rect 1500 4176 1508 4184
rect 1276 4036 1284 4044
rect 1324 3936 1332 3944
rect 972 3916 980 3924
rect 1068 3916 1076 3924
rect 1116 3916 1124 3924
rect 1308 3916 1316 3924
rect 1372 3916 1380 3924
rect 1084 3896 1092 3904
rect 1180 3896 1188 3904
rect 1196 3896 1204 3904
rect 1388 3896 1396 3904
rect 988 3876 996 3884
rect 1148 3876 1156 3884
rect 940 3796 948 3804
rect 924 3776 932 3784
rect 892 3696 900 3704
rect 908 3656 916 3664
rect 908 3636 916 3644
rect 812 3516 820 3524
rect 908 3516 916 3524
rect 940 3536 948 3544
rect 972 3536 980 3544
rect 508 3476 516 3484
rect 556 3476 564 3484
rect 860 3476 868 3484
rect 524 3456 532 3464
rect 508 3356 516 3364
rect 412 3316 420 3324
rect 124 3236 132 3244
rect 172 3236 180 3244
rect 316 3236 324 3244
rect 12 3196 20 3204
rect 140 2936 148 2944
rect 172 2936 180 2944
rect 140 2676 148 2684
rect 284 3076 292 3084
rect 380 3196 388 3204
rect 444 3176 452 3184
rect 476 3176 484 3184
rect 556 3356 564 3364
rect 540 3316 548 3324
rect 524 3216 532 3224
rect 572 3096 580 3104
rect 492 3076 500 3084
rect 316 3056 324 3064
rect 604 3416 612 3424
rect 812 3416 820 3424
rect 1116 3856 1124 3864
rect 1084 3816 1092 3824
rect 1116 3796 1124 3804
rect 1196 3856 1204 3864
rect 1212 3856 1220 3864
rect 1276 3836 1284 3844
rect 1212 3816 1220 3824
rect 1212 3736 1220 3744
rect 1244 3736 1252 3744
rect 1036 3716 1044 3724
rect 1020 3696 1028 3704
rect 1004 3676 1012 3684
rect 1212 3716 1220 3724
rect 1228 3716 1236 3724
rect 1196 3576 1204 3584
rect 1052 3516 1060 3524
rect 1132 3516 1140 3524
rect 1196 3516 1204 3524
rect 1036 3496 1044 3504
rect 924 3476 932 3484
rect 988 3476 996 3484
rect 1132 3476 1140 3484
rect 940 3416 948 3424
rect 908 3396 916 3404
rect 684 3356 692 3364
rect 764 3356 772 3364
rect 604 3216 612 3224
rect 284 2956 292 2964
rect 572 2956 580 2964
rect 588 2956 596 2964
rect 316 2936 324 2944
rect 796 3336 804 3344
rect 972 3336 980 3344
rect 956 3316 964 3324
rect 796 3116 804 3124
rect 1084 3356 1092 3364
rect 1228 3516 1236 3524
rect 1340 3836 1348 3844
rect 1388 3836 1396 3844
rect 1324 3796 1332 3804
rect 1292 3756 1300 3764
rect 1372 3736 1380 3744
rect 1420 3776 1428 3784
rect 1420 3756 1428 3764
rect 1372 3716 1380 3724
rect 1420 3716 1428 3724
rect 1260 3636 1268 3644
rect 1260 3516 1268 3524
rect 1388 3696 1396 3704
rect 1324 3676 1332 3684
rect 1452 3676 1460 3684
rect 1308 3656 1316 3664
rect 1436 3656 1444 3664
rect 1276 3496 1284 3504
rect 1196 3416 1204 3424
rect 1244 3416 1252 3424
rect 1420 3636 1428 3644
rect 1340 3536 1348 3544
rect 1564 4156 1572 4164
rect 1564 4116 1572 4124
rect 1628 4516 1636 4524
rect 1612 4496 1620 4504
rect 1628 4496 1636 4504
rect 1660 4636 1668 4644
rect 1676 4616 1684 4624
rect 1676 4556 1684 4564
rect 1724 4676 1732 4684
rect 1788 4756 1796 4764
rect 1772 4696 1780 4704
rect 2012 4956 2020 4964
rect 1948 4936 1956 4944
rect 1836 4916 1844 4924
rect 1852 4716 1860 4724
rect 1772 4676 1780 4684
rect 1804 4656 1812 4664
rect 1836 4656 1844 4664
rect 2044 4696 2052 4704
rect 2268 5236 2276 5244
rect 2332 5236 2340 5244
rect 3452 5496 3460 5504
rect 2700 5396 2708 5404
rect 2924 5416 2932 5424
rect 2988 5416 2996 5424
rect 2652 5356 2660 5364
rect 2732 5356 2740 5364
rect 2764 5356 2772 5364
rect 2892 5356 2900 5364
rect 2956 5356 2964 5364
rect 2988 5356 2996 5364
rect 2364 5096 2372 5104
rect 2412 5096 2420 5104
rect 2396 5076 2404 5084
rect 2380 5056 2388 5064
rect 2412 5056 2420 5064
rect 2252 5036 2260 5044
rect 2316 5036 2324 5044
rect 2364 5036 2372 5044
rect 2236 5016 2244 5024
rect 2156 4996 2164 5004
rect 2268 4956 2276 4964
rect 2140 4936 2148 4944
rect 2124 4836 2132 4844
rect 2252 4836 2260 4844
rect 2108 4716 2116 4724
rect 2236 4716 2244 4724
rect 2188 4696 2196 4704
rect 1964 4676 1972 4684
rect 2124 4676 2132 4684
rect 1836 4596 1844 4604
rect 1852 4596 1860 4604
rect 1964 4596 1972 4604
rect 1756 4556 1764 4564
rect 1772 4536 1780 4544
rect 1852 4536 1860 4544
rect 1932 4536 1940 4544
rect 1692 4516 1700 4524
rect 1692 4496 1700 4504
rect 1660 4476 1668 4484
rect 1644 4456 1652 4464
rect 1676 4376 1684 4384
rect 1676 4336 1684 4344
rect 1676 4316 1684 4324
rect 1756 4516 1764 4524
rect 1804 4516 1812 4524
rect 1884 4516 1892 4524
rect 1836 4496 1844 4504
rect 1724 4296 1732 4304
rect 1708 4276 1716 4284
rect 1692 4256 1700 4264
rect 1644 4216 1652 4224
rect 1612 4156 1620 4164
rect 1484 4096 1492 4104
rect 1502 4006 1510 4014
rect 1516 4006 1524 4014
rect 1530 4006 1538 4014
rect 1612 4096 1620 4104
rect 1612 4076 1620 4084
rect 1580 4056 1588 4064
rect 1676 4136 1684 4144
rect 1692 4116 1700 4124
rect 1676 4096 1684 4104
rect 1724 4256 1732 4264
rect 1980 4556 1988 4564
rect 2076 4636 2084 4644
rect 1980 4516 1988 4524
rect 2028 4516 2036 4524
rect 1996 4476 2004 4484
rect 1948 4336 1956 4344
rect 2012 4336 2020 4344
rect 2076 4576 2084 4584
rect 2108 4496 2116 4504
rect 2092 4476 2100 4484
rect 2220 4676 2228 4684
rect 2140 4636 2148 4644
rect 2380 4716 2388 4724
rect 2460 5076 2468 5084
rect 2476 5076 2484 5084
rect 2476 5056 2484 5064
rect 2524 5056 2532 5064
rect 2444 4976 2452 4984
rect 2348 4676 2356 4684
rect 2284 4656 2292 4664
rect 2300 4636 2308 4644
rect 2220 4536 2228 4544
rect 2284 4536 2292 4544
rect 2428 4676 2436 4684
rect 2412 4656 2420 4664
rect 2364 4536 2372 4544
rect 2396 4536 2404 4544
rect 2140 4376 2148 4384
rect 2076 4336 2084 4344
rect 2124 4336 2132 4344
rect 2252 4356 2260 4364
rect 2204 4336 2212 4344
rect 2332 4436 2340 4444
rect 2156 4316 2164 4324
rect 2188 4316 2196 4324
rect 2300 4316 2308 4324
rect 2108 4296 2116 4304
rect 2236 4296 2244 4304
rect 2268 4296 2276 4304
rect 2028 4276 2036 4284
rect 1820 4256 1828 4264
rect 1804 4236 1812 4244
rect 2188 4276 2196 4284
rect 2252 4256 2260 4264
rect 2172 4236 2180 4244
rect 2044 4216 2052 4224
rect 1932 4196 1940 4204
rect 1980 4196 1988 4204
rect 2140 4196 2148 4204
rect 1740 4156 1748 4164
rect 2476 5016 2484 5024
rect 2508 4956 2516 4964
rect 2460 4876 2468 4884
rect 2508 4716 2516 4724
rect 2460 4656 2468 4664
rect 2444 4636 2452 4644
rect 2476 4636 2484 4644
rect 2620 5076 2628 5084
rect 3038 5406 3046 5414
rect 3052 5406 3060 5414
rect 3066 5406 3074 5414
rect 3020 5376 3028 5384
rect 3436 5476 3444 5484
rect 3420 5396 3428 5404
rect 3100 5356 3108 5364
rect 3196 5356 3204 5364
rect 3324 5356 3332 5364
rect 3356 5356 3364 5364
rect 3180 5296 3188 5304
rect 2732 5216 2740 5224
rect 2812 5216 2820 5224
rect 3004 5216 3012 5224
rect 3452 5316 3460 5324
rect 3500 5476 3508 5484
rect 3516 5456 3524 5464
rect 3532 5396 3540 5404
rect 3500 5356 3508 5364
rect 3500 5336 3508 5344
rect 3612 5516 3620 5524
rect 3644 5516 3652 5524
rect 3628 5496 3636 5504
rect 3644 5476 3652 5484
rect 3628 5456 3636 5464
rect 3580 5396 3588 5404
rect 3580 5336 3588 5344
rect 3660 5456 3668 5464
rect 3708 5376 3716 5384
rect 4574 5606 4582 5614
rect 4588 5606 4596 5614
rect 4602 5606 4610 5614
rect 4060 5536 4068 5544
rect 4252 5536 4260 5544
rect 4204 5516 4212 5524
rect 3900 5496 3908 5504
rect 3996 5496 4004 5504
rect 4124 5496 4132 5504
rect 3772 5396 3780 5404
rect 3676 5356 3684 5364
rect 3596 5296 3604 5304
rect 3564 5276 3572 5284
rect 3292 5216 3300 5224
rect 3468 5216 3476 5224
rect 3660 5216 3668 5224
rect 3196 5116 3204 5124
rect 3356 5116 3364 5124
rect 2796 5096 2804 5104
rect 3132 5096 3140 5104
rect 3164 5096 3166 5104
rect 3166 5096 3172 5104
rect 2652 5056 2660 5064
rect 2636 4936 2644 4944
rect 2780 4936 2788 4944
rect 2812 4976 2820 4984
rect 2812 4936 2820 4944
rect 2860 4936 2868 4944
rect 2572 4716 2580 4724
rect 2540 4696 2548 4704
rect 2524 4656 2532 4664
rect 2460 4596 2468 4604
rect 2508 4596 2516 4604
rect 2700 4656 2708 4664
rect 2780 4636 2788 4644
rect 2572 4516 2580 4524
rect 2748 4556 2756 4564
rect 2764 4536 2772 4544
rect 2812 4556 2820 4564
rect 2844 4876 2852 4884
rect 2844 4856 2852 4864
rect 2828 4536 2836 4544
rect 2732 4516 2740 4524
rect 2460 4476 2468 4484
rect 2652 4476 2660 4484
rect 2428 4376 2436 4384
rect 2412 4316 2420 4324
rect 2380 4276 2388 4284
rect 2316 4256 2324 4264
rect 2300 4236 2308 4244
rect 2332 4236 2340 4244
rect 1756 4136 1764 4144
rect 1948 4136 1956 4144
rect 2156 4136 2164 4144
rect 2300 4136 2308 4144
rect 2348 4136 2356 4144
rect 2380 4136 2388 4144
rect 1804 4116 1812 4124
rect 2348 4116 2356 4124
rect 1708 4076 1716 4084
rect 1628 4056 1636 4064
rect 1772 3996 1780 4004
rect 1868 3996 1876 4004
rect 1676 3976 1684 3984
rect 2236 4096 2244 4104
rect 2396 4116 2404 4124
rect 2492 4416 2500 4424
rect 2428 4296 2436 4304
rect 2476 4236 2484 4244
rect 2476 4136 2484 4144
rect 2428 4096 2436 4104
rect 2188 4076 2196 4084
rect 2332 4076 2340 4084
rect 2028 4016 2036 4024
rect 2220 3996 2228 4004
rect 2044 3976 2052 3984
rect 2092 3936 2100 3944
rect 2124 3916 2132 3924
rect 2780 4376 2788 4384
rect 2780 4356 2788 4364
rect 2684 4336 2692 4344
rect 2716 4336 2724 4344
rect 2556 4316 2564 4324
rect 2764 4316 2772 4324
rect 2540 4296 2548 4304
rect 2604 4296 2612 4304
rect 2652 4296 2660 4304
rect 2748 4296 2756 4304
rect 2572 4276 2580 4284
rect 2668 4276 2676 4284
rect 2588 4256 2596 4264
rect 2524 4236 2532 4244
rect 2540 4236 2548 4244
rect 2588 4116 2596 4124
rect 2732 4276 2740 4284
rect 2700 4236 2708 4244
rect 2620 4156 2628 4164
rect 2668 4156 2676 4164
rect 2892 5076 2900 5084
rect 2972 5076 2980 5084
rect 3292 5096 3300 5104
rect 3276 5076 3284 5084
rect 3004 5056 3012 5064
rect 3196 5056 3204 5064
rect 3148 5016 3156 5024
rect 3038 5006 3046 5014
rect 3052 5006 3060 5014
rect 3066 5006 3074 5014
rect 2940 4976 2948 4984
rect 3020 4976 3028 4984
rect 2908 4936 2916 4944
rect 2924 4856 2932 4864
rect 2892 4736 2900 4744
rect 2924 4736 2932 4744
rect 2876 4716 2884 4724
rect 2956 4956 2964 4964
rect 2972 4936 2980 4944
rect 2988 4916 2996 4924
rect 3868 5356 3876 5364
rect 3996 5356 4004 5364
rect 3820 5336 3828 5344
rect 4028 5336 4036 5344
rect 4172 5456 4180 5464
rect 4444 5516 4452 5524
rect 4636 5516 4644 5524
rect 4876 5516 4884 5524
rect 4940 5516 4948 5524
rect 5180 5516 5188 5524
rect 5212 5516 5220 5524
rect 4316 5502 4324 5504
rect 4316 5496 4324 5502
rect 4412 5496 4420 5504
rect 4300 5456 4308 5464
rect 4172 5356 4180 5364
rect 4188 5336 4196 5344
rect 3916 5316 3924 5324
rect 3724 5296 3732 5304
rect 3804 5296 3812 5304
rect 3708 5276 3716 5284
rect 3836 5276 3844 5284
rect 4172 5276 4180 5284
rect 4124 5236 4132 5244
rect 3692 5216 3700 5224
rect 4060 5216 4068 5224
rect 3388 5102 3396 5104
rect 3388 5096 3396 5102
rect 3644 5096 3652 5104
rect 3324 5076 3332 5084
rect 3532 5076 3540 5084
rect 3356 5056 3364 5064
rect 3196 4976 3204 4984
rect 3308 4976 3316 4984
rect 3148 4956 3156 4964
rect 3196 4956 3204 4964
rect 3244 4956 3252 4964
rect 3116 4916 3124 4924
rect 3260 4916 3268 4924
rect 2956 4896 2964 4904
rect 3100 4896 3108 4904
rect 3004 4876 3012 4884
rect 2988 4816 2996 4824
rect 3164 4756 3172 4764
rect 2860 4636 2868 4644
rect 2860 4556 2868 4564
rect 2956 4556 2964 4564
rect 2860 4536 2868 4544
rect 2924 4536 2932 4544
rect 2812 4296 2820 4304
rect 2844 4296 2852 4304
rect 2796 4176 2804 4184
rect 2780 4156 2788 4164
rect 2828 4216 2836 4224
rect 2828 4176 2836 4184
rect 2636 4136 2644 4144
rect 2652 4116 2660 4124
rect 2780 4116 2788 4124
rect 2796 4116 2804 4124
rect 2844 4156 2852 4164
rect 3036 4636 3044 4644
rect 3038 4606 3046 4614
rect 3052 4606 3060 4614
rect 3066 4606 3074 4614
rect 3292 4876 3300 4884
rect 3228 4856 3236 4864
rect 3340 4936 3348 4944
rect 3548 5036 3556 5044
rect 3420 4996 3428 5004
rect 3516 4996 3524 5004
rect 3324 4916 3332 4924
rect 3356 4916 3364 4924
rect 3404 4916 3412 4924
rect 3308 4836 3316 4844
rect 3276 4736 3284 4744
rect 3292 4716 3300 4724
rect 3580 4956 3588 4964
rect 3932 5136 3940 5144
rect 4092 5136 4100 5144
rect 3468 4936 3476 4944
rect 3692 4936 3700 4944
rect 3452 4916 3460 4924
rect 3420 4896 3428 4904
rect 3372 4856 3380 4864
rect 3356 4836 3364 4844
rect 3308 4696 3316 4704
rect 3276 4676 3284 4684
rect 3324 4676 3332 4684
rect 3180 4596 3188 4604
rect 2972 4456 2980 4464
rect 2956 4436 2964 4444
rect 3052 4436 3060 4444
rect 2876 4316 2884 4324
rect 2972 4396 2980 4404
rect 2940 4196 2948 4204
rect 2892 4156 2900 4164
rect 2860 4116 2868 4124
rect 2780 4096 2788 4104
rect 2828 4096 2836 4104
rect 2572 4036 2580 4044
rect 2636 4036 2644 4044
rect 2460 3936 2468 3944
rect 2492 3936 2500 3944
rect 2540 3936 2548 3944
rect 1980 3896 1988 3904
rect 1564 3876 1572 3884
rect 1660 3856 1668 3864
rect 1836 3856 1844 3864
rect 1484 3776 1492 3784
rect 1724 3836 1732 3844
rect 1724 3756 1732 3764
rect 1900 3756 1908 3764
rect 1612 3736 1620 3744
rect 1868 3736 1876 3744
rect 1532 3716 1540 3724
rect 1516 3636 1524 3644
rect 1502 3606 1510 3614
rect 1516 3606 1524 3614
rect 1530 3606 1538 3614
rect 1596 3718 1604 3724
rect 1596 3716 1604 3718
rect 1532 3576 1540 3584
rect 1564 3576 1572 3584
rect 2076 3856 2084 3864
rect 2012 3836 2020 3844
rect 2044 3736 2052 3744
rect 2524 3916 2532 3924
rect 2172 3896 2180 3904
rect 2524 3896 2532 3904
rect 2636 3896 2644 3904
rect 2108 3876 2116 3884
rect 2268 3876 2276 3884
rect 2140 3856 2148 3864
rect 2284 3816 2292 3824
rect 2188 3776 2196 3784
rect 2268 3776 2276 3784
rect 2124 3736 2132 3744
rect 2204 3736 2212 3744
rect 2268 3736 2276 3744
rect 2316 3796 2324 3804
rect 2492 3796 2500 3804
rect 2508 3796 2516 3804
rect 2572 3816 2580 3824
rect 2300 3756 2308 3764
rect 2188 3716 2196 3724
rect 2284 3716 2292 3724
rect 2060 3696 2068 3704
rect 2124 3696 2132 3704
rect 1980 3616 1988 3624
rect 2028 3616 2036 3624
rect 1916 3596 1924 3604
rect 1468 3536 1476 3544
rect 1612 3536 1620 3544
rect 1324 3496 1332 3504
rect 1308 3476 1316 3484
rect 1292 3436 1300 3444
rect 1356 3436 1364 3444
rect 1340 3356 1348 3364
rect 1052 3316 1060 3324
rect 1276 3316 1284 3324
rect 1308 3318 1316 3324
rect 1308 3316 1316 3318
rect 1036 3216 1044 3224
rect 1580 3496 1588 3504
rect 1708 3496 1716 3504
rect 1452 3396 1460 3404
rect 1532 3356 1540 3364
rect 1502 3206 1510 3214
rect 1516 3206 1524 3214
rect 1530 3206 1538 3214
rect 1420 3196 1428 3204
rect 1020 3176 1028 3184
rect 1100 3176 1108 3184
rect 1180 3116 1188 3124
rect 1372 3116 1380 3124
rect 1692 3416 1700 3424
rect 2188 3616 2196 3624
rect 2108 3596 2116 3604
rect 2108 3576 2116 3584
rect 2220 3616 2228 3624
rect 2204 3576 2212 3584
rect 2028 3496 2036 3504
rect 2124 3496 2132 3504
rect 1740 3436 1748 3444
rect 1740 3416 1748 3424
rect 1948 3416 1956 3424
rect 2108 3416 2116 3424
rect 1724 3396 1732 3404
rect 1708 3356 1716 3364
rect 1964 3396 1972 3404
rect 1836 3316 1844 3324
rect 1916 3316 1924 3324
rect 1612 3176 1620 3184
rect 1692 3116 1700 3124
rect 1884 3296 1892 3304
rect 2076 3236 2084 3244
rect 2284 3496 2292 3504
rect 2268 3476 2276 3484
rect 2300 3476 2308 3484
rect 2268 3416 2276 3424
rect 2204 3316 2212 3324
rect 2348 3596 2356 3604
rect 2332 3496 2340 3504
rect 2380 3496 2388 3504
rect 2476 3476 2484 3484
rect 2604 3736 2612 3744
rect 2828 3976 2836 3984
rect 3068 4276 3076 4284
rect 3164 4536 3172 4544
rect 3356 4636 3364 4644
rect 3404 4616 3412 4624
rect 3452 4876 3460 4884
rect 3436 4836 3444 4844
rect 3516 4916 3524 4924
rect 3452 4676 3460 4684
rect 3420 4556 3428 4564
rect 3436 4518 3444 4524
rect 3436 4516 3444 4518
rect 3308 4496 3316 4504
rect 3564 4896 3572 4904
rect 3548 4876 3556 4884
rect 3564 4796 3572 4804
rect 3548 4756 3556 4764
rect 3548 4736 3556 4744
rect 3500 4716 3508 4724
rect 3564 4696 3572 4704
rect 3484 4636 3492 4644
rect 3532 4616 3540 4624
rect 3500 4556 3508 4564
rect 3516 4476 3524 4484
rect 3484 4436 3492 4444
rect 3468 4356 3476 4364
rect 3468 4316 3476 4324
rect 3596 4916 3604 4924
rect 3644 4876 3652 4884
rect 3660 4776 3668 4784
rect 3644 4756 3652 4764
rect 3612 4736 3620 4744
rect 3644 4716 3652 4724
rect 3756 5116 3764 5124
rect 3788 5116 3796 5124
rect 3980 5116 3988 5124
rect 4108 5116 4116 5124
rect 3740 4916 3748 4924
rect 3724 4836 3732 4844
rect 3708 4796 3716 4804
rect 3676 4736 3684 4744
rect 3900 5096 3908 5104
rect 3916 5096 3924 5104
rect 3964 5096 3972 5104
rect 3788 5036 3796 5044
rect 3964 5076 3972 5084
rect 3836 5016 3844 5024
rect 3836 4976 3844 4984
rect 3916 5016 3924 5024
rect 3868 4956 3876 4964
rect 3932 4996 3940 5004
rect 3932 4956 3940 4964
rect 3964 4936 3972 4944
rect 3788 4896 3796 4904
rect 3868 4896 3876 4904
rect 3772 4876 3780 4884
rect 3756 4776 3764 4784
rect 3724 4716 3732 4724
rect 3596 4696 3604 4704
rect 3644 4656 3652 4664
rect 3644 4556 3652 4564
rect 3612 4536 3620 4544
rect 3500 4376 3508 4384
rect 3564 4376 3572 4384
rect 3564 4356 3572 4364
rect 3548 4316 3556 4324
rect 3356 4296 3364 4304
rect 3548 4276 3556 4284
rect 3036 4256 3044 4264
rect 3132 4256 3140 4264
rect 3164 4256 3172 4264
rect 3038 4206 3046 4214
rect 3052 4206 3060 4214
rect 3066 4206 3074 4214
rect 2956 4156 2964 4164
rect 3036 4156 3044 4164
rect 2988 4136 2996 4144
rect 3132 4136 3140 4144
rect 3004 4116 3012 4124
rect 3164 4116 3172 4124
rect 2908 4076 2916 4084
rect 2972 3976 2980 3984
rect 2812 3856 2820 3864
rect 2844 3816 2852 3824
rect 2812 3796 2820 3804
rect 2812 3776 2820 3784
rect 2700 3736 2708 3744
rect 2748 3736 2756 3744
rect 2636 3716 2644 3724
rect 2668 3716 2676 3724
rect 2700 3696 2708 3704
rect 2668 3576 2676 3584
rect 2588 3516 2596 3524
rect 2732 3676 2740 3684
rect 2860 3796 2868 3804
rect 3420 4156 3428 4164
rect 3372 4116 3380 4124
rect 3548 4136 3556 4144
rect 3628 4516 3636 4524
rect 3804 4876 3812 4884
rect 3916 4796 3924 4804
rect 3852 4756 3860 4764
rect 3932 4756 3940 4764
rect 4012 4916 4020 4924
rect 3996 4896 4004 4904
rect 4156 5096 4164 5104
rect 4140 5076 4148 5084
rect 4044 5016 4052 5024
rect 4348 5436 4356 5444
rect 4380 5376 4388 5384
rect 4348 5336 4356 5344
rect 4380 5336 4388 5344
rect 4332 5316 4340 5324
rect 4300 5216 4308 5224
rect 4316 5196 4324 5204
rect 4236 5076 4244 5084
rect 4220 5036 4228 5044
rect 4220 5016 4228 5024
rect 4188 4956 4196 4964
rect 4204 4956 4212 4964
rect 4092 4916 4100 4924
rect 4060 4876 4068 4884
rect 4060 4836 4068 4844
rect 4076 4776 4084 4784
rect 4028 4736 4036 4744
rect 3740 4696 3748 4704
rect 3788 4696 3796 4704
rect 3756 4596 3764 4604
rect 3724 4576 3732 4584
rect 3692 4536 3700 4544
rect 3772 4576 3780 4584
rect 3676 4516 3684 4524
rect 3676 4496 3684 4504
rect 3756 4436 3764 4444
rect 3724 4376 3732 4384
rect 3676 4356 3684 4364
rect 3644 4316 3652 4324
rect 3612 4296 3620 4304
rect 3884 4676 3892 4684
rect 3932 4636 3940 4644
rect 3820 4536 3828 4544
rect 3868 4536 3876 4544
rect 3820 4496 3828 4504
rect 3820 4356 3828 4364
rect 3692 4276 3700 4284
rect 3644 4196 3652 4204
rect 3676 4196 3684 4204
rect 3580 4176 3588 4184
rect 3660 4176 3668 4184
rect 3612 4156 3620 4164
rect 3644 4156 3652 4164
rect 3804 4276 3812 4284
rect 3772 4196 3780 4204
rect 3740 4156 3748 4164
rect 3708 4136 3716 4144
rect 3724 4136 3732 4144
rect 3564 4116 3572 4124
rect 3532 4096 3540 4104
rect 3596 4096 3604 4104
rect 3324 4076 3332 4084
rect 3260 3996 3268 4004
rect 3372 3996 3380 4004
rect 3292 3976 3300 3984
rect 3420 3976 3428 3984
rect 3038 3806 3046 3814
rect 3052 3806 3060 3814
rect 3066 3806 3074 3814
rect 2892 3736 2900 3744
rect 3212 3856 3220 3864
rect 3212 3836 3220 3844
rect 3132 3816 3140 3824
rect 3180 3816 3188 3824
rect 3724 4116 3732 4124
rect 3756 4116 3764 4124
rect 3820 4176 3828 4184
rect 3852 4436 3860 4444
rect 3804 4156 3812 4164
rect 3900 4536 3908 4544
rect 3900 4496 3908 4504
rect 4044 4716 4052 4724
rect 3996 4676 4004 4684
rect 3980 4656 3988 4664
rect 4044 4656 4052 4664
rect 3964 4616 3972 4624
rect 3964 4596 3972 4604
rect 3996 4536 4004 4544
rect 4012 4496 4020 4504
rect 4060 4336 4068 4344
rect 3980 4316 3988 4324
rect 4092 4756 4100 4764
rect 4140 4736 4148 4744
rect 4108 4716 4116 4724
rect 4108 4616 4116 4624
rect 4108 4556 4116 4564
rect 4124 4556 4132 4564
rect 4108 4516 4116 4524
rect 4284 5076 4292 5084
rect 4380 5296 4388 5304
rect 4572 5476 4580 5484
rect 4492 5456 4500 5464
rect 4556 5456 4564 5464
rect 4508 5396 4516 5404
rect 4508 5376 4516 5384
rect 4556 5356 4564 5364
rect 4476 5336 4484 5344
rect 4524 5316 4532 5324
rect 4540 5316 4548 5324
rect 4396 5276 4404 5284
rect 4444 5276 4452 5284
rect 4524 5276 4532 5284
rect 4524 5256 4532 5264
rect 4380 5196 4388 5204
rect 4364 5116 4372 5124
rect 4348 5096 4356 5104
rect 4364 5076 4372 5084
rect 4348 5056 4356 5064
rect 4252 4836 4260 4844
rect 4268 4836 4276 4844
rect 4268 4796 4276 4804
rect 4204 4656 4212 4664
rect 4156 4616 4164 4624
rect 4156 4536 4164 4544
rect 4220 4536 4228 4544
rect 4140 4516 4148 4524
rect 4204 4516 4212 4524
rect 4300 4876 4308 4884
rect 4300 4856 4308 4864
rect 4300 4796 4308 4804
rect 4332 4976 4340 4984
rect 4588 5316 4596 5324
rect 4620 5296 4628 5304
rect 4572 5276 4580 5284
rect 4574 5206 4582 5214
rect 4588 5206 4596 5214
rect 4602 5206 4610 5214
rect 4412 5096 4420 5104
rect 4396 5076 4404 5084
rect 4332 4796 4340 4804
rect 4316 4736 4324 4744
rect 4348 4756 4356 4764
rect 4380 4756 4388 4764
rect 4540 5076 4548 5084
rect 4492 5036 4500 5044
rect 4476 4976 4484 4984
rect 4476 4956 4484 4964
rect 4444 4916 4452 4924
rect 4412 4736 4420 4744
rect 4460 4876 4468 4884
rect 4476 4796 4484 4804
rect 4748 5502 4756 5504
rect 4748 5496 4756 5502
rect 4780 5496 4788 5504
rect 4860 5496 4868 5504
rect 5052 5496 5060 5504
rect 4684 5436 4692 5444
rect 4748 5376 4756 5384
rect 4668 5356 4676 5364
rect 4812 5376 4820 5384
rect 4652 5336 4660 5344
rect 4716 5336 4724 5344
rect 4860 5436 4868 5444
rect 4876 5376 4884 5384
rect 4924 5436 4932 5444
rect 5132 5436 5140 5444
rect 5020 5416 5028 5424
rect 5100 5416 5108 5424
rect 4924 5356 4932 5364
rect 4988 5356 4996 5364
rect 5180 5476 5188 5484
rect 4844 5336 4852 5344
rect 4908 5336 4916 5344
rect 4972 5336 4980 5344
rect 5148 5336 5156 5344
rect 5324 5516 5332 5524
rect 5276 5496 5284 5504
rect 5228 5456 5236 5464
rect 5324 5496 5332 5504
rect 5292 5476 5300 5484
rect 5276 5436 5284 5444
rect 5324 5416 5332 5424
rect 5260 5356 5268 5364
rect 4748 5316 4756 5324
rect 4828 5316 4836 5324
rect 4924 5316 4932 5324
rect 5052 5318 5060 5324
rect 5052 5316 5060 5318
rect 5196 5316 5204 5324
rect 4652 5216 4660 5224
rect 4652 5116 4660 5124
rect 4732 5256 4740 5264
rect 4812 5296 4820 5304
rect 4876 5276 4884 5284
rect 4828 5156 4836 5164
rect 4844 5136 4852 5144
rect 4684 5116 4692 5124
rect 4668 5096 4676 5104
rect 4764 5096 4772 5104
rect 4636 5056 4644 5064
rect 4716 5056 4724 5064
rect 4796 5056 4804 5064
rect 4700 5036 4708 5044
rect 4556 5016 4564 5024
rect 4524 4976 4532 4984
rect 4540 4956 4548 4964
rect 4492 4776 4500 4784
rect 4476 4756 4484 4764
rect 4460 4736 4468 4744
rect 4428 4716 4436 4724
rect 4396 4696 4404 4704
rect 4316 4676 4324 4684
rect 4380 4676 4388 4684
rect 4444 4696 4452 4704
rect 4460 4676 4468 4684
rect 4300 4616 4308 4624
rect 4348 4616 4356 4624
rect 4412 4616 4420 4624
rect 4284 4536 4292 4544
rect 4092 4436 4100 4444
rect 4140 4376 4148 4384
rect 4124 4336 4132 4344
rect 3932 4296 3940 4304
rect 4012 4296 4020 4304
rect 4028 4296 4036 4304
rect 4108 4296 4116 4304
rect 3884 4276 3892 4284
rect 3980 4276 3988 4284
rect 3884 4236 3892 4244
rect 3964 4216 3972 4224
rect 3900 4156 3908 4164
rect 3916 4156 3924 4164
rect 3836 4116 3844 4124
rect 3964 4116 3972 4124
rect 3772 4096 3780 4104
rect 3708 3996 3716 4004
rect 3820 3996 3828 4004
rect 3500 3856 3508 3864
rect 3580 3856 3588 3864
rect 3612 3836 3620 3844
rect 3596 3816 3604 3824
rect 3420 3796 3428 3804
rect 3196 3756 3204 3764
rect 3372 3756 3380 3764
rect 3388 3736 3396 3744
rect 3564 3736 3572 3744
rect 3756 3796 3764 3804
rect 3116 3716 3124 3724
rect 3436 3716 3444 3724
rect 3468 3716 3476 3724
rect 3084 3696 3092 3704
rect 3100 3656 3108 3664
rect 3212 3696 3220 3704
rect 2812 3576 2820 3584
rect 2732 3556 2740 3564
rect 2364 3456 2372 3464
rect 2316 3296 2324 3304
rect 2300 3276 2308 3284
rect 2188 3256 2196 3264
rect 2108 3216 2116 3224
rect 2172 3216 2180 3224
rect 1916 3116 1924 3124
rect 2044 3116 2052 3124
rect 876 3096 884 3104
rect 1036 3096 1044 3104
rect 1292 3096 1300 3104
rect 1468 3096 1476 3104
rect 1564 3096 1572 3104
rect 716 3076 724 3084
rect 860 3076 868 3084
rect 684 3056 692 3064
rect 924 3056 932 3064
rect 860 2956 868 2964
rect 780 2936 788 2944
rect 748 2916 756 2924
rect 540 2896 548 2904
rect 588 2896 596 2904
rect 396 2836 404 2844
rect 476 2836 484 2844
rect 252 2696 260 2704
rect 284 2696 292 2704
rect 172 2656 180 2664
rect 332 2636 340 2644
rect 380 2556 388 2564
rect 12 2336 20 2344
rect 124 2336 132 2344
rect 92 2316 100 2324
rect 252 2516 260 2524
rect 220 2396 228 2404
rect 188 2356 196 2364
rect 300 2356 308 2364
rect 332 2356 340 2364
rect 156 2336 164 2344
rect 220 2316 228 2324
rect 252 2316 260 2324
rect 332 2316 340 2324
rect 44 2296 52 2304
rect 156 2296 164 2304
rect 188 2296 196 2304
rect 236 2296 244 2304
rect 268 2296 276 2304
rect 28 2276 36 2284
rect 76 2276 84 2284
rect 60 2256 68 2264
rect 188 2276 196 2284
rect 156 2156 164 2164
rect 204 2256 212 2264
rect 220 2256 228 2264
rect 332 2276 340 2284
rect 236 2136 244 2144
rect 60 2116 68 2124
rect 92 2116 100 2124
rect 140 2116 148 2124
rect 188 2116 196 2124
rect 12 2096 20 2104
rect 92 2096 100 2104
rect 316 2156 324 2164
rect 188 2096 196 2104
rect 220 2096 228 2104
rect 268 2096 276 2104
rect 252 2076 260 2084
rect 252 1916 260 1924
rect 140 1896 148 1904
rect 60 1876 68 1884
rect 140 1876 148 1884
rect 60 1856 68 1864
rect 172 1856 180 1864
rect 332 2136 340 2144
rect 364 2416 372 2424
rect 812 2796 820 2804
rect 652 2716 660 2724
rect 684 2716 692 2724
rect 892 2836 900 2844
rect 844 2736 852 2744
rect 460 2696 468 2704
rect 540 2696 548 2704
rect 748 2696 756 2704
rect 780 2696 788 2704
rect 748 2676 756 2684
rect 540 2656 548 2664
rect 572 2656 580 2664
rect 716 2636 724 2644
rect 748 2556 756 2564
rect 412 2516 420 2524
rect 508 2436 516 2444
rect 428 2276 436 2284
rect 412 2256 420 2264
rect 396 2136 404 2144
rect 460 2136 468 2144
rect 332 2096 340 2104
rect 348 2076 356 2084
rect 380 1936 388 1944
rect 332 1876 340 1884
rect 380 1876 388 1884
rect 316 1816 324 1824
rect 300 1776 308 1784
rect 252 1756 260 1764
rect 300 1756 308 1764
rect 92 1716 100 1724
rect 204 1716 212 1724
rect 236 1716 244 1724
rect 204 1696 212 1704
rect 236 1696 244 1704
rect 188 1676 196 1684
rect 204 1676 212 1684
rect 76 1496 84 1504
rect 188 1476 196 1484
rect 284 1676 292 1684
rect 268 1596 276 1604
rect 284 1576 292 1584
rect 268 1536 276 1544
rect 252 1436 260 1444
rect 60 1356 68 1364
rect 188 1356 196 1364
rect 220 1356 228 1364
rect 28 1296 36 1304
rect 12 876 20 884
rect 12 696 20 704
rect 92 1096 100 1104
rect 236 1156 244 1164
rect 188 1136 196 1144
rect 268 1136 276 1144
rect 412 1856 420 1864
rect 380 1836 388 1844
rect 316 1716 324 1724
rect 380 1816 388 1824
rect 396 1776 404 1784
rect 380 1536 388 1544
rect 364 1516 372 1524
rect 476 1916 484 1924
rect 476 1896 484 1904
rect 492 1856 500 1864
rect 412 1676 420 1684
rect 332 1496 340 1504
rect 396 1496 404 1504
rect 316 1476 324 1484
rect 364 1456 372 1464
rect 396 1456 404 1464
rect 380 1436 388 1444
rect 380 1416 388 1424
rect 412 1416 420 1424
rect 332 1316 340 1324
rect 300 1116 308 1124
rect 220 1096 228 1104
rect 204 1076 212 1084
rect 268 1076 276 1084
rect 252 1056 260 1064
rect 268 1056 276 1064
rect 204 1036 212 1044
rect 236 956 244 964
rect 220 936 228 944
rect 76 736 84 744
rect 108 736 116 744
rect 60 696 68 704
rect 28 636 36 644
rect 108 716 116 724
rect 92 616 100 624
rect 140 896 148 904
rect 172 716 180 724
rect 140 636 148 644
rect 316 976 324 984
rect 252 936 260 944
rect 284 916 292 924
rect 364 1336 372 1344
rect 412 1356 420 1364
rect 396 1296 404 1304
rect 460 1516 468 1524
rect 796 2676 804 2684
rect 828 2676 836 2684
rect 812 2656 820 2664
rect 876 2676 884 2684
rect 972 3076 980 3084
rect 956 2896 964 2904
rect 940 2836 948 2844
rect 1228 3016 1236 3024
rect 1436 3016 1444 3024
rect 1084 2956 1092 2964
rect 1260 2956 1268 2964
rect 1388 2956 1396 2964
rect 1004 2936 1012 2944
rect 1052 2936 1060 2944
rect 1020 2916 1028 2924
rect 1100 2916 1108 2924
rect 1180 2916 1188 2924
rect 1212 2916 1220 2924
rect 972 2796 980 2804
rect 924 2736 932 2744
rect 924 2716 932 2724
rect 1116 2896 1124 2904
rect 1068 2856 1076 2864
rect 1132 2856 1140 2864
rect 1036 2696 1044 2704
rect 1148 2696 1156 2704
rect 1420 2936 1428 2944
rect 1548 2936 1556 2944
rect 1692 3036 1700 3044
rect 1580 3016 1588 3024
rect 1804 3036 1812 3044
rect 1868 3036 1876 3044
rect 1772 2956 1780 2964
rect 1836 2936 1844 2944
rect 1564 2916 1572 2924
rect 1644 2916 1652 2924
rect 1516 2876 1524 2884
rect 1436 2836 1444 2844
rect 1228 2756 1236 2764
rect 1308 2756 1316 2764
rect 1228 2736 1236 2744
rect 1004 2676 1012 2684
rect 1132 2676 1140 2684
rect 1244 2676 1252 2684
rect 908 2656 916 2664
rect 1180 2656 1188 2664
rect 1148 2596 1156 2604
rect 1196 2596 1204 2604
rect 1004 2556 1012 2564
rect 1116 2556 1124 2564
rect 1388 2676 1396 2684
rect 1260 2556 1268 2564
rect 636 2516 644 2524
rect 684 2516 692 2524
rect 1244 2516 1252 2524
rect 1308 2516 1316 2524
rect 1372 2516 1380 2524
rect 524 2396 532 2404
rect 956 2436 964 2444
rect 1356 2436 1364 2444
rect 716 2416 724 2424
rect 780 2416 788 2424
rect 828 2336 836 2344
rect 764 2296 766 2304
rect 766 2296 772 2304
rect 828 2296 836 2304
rect 572 2276 580 2284
rect 844 2276 852 2284
rect 684 2256 692 2264
rect 556 2216 564 2224
rect 844 2216 852 2224
rect 604 2196 612 2204
rect 668 2196 676 2204
rect 748 2156 756 2164
rect 828 2116 836 2124
rect 572 1956 580 1964
rect 588 1916 596 1924
rect 668 1916 676 1924
rect 588 1896 596 1904
rect 620 1896 628 1904
rect 524 1776 532 1784
rect 700 1956 708 1964
rect 764 2076 772 2084
rect 796 2076 804 2084
rect 780 2016 788 2024
rect 844 2016 852 2024
rect 716 1936 724 1944
rect 732 1936 740 1944
rect 700 1916 708 1924
rect 780 1916 788 1924
rect 716 1896 724 1904
rect 684 1876 692 1884
rect 652 1816 660 1824
rect 668 1816 676 1824
rect 636 1756 644 1764
rect 796 1856 804 1864
rect 828 1816 836 1824
rect 780 1796 788 1804
rect 732 1776 740 1784
rect 652 1696 660 1704
rect 572 1596 580 1604
rect 556 1536 564 1544
rect 508 1516 516 1524
rect 812 1756 820 1764
rect 828 1756 836 1764
rect 1244 2336 1252 2344
rect 988 2316 996 2324
rect 1020 2276 1028 2284
rect 876 2236 884 2244
rect 860 1976 868 1984
rect 924 2176 932 2184
rect 956 2176 964 2184
rect 1068 2176 1076 2184
rect 1004 2156 1012 2164
rect 1180 2156 1188 2164
rect 1228 2156 1236 2164
rect 924 2136 932 2144
rect 1020 2136 1028 2144
rect 1100 2136 1108 2144
rect 1084 2116 1092 2124
rect 1052 2076 1060 2084
rect 988 1976 996 1984
rect 940 1916 948 1924
rect 1020 1896 1028 1904
rect 764 1736 772 1744
rect 828 1736 836 1744
rect 844 1736 852 1744
rect 796 1716 804 1724
rect 780 1656 788 1664
rect 684 1556 692 1564
rect 732 1556 740 1564
rect 636 1536 644 1544
rect 460 1476 468 1484
rect 460 1396 468 1404
rect 460 1336 468 1344
rect 636 1496 644 1504
rect 668 1496 676 1504
rect 540 1476 548 1484
rect 572 1336 580 1344
rect 444 1316 452 1324
rect 476 1316 484 1324
rect 556 1316 564 1324
rect 428 1276 436 1284
rect 412 1236 420 1244
rect 348 1076 356 1084
rect 332 936 340 944
rect 348 936 356 944
rect 364 916 372 924
rect 284 896 292 904
rect 396 1036 404 1044
rect 396 1016 404 1024
rect 460 1236 468 1244
rect 572 1296 580 1304
rect 540 1256 548 1264
rect 508 1156 516 1164
rect 540 1136 548 1144
rect 508 1116 516 1124
rect 620 1236 628 1244
rect 588 1116 596 1124
rect 780 1516 788 1524
rect 764 1502 772 1504
rect 764 1496 772 1502
rect 684 1476 692 1484
rect 684 1436 692 1444
rect 716 1416 724 1424
rect 684 1356 692 1364
rect 652 1316 660 1324
rect 668 1276 676 1284
rect 684 1236 692 1244
rect 540 1096 548 1104
rect 684 1096 692 1104
rect 780 1376 788 1384
rect 764 1336 772 1344
rect 748 1318 756 1324
rect 748 1316 756 1318
rect 732 1116 740 1124
rect 828 1696 836 1704
rect 828 1416 836 1424
rect 892 1876 900 1884
rect 924 1876 932 1884
rect 876 1776 884 1784
rect 908 1756 916 1764
rect 1132 2116 1140 2124
rect 1164 2116 1172 2124
rect 1244 2136 1252 2144
rect 1212 2096 1220 2104
rect 1068 1976 1076 1984
rect 1116 1976 1124 1984
rect 1148 1936 1156 1944
rect 1084 1916 1092 1924
rect 1116 1916 1124 1924
rect 1084 1896 1092 1904
rect 940 1776 948 1784
rect 1036 1776 1044 1784
rect 1132 1836 1140 1844
rect 1100 1796 1108 1804
rect 1052 1736 1060 1744
rect 1148 1776 1156 1784
rect 1212 1916 1220 1924
rect 1212 1836 1220 1844
rect 1308 2296 1316 2304
rect 1340 2296 1348 2304
rect 1324 2236 1332 2244
rect 1308 2076 1316 2084
rect 1340 2096 1348 2104
rect 1372 2076 1380 2084
rect 1356 1976 1364 1984
rect 1276 1896 1284 1904
rect 1356 1896 1364 1904
rect 1244 1876 1252 1884
rect 1276 1876 1284 1884
rect 1228 1776 1236 1784
rect 1324 1876 1332 1884
rect 1340 1856 1348 1864
rect 1260 1756 1268 1764
rect 1292 1736 1300 1744
rect 1132 1716 1140 1724
rect 1212 1716 1220 1724
rect 1292 1716 1300 1724
rect 940 1556 948 1564
rect 892 1536 900 1544
rect 924 1496 932 1504
rect 860 1376 868 1384
rect 812 1356 820 1364
rect 892 1356 900 1364
rect 844 1216 852 1224
rect 876 1216 884 1224
rect 828 1116 836 1124
rect 476 1076 484 1084
rect 492 1076 500 1084
rect 444 1036 452 1044
rect 428 976 436 984
rect 604 1056 612 1064
rect 604 976 612 984
rect 588 956 596 964
rect 412 916 420 924
rect 396 896 404 904
rect 380 816 388 824
rect 428 896 436 904
rect 300 756 308 764
rect 412 756 420 764
rect 284 736 292 744
rect 268 716 276 724
rect 380 736 388 744
rect 316 716 324 724
rect 364 716 372 724
rect 252 696 260 704
rect 220 676 228 684
rect 172 656 180 664
rect 140 616 148 624
rect 156 616 164 624
rect 124 596 132 604
rect 332 696 340 704
rect 492 716 500 724
rect 412 696 420 704
rect 460 696 468 704
rect 684 956 692 964
rect 636 936 644 944
rect 620 836 628 844
rect 668 896 676 904
rect 652 876 660 884
rect 684 876 692 884
rect 620 736 628 744
rect 636 736 644 744
rect 732 976 740 984
rect 716 956 724 964
rect 748 916 756 924
rect 764 896 772 904
rect 732 856 740 864
rect 700 716 708 724
rect 524 696 532 704
rect 652 696 660 704
rect 716 696 724 704
rect 460 676 468 684
rect 332 656 340 664
rect 364 656 372 664
rect 428 656 436 664
rect 172 596 180 604
rect 236 596 244 604
rect 348 636 356 644
rect 172 556 180 564
rect 12 296 20 304
rect 60 296 68 304
rect 444 636 452 644
rect 364 616 372 624
rect 492 556 500 564
rect 460 536 468 544
rect 172 376 180 384
rect 220 376 228 384
rect 188 276 196 284
rect 300 216 308 224
rect 172 196 180 204
rect 220 196 228 204
rect 332 156 340 164
rect 140 136 148 144
rect 380 396 388 404
rect 412 496 420 504
rect 412 396 420 404
rect 396 276 404 284
rect 364 176 372 184
rect 412 156 420 164
rect 716 676 724 684
rect 636 656 644 664
rect 700 656 708 664
rect 684 636 692 644
rect 636 596 644 604
rect 604 556 612 564
rect 876 1156 884 1164
rect 860 1136 868 1144
rect 956 1516 964 1524
rect 988 1656 996 1664
rect 1068 1656 1076 1664
rect 1036 1576 1044 1584
rect 1068 1556 1076 1564
rect 1020 1516 1028 1524
rect 1084 1516 1092 1524
rect 1052 1496 1060 1504
rect 1116 1556 1124 1564
rect 1116 1536 1124 1544
rect 1116 1476 1124 1484
rect 988 1456 996 1464
rect 956 1376 964 1384
rect 1020 1436 1028 1444
rect 1036 1336 1044 1344
rect 940 1316 948 1324
rect 1004 1316 1012 1324
rect 1100 1316 1108 1324
rect 1068 1296 1076 1304
rect 988 1216 996 1224
rect 1036 1216 1044 1224
rect 892 1016 900 1024
rect 796 976 804 984
rect 796 956 804 964
rect 780 816 788 824
rect 780 736 788 744
rect 796 736 804 744
rect 748 676 756 684
rect 748 616 756 624
rect 748 536 756 544
rect 764 536 772 544
rect 924 956 932 964
rect 828 936 836 944
rect 876 916 884 924
rect 844 856 852 864
rect 828 716 836 724
rect 796 656 804 664
rect 860 656 868 664
rect 844 596 852 604
rect 828 536 836 544
rect 860 536 868 544
rect 956 1136 964 1144
rect 1068 1136 1076 1144
rect 1148 1556 1156 1564
rect 1164 1556 1172 1564
rect 1164 1516 1172 1524
rect 1502 2806 1510 2814
rect 1516 2806 1524 2814
rect 1530 2806 1538 2814
rect 1644 2716 1652 2724
rect 1628 2696 1636 2704
rect 1500 2636 1508 2644
rect 1692 2896 1700 2904
rect 1756 2876 1764 2884
rect 1740 2756 1748 2764
rect 1692 2716 1700 2724
rect 1676 2656 1684 2664
rect 1692 2616 1700 2624
rect 1660 2596 1668 2604
rect 1868 2816 1876 2824
rect 1916 2816 1924 2824
rect 1756 2696 1764 2704
rect 1788 2696 1796 2704
rect 1612 2556 1620 2564
rect 1644 2536 1652 2544
rect 1532 2516 1540 2524
rect 1884 2676 1892 2684
rect 1964 3096 1972 3104
rect 2380 3416 2388 3424
rect 2508 3396 2516 3404
rect 2572 3396 2580 3404
rect 2540 3336 2548 3344
rect 2684 3336 2692 3344
rect 2540 3256 2548 3264
rect 2396 3116 2404 3124
rect 2332 3096 2334 3104
rect 2334 3096 2340 3104
rect 2380 3096 2388 3104
rect 2076 3056 2084 3064
rect 2140 3056 2148 3064
rect 2172 3036 2180 3044
rect 2348 3036 2356 3044
rect 2044 2936 2052 2944
rect 2060 2936 2068 2944
rect 2092 2936 2100 2944
rect 2316 2936 2324 2944
rect 1996 2916 2004 2924
rect 2220 2916 2228 2924
rect 1964 2896 1972 2904
rect 1948 2796 1956 2804
rect 2476 3096 2484 3104
rect 2460 3056 2468 3064
rect 2476 2956 2484 2964
rect 2140 2896 2148 2904
rect 2428 2896 2436 2904
rect 2076 2836 2084 2844
rect 2124 2736 2132 2744
rect 2124 2696 2132 2704
rect 1884 2656 1892 2664
rect 1916 2636 1924 2644
rect 1868 2616 1876 2624
rect 1884 2616 1892 2624
rect 1852 2596 1860 2604
rect 1820 2536 1828 2544
rect 1452 2436 1460 2444
rect 1628 2416 1636 2424
rect 1502 2406 1510 2414
rect 1516 2406 1524 2414
rect 1530 2406 1538 2414
rect 1788 2436 1796 2444
rect 1820 2416 1828 2424
rect 1820 2376 1828 2384
rect 1932 2596 1940 2604
rect 1868 2416 1876 2424
rect 2076 2676 2078 2684
rect 2078 2676 2084 2684
rect 2124 2676 2132 2684
rect 2108 2636 2116 2644
rect 2364 2836 2372 2844
rect 2284 2816 2292 2824
rect 2300 2776 2308 2784
rect 2172 2736 2180 2744
rect 2220 2716 2228 2724
rect 2204 2656 2212 2664
rect 2140 2616 2148 2624
rect 2172 2616 2180 2624
rect 2076 2536 2084 2544
rect 2252 2516 2260 2524
rect 2204 2416 2212 2424
rect 1932 2376 1940 2384
rect 2268 2376 2276 2384
rect 1852 2276 1860 2284
rect 2012 2216 2020 2224
rect 1500 2176 1508 2184
rect 1660 2176 1668 2184
rect 1724 2176 1732 2184
rect 1980 2176 1988 2184
rect 1948 2156 1956 2164
rect 1436 2136 1444 2144
rect 1484 2096 1492 2104
rect 1452 2076 1460 2084
rect 1502 2006 1510 2014
rect 1516 2006 1524 2014
rect 1530 2006 1538 2014
rect 2092 2216 2100 2224
rect 2044 2156 2052 2164
rect 1644 2136 1652 2144
rect 1756 2136 1764 2144
rect 2044 2116 2052 2124
rect 1660 2076 1668 2084
rect 1420 1976 1428 1984
rect 1612 1976 1620 1984
rect 1644 1976 1652 1984
rect 1516 1896 1524 1904
rect 1596 1896 1604 1904
rect 1708 1896 1716 1904
rect 1724 1876 1732 1884
rect 1500 1856 1508 1864
rect 1772 1856 1780 1864
rect 1388 1796 1396 1804
rect 1468 1756 1476 1764
rect 1404 1716 1412 1724
rect 1564 1716 1572 1724
rect 1372 1696 1380 1704
rect 1356 1676 1364 1684
rect 1676 1676 1684 1684
rect 1420 1656 1428 1664
rect 1516 1656 1524 1664
rect 1228 1556 1236 1564
rect 1340 1556 1348 1564
rect 1180 1496 1188 1504
rect 1292 1536 1300 1544
rect 1244 1476 1252 1484
rect 1196 1456 1204 1464
rect 1228 1456 1236 1464
rect 1132 1296 1140 1304
rect 1276 1496 1284 1504
rect 1308 1516 1316 1524
rect 1276 1476 1284 1484
rect 1372 1476 1380 1484
rect 1260 1456 1268 1464
rect 1340 1456 1348 1464
rect 1356 1436 1364 1444
rect 1292 1396 1300 1404
rect 1244 1316 1252 1324
rect 1244 1296 1252 1304
rect 1212 1256 1220 1264
rect 1404 1596 1412 1604
rect 1404 1556 1412 1564
rect 1612 1616 1620 1624
rect 1502 1606 1510 1614
rect 1516 1606 1524 1614
rect 1530 1606 1538 1614
rect 1516 1576 1524 1584
rect 1404 1456 1412 1464
rect 1388 1356 1396 1364
rect 1484 1456 1492 1464
rect 1436 1396 1444 1404
rect 1276 1336 1284 1344
rect 1340 1336 1348 1344
rect 1420 1336 1428 1344
rect 1500 1336 1508 1344
rect 1356 1316 1364 1324
rect 1420 1316 1428 1324
rect 1452 1316 1460 1324
rect 1324 1296 1332 1304
rect 1340 1296 1348 1304
rect 1308 1276 1316 1284
rect 1196 1236 1204 1244
rect 1260 1236 1268 1244
rect 1132 1156 1140 1164
rect 1180 1156 1188 1164
rect 988 1096 996 1104
rect 1100 1096 1108 1104
rect 1196 1136 1204 1144
rect 1212 1116 1220 1124
rect 972 1076 980 1084
rect 972 936 980 944
rect 940 896 948 904
rect 908 836 916 844
rect 908 696 916 704
rect 924 676 932 684
rect 892 616 900 624
rect 716 516 724 524
rect 636 356 644 364
rect 620 336 628 344
rect 556 316 564 324
rect 444 296 452 304
rect 44 116 52 124
rect 348 116 356 124
rect 380 116 388 124
rect 428 136 436 144
rect 604 296 612 304
rect 716 496 724 504
rect 700 316 708 324
rect 764 316 772 324
rect 652 296 660 304
rect 540 196 548 204
rect 508 176 516 184
rect 764 196 772 204
rect 732 176 740 184
rect 780 156 788 164
rect 828 336 836 344
rect 844 316 852 324
rect 844 296 852 304
rect 876 496 884 504
rect 924 656 932 664
rect 1020 1076 1028 1084
rect 1132 1076 1140 1084
rect 1212 1076 1220 1084
rect 1084 1056 1092 1064
rect 1052 956 1060 964
rect 1132 956 1140 964
rect 1004 916 1012 924
rect 988 816 996 824
rect 1196 936 1204 944
rect 1180 916 1188 924
rect 1068 896 1076 904
rect 1100 896 1108 904
rect 1116 896 1124 904
rect 1212 896 1220 904
rect 1036 876 1044 884
rect 1084 876 1092 884
rect 1148 876 1156 884
rect 1068 856 1076 864
rect 1276 1076 1284 1084
rect 1244 1056 1252 1064
rect 1276 936 1284 944
rect 1244 876 1252 884
rect 1228 816 1236 824
rect 1196 736 1204 744
rect 1212 716 1220 724
rect 988 696 996 704
rect 1004 676 1012 684
rect 1180 676 1188 684
rect 988 636 996 644
rect 1020 656 1028 664
rect 1084 656 1092 664
rect 924 576 932 584
rect 1052 576 1060 584
rect 1116 556 1124 564
rect 1196 556 1204 564
rect 956 536 964 544
rect 1116 536 1124 544
rect 1292 916 1300 924
rect 1388 1276 1396 1284
rect 1356 1256 1364 1264
rect 1356 1136 1364 1144
rect 1324 1116 1332 1124
rect 1420 1116 1428 1124
rect 1420 1096 1428 1104
rect 1372 996 1380 1004
rect 1468 1296 1476 1304
rect 1996 1916 2004 1924
rect 1788 1756 1796 1764
rect 1932 1876 1940 1884
rect 1900 1856 1908 1864
rect 1900 1816 1908 1824
rect 1932 1776 1940 1784
rect 1948 1756 1956 1764
rect 1932 1736 1940 1744
rect 1804 1716 1812 1724
rect 1820 1716 1828 1724
rect 1852 1716 1860 1724
rect 1772 1676 1780 1684
rect 1708 1596 1716 1604
rect 1740 1476 1748 1484
rect 1772 1416 1780 1424
rect 1804 1416 1812 1424
rect 1564 1376 1572 1384
rect 1852 1396 1860 1404
rect 1916 1616 1924 1624
rect 2444 2676 2452 2684
rect 2588 3236 2596 3244
rect 2732 3476 2740 3484
rect 2892 3516 2900 3524
rect 2860 3496 2868 3504
rect 3020 3496 3028 3504
rect 3180 3496 3182 3504
rect 3182 3496 3188 3504
rect 2988 3476 2996 3484
rect 2716 3396 2724 3404
rect 3212 3436 3220 3444
rect 3038 3406 3046 3414
rect 3052 3406 3060 3414
rect 3066 3406 3074 3414
rect 2940 3396 2948 3404
rect 2924 3376 2932 3384
rect 2732 3356 2740 3364
rect 2780 3356 2788 3364
rect 2828 3356 2836 3364
rect 2876 3316 2884 3324
rect 2908 3316 2916 3324
rect 2812 3296 2820 3304
rect 2844 3296 2852 3304
rect 2908 3296 2916 3304
rect 2652 3136 2660 3144
rect 2700 3136 2708 3144
rect 2572 3116 2580 3124
rect 2716 3116 2724 3124
rect 2620 3096 2628 3104
rect 2636 3036 2644 3044
rect 2636 3016 2644 3024
rect 2572 2936 2580 2944
rect 2556 2916 2564 2924
rect 2508 2836 2516 2844
rect 2492 2816 2500 2824
rect 2748 3116 2756 3124
rect 2892 3136 2900 3144
rect 2844 3116 2852 3124
rect 2972 3316 2980 3324
rect 3052 3316 3060 3324
rect 3164 3316 3172 3324
rect 3004 3276 3012 3284
rect 2844 3096 2852 3104
rect 2684 3076 2692 3084
rect 2668 2856 2676 2864
rect 2668 2816 2676 2824
rect 2796 3076 2804 3084
rect 2828 3076 2836 3084
rect 2876 3076 2884 3084
rect 2908 3056 2916 3064
rect 2892 3036 2900 3044
rect 2780 3016 2788 3024
rect 2828 2956 2836 2964
rect 2940 2976 2948 2984
rect 2940 2936 2948 2944
rect 2700 2916 2708 2924
rect 2796 2916 2804 2924
rect 2924 2896 2932 2904
rect 2908 2876 2916 2884
rect 2764 2816 2772 2824
rect 2796 2796 2804 2804
rect 2892 2796 2900 2804
rect 2780 2716 2788 2724
rect 2684 2696 2692 2704
rect 2764 2696 2772 2704
rect 2636 2656 2644 2664
rect 2428 2576 2436 2584
rect 2332 2536 2340 2544
rect 2364 2536 2372 2544
rect 2396 2536 2404 2544
rect 2700 2676 2708 2684
rect 2668 2636 2676 2644
rect 2668 2576 2676 2584
rect 2700 2576 2708 2584
rect 2476 2556 2484 2564
rect 2668 2556 2676 2564
rect 2476 2516 2484 2524
rect 2444 2476 2452 2484
rect 2588 2476 2596 2484
rect 2508 2436 2516 2444
rect 2716 2316 2724 2324
rect 2860 2676 2868 2684
rect 2780 2656 2788 2664
rect 2844 2656 2852 2664
rect 2812 2636 2820 2644
rect 2860 2576 2868 2584
rect 2844 2556 2852 2564
rect 2876 2556 2884 2564
rect 2780 2396 2788 2404
rect 2652 2296 2660 2304
rect 2668 2296 2676 2304
rect 2860 2496 2868 2504
rect 2972 3096 2980 3104
rect 2956 2736 2964 2744
rect 2988 3076 2994 3084
rect 2994 3076 2996 3084
rect 3308 3696 3316 3704
rect 3292 3476 3300 3484
rect 3276 3456 3284 3464
rect 3260 3436 3268 3444
rect 3244 3416 3252 3424
rect 3804 3696 3812 3704
rect 3676 3596 3684 3604
rect 3372 3476 3380 3484
rect 3452 3456 3460 3464
rect 3516 3456 3524 3464
rect 3356 3416 3364 3424
rect 3324 3376 3332 3384
rect 3260 3336 3268 3344
rect 3260 3316 3268 3324
rect 3292 3316 3300 3324
rect 3324 3316 3332 3324
rect 3292 3296 3300 3304
rect 3276 3276 3284 3284
rect 3212 3256 3220 3264
rect 3148 3216 3156 3224
rect 3340 3136 3348 3144
rect 3324 3076 3332 3084
rect 3068 3056 3076 3064
rect 3244 3056 3252 3064
rect 2988 2976 2996 2984
rect 2988 2736 2996 2744
rect 2908 2576 2916 2584
rect 2908 2536 2916 2544
rect 2956 2636 2964 2644
rect 3148 3036 3156 3044
rect 3180 3036 3188 3044
rect 3038 3006 3046 3014
rect 3052 3006 3060 3014
rect 3066 3006 3074 3014
rect 3164 2976 3172 2984
rect 3052 2916 3060 2924
rect 3228 2916 3236 2924
rect 3052 2896 3060 2904
rect 3148 2896 3156 2904
rect 3228 2896 3236 2904
rect 3132 2856 3140 2864
rect 3020 2736 3028 2744
rect 3004 2676 3012 2684
rect 3084 2676 3092 2684
rect 3004 2656 3012 2664
rect 3038 2606 3046 2614
rect 3052 2606 3060 2614
rect 3066 2606 3074 2614
rect 3148 2836 3156 2844
rect 3196 2836 3204 2844
rect 3372 3296 3380 3304
rect 3372 3276 3380 3284
rect 3404 3256 3412 3264
rect 3372 3236 3380 3244
rect 3404 3216 3412 3224
rect 3324 2976 3332 2984
rect 3276 2936 3284 2944
rect 3292 2936 3300 2944
rect 3308 2916 3316 2924
rect 3260 2896 3268 2904
rect 3340 2896 3348 2904
rect 3292 2856 3300 2864
rect 3340 2856 3348 2864
rect 3356 2816 3364 2824
rect 3260 2796 3268 2804
rect 3340 2796 3348 2804
rect 3132 2556 3140 2564
rect 3036 2536 3044 2544
rect 3084 2536 3092 2544
rect 3148 2536 3156 2544
rect 2876 2296 2884 2304
rect 2300 2276 2308 2284
rect 2444 2276 2452 2284
rect 2252 2256 2260 2264
rect 2172 2236 2180 2244
rect 2204 2236 2212 2244
rect 2444 2236 2452 2244
rect 2124 2116 2132 2124
rect 2156 2116 2164 2124
rect 2492 2216 2500 2224
rect 2284 2176 2292 2184
rect 2476 2176 2484 2184
rect 2252 2136 2260 2144
rect 2076 1896 2084 1904
rect 2108 1876 2116 1884
rect 2060 1856 2068 1864
rect 2124 1856 2132 1864
rect 2044 1836 2052 1844
rect 2156 1876 2164 1884
rect 2140 1836 2148 1844
rect 2236 1876 2244 1884
rect 2252 1816 2260 1824
rect 2076 1796 2084 1804
rect 2188 1796 2196 1804
rect 2012 1716 2020 1724
rect 1964 1696 1972 1704
rect 1996 1696 2004 1704
rect 2012 1696 2020 1704
rect 2300 2036 2308 2044
rect 2364 2036 2372 2044
rect 2444 2036 2452 2044
rect 2444 1936 2452 1944
rect 2348 1896 2356 1904
rect 2316 1876 2324 1884
rect 2380 1876 2388 1884
rect 2332 1836 2340 1844
rect 2396 1836 2404 1844
rect 2252 1776 2260 1784
rect 2284 1776 2292 1784
rect 2124 1756 2132 1764
rect 2092 1696 2100 1704
rect 2012 1496 2020 1504
rect 2044 1496 2052 1504
rect 1980 1476 1988 1484
rect 1932 1396 1940 1404
rect 1580 1356 1588 1364
rect 1900 1356 1908 1364
rect 1564 1316 1572 1324
rect 1548 1276 1556 1284
rect 1468 1236 1476 1244
rect 1500 1236 1508 1244
rect 1532 1236 1540 1244
rect 1502 1206 1510 1214
rect 1516 1206 1524 1214
rect 1530 1206 1538 1214
rect 1612 1276 1620 1284
rect 1580 1236 1588 1244
rect 1500 1116 1508 1124
rect 1468 1076 1476 1084
rect 1452 1036 1460 1044
rect 1324 956 1332 964
rect 1308 896 1316 904
rect 1324 876 1332 884
rect 1372 916 1380 924
rect 1420 896 1428 904
rect 1356 876 1364 884
rect 1404 876 1412 884
rect 1308 756 1316 764
rect 1340 696 1348 704
rect 940 516 948 524
rect 876 456 884 464
rect 908 456 916 464
rect 828 156 836 164
rect 828 136 836 144
rect 780 116 788 124
rect 860 236 868 244
rect 892 356 900 364
rect 892 316 900 324
rect 924 316 932 324
rect 908 296 916 304
rect 924 296 932 304
rect 1244 496 1252 504
rect 1132 356 1140 364
rect 1148 336 1156 344
rect 1020 316 1028 324
rect 1164 316 1172 324
rect 1212 356 1220 364
rect 1276 336 1284 344
rect 1244 296 1252 304
rect 1436 856 1444 864
rect 1388 816 1396 824
rect 1356 516 1364 524
rect 1836 1336 1844 1344
rect 2044 1456 2052 1464
rect 2076 1356 2084 1364
rect 1964 1336 1972 1344
rect 2012 1336 2020 1344
rect 2028 1336 2036 1344
rect 2636 2276 2638 2284
rect 2638 2276 2644 2284
rect 2748 2276 2756 2284
rect 2972 2516 2980 2524
rect 3004 2456 3012 2464
rect 2924 2436 2932 2444
rect 3020 2356 3028 2364
rect 3148 2496 3156 2504
rect 3100 2436 3108 2444
rect 3020 2316 3028 2324
rect 3036 2316 3044 2324
rect 2972 2296 2980 2304
rect 2828 2256 2836 2264
rect 2668 2156 2676 2164
rect 2748 2156 2756 2164
rect 2636 2136 2644 2144
rect 2796 2136 2804 2144
rect 2828 2056 2836 2064
rect 2716 1956 2724 1964
rect 2476 1916 2484 1924
rect 2492 1896 2500 1904
rect 2588 1896 2596 1904
rect 2476 1876 2484 1884
rect 2460 1736 2468 1744
rect 2684 1876 2692 1884
rect 2876 2056 2884 2064
rect 2860 1936 2868 1944
rect 2876 1936 2884 1944
rect 2940 2276 2948 2284
rect 3036 2276 3044 2284
rect 3052 2276 3060 2284
rect 2956 2216 2964 2224
rect 3038 2206 3046 2214
rect 3052 2206 3060 2214
rect 3066 2206 3074 2214
rect 3132 2316 3140 2324
rect 3228 2676 3236 2684
rect 3260 2656 3268 2664
rect 3180 2576 3188 2584
rect 3276 2556 3284 2564
rect 3196 2516 3204 2524
rect 3180 2496 3188 2504
rect 3244 2496 3252 2504
rect 3164 2476 3172 2484
rect 3196 2476 3204 2484
rect 3164 2456 3172 2464
rect 3244 2476 3252 2484
rect 3292 2476 3300 2484
rect 3212 2436 3220 2444
rect 3260 2436 3268 2444
rect 3212 2336 3220 2344
rect 3116 2296 3124 2304
rect 3196 2296 3204 2304
rect 3116 2216 3124 2224
rect 3004 2176 3012 2184
rect 2972 2136 2980 2144
rect 2908 1956 2916 1964
rect 2540 1816 2548 1824
rect 2956 1896 2964 1904
rect 2924 1856 2932 1864
rect 2748 1776 2756 1784
rect 2892 1776 2900 1784
rect 2556 1736 2564 1744
rect 2284 1716 2292 1724
rect 2252 1676 2260 1684
rect 2236 1556 2244 1564
rect 2140 1516 2148 1524
rect 2412 1596 2420 1604
rect 2140 1496 2148 1504
rect 2204 1496 2212 1504
rect 2172 1476 2180 1484
rect 2220 1476 2228 1484
rect 2188 1456 2196 1464
rect 2764 1736 2772 1744
rect 2812 1736 2820 1744
rect 2908 1736 2916 1744
rect 2588 1596 2596 1604
rect 2572 1556 2580 1564
rect 2812 1596 2820 1604
rect 2844 1596 2852 1604
rect 2716 1536 2724 1544
rect 2780 1536 2788 1544
rect 2604 1516 2612 1524
rect 2524 1496 2532 1504
rect 2492 1456 2500 1464
rect 2156 1436 2164 1444
rect 2380 1436 2388 1444
rect 1932 1316 1940 1324
rect 2028 1316 2036 1324
rect 2092 1316 2100 1324
rect 1708 1196 1716 1204
rect 1804 1196 1812 1204
rect 2092 1296 2100 1304
rect 1932 1176 1940 1184
rect 1644 1116 1652 1124
rect 1532 1096 1540 1104
rect 1756 1096 1764 1104
rect 1564 1056 1572 1064
rect 1468 876 1476 884
rect 1502 806 1510 814
rect 1516 806 1524 814
rect 1530 806 1538 814
rect 1500 756 1508 764
rect 1452 736 1460 744
rect 1484 736 1492 744
rect 1468 696 1476 704
rect 1404 676 1412 684
rect 1404 556 1412 564
rect 1468 556 1476 564
rect 1468 516 1476 524
rect 1372 496 1380 504
rect 1340 456 1348 464
rect 1308 356 1316 364
rect 1340 336 1348 344
rect 1292 316 1300 324
rect 1340 316 1348 324
rect 892 276 900 284
rect 940 276 948 284
rect 1260 276 1268 284
rect 908 236 916 244
rect 1292 256 1300 264
rect 1004 196 1012 204
rect 1260 196 1268 204
rect 1100 176 1108 184
rect 1308 196 1316 204
rect 1020 136 1028 144
rect 1580 1036 1588 1044
rect 1580 776 1588 784
rect 1564 736 1572 744
rect 1548 556 1556 564
rect 1452 476 1460 484
rect 1484 476 1492 484
rect 1804 1076 1812 1084
rect 1740 1036 1748 1044
rect 1788 936 1796 944
rect 1628 702 1636 704
rect 1628 696 1636 702
rect 1644 676 1652 684
rect 1596 536 1604 544
rect 1532 456 1540 464
rect 1502 406 1510 414
rect 1516 406 1524 414
rect 1530 406 1538 414
rect 1404 376 1412 384
rect 1452 376 1460 384
rect 1596 476 1604 484
rect 1372 296 1380 304
rect 1532 302 1540 304
rect 1532 296 1540 302
rect 1564 296 1572 304
rect 1628 596 1636 604
rect 1852 1096 1860 1104
rect 1868 1076 1876 1084
rect 1916 1076 1924 1084
rect 1836 1056 1844 1064
rect 1980 1156 1988 1164
rect 1980 1096 1988 1104
rect 2028 1096 2036 1104
rect 2188 1336 2196 1344
rect 2236 1196 2244 1204
rect 2300 1336 2308 1344
rect 2444 1336 2452 1344
rect 2380 1276 2388 1284
rect 2284 1216 2292 1224
rect 2268 1176 2276 1184
rect 2204 1136 2212 1144
rect 2236 1136 2244 1144
rect 2268 1136 2276 1144
rect 2140 1116 2148 1124
rect 2188 1116 2196 1124
rect 2092 1076 2100 1084
rect 2044 1036 2052 1044
rect 1900 936 1908 944
rect 1756 856 1764 864
rect 1708 816 1716 824
rect 1868 816 1876 824
rect 1900 796 1908 804
rect 1820 776 1828 784
rect 1884 736 1892 744
rect 1820 696 1828 704
rect 1772 676 1780 684
rect 1740 616 1748 624
rect 1660 536 1668 544
rect 1692 536 1700 544
rect 1628 496 1636 504
rect 1468 256 1476 264
rect 1468 236 1476 244
rect 1628 236 1636 244
rect 1388 196 1396 204
rect 1548 216 1556 224
rect 1340 176 1348 184
rect 1340 156 1348 164
rect 1996 736 2004 744
rect 1964 716 1972 724
rect 2044 896 2052 904
rect 2108 1056 2116 1064
rect 2188 1096 2196 1104
rect 2220 1096 2228 1104
rect 2252 1096 2260 1104
rect 2172 1076 2180 1084
rect 2188 1076 2196 1084
rect 2156 1036 2164 1044
rect 2268 1076 2276 1084
rect 2236 1036 2244 1044
rect 2268 976 2276 984
rect 2268 956 2276 964
rect 2220 936 2228 944
rect 2124 916 2132 924
rect 2156 916 2164 924
rect 2172 916 2180 924
rect 2268 916 2276 924
rect 2124 896 2132 904
rect 2156 896 2164 904
rect 2076 796 2084 804
rect 2028 716 2036 724
rect 1916 696 1924 704
rect 2012 696 2020 704
rect 2076 696 2084 704
rect 1868 676 1876 684
rect 1932 676 1940 684
rect 2012 676 2020 684
rect 2172 676 2180 684
rect 1964 656 1972 664
rect 2204 656 2212 664
rect 1788 596 1796 604
rect 2124 576 2132 584
rect 2220 576 2228 584
rect 1932 556 1940 564
rect 2204 556 2212 564
rect 2380 1156 2388 1164
rect 2492 1336 2500 1344
rect 2540 1356 2548 1364
rect 2604 1336 2612 1344
rect 2620 1336 2628 1344
rect 2524 1316 2532 1324
rect 2620 1316 2628 1324
rect 2572 1296 2580 1304
rect 2476 1196 2484 1204
rect 2492 1176 2500 1184
rect 2332 1096 2340 1104
rect 2364 1096 2372 1104
rect 2444 1096 2452 1104
rect 2348 1056 2356 1064
rect 2364 1056 2372 1064
rect 2412 1056 2420 1064
rect 2316 956 2324 964
rect 2428 1036 2436 1044
rect 2476 1036 2484 1044
rect 2396 976 2404 984
rect 2444 956 2452 964
rect 2412 936 2420 944
rect 2396 916 2404 924
rect 2348 896 2356 904
rect 2460 796 2468 804
rect 2380 716 2388 724
rect 2508 1156 2516 1164
rect 2652 1216 2660 1224
rect 2668 1196 2676 1204
rect 2620 1176 2628 1184
rect 2604 1136 2612 1144
rect 2508 1120 2516 1124
rect 2508 1116 2516 1120
rect 2572 1116 2580 1124
rect 2604 1096 2612 1104
rect 2572 1056 2580 1064
rect 2780 1476 2788 1484
rect 2956 1876 2964 1884
rect 2940 1836 2948 1844
rect 3180 2156 3188 2164
rect 3020 2136 3028 2144
rect 3388 3036 3396 3044
rect 3388 2956 3396 2964
rect 3532 3376 3540 3384
rect 3564 3336 3572 3344
rect 3644 3316 3652 3324
rect 3596 3176 3604 3184
rect 3580 3136 3588 3144
rect 3484 3116 3492 3124
rect 3468 3076 3476 3084
rect 3484 2956 3492 2964
rect 3564 3056 3572 3064
rect 3516 2936 3524 2944
rect 3452 2916 3460 2924
rect 3516 2896 3524 2904
rect 3420 2856 3428 2864
rect 3468 2856 3476 2864
rect 3404 2796 3412 2804
rect 3388 2756 3396 2764
rect 3436 2736 3444 2744
rect 3452 2736 3460 2744
rect 3404 2676 3412 2684
rect 3436 2676 3444 2684
rect 3372 2556 3380 2564
rect 3388 2556 3396 2564
rect 3372 2476 3380 2484
rect 3356 2336 3364 2344
rect 3420 2536 3428 2544
rect 3436 2496 3444 2504
rect 3484 2716 3492 2724
rect 3516 2716 3524 2724
rect 3548 2936 3556 2944
rect 3596 2976 3604 2984
rect 3612 2916 3620 2924
rect 3596 2896 3604 2904
rect 3548 2876 3556 2884
rect 3612 2776 3620 2784
rect 3596 2756 3604 2764
rect 3564 2736 3572 2744
rect 3564 2716 3572 2724
rect 3500 2696 3508 2704
rect 3548 2696 3556 2704
rect 3596 2696 3604 2704
rect 3932 4096 3940 4104
rect 3948 4096 3956 4104
rect 3916 4076 3924 4084
rect 3948 4076 3956 4084
rect 4076 4216 4084 4224
rect 3996 4196 4004 4204
rect 4012 4136 4020 4144
rect 4028 4136 4036 4144
rect 4092 4176 4100 4184
rect 4108 4176 4116 4184
rect 4156 4336 4164 4344
rect 4204 4376 4212 4384
rect 4140 4296 4148 4304
rect 4156 4156 4164 4164
rect 4172 4156 4180 4164
rect 4300 4496 4308 4504
rect 4028 4116 4036 4124
rect 4060 4116 4068 4124
rect 4108 4116 4116 4124
rect 4156 4116 4164 4124
rect 4012 4096 4020 4104
rect 4220 4116 4228 4124
rect 4396 4536 4404 4544
rect 4444 4516 4452 4524
rect 4364 4476 4372 4484
rect 4316 4456 4324 4464
rect 4348 4436 4356 4444
rect 4252 4296 4260 4304
rect 4252 4276 4260 4284
rect 4236 4076 4244 4084
rect 3996 4056 4004 4064
rect 4236 4036 4244 4044
rect 3836 3976 3844 3984
rect 3932 3976 3940 3984
rect 4092 3936 4100 3944
rect 4012 3896 4020 3904
rect 4268 4196 4276 4204
rect 4284 4176 4292 4184
rect 4572 4956 4580 4964
rect 4764 4976 4772 4984
rect 4716 4956 4724 4964
rect 4732 4936 4740 4944
rect 4796 4936 4804 4944
rect 4556 4896 4564 4904
rect 4540 4836 4548 4844
rect 4556 4836 4564 4844
rect 4508 4516 4516 4524
rect 4460 4476 4468 4484
rect 4412 4436 4420 4444
rect 4396 4296 4404 4304
rect 4460 4276 4468 4284
rect 4380 4216 4388 4224
rect 4364 4156 4372 4164
rect 4412 4156 4420 4164
rect 4348 4136 4356 4144
rect 4364 4116 4372 4124
rect 4444 4176 4452 4184
rect 4524 4476 4532 4484
rect 4508 4436 4516 4444
rect 4574 4806 4582 4814
rect 4588 4806 4596 4814
rect 4602 4806 4610 4814
rect 4668 4916 4676 4924
rect 4668 4896 4676 4904
rect 4700 4876 4708 4884
rect 4716 4816 4724 4824
rect 4668 4776 4676 4784
rect 4652 4716 4660 4724
rect 4684 4736 4692 4744
rect 4652 4676 4660 4684
rect 4684 4676 4692 4684
rect 4748 4896 4756 4904
rect 4716 4656 4724 4664
rect 4604 4636 4612 4644
rect 4604 4576 4612 4584
rect 4556 4556 4564 4564
rect 4716 4616 4724 4624
rect 4700 4536 4708 4544
rect 4780 4876 4788 4884
rect 4780 4816 4788 4824
rect 4780 4736 4788 4744
rect 4812 4736 4820 4744
rect 4812 4716 4820 4724
rect 4988 5296 4996 5304
rect 4908 5276 4916 5284
rect 4940 5276 4948 5284
rect 5180 5276 5188 5284
rect 5196 5216 5204 5224
rect 5164 5196 5172 5204
rect 5212 5196 5220 5204
rect 4988 5176 4996 5184
rect 5036 5176 5044 5184
rect 4908 5116 4916 5124
rect 5052 5136 5060 5144
rect 5308 5296 5316 5304
rect 5228 5136 5236 5144
rect 5116 5116 5124 5124
rect 5180 5116 5188 5124
rect 5228 5116 5236 5124
rect 4860 5096 4868 5104
rect 4876 5096 4884 5104
rect 4908 5016 4916 5024
rect 4892 4956 4900 4964
rect 4892 4896 4900 4904
rect 5004 5056 5012 5064
rect 4956 4976 4964 4984
rect 5068 5036 5076 5044
rect 5084 4996 5092 5004
rect 5068 4976 5076 4984
rect 5036 4956 5044 4964
rect 5004 4936 5012 4944
rect 4972 4896 4980 4904
rect 4924 4836 4932 4844
rect 4940 4836 4948 4844
rect 4860 4756 4868 4764
rect 4876 4756 4884 4764
rect 4860 4716 4868 4724
rect 4828 4696 4836 4704
rect 4780 4636 4788 4644
rect 4764 4556 4772 4564
rect 4812 4556 4820 4564
rect 4748 4536 4756 4544
rect 4796 4536 4804 4544
rect 4748 4516 4756 4524
rect 4716 4496 4724 4504
rect 4540 4456 4548 4464
rect 4636 4456 4644 4464
rect 4574 4406 4582 4414
rect 4588 4406 4596 4414
rect 4602 4406 4610 4414
rect 4540 4376 4548 4384
rect 4524 4356 4532 4364
rect 4508 4296 4516 4304
rect 4492 4156 4500 4164
rect 4620 4336 4628 4344
rect 4572 4156 4580 4164
rect 4524 4136 4532 4144
rect 4604 4136 4612 4144
rect 4700 4356 4708 4364
rect 4860 4596 4868 4604
rect 4844 4556 4852 4564
rect 4860 4536 4868 4544
rect 4956 4816 4964 4824
rect 4940 4776 4948 4784
rect 4988 4876 4996 4884
rect 4972 4716 4980 4724
rect 5068 4896 5076 4904
rect 5020 4876 5028 4884
rect 5036 4876 5044 4884
rect 5036 4716 5044 4724
rect 5084 4716 5092 4724
rect 5004 4676 5012 4684
rect 5020 4676 5028 4684
rect 5068 4656 5076 4664
rect 5052 4576 5060 4584
rect 4940 4536 4948 4544
rect 4988 4536 4996 4544
rect 5052 4536 5060 4544
rect 4844 4516 4852 4524
rect 4924 4516 4932 4524
rect 5004 4516 5012 4524
rect 5084 4516 5092 4524
rect 4924 4496 4932 4504
rect 5036 4496 5044 4504
rect 4956 4436 4964 4444
rect 4764 4376 4772 4384
rect 4748 4336 4756 4344
rect 4956 4296 4964 4304
rect 4652 4176 4660 4184
rect 4812 4276 4820 4284
rect 4956 4276 4964 4284
rect 4924 4256 4932 4264
rect 4988 4196 4996 4204
rect 4716 4156 4724 4164
rect 4908 4156 4916 4164
rect 4668 4136 4676 4144
rect 4748 4136 4756 4144
rect 4636 4116 4644 4124
rect 4716 4116 4724 4124
rect 4412 4096 4420 4104
rect 4476 4096 4484 4104
rect 4268 4076 4276 4084
rect 4332 4076 4340 4084
rect 4652 4076 4660 4084
rect 4892 4116 4900 4124
rect 4844 4096 4852 4104
rect 4732 4076 4740 4084
rect 4300 3976 4308 3984
rect 4428 3976 4436 3984
rect 4284 3876 4292 3884
rect 3868 3816 3876 3824
rect 3964 3816 3972 3824
rect 3948 3796 3956 3804
rect 4252 3836 4260 3844
rect 3980 3796 3988 3804
rect 4044 3796 4052 3804
rect 4076 3776 4084 3784
rect 3996 3736 4004 3744
rect 3932 3536 3940 3544
rect 3948 3516 3956 3524
rect 4012 3516 4020 3524
rect 4076 3516 4084 3524
rect 4316 3816 4324 3824
rect 4172 3756 4180 3764
rect 4428 3876 4436 3884
rect 4574 4006 4582 4014
rect 4588 4006 4596 4014
rect 4602 4006 4610 4014
rect 4460 3936 4468 3944
rect 4508 3896 4516 3904
rect 4444 3856 4452 3864
rect 4380 3776 4388 3784
rect 4188 3736 4196 3744
rect 4204 3716 4212 3724
rect 4332 3716 4340 3724
rect 4476 3736 4484 3744
rect 4860 4076 4868 4084
rect 4844 3996 4852 4004
rect 4956 4140 4964 4144
rect 4956 4136 4964 4140
rect 4988 4116 4996 4124
rect 5020 4096 5028 4104
rect 5052 4476 5060 4484
rect 5052 4356 5060 4364
rect 5052 4296 5060 4304
rect 5212 5076 5220 5084
rect 5196 5056 5204 5064
rect 5180 4996 5188 5004
rect 5164 4976 5172 4984
rect 5116 4956 5124 4964
rect 5164 4916 5172 4924
rect 5276 5076 5284 5084
rect 5228 5056 5236 5064
rect 5292 5036 5300 5044
rect 5116 4896 5124 4904
rect 5212 4896 5220 4904
rect 5132 4876 5140 4884
rect 5196 4876 5204 4884
rect 5164 4836 5172 4844
rect 5180 4736 5188 4744
rect 5196 4696 5204 4704
rect 5212 4596 5220 4604
rect 5148 4576 5156 4584
rect 5244 4836 5252 4844
rect 5276 4976 5284 4984
rect 5260 4676 5268 4684
rect 5132 4516 5140 4524
rect 5148 4516 5156 4524
rect 5180 4516 5188 4524
rect 5292 4956 5300 4964
rect 5292 4716 5300 4724
rect 5500 5516 5508 5524
rect 5916 5556 5924 5564
rect 5788 5476 5796 5484
rect 5388 5456 5396 5464
rect 5340 5376 5348 5384
rect 5548 5456 5556 5464
rect 5612 5456 5620 5464
rect 5756 5456 5764 5464
rect 5868 5456 5876 5464
rect 5596 5436 5604 5444
rect 5452 5416 5460 5424
rect 5388 5396 5396 5404
rect 5436 5356 5444 5364
rect 5644 5356 5652 5364
rect 5788 5336 5796 5344
rect 5420 5156 5428 5164
rect 5356 5136 5364 5144
rect 5724 5236 5732 5244
rect 5756 5176 5764 5184
rect 5452 5156 5460 5164
rect 5452 5136 5460 5144
rect 5484 5116 5492 5124
rect 5692 5116 5700 5124
rect 5788 5116 5796 5124
rect 5388 5096 5396 5104
rect 5436 5076 5444 5084
rect 5356 5056 5364 5064
rect 5324 5016 5332 5024
rect 5388 5036 5396 5044
rect 5372 4996 5380 5004
rect 5436 4996 5444 5004
rect 5436 4956 5444 4964
rect 5436 4896 5444 4904
rect 5404 4836 5412 4844
rect 5724 5076 5732 5084
rect 5756 5076 5764 5084
rect 5612 5056 5620 5064
rect 5676 4996 5684 5004
rect 5628 4956 5636 4964
rect 5468 4916 5476 4924
rect 5740 4936 5748 4944
rect 5724 4916 5732 4924
rect 5468 4896 5476 4904
rect 5788 4836 5796 4844
rect 5452 4756 5460 4764
rect 5308 4696 5316 4704
rect 5484 4676 5492 4684
rect 5356 4576 5364 4584
rect 5404 4576 5412 4584
rect 5436 4576 5444 4584
rect 5308 4516 5316 4524
rect 5420 4516 5428 4524
rect 5116 4476 5124 4484
rect 5132 4476 5140 4484
rect 5164 4476 5172 4484
rect 5100 4456 5108 4464
rect 5260 4496 5268 4504
rect 5196 4436 5204 4444
rect 5356 4396 5364 4404
rect 5116 4376 5124 4384
rect 5292 4376 5300 4384
rect 5548 4736 5556 4744
rect 5532 4716 5540 4724
rect 5548 4696 5556 4704
rect 5772 4696 5780 4704
rect 5676 4676 5684 4684
rect 5788 4676 5796 4684
rect 5564 4656 5572 4664
rect 5516 4596 5524 4604
rect 5628 4596 5636 4604
rect 5596 4576 5604 4584
rect 5564 4556 5572 4564
rect 5596 4516 5604 4524
rect 5596 4496 5604 4504
rect 5452 4396 5460 4404
rect 5484 4396 5492 4404
rect 5516 4396 5524 4404
rect 5724 4536 5732 4544
rect 5660 4416 5668 4424
rect 5196 4296 5204 4304
rect 5468 4296 5476 4304
rect 5564 4296 5572 4304
rect 5084 4156 5092 4164
rect 5052 4136 5060 4144
rect 5100 4136 5108 4144
rect 5148 4136 5156 4144
rect 5052 4116 5060 4124
rect 5132 4116 5140 4124
rect 5164 4116 5172 4124
rect 5164 4096 5172 4104
rect 5180 4096 5188 4104
rect 5084 4016 5092 4024
rect 5036 3996 5044 4004
rect 5068 3956 5076 3964
rect 4892 3916 4900 3924
rect 4748 3876 4756 3884
rect 4748 3836 4756 3844
rect 4524 3816 4532 3824
rect 4572 3776 4580 3784
rect 5100 3996 5108 4004
rect 5164 3936 5172 3944
rect 5132 3916 5140 3924
rect 5084 3896 5092 3904
rect 5276 4256 5284 4264
rect 5260 4216 5268 4224
rect 5308 4216 5316 4224
rect 5452 4196 5460 4204
rect 5420 4176 5428 4184
rect 5468 4176 5476 4184
rect 5212 4156 5220 4164
rect 5500 4156 5508 4164
rect 5356 4136 5364 4144
rect 5468 4136 5476 4144
rect 5324 4116 5332 4124
rect 5452 4116 5460 4124
rect 5212 4096 5220 4104
rect 5532 4276 5540 4284
rect 5532 4236 5540 4244
rect 5612 4276 5620 4284
rect 5708 4276 5716 4284
rect 5660 4236 5668 4244
rect 5692 4236 5700 4244
rect 5660 4216 5668 4224
rect 5580 4196 5588 4204
rect 5516 4136 5524 4144
rect 5292 3976 5300 3984
rect 5484 3916 5492 3924
rect 5516 3976 5524 3984
rect 5500 3896 5502 3904
rect 5502 3896 5508 3904
rect 4940 3876 4948 3884
rect 5148 3876 5156 3884
rect 4844 3836 4852 3844
rect 4844 3816 4852 3824
rect 5116 3836 5124 3844
rect 5148 3836 5156 3844
rect 5084 3816 5092 3824
rect 5308 3876 5316 3884
rect 5212 3816 5220 3824
rect 5340 3816 5348 3824
rect 5372 3816 5380 3824
rect 5692 4116 5700 4124
rect 5804 4416 5812 4424
rect 5756 4396 5764 4404
rect 5836 5256 5844 5264
rect 5836 5236 5844 5244
rect 5884 5236 5892 5244
rect 6092 5596 6100 5604
rect 6076 5556 6084 5564
rect 5932 5476 5940 5484
rect 5948 5396 5956 5404
rect 6028 5396 6036 5404
rect 5980 5336 5988 5344
rect 6124 5336 6132 5344
rect 5996 5296 6004 5304
rect 5948 5196 5956 5204
rect 5980 5196 5988 5204
rect 5916 4996 5924 5004
rect 5948 4996 5956 5004
rect 5980 4916 5988 4924
rect 5996 4676 6004 4684
rect 5836 4656 5844 4664
rect 5884 4656 5892 4664
rect 5916 4596 5924 4604
rect 5964 4596 5972 4604
rect 5916 4556 5924 4564
rect 5948 4496 5956 4504
rect 5996 4416 6004 4424
rect 6060 4416 6068 4424
rect 5820 4276 5828 4284
rect 5820 4256 5828 4264
rect 5852 4216 5860 4224
rect 5564 4076 5572 4084
rect 5676 4076 5684 4084
rect 5548 4016 5556 4024
rect 5580 3996 5588 4004
rect 5612 3936 5620 3944
rect 5660 3916 5668 3924
rect 5564 3896 5572 3904
rect 5580 3896 5588 3904
rect 5612 3896 5620 3904
rect 5548 3876 5556 3884
rect 5596 3876 5604 3884
rect 5532 3836 5540 3844
rect 5420 3796 5428 3804
rect 5468 3796 5476 3804
rect 4988 3756 4996 3764
rect 5068 3756 5076 3764
rect 4684 3736 4692 3744
rect 4780 3736 4788 3744
rect 4828 3736 4836 3744
rect 5004 3736 5012 3744
rect 4508 3716 4516 3724
rect 4652 3716 4660 3724
rect 4764 3716 4772 3724
rect 4860 3716 4868 3724
rect 4236 3696 4244 3704
rect 4380 3696 4388 3704
rect 4492 3696 4500 3704
rect 4140 3676 4148 3684
rect 4380 3596 4388 3604
rect 4574 3606 4582 3614
rect 4588 3606 4596 3614
rect 4602 3606 4610 3614
rect 4140 3536 4148 3544
rect 4124 3516 4132 3524
rect 4348 3516 4356 3524
rect 4460 3516 4468 3524
rect 3884 3496 3892 3504
rect 3900 3496 3908 3504
rect 3996 3496 4004 3504
rect 4092 3496 4100 3504
rect 3740 3476 3748 3484
rect 3788 3456 3796 3464
rect 3708 3436 3716 3444
rect 3820 3396 3828 3404
rect 3804 3356 3812 3364
rect 3756 3336 3764 3344
rect 3740 3316 3748 3324
rect 3724 3296 3732 3304
rect 3740 3276 3748 3284
rect 3788 3276 3796 3284
rect 3772 3236 3780 3244
rect 3724 3136 3732 3144
rect 3708 3116 3716 3124
rect 3708 3096 3716 3104
rect 3692 3076 3700 3084
rect 3676 2936 3684 2944
rect 3756 3176 3764 3184
rect 3756 3136 3764 3144
rect 3916 3336 3924 3344
rect 3980 3316 3988 3324
rect 3852 3296 3860 3304
rect 3916 3296 3924 3304
rect 4044 3476 4052 3484
rect 4092 3476 4100 3484
rect 4012 3456 4020 3464
rect 4028 3396 4036 3404
rect 4012 3336 4020 3344
rect 3996 3276 4004 3284
rect 3836 3216 3844 3224
rect 3980 3196 3988 3204
rect 3996 3176 4004 3184
rect 3884 3156 3892 3164
rect 3852 3116 3860 3124
rect 3788 3096 3796 3104
rect 3836 3096 3844 3104
rect 3740 2936 3748 2944
rect 3708 2916 3716 2924
rect 3644 2816 3652 2824
rect 3644 2716 3652 2724
rect 3532 2616 3540 2624
rect 3628 2596 3636 2604
rect 3500 2556 3508 2564
rect 3468 2536 3476 2544
rect 3468 2516 3476 2524
rect 3452 2476 3460 2484
rect 3468 2456 3476 2464
rect 3452 2436 3460 2444
rect 3420 2336 3428 2344
rect 3772 3076 3780 3084
rect 3804 3076 3812 3084
rect 3772 2976 3780 2984
rect 3804 2936 3812 2944
rect 3964 3116 3972 3124
rect 3916 3096 3924 3104
rect 3900 3076 3908 3084
rect 3900 3016 3908 3024
rect 3884 2976 3892 2984
rect 3868 2936 3876 2944
rect 3804 2876 3812 2884
rect 3820 2876 3828 2884
rect 3692 2836 3700 2844
rect 3724 2756 3732 2764
rect 3788 2816 3796 2824
rect 3852 2856 3860 2864
rect 3836 2836 3844 2844
rect 3852 2816 3860 2824
rect 3820 2736 3828 2744
rect 3692 2716 3700 2724
rect 3756 2716 3764 2724
rect 3772 2716 3780 2724
rect 3676 2696 3684 2704
rect 3724 2696 3732 2704
rect 3756 2696 3764 2704
rect 3820 2696 3828 2704
rect 3836 2696 3844 2704
rect 3660 2616 3668 2624
rect 3676 2616 3684 2624
rect 3676 2596 3684 2604
rect 3932 3076 3940 3084
rect 3980 3076 3988 3084
rect 3948 3056 3956 3064
rect 3964 3056 3972 3064
rect 4076 3456 4084 3464
rect 4156 3456 4164 3464
rect 4108 3416 4116 3424
rect 4140 3416 4148 3424
rect 4140 3376 4148 3384
rect 4060 3316 4068 3324
rect 4044 3176 4052 3184
rect 4028 3156 4036 3164
rect 4012 3116 4020 3124
rect 4044 3076 4052 3084
rect 4028 3056 4036 3064
rect 4012 2976 4020 2984
rect 3996 2956 4004 2964
rect 3900 2856 3908 2864
rect 3900 2776 3908 2784
rect 3964 2856 3972 2864
rect 3916 2736 3924 2744
rect 3868 2656 3876 2664
rect 3772 2636 3780 2644
rect 3868 2616 3876 2624
rect 3900 2576 3908 2584
rect 3916 2576 3924 2584
rect 3756 2556 3764 2564
rect 3516 2376 3524 2384
rect 3532 2356 3540 2364
rect 3484 2336 3492 2344
rect 3516 2336 3524 2344
rect 3404 2316 3412 2324
rect 3468 2316 3476 2324
rect 3516 2316 3524 2324
rect 3548 2316 3556 2324
rect 3404 2296 3412 2304
rect 3340 2256 3348 2264
rect 3372 2216 3380 2224
rect 3484 2276 3492 2284
rect 3468 2196 3476 2204
rect 3516 2196 3524 2204
rect 3404 2156 3412 2164
rect 3372 2136 3380 2144
rect 3500 2136 3508 2144
rect 3100 2016 3108 2024
rect 3004 1876 3012 1884
rect 3244 2036 3252 2044
rect 3404 1956 3412 1964
rect 3132 1896 3140 1904
rect 3180 1896 3188 1904
rect 3084 1856 3092 1864
rect 3038 1806 3046 1814
rect 3052 1806 3060 1814
rect 3066 1806 3074 1814
rect 3164 1816 3172 1824
rect 3212 1796 3220 1804
rect 2988 1756 2996 1764
rect 3148 1756 3156 1764
rect 3180 1756 3188 1764
rect 2972 1596 2980 1604
rect 2924 1556 2932 1564
rect 3148 1736 3156 1744
rect 3452 2036 3460 2044
rect 3436 1936 3444 1944
rect 3948 2696 3956 2704
rect 3964 2676 3972 2684
rect 3996 2836 4004 2844
rect 3996 2756 4004 2764
rect 4028 2916 4036 2924
rect 3980 2556 3988 2564
rect 4012 2656 4020 2664
rect 4076 3116 4084 3124
rect 4124 3116 4132 3124
rect 4076 3096 4084 3104
rect 4092 3076 4100 3084
rect 4108 3076 4116 3084
rect 4316 3416 4324 3424
rect 4316 3376 4324 3384
rect 4348 3376 4356 3384
rect 4172 3316 4180 3324
rect 4396 3336 4404 3344
rect 4364 3296 4372 3304
rect 4412 3296 4420 3304
rect 4348 3276 4356 3284
rect 4236 3196 4244 3204
rect 4332 3196 4340 3204
rect 4188 3156 4196 3164
rect 4172 3096 4180 3104
rect 4140 3056 4148 3064
rect 4124 3016 4132 3024
rect 4604 3476 4610 3484
rect 4610 3476 4612 3484
rect 5052 3656 5060 3664
rect 5116 3656 5124 3664
rect 4796 3596 4804 3604
rect 4828 3596 4836 3604
rect 5324 3596 5332 3604
rect 5324 3536 5332 3544
rect 5340 3536 5348 3544
rect 5212 3516 5220 3524
rect 4892 3496 4900 3504
rect 4956 3496 4964 3504
rect 5180 3496 5188 3504
rect 5068 3476 5076 3484
rect 4764 3456 4772 3464
rect 5100 3456 5108 3464
rect 5228 3456 5236 3464
rect 5292 3456 5300 3464
rect 4492 3436 4500 3444
rect 4524 3396 4532 3404
rect 4620 3396 4628 3404
rect 4556 3356 4564 3364
rect 4508 3336 4516 3344
rect 5260 3416 5268 3424
rect 5260 3396 5268 3404
rect 5308 3396 5316 3404
rect 4668 3356 4676 3364
rect 4908 3356 4916 3364
rect 5228 3356 5236 3364
rect 4652 3336 4660 3344
rect 4684 3336 4692 3344
rect 4892 3336 4900 3344
rect 4476 3296 4484 3304
rect 4508 3296 4516 3304
rect 4428 3236 4436 3244
rect 4540 3276 4548 3284
rect 4492 3236 4500 3244
rect 4444 3196 4452 3204
rect 4364 3176 4372 3184
rect 4508 3196 4516 3204
rect 4236 3096 4244 3104
rect 4380 3096 4388 3104
rect 4188 3016 4196 3024
rect 4204 3016 4212 3024
rect 4156 2996 4164 3004
rect 4156 2956 4164 2964
rect 4412 3056 4420 3064
rect 4604 3256 4612 3264
rect 4574 3206 4582 3214
rect 4588 3206 4596 3214
rect 4602 3206 4610 3214
rect 4604 3176 4612 3184
rect 4540 3156 4548 3164
rect 4572 3156 4580 3164
rect 4588 3156 4596 3164
rect 4492 3036 4500 3044
rect 4508 3036 4516 3044
rect 4428 3016 4436 3024
rect 4348 2996 4356 3004
rect 4380 2936 4388 2944
rect 4476 2936 4484 2944
rect 4060 2856 4068 2864
rect 4396 2916 4404 2924
rect 4348 2876 4356 2884
rect 4396 2856 4404 2864
rect 4204 2776 4212 2784
rect 4076 2736 4084 2744
rect 4108 2736 4116 2744
rect 4140 2736 4148 2744
rect 4172 2736 4180 2744
rect 4092 2696 4100 2704
rect 4124 2696 4132 2704
rect 4044 2676 4052 2684
rect 4028 2596 4036 2604
rect 3996 2516 4004 2524
rect 4076 2656 4084 2664
rect 4060 2636 4068 2644
rect 4060 2556 4068 2564
rect 4332 2756 4340 2764
rect 4476 2916 4484 2924
rect 4428 2776 4436 2784
rect 4348 2736 4356 2744
rect 4396 2736 4404 2744
rect 4444 2716 4452 2724
rect 4268 2696 4276 2704
rect 4316 2696 4324 2704
rect 4428 2696 4436 2704
rect 4460 2696 4468 2704
rect 4156 2676 4164 2684
rect 4172 2636 4180 2644
rect 4140 2596 4148 2604
rect 4156 2596 4164 2604
rect 4204 2596 4212 2604
rect 4140 2536 4148 2544
rect 4044 2516 4052 2524
rect 4076 2516 4084 2524
rect 4012 2456 4020 2464
rect 4092 2456 4100 2464
rect 4060 2436 4068 2444
rect 4108 2436 4116 2444
rect 3836 2396 3844 2404
rect 3884 2396 3892 2404
rect 3596 2376 3604 2384
rect 3996 2336 4004 2344
rect 4044 2336 4052 2344
rect 3580 2296 3588 2304
rect 3644 2296 3652 2304
rect 4012 2296 4020 2304
rect 3564 2276 3572 2284
rect 3708 2276 3716 2284
rect 3724 2276 3732 2284
rect 3804 2276 3812 2284
rect 3548 2256 3556 2264
rect 4108 2416 4116 2424
rect 4092 2356 4100 2364
rect 4076 2316 4084 2324
rect 4108 2296 4116 2304
rect 4108 2256 4116 2264
rect 4012 2216 4020 2224
rect 3676 2196 3684 2204
rect 3836 2196 3844 2204
rect 3564 2156 3572 2164
rect 3708 2156 3716 2164
rect 3868 2156 3876 2164
rect 3852 2136 3860 2144
rect 4108 2136 4116 2144
rect 3900 2116 3908 2124
rect 3884 2096 3892 2104
rect 3900 2036 3908 2044
rect 3740 2016 3748 2024
rect 3788 2016 3796 2024
rect 3676 1956 3684 1964
rect 3532 1936 3540 1944
rect 3580 1936 3588 1944
rect 3660 1936 3668 1944
rect 3820 1956 3828 1964
rect 3612 1896 3620 1904
rect 3660 1896 3668 1904
rect 3628 1876 3636 1884
rect 3404 1836 3412 1844
rect 3436 1836 3444 1844
rect 3372 1796 3380 1804
rect 3468 1816 3476 1824
rect 3532 1796 3540 1804
rect 3468 1776 3476 1784
rect 3500 1756 3508 1764
rect 3436 1736 3444 1744
rect 3484 1736 3492 1744
rect 3564 1776 3572 1784
rect 3564 1736 3572 1744
rect 3644 1736 3652 1744
rect 3852 1876 3860 1884
rect 3820 1856 3828 1864
rect 3804 1816 3812 1824
rect 3964 1876 3972 1884
rect 4188 2556 4196 2564
rect 4204 2516 4212 2524
rect 4140 2496 4148 2504
rect 4172 2496 4180 2504
rect 4252 2636 4260 2644
rect 4268 2616 4276 2624
rect 4236 2556 4244 2564
rect 4332 2676 4340 2684
rect 4412 2676 4420 2684
rect 4316 2636 4324 2644
rect 4300 2616 4308 2624
rect 4284 2596 4292 2604
rect 4300 2556 4308 2564
rect 4268 2536 4276 2544
rect 4236 2516 4244 2524
rect 4236 2496 4244 2504
rect 4284 2496 4292 2504
rect 4412 2596 4420 2604
rect 4364 2556 4372 2564
rect 4412 2556 4420 2564
rect 4396 2536 4404 2544
rect 4332 2496 4340 2504
rect 4220 2436 4228 2444
rect 4188 2416 4196 2424
rect 4284 2316 4292 2324
rect 4140 2296 4148 2304
rect 4156 2276 4164 2284
rect 4284 2276 4292 2284
rect 4300 2276 4308 2284
rect 4204 2136 4212 2144
rect 4252 2136 4260 2144
rect 4108 2096 4116 2104
rect 4124 2096 4132 2104
rect 4268 2096 4276 2104
rect 4172 1976 4180 1984
rect 4124 1936 4132 1944
rect 4028 1896 4036 1904
rect 4044 1876 4052 1884
rect 4044 1836 4052 1844
rect 3980 1796 3988 1804
rect 3708 1776 3716 1784
rect 3916 1776 3924 1784
rect 3692 1736 3700 1744
rect 3772 1736 3780 1744
rect 3260 1716 3268 1724
rect 3324 1716 3332 1724
rect 3452 1716 3460 1724
rect 3644 1716 3652 1724
rect 3692 1716 3700 1724
rect 3180 1656 3188 1664
rect 3196 1596 3204 1604
rect 3100 1496 3108 1504
rect 2988 1476 2996 1484
rect 2892 1456 2900 1464
rect 3084 1436 3092 1444
rect 2812 1396 2820 1404
rect 3038 1406 3046 1414
rect 3052 1406 3060 1414
rect 3066 1406 3074 1414
rect 2876 1336 2884 1344
rect 2972 1336 2980 1344
rect 2844 1316 2852 1324
rect 3068 1316 3076 1324
rect 2764 1296 2772 1304
rect 2828 1176 2836 1184
rect 2764 1136 2772 1144
rect 2844 1096 2852 1104
rect 2796 1076 2804 1084
rect 2812 1076 2820 1084
rect 2716 1016 2724 1024
rect 2556 996 2564 1004
rect 2604 996 2612 1004
rect 2668 996 2676 1004
rect 2508 956 2516 964
rect 2524 736 2532 744
rect 2588 736 2596 744
rect 2572 676 2580 684
rect 2700 916 2708 924
rect 2796 916 2804 924
rect 2908 1136 2916 1144
rect 3340 1696 3348 1704
rect 3420 1696 3428 1704
rect 3516 1676 3524 1684
rect 3404 1656 3412 1664
rect 3516 1536 3524 1544
rect 3436 1496 3444 1504
rect 3324 1476 3332 1484
rect 3228 1456 3236 1464
rect 3356 1456 3364 1464
rect 3484 1456 3492 1464
rect 3372 1376 3380 1384
rect 3340 1336 3348 1344
rect 3452 1236 3460 1244
rect 3308 1196 3316 1204
rect 3372 1196 3380 1204
rect 2924 1076 2932 1084
rect 3020 1076 3028 1084
rect 3180 1076 3188 1084
rect 2892 1056 2900 1064
rect 3084 1056 3092 1064
rect 2876 916 2884 924
rect 2844 796 2852 804
rect 3038 1006 3046 1014
rect 3052 1006 3060 1014
rect 3066 1006 3074 1014
rect 3004 956 3012 964
rect 3036 736 3044 744
rect 2780 676 2788 684
rect 2892 676 2900 684
rect 2924 676 2932 684
rect 2668 656 2676 664
rect 2748 656 2756 664
rect 2844 636 2852 644
rect 2524 616 2532 624
rect 2460 576 2468 584
rect 1788 536 1796 544
rect 1964 536 1972 544
rect 2156 536 2164 544
rect 2188 536 2196 544
rect 2236 536 2244 544
rect 1676 316 1684 324
rect 1802 316 1810 324
rect 1644 196 1652 204
rect 1628 156 1636 164
rect 2044 516 2052 524
rect 2316 556 2324 564
rect 2364 556 2372 564
rect 2412 556 2420 564
rect 2748 556 2756 564
rect 2284 536 2292 544
rect 2220 316 2228 324
rect 2172 296 2180 304
rect 2204 296 2212 304
rect 2380 536 2388 544
rect 2460 516 2468 524
rect 2364 496 2372 504
rect 2556 496 2564 504
rect 2460 396 2468 404
rect 2572 296 2580 304
rect 1996 276 2004 284
rect 2220 276 2228 284
rect 2284 276 2292 284
rect 1836 196 1844 204
rect 1852 196 1860 204
rect 1884 196 1892 204
rect 1660 136 1668 144
rect 1724 136 1732 144
rect 1964 156 1972 164
rect 1932 136 1940 144
rect 2316 216 2324 224
rect 2524 216 2532 224
rect 2780 536 2788 544
rect 2700 516 2708 524
rect 2796 516 2804 524
rect 3164 936 3166 944
rect 3166 936 3172 944
rect 3436 1096 3444 1104
rect 3340 1076 3348 1084
rect 3548 1696 3556 1704
rect 3628 1696 3636 1704
rect 3612 1676 3620 1684
rect 3564 1556 3572 1564
rect 3548 1476 3556 1484
rect 3548 1456 3556 1464
rect 3580 1536 3588 1544
rect 3596 1496 3604 1504
rect 3596 1356 3604 1364
rect 3532 1316 3540 1324
rect 3500 1096 3508 1104
rect 3532 1076 3540 1084
rect 3484 996 3492 1004
rect 3324 976 3332 984
rect 3308 956 3316 964
rect 3516 936 3524 944
rect 3580 916 3588 924
rect 3260 796 3268 804
rect 3372 796 3380 804
rect 3596 796 3604 804
rect 3100 636 3108 644
rect 2892 536 2900 544
rect 2828 496 2836 504
rect 3038 606 3046 614
rect 3052 606 3060 614
rect 3066 606 3074 614
rect 3548 736 3556 744
rect 3388 696 3396 704
rect 3196 656 3204 664
rect 3228 656 3236 664
rect 3388 636 3396 644
rect 3116 576 3124 584
rect 3196 576 3204 584
rect 3260 576 3268 584
rect 3084 536 3092 544
rect 2940 496 2948 504
rect 2892 436 2900 444
rect 2732 296 2740 304
rect 2604 196 2612 204
rect 2364 176 2372 184
rect 2492 176 2500 184
rect 2588 176 2596 184
rect 2172 136 2180 144
rect 2236 136 2244 144
rect 2332 136 2340 144
rect 2796 396 2804 404
rect 2844 296 2852 304
rect 2876 276 2884 284
rect 2748 196 2756 204
rect 2860 176 2868 184
rect 2828 136 2836 144
rect 3036 276 3038 284
rect 3038 276 3044 284
rect 3038 206 3046 214
rect 3052 206 3060 214
rect 3066 206 3074 214
rect 3132 436 3140 444
rect 3580 696 3588 704
rect 3980 1756 3988 1764
rect 4156 1856 4164 1864
rect 4124 1816 4132 1824
rect 4108 1756 4116 1764
rect 4140 1756 4148 1764
rect 4172 1756 4180 1764
rect 4012 1736 4020 1744
rect 3740 1696 3748 1704
rect 3804 1696 3812 1704
rect 3852 1696 3860 1704
rect 3804 1656 3812 1664
rect 3708 1556 3716 1564
rect 3660 1536 3668 1544
rect 3708 1516 3716 1524
rect 3772 1516 3780 1524
rect 3692 1456 3700 1464
rect 3644 1436 3652 1444
rect 3628 1376 3636 1384
rect 3692 1396 3700 1404
rect 3692 1376 3700 1384
rect 3628 1336 3636 1344
rect 3644 1336 3652 1344
rect 3676 1336 3684 1344
rect 3660 1316 3668 1324
rect 3660 1156 3668 1164
rect 3692 1156 3700 1164
rect 3644 1076 3652 1084
rect 3628 1016 3636 1024
rect 3612 776 3620 784
rect 3644 776 3652 784
rect 3692 1136 3700 1144
rect 3692 1076 3700 1084
rect 3692 916 3700 924
rect 3676 796 3684 804
rect 3660 696 3668 704
rect 3436 676 3444 684
rect 3532 676 3540 684
rect 3564 676 3572 684
rect 3612 676 3620 684
rect 3420 576 3428 584
rect 3276 496 3284 504
rect 3276 316 3284 324
rect 3148 296 3156 304
rect 3148 276 3156 284
rect 3756 1496 3764 1504
rect 3740 1436 3748 1444
rect 4092 1696 4100 1704
rect 4172 1696 4180 1704
rect 4156 1676 4164 1684
rect 4204 1676 4212 1684
rect 4076 1636 4084 1644
rect 4060 1616 4068 1624
rect 4044 1576 4052 1584
rect 3900 1556 3908 1564
rect 4028 1556 4036 1564
rect 3980 1536 3988 1544
rect 4044 1536 4052 1544
rect 3852 1516 3860 1524
rect 3884 1516 3892 1524
rect 3964 1516 3972 1524
rect 4012 1516 4020 1524
rect 3852 1496 3860 1504
rect 3932 1496 3940 1504
rect 3996 1496 4004 1504
rect 3820 1476 3828 1484
rect 3900 1476 3908 1484
rect 3804 1416 3812 1424
rect 3948 1476 3956 1484
rect 3932 1396 3940 1404
rect 3820 1356 3828 1364
rect 3948 1356 3956 1364
rect 3772 1336 3780 1344
rect 3916 1336 3924 1344
rect 3740 1276 3748 1284
rect 3948 1236 3956 1244
rect 3772 1216 3780 1224
rect 4012 1216 4020 1224
rect 3868 1096 3876 1104
rect 3836 1076 3844 1084
rect 3820 996 3828 1004
rect 3868 996 3876 1004
rect 4108 1616 4116 1624
rect 4092 1576 4100 1584
rect 4060 1496 4068 1504
rect 4124 1576 4132 1584
rect 4140 1516 4148 1524
rect 4124 1476 4132 1484
rect 4172 1476 4180 1484
rect 4124 1396 4132 1404
rect 4108 1376 4116 1384
rect 4092 1336 4100 1344
rect 4060 1316 4068 1324
rect 4108 1276 4116 1284
rect 4060 1216 4068 1224
rect 4044 1036 4052 1044
rect 4028 1016 4036 1024
rect 3980 836 3988 844
rect 3788 816 3796 824
rect 3980 816 3988 824
rect 3868 736 3876 744
rect 3900 736 3908 744
rect 4076 936 4084 944
rect 4140 1356 4148 1364
rect 4236 1776 4244 1784
rect 4508 2996 4516 3004
rect 4572 2956 4580 2964
rect 4508 2936 4516 2944
rect 4780 3316 4788 3324
rect 4684 3296 4692 3304
rect 4700 3296 4708 3304
rect 4668 3276 4676 3284
rect 4652 3156 4660 3164
rect 4668 3096 4676 3104
rect 4636 2936 4644 2944
rect 4620 2916 4628 2924
rect 4524 2876 4532 2884
rect 4636 2876 4644 2884
rect 4716 3256 4724 3264
rect 4844 3316 4852 3324
rect 4828 3296 4836 3304
rect 4876 3256 4884 3264
rect 4812 3176 4820 3184
rect 4780 3136 4788 3144
rect 4812 3136 4820 3144
rect 4844 3136 4852 3144
rect 4748 3116 4756 3124
rect 4796 3116 4804 3124
rect 4876 3156 4884 3164
rect 4860 3116 4868 3124
rect 4716 3096 4724 3104
rect 4764 3096 4772 3104
rect 4796 3056 4804 3064
rect 4812 3036 4820 3044
rect 4764 3016 4772 3024
rect 4860 3016 4868 3024
rect 4700 2996 4708 3004
rect 4716 2996 4724 3004
rect 4668 2956 4676 2964
rect 4684 2916 4692 2924
rect 4668 2876 4676 2884
rect 4636 2836 4644 2844
rect 4652 2836 4660 2844
rect 4574 2806 4582 2814
rect 4588 2806 4596 2814
rect 4602 2806 4610 2814
rect 4508 2736 4516 2744
rect 4540 2716 4548 2724
rect 4396 2496 4404 2504
rect 4364 2396 4372 2404
rect 4348 2236 4356 2244
rect 4476 2536 4484 2544
rect 4540 2596 4548 2604
rect 4508 2556 4516 2564
rect 4652 2776 4660 2784
rect 4732 2936 4740 2944
rect 4748 2936 4756 2944
rect 4796 2936 4804 2944
rect 4828 2936 4836 2944
rect 4780 2916 4788 2924
rect 4716 2856 4724 2864
rect 4684 2776 4692 2784
rect 4668 2756 4676 2764
rect 4636 2616 4644 2624
rect 4524 2536 4532 2544
rect 4556 2536 4564 2544
rect 4572 2536 4580 2544
rect 4524 2516 4532 2524
rect 4588 2516 4596 2524
rect 4476 2456 4484 2464
rect 4444 2256 4452 2264
rect 4524 2496 4532 2504
rect 4556 2496 4564 2504
rect 4524 2456 4532 2464
rect 4652 2596 4660 2604
rect 4812 2836 4820 2844
rect 4796 2816 4804 2824
rect 4748 2796 4756 2804
rect 4748 2756 4756 2764
rect 4780 2716 4788 2724
rect 4748 2696 4756 2704
rect 4716 2616 4724 2624
rect 4668 2576 4676 2584
rect 4716 2576 4724 2584
rect 4652 2496 4660 2504
rect 4700 2536 4708 2544
rect 4780 2696 4788 2704
rect 4764 2676 4772 2684
rect 4764 2656 4772 2664
rect 4796 2656 4804 2664
rect 4716 2516 4724 2524
rect 4652 2476 4660 2484
rect 4668 2476 4676 2484
rect 4636 2416 4644 2424
rect 4574 2406 4582 2414
rect 4588 2406 4596 2414
rect 4602 2406 4610 2414
rect 4540 2396 4548 2404
rect 4508 2316 4516 2324
rect 4636 2376 4644 2384
rect 4524 2296 4532 2304
rect 4476 2276 4484 2284
rect 4556 2276 4564 2284
rect 4460 2236 4468 2244
rect 4412 2196 4420 2204
rect 4588 2236 4596 2244
rect 4604 2196 4612 2204
rect 4636 2196 4644 2204
rect 4780 2616 4788 2624
rect 4828 2736 4836 2744
rect 4828 2716 4836 2724
rect 4956 3316 4964 3324
rect 5004 3316 5012 3324
rect 4940 3276 4948 3284
rect 4908 3216 4916 3224
rect 4908 3176 4916 3184
rect 5100 3316 5108 3324
rect 5260 3316 5268 3324
rect 5052 3296 5060 3304
rect 5020 3176 5028 3184
rect 5068 3196 5076 3204
rect 5004 3156 5012 3164
rect 5020 3136 5028 3144
rect 4956 3096 4964 3104
rect 4988 3096 4996 3104
rect 5004 3096 5012 3104
rect 5052 3096 5060 3104
rect 4908 3076 4916 3084
rect 4924 3056 4932 3064
rect 4892 2996 4900 3004
rect 4972 3016 4980 3024
rect 4892 2976 4900 2984
rect 4940 2976 4948 2984
rect 4892 2936 4900 2944
rect 4876 2816 4884 2824
rect 4956 2936 4964 2944
rect 5004 3076 5012 3084
rect 5084 3136 5092 3144
rect 5180 3216 5188 3224
rect 5244 3216 5252 3224
rect 5132 3176 5140 3184
rect 5212 3196 5220 3204
rect 5228 3176 5236 3184
rect 5116 3116 5124 3124
rect 5212 3116 5220 3124
rect 5116 3096 5124 3104
rect 5020 2996 5028 3004
rect 5004 2956 5012 2964
rect 4924 2916 4932 2924
rect 4940 2916 4948 2924
rect 4988 2916 4996 2924
rect 4908 2796 4916 2804
rect 4956 2896 4964 2904
rect 4972 2816 4980 2824
rect 4876 2756 4884 2764
rect 4860 2696 4868 2704
rect 4892 2736 4900 2744
rect 4860 2676 4868 2684
rect 4844 2656 4852 2664
rect 4844 2616 4852 2624
rect 4796 2556 4804 2564
rect 4828 2556 4836 2564
rect 4956 2696 4964 2704
rect 5004 2856 5012 2864
rect 5004 2776 5012 2784
rect 5068 2956 5076 2964
rect 5068 2816 5076 2824
rect 5052 2796 5060 2804
rect 5020 2716 5028 2724
rect 4972 2676 4980 2684
rect 4956 2656 4964 2664
rect 4940 2636 4948 2644
rect 4924 2576 4932 2584
rect 4956 2616 4964 2624
rect 4844 2516 4852 2524
rect 4828 2496 4836 2504
rect 4844 2456 4852 2464
rect 4812 2416 4820 2424
rect 4828 2416 4836 2424
rect 4748 2396 4756 2404
rect 4764 2336 4772 2344
rect 4700 2316 4708 2324
rect 4748 2316 4756 2324
rect 4716 2276 4724 2284
rect 4668 2256 4676 2264
rect 4684 2236 4692 2244
rect 4780 2316 4788 2324
rect 4812 2316 4820 2324
rect 4844 2316 4852 2324
rect 4780 2296 4788 2304
rect 4828 2276 4836 2284
rect 4748 2196 4756 2204
rect 4828 2176 4836 2184
rect 4556 2156 4564 2164
rect 4812 2156 4820 2164
rect 4332 1996 4340 2004
rect 4316 1836 4324 1844
rect 4892 2556 4900 2564
rect 4892 2536 4900 2544
rect 4876 2336 4884 2344
rect 4876 2316 4884 2324
rect 4972 2536 4980 2544
rect 4956 2496 4964 2504
rect 4908 2436 4916 2444
rect 4908 2396 4916 2404
rect 4956 2376 4964 2384
rect 4924 2336 4932 2344
rect 4956 2316 4964 2324
rect 4940 2296 4948 2304
rect 4972 2296 4980 2304
rect 4972 2196 4980 2204
rect 5036 2696 5044 2704
rect 5004 2656 5012 2664
rect 5020 2636 5028 2644
rect 5020 2616 5028 2624
rect 5052 2636 5060 2644
rect 5004 2596 5012 2604
rect 5036 2596 5044 2604
rect 5164 3076 5172 3084
rect 5116 3056 5124 3064
rect 5212 3016 5220 3024
rect 5212 2976 5220 2984
rect 5100 2736 5108 2744
rect 5132 2936 5140 2944
rect 5180 2936 5188 2944
rect 5212 2916 5220 2924
rect 5180 2896 5188 2904
rect 5132 2816 5140 2824
rect 5084 2696 5092 2704
rect 5084 2636 5092 2644
rect 5020 2576 5028 2584
rect 5068 2576 5076 2584
rect 5052 2556 5060 2564
rect 5212 2856 5220 2864
rect 5196 2776 5204 2784
rect 5164 2736 5172 2744
rect 5164 2696 5172 2704
rect 5228 2796 5236 2804
rect 5276 3136 5284 3144
rect 5324 3136 5332 3144
rect 5260 3096 5268 3104
rect 5292 3116 5300 3124
rect 5404 3736 5412 3744
rect 5548 3736 5556 3744
rect 5580 3716 5588 3724
rect 5516 3656 5524 3664
rect 5548 3656 5556 3664
rect 5548 3596 5556 3604
rect 5420 3576 5428 3584
rect 5388 3556 5396 3564
rect 5404 3516 5412 3524
rect 5372 3356 5380 3364
rect 5372 3336 5380 3344
rect 5356 3316 5364 3324
rect 5388 3116 5396 3124
rect 5340 3096 5348 3104
rect 5292 3076 5300 3084
rect 5260 3036 5268 3044
rect 5260 3016 5268 3024
rect 5260 2916 5268 2924
rect 5516 3556 5524 3564
rect 5724 3896 5732 3904
rect 5676 3876 5684 3884
rect 5724 3876 5732 3884
rect 5612 3856 5620 3864
rect 5660 3836 5668 3844
rect 5628 3756 5636 3764
rect 5644 3736 5652 3744
rect 5596 3536 5604 3544
rect 5580 3516 5588 3524
rect 5612 3516 5620 3524
rect 5436 3476 5444 3484
rect 5596 3476 5604 3484
rect 5452 3396 5460 3404
rect 5436 3316 5444 3324
rect 5708 3836 5716 3844
rect 5692 3736 5700 3744
rect 5676 3496 5684 3504
rect 5660 3476 5668 3484
rect 5644 3376 5652 3384
rect 5564 3356 5572 3364
rect 5820 4156 5828 4164
rect 5916 4156 5924 4164
rect 5884 4136 5892 4144
rect 5772 3716 5780 3724
rect 5740 3616 5748 3624
rect 6012 4156 6020 4164
rect 6044 3996 6052 4004
rect 6060 3996 6068 4004
rect 5868 3896 5876 3904
rect 5932 3756 5940 3764
rect 5820 3716 5828 3724
rect 5932 3716 5940 3724
rect 5900 3476 5908 3484
rect 5724 3376 5732 3384
rect 5708 3336 5716 3344
rect 5788 3316 5796 3324
rect 5852 3416 5860 3424
rect 5884 3356 5892 3364
rect 6124 3956 6132 3964
rect 5980 3496 5982 3504
rect 5982 3496 5988 3504
rect 6044 3496 6052 3504
rect 5948 3376 5956 3384
rect 5900 3336 5908 3344
rect 5852 3316 5860 3324
rect 5932 3316 5940 3324
rect 6012 3476 6020 3484
rect 6060 3476 6068 3484
rect 5980 3356 5988 3364
rect 5996 3316 6004 3324
rect 5468 3236 5476 3244
rect 5756 3116 5764 3124
rect 5628 3076 5636 3084
rect 5420 3056 5428 3064
rect 5340 3036 5348 3044
rect 5372 2956 5380 2964
rect 5356 2936 5364 2944
rect 5420 2936 5428 2944
rect 5308 2896 5316 2904
rect 5308 2816 5316 2824
rect 5292 2796 5300 2804
rect 5324 2776 5332 2784
rect 5276 2756 5284 2764
rect 5276 2696 5284 2704
rect 5148 2656 5156 2664
rect 5164 2656 5172 2664
rect 5244 2656 5252 2664
rect 5212 2636 5220 2644
rect 5196 2616 5204 2624
rect 5148 2596 5156 2604
rect 5228 2596 5236 2604
rect 5116 2576 5124 2584
rect 5180 2576 5188 2584
rect 5100 2556 5108 2564
rect 5084 2516 5092 2524
rect 5116 2516 5124 2524
rect 5020 2496 5028 2504
rect 5004 2456 5012 2464
rect 5004 2416 5012 2424
rect 5052 2456 5060 2464
rect 5036 2416 5044 2424
rect 5068 2376 5076 2384
rect 5052 2356 5060 2364
rect 5068 2356 5076 2364
rect 5004 2296 5012 2304
rect 5004 2216 5012 2224
rect 5100 2456 5108 2464
rect 5084 2336 5092 2344
rect 5068 2296 5076 2304
rect 5084 2276 5092 2284
rect 5180 2516 5188 2524
rect 5196 2516 5204 2524
rect 5164 2496 5172 2504
rect 5148 2396 5156 2404
rect 5116 2356 5124 2364
rect 5228 2396 5236 2404
rect 5196 2336 5204 2344
rect 5308 2596 5316 2604
rect 5292 2576 5300 2584
rect 5276 2516 5284 2524
rect 5260 2356 5268 2364
rect 5244 2316 5252 2324
rect 5132 2276 5140 2284
rect 5052 2196 5060 2204
rect 5116 2156 5124 2164
rect 4460 2136 4468 2144
rect 4844 2116 4852 2124
rect 4892 2096 4900 2104
rect 5196 2276 5204 2284
rect 5196 2256 5204 2264
rect 5260 2256 5268 2264
rect 5180 2216 5188 2224
rect 5228 2216 5236 2224
rect 5164 2136 5172 2144
rect 5308 2356 5316 2364
rect 5308 2336 5316 2344
rect 5308 2316 5316 2324
rect 5308 2296 5316 2304
rect 5308 2236 5316 2244
rect 5292 2216 5300 2224
rect 5196 2116 5204 2124
rect 5388 2896 5396 2904
rect 5740 3056 5748 3064
rect 5548 3036 5556 3044
rect 5660 3036 5668 3044
rect 5452 2836 5460 2844
rect 5372 2796 5380 2804
rect 5340 2756 5348 2764
rect 5340 2736 5348 2744
rect 5404 2716 5412 2724
rect 5452 2716 5460 2724
rect 5340 2696 5348 2704
rect 5356 2616 5364 2624
rect 5340 2556 5348 2564
rect 5356 2556 5364 2564
rect 5388 2696 5396 2704
rect 5436 2656 5444 2664
rect 5372 2536 5380 2544
rect 5420 2616 5428 2624
rect 5420 2556 5428 2564
rect 5724 3016 5732 3024
rect 5580 2956 5588 2964
rect 5788 3056 5796 3064
rect 5548 2936 5556 2944
rect 5500 2716 5508 2724
rect 5484 2676 5492 2684
rect 5468 2596 5476 2604
rect 5468 2576 5476 2584
rect 5452 2556 5460 2564
rect 5852 3116 5860 3124
rect 5852 3076 5860 3084
rect 5900 3076 5908 3084
rect 5996 3076 6004 3084
rect 5820 3056 5828 3064
rect 5804 3036 5812 3044
rect 5932 3056 5940 3064
rect 5932 3036 5940 3044
rect 5900 3016 5908 3024
rect 5900 2996 5908 3004
rect 5948 2996 5956 3004
rect 5580 2916 5588 2924
rect 5564 2756 5572 2764
rect 5676 2756 5684 2764
rect 5644 2736 5652 2744
rect 5548 2676 5556 2684
rect 5580 2636 5588 2644
rect 5388 2516 5396 2524
rect 5388 2496 5396 2504
rect 5452 2456 5460 2464
rect 5356 2436 5364 2444
rect 5372 2416 5380 2424
rect 5404 2376 5412 2384
rect 5436 2336 5444 2344
rect 5452 2316 5460 2324
rect 5484 2316 5492 2324
rect 5500 2316 5508 2324
rect 5388 2296 5396 2304
rect 5420 2296 5428 2304
rect 5340 2276 5348 2284
rect 5548 2376 5556 2384
rect 5516 2256 5524 2264
rect 5484 2236 5492 2244
rect 5468 2216 5476 2224
rect 5388 2196 5396 2204
rect 5324 2176 5332 2184
rect 6028 3376 6036 3384
rect 6124 3696 6132 3704
rect 6124 3496 6132 3504
rect 6108 3396 6116 3404
rect 6028 3356 6036 3364
rect 6076 3356 6084 3364
rect 6076 3336 6084 3344
rect 6108 3336 6116 3344
rect 6044 3056 6052 3064
rect 5724 2756 5732 2764
rect 5756 2756 5764 2764
rect 5788 2756 5796 2764
rect 5756 2736 5764 2744
rect 5692 2696 5700 2704
rect 5788 2696 5796 2704
rect 5868 2696 5876 2704
rect 5644 2676 5652 2684
rect 5772 2676 5780 2684
rect 5612 2576 5620 2584
rect 5772 2596 5780 2604
rect 5708 2576 5716 2584
rect 5644 2536 5652 2544
rect 5612 2476 5620 2484
rect 5660 2376 5668 2384
rect 5660 2356 5668 2364
rect 5580 2296 5588 2304
rect 5628 2316 5636 2324
rect 5628 2296 5636 2304
rect 6028 2816 6036 2824
rect 6060 2816 6068 2824
rect 5980 2676 5988 2684
rect 6044 2676 6052 2684
rect 5868 2656 5876 2664
rect 5948 2656 5956 2664
rect 5900 2536 5908 2544
rect 5596 2276 5604 2284
rect 5724 2276 5732 2284
rect 5692 2216 5700 2224
rect 5532 2196 5540 2204
rect 5564 2196 5572 2204
rect 5580 2176 5588 2184
rect 5676 2156 5684 2164
rect 5356 2136 5364 2144
rect 5468 2136 5476 2144
rect 5548 2136 5556 2144
rect 4574 2006 4582 2014
rect 4588 2006 4596 2014
rect 4602 2006 4610 2014
rect 4428 1996 4436 2004
rect 4508 1996 4516 2004
rect 4668 1896 4676 1904
rect 4348 1876 4356 1884
rect 4380 1876 4388 1884
rect 4508 1876 4516 1884
rect 4380 1856 4388 1864
rect 4332 1736 4340 1744
rect 4316 1716 4324 1724
rect 4332 1716 4340 1724
rect 4284 1556 4292 1564
rect 4284 1516 4292 1524
rect 4316 1516 4324 1524
rect 4300 1496 4308 1504
rect 4316 1436 4324 1444
rect 4316 1376 4324 1384
rect 4332 1336 4340 1344
rect 4332 1296 4340 1304
rect 4268 1256 4276 1264
rect 4252 1196 4260 1204
rect 4332 1276 4340 1284
rect 4284 1216 4292 1224
rect 4220 1176 4228 1184
rect 4284 1156 4292 1164
rect 4316 1156 4324 1164
rect 4220 1116 4228 1124
rect 4156 1096 4164 1104
rect 4188 1102 4196 1104
rect 4188 1096 4196 1102
rect 4188 996 4196 1004
rect 4140 936 4148 944
rect 4284 1096 4292 1104
rect 4204 956 4212 964
rect 4060 836 4068 844
rect 3708 716 3716 724
rect 3740 716 3748 724
rect 3820 716 3828 724
rect 3948 716 3956 724
rect 4012 716 4020 724
rect 3756 696 3764 704
rect 3628 656 3636 664
rect 3676 656 3684 664
rect 3724 656 3732 664
rect 3708 636 3716 644
rect 3708 616 3716 624
rect 3772 616 3780 624
rect 3532 596 3540 604
rect 3548 576 3556 584
rect 3628 576 3636 584
rect 3676 576 3684 584
rect 3612 556 3620 564
rect 3692 556 3700 564
rect 4108 736 4116 744
rect 4108 696 4116 704
rect 4076 676 4084 684
rect 4156 876 4164 884
rect 4476 1816 4484 1824
rect 4508 1816 4516 1824
rect 4460 1736 4468 1744
rect 4444 1696 4452 1704
rect 4492 1716 4500 1724
rect 4460 1676 4468 1684
rect 4524 1696 4532 1704
rect 4524 1676 4532 1684
rect 4572 1676 4580 1684
rect 4508 1536 4516 1544
rect 4476 1516 4484 1524
rect 4508 1516 4516 1524
rect 4412 1496 4420 1504
rect 4476 1496 4484 1504
rect 4380 1456 4388 1464
rect 4396 1396 4404 1404
rect 4412 1356 4420 1364
rect 4380 1336 4388 1344
rect 4364 1216 4372 1224
rect 4444 1316 4452 1324
rect 4412 1136 4420 1144
rect 4396 1116 4404 1124
rect 4348 1016 4356 1024
rect 4284 976 4292 984
rect 4252 916 4260 924
rect 4252 896 4260 904
rect 4252 836 4260 844
rect 4236 796 4244 804
rect 4140 716 4148 724
rect 4172 716 4180 724
rect 4204 716 4212 724
rect 4156 676 4164 684
rect 4124 656 4132 664
rect 3932 636 3940 644
rect 4092 636 4100 644
rect 4172 636 4180 644
rect 3996 616 4004 624
rect 4188 616 4196 624
rect 3900 596 3908 604
rect 3884 576 3892 584
rect 3852 556 3860 564
rect 3884 556 3892 564
rect 3468 536 3476 544
rect 3564 536 3572 544
rect 3788 536 3796 544
rect 3852 536 3860 544
rect 3484 516 3492 524
rect 3452 496 3460 504
rect 3404 456 3412 464
rect 3388 316 3396 324
rect 3468 456 3476 464
rect 3548 456 3556 464
rect 3612 516 3620 524
rect 3644 516 3652 524
rect 3756 516 3764 524
rect 3580 496 3588 504
rect 3628 496 3636 504
rect 3452 276 3460 284
rect 3484 276 3492 284
rect 3356 256 3364 264
rect 3468 256 3476 264
rect 3276 196 3284 204
rect 3340 196 3348 204
rect 3116 176 3124 184
rect 3308 176 3316 184
rect 3532 256 3540 264
rect 3596 256 3604 264
rect 3612 256 3620 264
rect 3628 256 3636 264
rect 3500 156 3508 164
rect 3596 156 3604 164
rect 3596 136 3604 144
rect 3788 276 3796 284
rect 3756 216 3764 224
rect 3804 216 3812 224
rect 3948 176 3956 184
rect 3964 176 3972 184
rect 3804 156 3812 164
rect 3772 136 3780 144
rect 4044 596 4052 604
rect 4092 556 4100 564
rect 4140 536 4148 544
rect 4076 276 4084 284
rect 4284 876 4292 884
rect 4332 936 4340 944
rect 4380 936 4388 944
rect 4412 1096 4420 1104
rect 4540 1656 4548 1664
rect 4574 1606 4582 1614
rect 4588 1606 4596 1614
rect 4602 1606 4610 1614
rect 4604 1556 4612 1564
rect 4556 1536 4564 1544
rect 4652 1696 4660 1704
rect 4700 1756 4708 1764
rect 4700 1736 4708 1744
rect 4684 1656 4692 1664
rect 4716 1716 4724 1724
rect 4700 1596 4708 1604
rect 4668 1556 4676 1564
rect 4700 1556 4708 1564
rect 4668 1496 4676 1504
rect 4636 1436 4644 1444
rect 4636 1376 4644 1384
rect 4524 1336 4532 1344
rect 4492 1316 4500 1324
rect 4508 1316 4516 1324
rect 4476 1256 4484 1264
rect 4460 1196 4468 1204
rect 4444 1156 4452 1164
rect 4460 1136 4468 1144
rect 4444 1116 4452 1124
rect 4428 1076 4436 1084
rect 4412 996 4420 1004
rect 4332 916 4340 924
rect 4364 916 4372 924
rect 4412 916 4420 924
rect 4524 1296 4532 1304
rect 4508 1276 4516 1284
rect 4508 1156 4516 1164
rect 4444 1056 4452 1064
rect 4476 1056 4484 1064
rect 4492 1056 4500 1064
rect 4492 1036 4500 1044
rect 4574 1206 4582 1214
rect 4588 1206 4596 1214
rect 4602 1206 4610 1214
rect 4556 1096 4564 1104
rect 4524 1036 4532 1044
rect 4508 996 4516 1004
rect 4476 956 4484 964
rect 4524 956 4532 964
rect 4476 936 4484 944
rect 4300 836 4308 844
rect 4268 756 4276 764
rect 4252 716 4260 724
rect 4236 696 4244 704
rect 4268 696 4276 704
rect 4220 676 4228 684
rect 4252 676 4260 684
rect 4284 676 4292 684
rect 4236 656 4244 664
rect 4204 596 4212 604
rect 4220 596 4228 604
rect 4268 556 4276 564
rect 4236 516 4244 524
rect 4220 496 4228 504
rect 4268 316 4276 324
rect 4316 516 4324 524
rect 4316 496 4324 504
rect 4300 336 4308 344
rect 4236 296 4244 304
rect 4268 296 4276 304
rect 4284 296 4292 304
rect 4316 296 4324 304
rect 4236 216 4244 224
rect 4092 156 4100 164
rect 4108 136 4116 144
rect 4380 776 4388 784
rect 4444 896 4452 904
rect 4396 696 4404 704
rect 4460 796 4468 804
rect 4444 736 4452 744
rect 4460 736 4468 744
rect 4444 716 4452 724
rect 4348 596 4356 604
rect 4492 916 4500 924
rect 4492 896 4500 904
rect 4524 716 4532 724
rect 4476 676 4484 684
rect 4412 636 4420 644
rect 4348 576 4356 584
rect 4396 576 4404 584
rect 4364 556 4372 564
rect 4444 556 4452 564
rect 4460 556 4468 564
rect 4396 536 4404 544
rect 4412 536 4420 544
rect 4348 496 4356 504
rect 4364 316 4372 324
rect 4332 216 4340 224
rect 4332 196 4340 204
rect 4252 136 4260 144
rect 1004 116 1012 124
rect 1164 116 1172 124
rect 1228 118 1236 124
rect 1228 116 1236 118
rect 1324 116 1332 124
rect 1772 116 1780 124
rect 1836 116 1844 124
rect 2044 116 2052 124
rect 2236 116 2244 124
rect 2972 116 2980 124
rect 3180 116 3188 124
rect 4300 116 4308 124
rect 4396 516 4404 524
rect 4396 496 4404 504
rect 4492 596 4500 604
rect 4620 1076 4628 1084
rect 4636 1016 4644 1024
rect 4716 1476 4724 1484
rect 4716 1456 4724 1464
rect 4684 1096 4692 1104
rect 4796 1956 4804 1964
rect 5036 2096 5044 2104
rect 5116 2096 5124 2104
rect 5164 2056 5172 2064
rect 5116 2036 5124 2044
rect 5036 1936 5044 1944
rect 4764 1916 4772 1924
rect 4956 1916 4964 1924
rect 4988 1916 4996 1924
rect 5020 1916 5028 1924
rect 5100 1916 5108 1924
rect 4764 1896 4772 1904
rect 4796 1902 4804 1904
rect 4796 1896 4804 1902
rect 4940 1896 4948 1904
rect 4748 1776 4756 1784
rect 4812 1876 4820 1884
rect 5004 1836 5012 1844
rect 4972 1796 4980 1804
rect 4828 1736 4836 1744
rect 4924 1736 4932 1744
rect 5132 1896 5140 1904
rect 5180 1936 5188 1944
rect 5260 1936 5268 1944
rect 5196 1876 5204 1884
rect 5372 1916 5380 1924
rect 5292 1896 5300 1904
rect 5036 1856 5044 1864
rect 5228 1856 5236 1864
rect 5452 1856 5460 1864
rect 5164 1836 5172 1844
rect 5148 1816 5156 1824
rect 5100 1796 5108 1804
rect 4988 1776 4996 1784
rect 5020 1776 5028 1784
rect 4780 1716 4788 1724
rect 4748 1696 4756 1704
rect 4764 1696 4772 1704
rect 4892 1696 4900 1704
rect 4844 1676 4852 1684
rect 4860 1676 4868 1684
rect 4924 1676 4932 1684
rect 4828 1656 4836 1664
rect 4796 1576 4804 1584
rect 4844 1556 4852 1564
rect 4876 1536 4884 1544
rect 4892 1516 4900 1524
rect 4908 1496 4916 1504
rect 4812 1476 4820 1484
rect 4892 1476 4900 1484
rect 4828 1456 4836 1464
rect 4860 1456 4868 1464
rect 4780 1436 4788 1444
rect 4732 1376 4740 1384
rect 4732 1356 4740 1364
rect 4796 1376 4804 1384
rect 4812 1376 4820 1384
rect 4764 1336 4772 1344
rect 4780 1336 4788 1344
rect 4748 1276 4756 1284
rect 4716 1136 4724 1144
rect 4764 1096 4772 1104
rect 4716 1076 4724 1084
rect 4780 1076 4788 1084
rect 4684 1056 4692 1064
rect 4636 956 4644 964
rect 4668 956 4676 964
rect 4556 936 4564 944
rect 4556 916 4564 924
rect 4572 896 4580 904
rect 4732 936 4740 944
rect 4652 916 4660 924
rect 4748 916 4756 924
rect 4588 856 4596 864
rect 4574 806 4582 814
rect 4588 806 4596 814
rect 4602 806 4610 814
rect 4556 756 4564 764
rect 4572 756 4580 764
rect 4636 736 4644 744
rect 4540 656 4548 664
rect 4524 556 4532 564
rect 4556 556 4564 564
rect 4508 536 4516 544
rect 4764 896 4772 904
rect 4828 1336 4836 1344
rect 4844 1336 4852 1344
rect 4844 1296 4852 1304
rect 4812 1216 4820 1224
rect 4812 1096 4820 1104
rect 4828 1096 4836 1104
rect 4828 996 4836 1004
rect 4892 1336 4900 1344
rect 4876 1296 4884 1304
rect 4876 1196 4884 1204
rect 4892 1176 4900 1184
rect 4892 1096 4900 1104
rect 4940 1316 4948 1324
rect 4924 1296 4932 1304
rect 4972 1416 4980 1424
rect 5676 2116 5684 2124
rect 5884 2376 5892 2384
rect 5964 2336 5972 2344
rect 5852 2256 5860 2264
rect 5916 2196 5924 2204
rect 5788 2136 5796 2144
rect 5772 2116 5780 2124
rect 5740 2096 5748 2104
rect 5724 2036 5732 2044
rect 5772 1976 5780 1984
rect 5756 1916 5764 1924
rect 5596 1896 5604 1904
rect 5660 1896 5668 1904
rect 5548 1856 5556 1864
rect 5452 1756 5460 1764
rect 5516 1756 5524 1764
rect 5068 1736 5076 1744
rect 5212 1736 5220 1744
rect 5292 1736 5300 1744
rect 5436 1736 5444 1744
rect 5020 1656 5028 1664
rect 5116 1696 5124 1704
rect 5276 1716 5284 1724
rect 5372 1716 5380 1724
rect 5068 1596 5076 1604
rect 5132 1596 5140 1604
rect 5052 1536 5060 1544
rect 5100 1516 5108 1524
rect 5084 1496 5092 1504
rect 5196 1696 5204 1704
rect 5244 1696 5252 1704
rect 5196 1656 5204 1664
rect 5180 1576 5188 1584
rect 5340 1696 5348 1704
rect 5292 1676 5300 1684
rect 5292 1636 5300 1644
rect 5244 1556 5252 1564
rect 5164 1516 5172 1524
rect 5388 1596 5396 1604
rect 5420 1676 5428 1684
rect 5276 1496 5284 1504
rect 5324 1496 5332 1504
rect 5372 1496 5380 1504
rect 5404 1496 5412 1504
rect 5036 1476 5044 1484
rect 5068 1476 5076 1484
rect 5324 1476 5332 1484
rect 5004 1456 5012 1464
rect 5020 1396 5028 1404
rect 5020 1376 5028 1384
rect 5244 1456 5252 1464
rect 5356 1456 5364 1464
rect 5180 1376 5188 1384
rect 5132 1356 5140 1364
rect 5148 1356 5156 1364
rect 5084 1336 5092 1344
rect 5116 1336 5124 1344
rect 5068 1256 5076 1264
rect 5036 1216 5044 1224
rect 5052 1196 5060 1204
rect 4956 1176 4964 1184
rect 5036 1156 5044 1164
rect 5036 1096 5044 1104
rect 4908 1076 4916 1084
rect 4940 1076 4948 1084
rect 5004 1076 5012 1084
rect 4860 1016 4868 1024
rect 4956 996 4964 1004
rect 4796 916 4804 924
rect 4908 916 4916 924
rect 4924 916 4932 924
rect 4972 976 4980 984
rect 5100 1316 5108 1324
rect 5100 1216 5108 1224
rect 5100 1116 5108 1124
rect 5084 1076 5092 1084
rect 5116 1076 5124 1084
rect 5148 1096 5156 1104
rect 5068 1056 5076 1064
rect 5084 1016 5092 1024
rect 5068 976 5076 984
rect 4988 916 4996 924
rect 4780 836 4788 844
rect 4716 736 4724 744
rect 4700 716 4708 724
rect 4844 716 4852 724
rect 4748 696 4756 704
rect 4796 696 4804 704
rect 4668 656 4676 664
rect 4732 616 4740 624
rect 4828 676 4836 684
rect 4924 796 4932 804
rect 4892 736 4900 744
rect 4924 696 4932 704
rect 4892 676 4900 684
rect 4844 616 4852 624
rect 4796 596 4804 604
rect 4716 556 4724 564
rect 4764 556 4772 564
rect 4796 556 4804 564
rect 4492 516 4500 524
rect 4428 496 4436 504
rect 4444 496 4452 504
rect 4476 496 4484 504
rect 4444 476 4452 484
rect 4428 336 4436 344
rect 4444 296 4452 304
rect 4460 276 4468 284
rect 4652 516 4660 524
rect 4732 516 4740 524
rect 4636 476 4644 484
rect 4556 436 4564 444
rect 4574 406 4582 414
rect 4588 406 4596 414
rect 4602 406 4610 414
rect 4652 296 4660 304
rect 4700 276 4708 284
rect 4476 196 4484 204
rect 4460 136 4468 144
rect 4572 256 4580 264
rect 4524 236 4532 244
rect 4636 216 4644 224
rect 4524 136 4532 144
rect 4556 136 4564 144
rect 4652 196 4660 204
rect 4668 136 4676 144
rect 4748 496 4756 504
rect 4748 436 4756 444
rect 4764 316 4772 324
rect 4844 316 4852 324
rect 4940 536 4948 544
rect 5036 936 5044 944
rect 5004 816 5012 824
rect 4988 756 4996 764
rect 5068 776 5076 784
rect 5052 716 5060 724
rect 5100 956 5108 964
rect 5148 1036 5156 1044
rect 5116 936 5124 944
rect 5228 1236 5236 1244
rect 5228 1136 5236 1144
rect 5212 1116 5220 1124
rect 5180 1096 5188 1104
rect 5212 1056 5220 1064
rect 5212 1016 5220 1024
rect 5180 916 5188 924
rect 5132 876 5140 884
rect 5116 796 5124 804
rect 5020 696 5028 704
rect 5052 696 5060 704
rect 5084 696 5092 704
rect 5004 676 5012 684
rect 5036 676 5044 684
rect 5084 676 5092 684
rect 4972 516 4980 524
rect 5052 516 5060 524
rect 5020 396 5028 404
rect 5148 756 5156 764
rect 5132 656 5140 664
rect 5132 636 5140 644
rect 5164 576 5172 584
rect 5164 536 5172 544
rect 5116 496 5124 504
rect 5084 396 5092 404
rect 5084 336 5092 344
rect 4812 296 4820 304
rect 4892 296 4900 304
rect 4924 296 4932 304
rect 4972 296 4980 304
rect 5132 296 5140 304
rect 4780 256 4788 264
rect 4828 256 4836 264
rect 4892 236 4900 244
rect 4780 136 4788 144
rect 4844 136 4852 144
rect 4892 136 4900 144
rect 4748 116 4756 124
rect 4812 116 4820 124
rect 4492 96 4500 104
rect 4524 96 4532 104
rect 4796 96 4804 104
rect 5020 276 5028 284
rect 5100 256 5108 264
rect 4940 136 4948 144
rect 5164 336 5172 344
rect 5196 896 5204 904
rect 5372 1436 5380 1444
rect 5356 1416 5364 1424
rect 5516 1736 5524 1744
rect 5452 1696 5460 1704
rect 5452 1556 5460 1564
rect 5452 1476 5460 1484
rect 5516 1596 5524 1604
rect 5500 1496 5508 1504
rect 5484 1376 5492 1384
rect 5452 1356 5460 1364
rect 5548 1776 5556 1784
rect 5756 1876 5764 1884
rect 5788 1856 5796 1864
rect 5724 1816 5732 1824
rect 5676 1756 5684 1764
rect 5580 1716 5588 1724
rect 5660 1716 5668 1724
rect 5564 1696 5572 1704
rect 5628 1696 5636 1704
rect 5644 1696 5652 1704
rect 5596 1676 5604 1684
rect 5628 1676 5636 1684
rect 5676 1676 5684 1684
rect 5628 1476 5636 1484
rect 5692 1476 5700 1484
rect 5596 1396 5604 1404
rect 5692 1436 5700 1444
rect 5564 1356 5572 1364
rect 5580 1356 5588 1364
rect 5628 1356 5636 1364
rect 5388 1336 5396 1344
rect 5436 1336 5444 1344
rect 5404 1316 5412 1324
rect 5516 1316 5524 1324
rect 5292 1296 5300 1304
rect 5644 1316 5652 1324
rect 5676 1316 5684 1324
rect 5532 1296 5540 1304
rect 5564 1296 5572 1304
rect 5612 1296 5620 1304
rect 5676 1296 5684 1304
rect 5468 1276 5476 1284
rect 5340 1136 5348 1144
rect 5500 1136 5508 1144
rect 5308 1116 5316 1124
rect 5372 1116 5380 1124
rect 5708 1296 5716 1304
rect 5692 1236 5700 1244
rect 5676 1156 5684 1164
rect 5692 1116 5700 1124
rect 5260 1096 5268 1104
rect 5292 1096 5300 1104
rect 5484 1096 5492 1104
rect 5644 1096 5652 1104
rect 5708 1096 5716 1104
rect 5356 1076 5364 1084
rect 5388 1076 5396 1084
rect 5244 956 5252 964
rect 5276 956 5284 964
rect 5340 956 5348 964
rect 5372 956 5380 964
rect 5228 916 5236 924
rect 5244 876 5252 884
rect 5228 816 5236 824
rect 5260 716 5268 724
rect 5196 316 5204 324
rect 5244 496 5252 504
rect 5532 1056 5540 1064
rect 5628 1076 5636 1084
rect 5564 1016 5572 1024
rect 5420 996 5428 1004
rect 5660 1036 5668 1044
rect 5484 976 5492 984
rect 5628 976 5636 984
rect 5692 976 5700 984
rect 5404 936 5412 944
rect 5324 916 5332 924
rect 5340 896 5348 904
rect 5452 896 5460 904
rect 5436 756 5444 764
rect 5468 756 5476 764
rect 5356 736 5364 744
rect 5436 736 5444 744
rect 5356 696 5364 704
rect 5404 676 5412 684
rect 5436 676 5444 684
rect 5308 616 5316 624
rect 5276 596 5284 604
rect 5276 556 5284 564
rect 5308 536 5316 544
rect 5324 536 5332 544
rect 5292 516 5300 524
rect 5260 436 5268 444
rect 5244 396 5252 404
rect 5212 296 5220 304
rect 5228 276 5236 284
rect 5420 596 5428 604
rect 5388 576 5396 584
rect 5356 556 5364 564
rect 5340 476 5348 484
rect 5372 476 5380 484
rect 5356 456 5364 464
rect 5452 656 5460 664
rect 5436 556 5444 564
rect 5404 496 5412 504
rect 5404 476 5412 484
rect 5388 376 5396 384
rect 5356 356 5364 364
rect 5324 316 5332 324
rect 5260 276 5268 284
rect 5244 256 5252 264
rect 5212 236 5220 244
rect 5212 136 5220 144
rect 5308 136 5316 144
rect 4892 96 4900 104
rect 5180 116 5188 124
rect 5228 116 5236 124
rect 5292 116 5300 124
rect 5436 336 5444 344
rect 5612 956 5620 964
rect 5644 936 5652 944
rect 5788 1796 5796 1804
rect 5820 1796 5828 1804
rect 5948 1936 5956 1944
rect 5948 1896 5950 1904
rect 5950 1896 5956 1904
rect 5916 1756 5924 1764
rect 5740 1716 5748 1724
rect 5852 1736 5860 1744
rect 5820 1596 5828 1604
rect 5852 1596 5860 1604
rect 5756 1556 5764 1564
rect 5884 1476 5892 1484
rect 5788 1416 5796 1424
rect 5852 1416 5860 1424
rect 5868 1416 5876 1424
rect 5916 1416 5924 1424
rect 5852 1376 5860 1384
rect 5836 1316 5844 1324
rect 5852 1316 5860 1324
rect 5852 1176 5860 1184
rect 5724 1036 5732 1044
rect 5884 1336 5892 1344
rect 5948 1318 5956 1324
rect 5948 1316 5956 1318
rect 6044 2336 6052 2344
rect 6044 2316 6052 2324
rect 6044 2296 6052 2304
rect 6028 2276 6036 2284
rect 6044 2256 6052 2264
rect 5980 1916 5988 1924
rect 6028 1896 6036 1904
rect 6028 1876 6036 1884
rect 6012 1836 6020 1844
rect 5996 1736 6004 1744
rect 5996 1696 6004 1704
rect 5996 1676 6004 1684
rect 5980 1596 5988 1604
rect 5964 1196 5972 1204
rect 5996 1096 6004 1104
rect 5900 1076 5908 1084
rect 6028 1676 6036 1684
rect 6124 3096 6132 3104
rect 6092 2816 6100 2824
rect 6124 1896 6132 1904
rect 6076 1836 6084 1844
rect 6124 1696 6132 1704
rect 6124 1516 6132 1524
rect 6044 1476 6052 1484
rect 6028 1396 6036 1404
rect 6092 1396 6100 1404
rect 6076 1296 6084 1304
rect 6044 1116 6052 1124
rect 6060 1096 6068 1104
rect 6076 1096 6084 1104
rect 5868 1056 5876 1064
rect 5884 976 5892 984
rect 5916 956 5924 964
rect 5564 916 5572 924
rect 5708 916 5716 924
rect 5676 896 5684 904
rect 5740 896 5748 904
rect 5612 856 5620 864
rect 5580 736 5588 744
rect 5628 816 5636 824
rect 5612 716 5620 724
rect 5612 696 5620 704
rect 5484 676 5492 684
rect 5516 476 5524 484
rect 5500 436 5508 444
rect 5596 636 5604 644
rect 5564 616 5572 624
rect 5548 536 5556 544
rect 5532 396 5540 404
rect 5516 356 5524 364
rect 5532 336 5540 344
rect 5644 716 5652 724
rect 5692 876 5700 884
rect 5708 756 5716 764
rect 5724 736 5732 744
rect 5756 736 5764 744
rect 5836 736 5844 744
rect 5708 696 5716 704
rect 5756 696 5764 704
rect 5804 636 5812 644
rect 5772 596 5780 604
rect 6044 1076 6052 1084
rect 6012 916 6020 924
rect 5916 776 5924 784
rect 5948 776 5956 784
rect 5676 576 5684 584
rect 5788 576 5796 584
rect 6076 976 6084 984
rect 6060 816 6068 824
rect 6028 756 6036 764
rect 5964 716 5972 724
rect 5980 676 5988 684
rect 6012 676 6020 684
rect 6060 676 6068 684
rect 5980 596 5988 604
rect 6028 596 6036 604
rect 5868 496 5876 504
rect 5948 496 5956 504
rect 5756 456 5764 464
rect 5468 316 5476 324
rect 5516 316 5524 324
rect 5564 316 5572 324
rect 5628 316 5636 324
rect 5420 296 5428 304
rect 5484 296 5492 304
rect 5388 276 5396 284
rect 5388 236 5396 244
rect 5436 276 5444 284
rect 5516 276 5524 284
rect 5596 276 5604 284
rect 5612 276 5620 284
rect 5580 256 5588 264
rect 5628 256 5636 264
rect 5452 236 5460 244
rect 5740 376 5748 384
rect 5708 356 5716 364
rect 5708 336 5716 344
rect 5596 176 5604 184
rect 5644 176 5652 184
rect 5532 156 5540 164
rect 5436 136 5444 144
rect 5548 116 5556 124
rect 5132 96 5140 104
rect 5180 96 5188 104
rect 5260 96 5268 104
rect 4220 76 4228 84
rect 4252 76 4260 84
rect 4348 76 4356 84
rect 4876 76 4884 84
rect 5004 76 5012 84
rect 1502 6 1510 14
rect 1516 6 1524 14
rect 1530 6 1538 14
rect 4574 6 4582 14
rect 4588 6 4596 14
rect 4602 6 4610 14
rect 6044 416 6052 424
rect 6060 296 6068 304
rect 5900 276 5908 284
rect 5868 256 5876 264
rect 5900 256 5908 264
rect 5900 176 5908 184
rect 5932 156 5940 164
rect 5660 136 5668 144
rect 5676 136 5684 144
rect 6060 276 6068 284
rect 6124 316 6132 324
rect 5676 116 5684 124
rect 5708 96 5716 104
rect 6108 96 6116 104
rect 5660 16 5668 24
<< metal3 >>
rect 1496 5614 1544 5616
rect 1496 5606 1500 5614
rect 1510 5606 1516 5614
rect 1524 5606 1530 5614
rect 1540 5606 1544 5614
rect 1496 5604 1544 5606
rect 4568 5614 4616 5616
rect 4568 5606 4572 5614
rect 4582 5606 4588 5614
rect 4596 5606 4602 5614
rect 4612 5606 4616 5614
rect 4568 5604 4616 5606
rect 5924 5557 6076 5563
rect 484 5537 636 5543
rect 1572 5537 1900 5543
rect 4068 5537 4252 5543
rect 580 5517 604 5523
rect 1876 5517 1932 5523
rect 3620 5517 3644 5523
rect 4212 5517 4444 5523
rect 4644 5517 4876 5523
rect 4884 5517 4940 5523
rect 5188 5517 5212 5523
rect 5332 5517 5500 5523
rect 340 5497 444 5503
rect 452 5497 604 5503
rect 1236 5497 1244 5503
rect 1684 5497 1772 5503
rect 1876 5497 1900 5503
rect 2164 5497 2444 5503
rect 3332 5497 3452 5503
rect 3636 5497 3900 5503
rect 4004 5497 4124 5503
rect 4324 5497 4412 5503
rect 4756 5497 4780 5503
rect 4868 5497 5052 5503
rect 5284 5497 5324 5503
rect 36 5477 172 5483
rect 580 5477 860 5483
rect 1124 5477 1212 5483
rect 1764 5477 1836 5483
rect 2276 5477 2620 5483
rect 3236 5477 3436 5483
rect 3508 5477 3644 5483
rect 3652 5477 4572 5483
rect 5188 5477 5292 5483
rect 5796 5477 5932 5483
rect 180 5457 204 5463
rect 292 5457 332 5463
rect 340 5457 748 5463
rect 964 5457 1452 5463
rect 2388 5457 2556 5463
rect 3524 5457 3628 5463
rect 3636 5457 3660 5463
rect 4180 5457 4300 5463
rect 4500 5457 4556 5463
rect 5236 5457 5388 5463
rect 5556 5457 5612 5463
rect 5620 5457 5756 5463
rect 5764 5457 5868 5463
rect 1108 5437 1180 5443
rect 4356 5437 4684 5443
rect 4868 5437 4924 5443
rect 4932 5437 5132 5443
rect 5140 5437 5276 5443
rect 5588 5437 5596 5443
rect 1188 5417 1228 5423
rect 1940 5417 2204 5423
rect 2212 5417 2412 5423
rect 2420 5417 2476 5423
rect 2484 5417 2924 5423
rect 2932 5417 2988 5423
rect 4685 5423 4691 5436
rect 4685 5417 5020 5423
rect 5108 5417 5324 5423
rect 5332 5417 5452 5423
rect 3032 5414 3080 5416
rect 3032 5406 3036 5414
rect 3046 5406 3052 5414
rect 3060 5406 3066 5414
rect 3076 5406 3080 5414
rect 3032 5404 3080 5406
rect 1172 5397 1372 5403
rect 1972 5397 2268 5403
rect 3428 5397 3532 5403
rect 3540 5397 3580 5403
rect 3588 5397 3772 5403
rect 3780 5397 4508 5403
rect 4516 5397 5388 5403
rect 5396 5397 5948 5403
rect 5956 5397 6028 5403
rect 2020 5377 2076 5383
rect 2701 5383 2707 5396
rect 2701 5377 3020 5383
rect 3716 5377 3724 5383
rect 4388 5377 4508 5383
rect 4516 5377 4748 5383
rect 4756 5377 4812 5383
rect 4820 5377 4876 5383
rect 4884 5377 5340 5383
rect 356 5357 428 5363
rect 1044 5357 1084 5363
rect 1892 5357 2172 5363
rect 2196 5357 2428 5363
rect 2436 5357 2444 5363
rect 2660 5357 2732 5363
rect 2740 5357 2764 5363
rect 2900 5357 2956 5363
rect 2996 5357 3100 5363
rect 3204 5357 3324 5363
rect 3364 5357 3500 5363
rect 3684 5357 3868 5363
rect 3876 5357 3996 5363
rect 4004 5357 4172 5363
rect 4564 5357 4668 5363
rect 4676 5357 4924 5363
rect 4932 5357 4988 5363
rect 5444 5357 5644 5363
rect 148 5337 364 5343
rect 420 5337 460 5343
rect 564 5337 844 5343
rect 980 5337 1052 5343
rect 1060 5337 1116 5343
rect 1476 5337 1580 5343
rect 1588 5337 1916 5343
rect 2148 5337 2204 5343
rect 2436 5337 2460 5343
rect 3508 5337 3580 5343
rect 3828 5337 4028 5343
rect 4196 5337 4348 5343
rect 4356 5337 4380 5343
rect 4484 5337 4652 5343
rect 4660 5337 4716 5343
rect 4724 5337 4844 5343
rect 4852 5337 4908 5343
rect 4916 5337 4972 5343
rect 4980 5337 5148 5343
rect 5620 5337 5788 5343
rect 5988 5337 6124 5343
rect 404 5317 444 5323
rect 452 5317 524 5323
rect 1060 5317 1132 5323
rect 1412 5317 1612 5323
rect 2004 5317 2044 5323
rect 3460 5317 3916 5323
rect 4340 5317 4524 5323
rect 4548 5317 4588 5323
rect 4596 5317 4739 5323
rect 340 5297 364 5303
rect 372 5297 428 5303
rect 564 5297 588 5303
rect 996 5297 1244 5303
rect 1252 5297 1724 5303
rect 3188 5297 3596 5303
rect 3732 5297 3804 5303
rect 4388 5297 4620 5303
rect 4733 5303 4739 5317
rect 4756 5317 4828 5323
rect 4932 5317 5052 5323
rect 4733 5297 4812 5303
rect 4996 5297 5308 5303
rect 5908 5297 5996 5303
rect 36 5277 524 5283
rect 1012 5277 1324 5283
rect 3572 5277 3708 5283
rect 3716 5277 3836 5283
rect 4180 5277 4396 5283
rect 4452 5277 4524 5283
rect 4580 5277 4876 5283
rect 4916 5277 4940 5283
rect 4948 5277 5180 5283
rect 4532 5257 4732 5263
rect 5844 5257 5996 5263
rect 1604 5237 1676 5243
rect 2276 5237 2332 5243
rect 4132 5237 5724 5243
rect 5732 5237 5836 5243
rect 5844 5237 5884 5243
rect 324 5217 412 5223
rect 420 5217 572 5223
rect 900 5217 1052 5223
rect 2740 5217 2812 5223
rect 3012 5217 3292 5223
rect 3300 5217 3468 5223
rect 3668 5217 3692 5223
rect 3700 5217 4060 5223
rect 4308 5217 4428 5223
rect 4660 5217 5196 5223
rect 1496 5214 1544 5216
rect 1496 5206 1500 5214
rect 1510 5206 1516 5214
rect 1524 5206 1530 5214
rect 1540 5206 1544 5214
rect 1496 5204 1544 5206
rect 4568 5214 4616 5216
rect 4568 5206 4572 5214
rect 4582 5206 4588 5214
rect 4596 5206 4602 5214
rect 4612 5206 4616 5214
rect 4568 5204 4616 5206
rect 4324 5197 4380 5203
rect 5172 5197 5212 5203
rect 5956 5197 5980 5203
rect 4116 5177 4988 5183
rect 5044 5177 5420 5183
rect 5428 5177 5756 5183
rect 4836 5157 5420 5163
rect 5428 5157 5452 5163
rect 445 5137 460 5143
rect 276 5097 428 5103
rect 445 5103 451 5137
rect 820 5137 860 5143
rect 868 5137 1020 5143
rect 1028 5137 1052 5143
rect 1060 5137 1532 5143
rect 3732 5137 3932 5143
rect 3988 5137 4092 5143
rect 4100 5137 4844 5143
rect 4852 5137 5052 5143
rect 5060 5137 5228 5143
rect 5364 5137 5452 5143
rect 468 5117 540 5123
rect 724 5117 796 5123
rect 1108 5117 1148 5123
rect 1156 5117 1308 5123
rect 3204 5117 3356 5123
rect 3764 5117 3788 5123
rect 3796 5117 3980 5123
rect 3988 5117 4108 5123
rect 4372 5117 4396 5123
rect 4404 5117 4652 5123
rect 4692 5117 4908 5123
rect 5124 5117 5180 5123
rect 5236 5117 5484 5123
rect 5700 5117 5788 5123
rect 445 5097 460 5103
rect 532 5097 1212 5103
rect 1716 5097 1836 5103
rect 2372 5097 2412 5103
rect 2804 5097 3132 5103
rect 3140 5097 3164 5103
rect 3300 5097 3388 5103
rect 3652 5097 3900 5103
rect 3924 5097 3964 5103
rect 4148 5097 4156 5103
rect 4356 5097 4412 5103
rect 4420 5097 4668 5103
rect 4772 5097 4860 5103
rect 4884 5097 5388 5103
rect 5693 5103 5699 5116
rect 5396 5097 5699 5103
rect 132 5077 172 5083
rect 180 5077 220 5083
rect 388 5077 476 5083
rect 484 5077 556 5083
rect 564 5077 796 5083
rect 1172 5077 1260 5083
rect 1652 5077 1852 5083
rect 1860 5077 1900 5083
rect 2404 5077 2460 5083
rect 2484 5077 2620 5083
rect 2900 5077 2972 5083
rect 3284 5077 3324 5083
rect 3332 5077 3532 5083
rect 3540 5077 3964 5083
rect 4148 5077 4236 5083
rect 4292 5077 4364 5083
rect 4404 5077 4540 5083
rect 4884 5077 5212 5083
rect 5268 5077 5276 5083
rect 5444 5077 5724 5083
rect 5732 5077 5756 5083
rect 420 5057 492 5063
rect 1204 5057 1308 5063
rect 1316 5057 1388 5063
rect 1396 5057 1660 5063
rect 1684 5057 1740 5063
rect 2388 5057 2412 5063
rect 2484 5057 2524 5063
rect 2660 5057 3004 5063
rect 3012 5057 3196 5063
rect 3364 5057 4348 5063
rect 4644 5057 4716 5063
rect 4804 5057 5004 5063
rect 5204 5057 5228 5063
rect 5364 5057 5612 5063
rect 20 5037 60 5043
rect 740 5037 908 5043
rect 948 5037 1004 5043
rect 1252 5037 1500 5043
rect 1508 5037 1692 5043
rect 2260 5037 2316 5043
rect 2324 5037 2364 5043
rect 2964 5037 3548 5043
rect 3796 5037 4220 5043
rect 4500 5037 4700 5043
rect 4708 5037 4876 5043
rect 5076 5037 5292 5043
rect 5300 5037 5388 5043
rect 196 5017 748 5023
rect 1716 5017 1724 5023
rect 2244 5017 2476 5023
rect 3156 5017 3836 5023
rect 3924 5017 4044 5023
rect 4228 5017 4556 5023
rect 4916 5017 5324 5023
rect 3032 5014 3080 5016
rect 3032 5006 3036 5014
rect 3046 5006 3052 5014
rect 3060 5006 3066 5014
rect 3076 5006 3080 5014
rect 3032 5004 3080 5006
rect 164 4997 460 5003
rect 676 4997 844 5003
rect 852 4997 924 5003
rect 1060 4997 1132 5003
rect 1300 4997 1404 5003
rect 1924 4997 1964 5003
rect 1972 4997 2156 5003
rect 3428 4997 3516 5003
rect 3924 4997 3932 5003
rect 5092 4997 5180 5003
rect 5188 4997 5372 5003
rect 5380 4997 5436 5003
rect 5684 4997 5916 5003
rect 5924 4997 5948 5003
rect 564 4977 1068 4983
rect 1828 4977 2252 4983
rect 2260 4977 2444 4983
rect 2820 4977 2940 4983
rect 3028 4977 3196 4983
rect 3844 4977 4332 4983
rect 4340 4977 4476 4983
rect 4532 4977 4764 4983
rect 4772 4977 4956 4983
rect 4964 4977 5068 4983
rect 5172 4977 5276 4983
rect 356 4957 652 4963
rect 660 4957 908 4963
rect 916 4957 1276 4963
rect 2020 4957 2268 4963
rect 2276 4957 2444 4963
rect 2452 4957 2508 4963
rect 2964 4957 3148 4963
rect 3204 4957 3244 4963
rect 3252 4957 3580 4963
rect 3588 4957 3868 4963
rect 3940 4957 4188 4963
rect 4212 4957 4476 4963
rect 4548 4957 4572 4963
rect 4724 4957 4892 4963
rect 5124 4957 5292 4963
rect 5444 4957 5628 4963
rect 452 4937 492 4943
rect 644 4937 876 4943
rect 884 4937 972 4943
rect 1028 4937 1116 4943
rect 1508 4937 1772 4943
rect 1956 4937 2140 4943
rect 2644 4937 2764 4943
rect 2772 4937 2780 4943
rect 2820 4937 2860 4943
rect 2916 4937 2972 4943
rect 2980 4937 3340 4943
rect 3476 4937 3692 4943
rect 3972 4937 4732 4943
rect 4740 4937 4796 4943
rect 5012 4937 5580 4943
rect 5588 4937 5740 4943
rect 20 4917 172 4923
rect 308 4917 460 4923
rect 484 4917 588 4923
rect 628 4917 876 4923
rect 884 4917 892 4923
rect 1044 4917 1164 4923
rect 1172 4917 1468 4923
rect 1604 4917 1836 4923
rect 2836 4917 2988 4923
rect 3124 4917 3260 4923
rect 3332 4917 3356 4923
rect 3412 4917 3452 4923
rect 3524 4917 3596 4923
rect 3748 4917 4012 4923
rect 4100 4917 4444 4923
rect 4452 4917 4668 4923
rect 4676 4917 5164 4923
rect 5172 4917 5468 4923
rect 5732 4917 5980 4923
rect 1037 4904 1043 4916
rect 148 4897 172 4903
rect 212 4897 300 4903
rect 420 4897 556 4903
rect 564 4897 588 4903
rect 660 4897 748 4903
rect 788 4897 828 4903
rect 852 4897 1004 4903
rect 3108 4897 3420 4903
rect 3572 4897 3788 4903
rect 3876 4897 3996 4903
rect 4004 4897 4268 4903
rect 4564 4897 4668 4903
rect 4756 4897 4892 4903
rect 4980 4897 5068 4903
rect 5124 4897 5212 4903
rect 5444 4897 5468 4903
rect 532 4877 652 4883
rect 820 4877 1132 4883
rect 2468 4877 2844 4883
rect 2852 4877 3004 4883
rect 3300 4877 3452 4883
rect 3556 4877 3644 4883
rect 3780 4877 3804 4883
rect 3812 4877 4060 4883
rect 4308 4877 4460 4883
rect 4708 4877 4780 4883
rect 4996 4877 5020 4883
rect 5044 4877 5132 4883
rect 5140 4877 5196 4883
rect 68 4857 204 4863
rect 212 4857 396 4863
rect 404 4857 428 4863
rect 436 4857 732 4863
rect 1044 4857 1964 4863
rect 2852 4857 2924 4863
rect 3236 4857 3372 4863
rect 3380 4857 4108 4863
rect 4308 4857 4396 4863
rect 164 4837 172 4843
rect 484 4837 716 4843
rect 884 4837 1212 4843
rect 2132 4837 2252 4843
rect 3316 4837 3356 4843
rect 3444 4837 3724 4843
rect 4068 4837 4252 4843
rect 4276 4837 4540 4843
rect 4564 4837 4924 4843
rect 4948 4837 5164 4843
rect 5172 4837 5196 4843
rect 5252 4837 5404 4843
rect 5796 4837 6028 4843
rect 580 4817 732 4823
rect 868 4817 915 4823
rect 228 4797 316 4803
rect 724 4797 860 4803
rect 909 4803 915 4817
rect 932 4817 1020 4823
rect 2996 4817 4492 4823
rect 4660 4817 4716 4823
rect 4788 4817 4956 4823
rect 1496 4814 1544 4816
rect 1496 4806 1500 4814
rect 1510 4806 1516 4814
rect 1524 4806 1530 4814
rect 1540 4806 1544 4814
rect 1496 4804 1544 4806
rect 4568 4814 4616 4816
rect 4568 4806 4572 4814
rect 4582 4806 4588 4814
rect 4596 4806 4602 4814
rect 4612 4806 4616 4814
rect 4568 4804 4616 4806
rect 909 4797 1155 4803
rect 836 4777 972 4783
rect 1149 4783 1155 4797
rect 1172 4797 1356 4803
rect 3572 4797 3708 4803
rect 3924 4797 3980 4803
rect 4276 4797 4300 4803
rect 4340 4797 4476 4803
rect 1149 4777 1452 4783
rect 3668 4777 3756 4783
rect 3764 4777 4076 4783
rect 4084 4777 4492 4783
rect 4676 4777 4940 4783
rect 516 4757 572 4763
rect 1124 4757 1212 4763
rect 1252 4757 1788 4763
rect 3172 4757 3548 4763
rect 3652 4757 3820 4763
rect 3828 4757 3852 4763
rect 3924 4757 3932 4763
rect 4100 4757 4348 4763
rect 4388 4757 4476 4763
rect 4500 4757 4860 4763
rect 4868 4757 4876 4763
rect 196 4737 268 4743
rect 276 4737 716 4743
rect 724 4737 1148 4743
rect 1204 4737 1276 4743
rect 1364 4737 2892 4743
rect 2900 4737 2924 4743
rect 3284 4737 3507 4743
rect 3501 4724 3507 4737
rect 3556 4737 3612 4743
rect 3684 4737 4028 4743
rect 4036 4737 4140 4743
rect 4148 4737 4316 4743
rect 4324 4737 4412 4743
rect 4468 4737 4684 4743
rect 4788 4737 4812 4743
rect 5188 4737 5548 4743
rect 404 4717 588 4723
rect 948 4717 1116 4723
rect 1124 4717 1548 4723
rect 1700 4717 1852 4723
rect 2116 4717 2236 4723
rect 2388 4717 2508 4723
rect 2516 4717 2572 4723
rect 2580 4717 2876 4723
rect 3300 4717 3308 4723
rect 3508 4717 3644 4723
rect 3732 4717 4044 4723
rect 4116 4717 4428 4723
rect 4436 4717 4652 4723
rect 4660 4717 4684 4723
rect 4692 4717 4812 4723
rect 4868 4717 4972 4723
rect 5092 4717 5292 4723
rect 5300 4717 5532 4723
rect 84 4697 236 4703
rect 308 4697 540 4703
rect 740 4697 1036 4703
rect 1140 4697 1260 4703
rect 1284 4697 1308 4703
rect 1668 4697 1724 4703
rect 1748 4697 1772 4703
rect 2052 4697 2188 4703
rect 2420 4697 2540 4703
rect 3316 4697 3564 4703
rect 3604 4697 3740 4703
rect 3796 4697 4396 4703
rect 4404 4697 4444 4703
rect 4452 4697 4828 4703
rect 4836 4697 5196 4703
rect 5204 4697 5308 4703
rect 5556 4697 5772 4703
rect 324 4677 412 4683
rect 420 4677 524 4683
rect 580 4677 812 4683
rect 1044 4677 1484 4683
rect 1636 4677 1708 4683
rect 1716 4677 1724 4683
rect 1780 4677 1964 4683
rect 2132 4677 2220 4683
rect 2356 4677 2428 4683
rect 3284 4677 3324 4683
rect 3460 4677 3884 4683
rect 3965 4677 3996 4683
rect 628 4657 796 4663
rect 813 4663 819 4676
rect 813 4657 1116 4663
rect 1284 4657 1340 4663
rect 1540 4657 1804 4663
rect 1844 4657 2284 4663
rect 2420 4657 2460 4663
rect 2532 4657 2700 4663
rect 3965 4663 3971 4677
rect 4276 4677 4316 4683
rect 4388 4677 4460 4683
rect 4660 4677 4684 4683
rect 4948 4677 5004 4683
rect 5028 4677 5260 4683
rect 5492 4677 5676 4683
rect 5796 4677 5996 4683
rect 3652 4657 3971 4663
rect 3988 4657 4044 4663
rect 4381 4663 4387 4676
rect 4212 4657 4387 4663
rect 4724 4657 5068 4663
rect 5204 4657 5564 4663
rect 5844 4657 5884 4663
rect 228 4637 684 4643
rect 1188 4637 1436 4643
rect 1444 4637 1660 4643
rect 2084 4637 2140 4643
rect 2308 4637 2444 4643
rect 2452 4637 2476 4643
rect 2788 4637 2860 4643
rect 2868 4637 3036 4643
rect 3364 4637 3404 4643
rect 3492 4637 3932 4643
rect 3940 4637 4140 4643
rect 4612 4637 4780 4643
rect 644 4617 812 4623
rect 820 4617 1068 4623
rect 1172 4617 1404 4623
rect 1412 4617 1676 4623
rect 3412 4617 3532 4623
rect 3972 4617 3980 4623
rect 4116 4617 4156 4623
rect 4308 4617 4348 4623
rect 4420 4617 4716 4623
rect 3032 4614 3080 4616
rect 3032 4606 3036 4614
rect 3046 4606 3052 4614
rect 3060 4606 3066 4614
rect 3076 4606 3080 4614
rect 3032 4604 3080 4606
rect 388 4597 1004 4603
rect 1364 4597 1388 4603
rect 1396 4597 1436 4603
rect 1444 4597 1772 4603
rect 1780 4597 1836 4603
rect 1860 4597 1964 4603
rect 2468 4597 2508 4603
rect 3188 4597 3756 4603
rect 3764 4597 3964 4603
rect 3972 4597 4860 4603
rect 5172 4597 5212 4603
rect 5220 4597 5516 4603
rect 5636 4597 5836 4603
rect 5924 4597 5964 4603
rect 900 4577 956 4583
rect 1476 4577 1596 4583
rect 1604 4577 2076 4583
rect 3732 4577 3772 4583
rect 3780 4577 4604 4583
rect 5060 4577 5148 4583
rect 5156 4577 5356 4583
rect 5364 4577 5404 4583
rect 5444 4577 5596 4583
rect 180 4557 540 4563
rect 1060 4557 1404 4563
rect 1684 4557 1756 4563
rect 1764 4557 1980 4563
rect 2756 4557 2812 4563
rect 2868 4557 2956 4563
rect 3428 4557 3500 4563
rect 3652 4557 4108 4563
rect 4132 4557 4556 4563
rect 4772 4557 4812 4563
rect 4852 4557 5068 4563
rect 5572 4557 5916 4563
rect 228 4537 268 4543
rect 340 4537 364 4543
rect 436 4537 508 4543
rect 516 4537 524 4543
rect 532 4537 780 4543
rect 804 4537 828 4543
rect 868 4537 1212 4543
rect 1268 4537 1452 4543
rect 1460 4537 1772 4543
rect 1789 4537 1852 4543
rect 148 4517 236 4523
rect 292 4517 796 4523
rect 1012 4517 1036 4523
rect 1092 4517 1148 4523
rect 1492 4517 1628 4523
rect 1636 4517 1692 4523
rect 1789 4523 1795 4537
rect 1940 4537 2220 4543
rect 2292 4537 2364 4543
rect 2404 4537 2764 4543
rect 2772 4537 2828 4543
rect 2836 4537 2860 4543
rect 2932 4537 3164 4543
rect 3620 4537 3692 4543
rect 3828 4537 3868 4543
rect 3908 4537 3996 4543
rect 4164 4537 4220 4543
rect 4292 4537 4396 4543
rect 4692 4537 4700 4543
rect 4804 4537 4860 4543
rect 4948 4537 4988 4543
rect 5060 4537 5724 4543
rect 1764 4517 1795 4523
rect 1812 4517 1884 4523
rect 1988 4517 2028 4523
rect 2580 4517 2732 4523
rect 3444 4517 3628 4523
rect 3684 4517 4108 4523
rect 4148 4517 4204 4523
rect 4452 4517 4508 4523
rect 4756 4517 4844 4523
rect 4932 4517 5004 4523
rect 5092 4517 5132 4523
rect 5156 4517 5164 4523
rect 5188 4517 5308 4523
rect 5428 4517 5596 4523
rect 5908 4517 5932 4523
rect 260 4497 284 4503
rect 596 4497 828 4503
rect 1028 4497 1132 4503
rect 1156 4497 1388 4503
rect 1428 4497 1484 4503
rect 1620 4497 1628 4503
rect 1636 4497 1692 4503
rect 1700 4497 1836 4503
rect 1908 4497 2108 4503
rect 2116 4497 2764 4503
rect 3316 4497 3676 4503
rect 3828 4497 3900 4503
rect 4020 4497 4300 4503
rect 4724 4497 4924 4503
rect 5044 4497 5260 4503
rect 5604 4497 5948 4503
rect 100 4477 268 4483
rect 468 4477 492 4483
rect 708 4477 732 4483
rect 740 4477 876 4483
rect 884 4477 1068 4483
rect 1108 4477 1164 4483
rect 1668 4477 1996 4483
rect 2004 4477 2092 4483
rect 2468 4477 2652 4483
rect 3524 4477 4364 4483
rect 4468 4477 4524 4483
rect 5060 4477 5116 4483
rect 5140 4477 5164 4483
rect 788 4457 940 4463
rect 1332 4457 1372 4463
rect 1380 4457 1644 4463
rect 2980 4457 2988 4463
rect 4324 4457 4540 4463
rect 4548 4457 4636 4463
rect 4644 4457 5100 4463
rect 452 4437 988 4443
rect 1556 4437 1612 4443
rect 2340 4437 2956 4443
rect 2964 4437 3052 4443
rect 3492 4437 3756 4443
rect 3860 4437 4092 4443
rect 4100 4437 4348 4443
rect 4420 4437 4508 4443
rect 4964 4437 5196 4443
rect 884 4417 1164 4423
rect 1348 4417 1356 4423
rect 2500 4417 2508 4423
rect 5236 4417 5660 4423
rect 5748 4417 5804 4423
rect 6004 4417 6060 4423
rect 1496 4414 1544 4416
rect 1496 4406 1500 4414
rect 1510 4406 1516 4414
rect 1524 4406 1530 4414
rect 1540 4406 1544 4414
rect 1496 4404 1544 4406
rect 4568 4414 4616 4416
rect 4568 4406 4572 4414
rect 4582 4406 4588 4414
rect 4596 4406 4602 4414
rect 4612 4406 4616 4414
rect 4568 4404 4616 4406
rect 132 4397 220 4403
rect 1300 4397 1340 4403
rect 2964 4397 2972 4403
rect 5364 4397 5452 4403
rect 5460 4397 5484 4403
rect 5524 4397 5756 4403
rect 2148 4377 2428 4383
rect 2676 4377 2780 4383
rect 3508 4377 3564 4383
rect 3572 4377 3724 4383
rect 4148 4377 4204 4383
rect 4548 4377 4764 4383
rect 5076 4377 5116 4383
rect 5300 4377 5356 4383
rect 180 4357 492 4363
rect 500 4357 716 4363
rect 724 4357 1276 4363
rect 1284 4357 1372 4363
rect 1412 4357 2252 4363
rect 2260 4357 2780 4363
rect 3476 4357 3564 4363
rect 3572 4357 3676 4363
rect 3684 4357 3820 4363
rect 4532 4357 4700 4363
rect 4708 4357 5052 4363
rect 708 4337 732 4343
rect 820 4337 1084 4343
rect 1188 4337 1292 4343
rect 1684 4337 1948 4343
rect 2020 4337 2076 4343
rect 2132 4337 2204 4343
rect 2212 4337 2684 4343
rect 2692 4337 2716 4343
rect 4068 4337 4124 4343
rect 4132 4337 4156 4343
rect 4628 4337 4748 4343
rect 20 4317 252 4323
rect 260 4317 332 4323
rect 740 4317 876 4323
rect 884 4317 940 4323
rect 1140 4317 1452 4323
rect 1476 4317 1564 4323
rect 1588 4317 1676 4323
rect 2164 4317 2188 4323
rect 2228 4317 2300 4323
rect 2420 4317 2556 4323
rect 2564 4317 2764 4323
rect 2772 4317 2876 4323
rect 3476 4317 3548 4323
rect 3556 4317 3644 4323
rect 3988 4317 4940 4323
rect -19 4297 12 4303
rect 36 4297 60 4303
rect 68 4297 364 4303
rect 452 4297 588 4303
rect 612 4297 844 4303
rect 900 4297 988 4303
rect 1076 4297 1148 4303
rect 1156 4297 1340 4303
rect 1572 4297 1724 4303
rect 1972 4297 2108 4303
rect 2244 4297 2268 4303
rect 2285 4297 2428 4303
rect 116 4277 140 4283
rect 340 4277 364 4283
rect 372 4277 396 4283
rect 516 4277 540 4283
rect 644 4277 1004 4283
rect 1076 4277 1100 4283
rect 1252 4277 1564 4283
rect 1588 4277 1708 4283
rect 2285 4283 2291 4297
rect 2548 4297 2604 4303
rect 2660 4297 2748 4303
rect 2820 4297 2844 4303
rect 3364 4297 3612 4303
rect 3940 4297 4012 4303
rect 4036 4297 4108 4303
rect 4148 4297 4252 4303
rect 4404 4297 4508 4303
rect 4516 4297 4956 4303
rect 5060 4297 5196 4303
rect 5476 4297 5564 4303
rect 2196 4277 2291 4283
rect 2388 4277 2572 4283
rect 2580 4277 2668 4283
rect 2740 4277 3068 4283
rect 3556 4277 3692 4283
rect 3700 4277 3804 4283
rect 3812 4277 3884 4283
rect 4260 4277 4460 4283
rect 4820 4277 4956 4283
rect 5540 4277 5612 4283
rect 5716 4277 5820 4283
rect 141 4263 147 4276
rect 141 4257 380 4263
rect 1012 4257 1052 4263
rect 1236 4257 1683 4263
rect 100 4237 364 4243
rect 532 4237 636 4243
rect 932 4237 1196 4243
rect 1268 4237 1356 4243
rect 1677 4243 1683 4257
rect 1700 4257 1724 4263
rect 1732 4257 1820 4263
rect 1828 4257 2252 4263
rect 2260 4257 2316 4263
rect 2324 4257 2588 4263
rect 3044 4257 3132 4263
rect 3140 4257 3164 4263
rect 4932 4257 5276 4263
rect 5284 4257 5820 4263
rect 1364 4237 1651 4243
rect 1677 4237 1804 4243
rect 1645 4224 1651 4237
rect 2180 4237 2300 4243
rect 2308 4237 2332 4243
rect 2340 4237 2476 4243
rect 2484 4237 2524 4243
rect 2548 4237 2700 4243
rect 3892 4237 4083 4243
rect 4077 4224 4083 4237
rect 5540 4237 5612 4243
rect 5668 4237 5692 4243
rect 324 4217 428 4223
rect 916 4217 1180 4223
rect 1188 4217 1244 4223
rect 1300 4217 1308 4223
rect 1652 4217 2044 4223
rect 2324 4217 2828 4223
rect 3380 4217 3964 4223
rect 4084 4217 4380 4223
rect 5268 4217 5308 4223
rect 5668 4217 5852 4223
rect 3032 4214 3080 4216
rect 3032 4206 3036 4214
rect 3046 4206 3052 4214
rect 3060 4206 3066 4214
rect 3076 4206 3080 4214
rect 3032 4204 3080 4206
rect 964 4197 1068 4203
rect 1508 4197 1900 4203
rect 1908 4197 1932 4203
rect 1940 4197 1980 4203
rect 2148 4197 2940 4203
rect 3652 4197 3676 4203
rect 3780 4197 3996 4203
rect 4212 4197 4268 4203
rect 4996 4197 5452 4203
rect 5460 4197 5580 4203
rect 980 4177 1036 4183
rect 1044 4177 1420 4183
rect 1428 4177 1500 4183
rect 2804 4177 2828 4183
rect 3588 4177 3660 4183
rect 3668 4177 3820 4183
rect 3828 4177 4092 4183
rect 4116 4177 4284 4183
rect 4452 4177 4652 4183
rect 5428 4177 5468 4183
rect 292 4157 444 4163
rect 452 4157 716 4163
rect 932 4157 956 4163
rect 1172 4157 1212 4163
rect 1300 4157 1564 4163
rect 1620 4157 1740 4163
rect 2628 4157 2668 4163
rect 2788 4157 2844 4163
rect 2900 4157 2956 4163
rect 2964 4157 3036 4163
rect 3428 4157 3612 4163
rect 3652 4157 3740 4163
rect 3812 4157 3900 4163
rect 3924 4157 4156 4163
rect 4180 4157 4364 4163
rect 4420 4157 4492 4163
rect 4500 4157 4572 4163
rect 4580 4157 4716 4163
rect 4724 4157 4908 4163
rect 4916 4157 5084 4163
rect 5108 4157 5212 4163
rect 5220 4157 5500 4163
rect 5828 4157 5916 4163
rect 5924 4157 6012 4163
rect 84 4137 140 4143
rect 564 4137 620 4143
rect 644 4137 812 4143
rect 820 4137 844 4143
rect 1092 4137 1324 4143
rect 1396 4137 1452 4143
rect 1684 4137 1756 4143
rect 1956 4137 2156 4143
rect 2308 4137 2348 4143
rect 2388 4137 2476 4143
rect 2644 4137 2803 4143
rect 2797 4124 2803 4137
rect 2996 4137 3132 4143
rect 3556 4137 3708 4143
rect 3732 4137 4012 4143
rect 4036 4137 4348 4143
rect 4356 4137 4524 4143
rect 4612 4137 4668 4143
rect 4676 4137 4748 4143
rect 4964 4137 5052 4143
rect 5108 4137 5148 4143
rect 5156 4137 5356 4143
rect 5364 4137 5468 4143
rect 5476 4137 5516 4143
rect 5892 4137 5900 4143
rect 260 4117 332 4123
rect 484 4117 588 4123
rect 612 4117 700 4123
rect 724 4117 940 4123
rect 948 4117 1100 4123
rect 1140 4117 1196 4123
rect 1572 4117 1612 4123
rect 1620 4117 1692 4123
rect 1780 4117 1804 4123
rect 2356 4117 2396 4123
rect 2404 4117 2588 4123
rect 2660 4117 2780 4123
rect 2804 4117 2860 4123
rect 3012 4117 3164 4123
rect 3172 4117 3372 4123
rect 3572 4117 3724 4123
rect 3764 4117 3836 4123
rect 3972 4117 4028 4123
rect 4068 4117 4108 4123
rect 4164 4117 4220 4123
rect 4372 4117 4636 4123
rect 4644 4117 4716 4123
rect 4900 4117 4988 4123
rect 5060 4117 5100 4123
rect 5140 4117 5164 4123
rect 5172 4117 5324 4123
rect 5332 4117 5452 4123
rect 5460 4117 5692 4123
rect 484 4097 508 4103
rect 516 4097 828 4103
rect 836 4097 972 4103
rect 1012 4097 1036 4103
rect 1492 4097 1612 4103
rect 2244 4097 2428 4103
rect 2788 4097 2828 4103
rect 3540 4097 3596 4103
rect 3604 4097 3772 4103
rect 3828 4097 3932 4103
rect 3956 4097 4012 4103
rect 4020 4097 4412 4103
rect 4484 4097 4844 4103
rect 5028 4097 5164 4103
rect 5188 4097 5212 4103
rect 1620 4077 1708 4083
rect 2196 4077 2332 4083
rect 2916 4077 3324 4083
rect 3332 4077 3436 4083
rect 3924 4077 3948 4083
rect 4244 4077 4268 4083
rect 4276 4077 4332 4083
rect 4477 4083 4483 4096
rect 4340 4077 4483 4083
rect 4660 4077 4732 4083
rect 4740 4077 4860 4083
rect 4868 4077 5564 4083
rect 5572 4077 5676 4083
rect 868 4057 924 4063
rect 1588 4057 1628 4063
rect 4004 4057 4748 4063
rect 660 4037 908 4043
rect 916 4037 956 4043
rect 964 4037 1276 4043
rect 2580 4037 2636 4043
rect 4244 4037 4908 4043
rect 564 4017 748 4023
rect 756 4017 796 4023
rect 5092 4017 5548 4023
rect 1496 4014 1544 4016
rect 1496 4006 1500 4014
rect 1510 4006 1516 4014
rect 1524 4006 1530 4014
rect 1540 4006 1544 4014
rect 1496 4004 1544 4006
rect 4568 4014 4616 4016
rect 4568 4006 4572 4014
rect 4582 4006 4588 4014
rect 4596 4006 4602 4014
rect 4612 4006 4616 4014
rect 4568 4004 4616 4006
rect 1780 3997 1859 4003
rect 676 3977 1676 3983
rect 1853 3983 1859 3997
rect 1876 3997 2220 4003
rect 3268 3997 3372 4003
rect 3716 3997 3820 4003
rect 4852 3997 5036 4003
rect 5044 3997 5100 4003
rect 5108 3997 5580 4003
rect 6004 3997 6044 4003
rect 6052 3997 6060 4003
rect 1853 3977 2044 3983
rect 2836 3977 2924 3983
rect 2932 3977 2972 3983
rect 3300 3977 3404 3983
rect 3412 3977 3420 3983
rect 3844 3977 3932 3983
rect 4308 3977 4428 3983
rect 5300 3977 5516 3983
rect 5076 3957 6124 3963
rect 1332 3937 2092 3943
rect 2468 3937 2492 3943
rect 2500 3937 2540 3943
rect 4100 3937 4460 3943
rect 5172 3937 5612 3943
rect 548 3917 860 3923
rect 916 3917 972 3923
rect 1076 3917 1116 3923
rect 1316 3917 1372 3923
rect 2132 3917 2195 3923
rect 372 3897 396 3903
rect 468 3897 588 3903
rect 596 3897 668 3903
rect 756 3897 860 3903
rect 1092 3897 1180 3903
rect 1204 3897 1388 3903
rect 1988 3897 2172 3903
rect 2189 3903 2195 3917
rect 2260 3917 2524 3923
rect 4900 3917 5132 3923
rect 5492 3917 5660 3923
rect 2189 3897 2524 3903
rect 2644 3897 2668 3903
rect 2676 3897 4012 3903
rect 4516 3897 5084 3903
rect 5508 3897 5564 3903
rect 5588 3897 5612 3903
rect 5732 3897 5868 3903
rect 404 3877 428 3883
rect 436 3877 556 3883
rect 564 3877 780 3883
rect 788 3877 988 3883
rect 1085 3883 1091 3896
rect 996 3877 1091 3883
rect 1156 3877 1564 3883
rect 2116 3877 2268 3883
rect 4292 3877 4428 3883
rect 4756 3877 4940 3883
rect 5156 3877 5308 3883
rect 5556 3877 5596 3883
rect 5604 3877 5676 3883
rect 5684 3877 5724 3883
rect 5732 3877 5740 3883
rect 1124 3857 1196 3863
rect 1220 3857 1660 3863
rect 1668 3857 1836 3863
rect 2084 3857 2140 3863
rect 2820 3857 3212 3863
rect 3508 3857 3580 3863
rect 4452 3857 5612 3863
rect 468 3837 476 3843
rect 900 3837 1276 3843
rect 1348 3837 1388 3843
rect 1732 3837 2012 3843
rect 3220 3837 3612 3843
rect 4260 3837 4748 3843
rect 4852 3837 5116 3843
rect 5124 3837 5148 3843
rect 5540 3837 5660 3843
rect 5668 3837 5708 3843
rect 276 3817 396 3823
rect 404 3817 1068 3823
rect 1092 3817 1212 3823
rect 2292 3817 2572 3823
rect 2836 3817 2844 3823
rect 3140 3817 3180 3823
rect 3604 3817 3868 3823
rect 3876 3817 3964 3823
rect 4253 3823 4259 3836
rect 3972 3817 4259 3823
rect 4324 3817 4524 3823
rect 4532 3817 4844 3823
rect 5092 3817 5212 3823
rect 5348 3817 5372 3823
rect 3032 3814 3080 3816
rect 3032 3806 3036 3814
rect 3046 3806 3052 3814
rect 3060 3806 3066 3814
rect 3076 3806 3080 3814
rect 3032 3804 3080 3806
rect 788 3797 940 3803
rect 948 3797 1116 3803
rect 1124 3797 1324 3803
rect 2324 3797 2492 3803
rect 2516 3797 2812 3803
rect 2820 3797 2860 3803
rect 3428 3797 3756 3803
rect 3764 3797 3948 3803
rect 3965 3797 3980 3803
rect 820 3777 844 3783
rect 852 3777 924 3783
rect 932 3777 1292 3783
rect 1428 3777 1484 3783
rect 2196 3777 2268 3783
rect 3965 3783 3971 3797
rect 4052 3797 4748 3803
rect 5428 3797 5468 3803
rect 2820 3777 3971 3783
rect 4084 3777 4380 3783
rect 4388 3777 4572 3783
rect 68 3757 92 3763
rect 132 3757 332 3763
rect 708 3757 780 3763
rect 836 3757 892 3763
rect 1076 3757 1292 3763
rect 1300 3757 1324 3763
rect 1428 3757 1724 3763
rect 1908 3757 2300 3763
rect 3204 3757 3372 3763
rect 4180 3757 4428 3763
rect 4436 3757 4988 3763
rect 4996 3757 5068 3763
rect 5636 3757 5932 3763
rect -19 3737 12 3743
rect 68 3737 140 3743
rect 276 3737 380 3743
rect 388 3737 428 3743
rect 452 3737 492 3743
rect 500 3737 556 3743
rect 580 3737 908 3743
rect 1220 3737 1244 3743
rect 1252 3737 1372 3743
rect 1380 3737 1612 3743
rect 1876 3737 2044 3743
rect 2132 3737 2204 3743
rect 2276 3737 2604 3743
rect 2708 3737 2748 3743
rect 2756 3737 2764 3743
rect 2772 3737 2892 3743
rect 3396 3737 3564 3743
rect 4004 3737 4188 3743
rect 4484 3737 4684 3743
rect 4788 3737 4828 3743
rect 4836 3737 5004 3743
rect 5412 3737 5548 3743
rect 5652 3737 5692 3743
rect 52 3717 76 3723
rect 100 3717 156 3723
rect 292 3717 364 3723
rect 436 3717 492 3723
rect 820 3717 1036 3723
rect 1044 3717 1212 3723
rect 1220 3717 1228 3723
rect 1380 3717 1420 3723
rect 1540 3717 1596 3723
rect 2196 3717 2284 3723
rect 2644 3717 2668 3723
rect 3124 3717 3436 3723
rect 3444 3717 3468 3723
rect 4340 3717 4508 3723
rect 4660 3717 4764 3723
rect 4772 3717 4860 3723
rect 5588 3717 5772 3723
rect 5780 3717 5820 3723
rect 5908 3717 5932 3723
rect -19 3697 28 3703
rect 340 3697 348 3703
rect 356 3697 460 3703
rect 596 3697 732 3703
rect 740 3697 780 3703
rect 900 3697 1020 3703
rect 1229 3703 1235 3716
rect 1229 3697 1388 3703
rect 2068 3697 2124 3703
rect 2132 3697 2380 3703
rect 2708 3697 3084 3703
rect 3092 3697 3212 3703
rect 3220 3697 3308 3703
rect 3796 3697 3804 3703
rect 3812 3697 4236 3703
rect 4388 3697 4492 3703
rect 6132 3697 6163 3703
rect 324 3677 348 3683
rect 788 3677 1004 3683
rect 1332 3677 1452 3683
rect 2740 3677 4140 3683
rect 676 3657 908 3663
rect 916 3657 1308 3663
rect 1316 3657 1436 3663
rect 2452 3657 3100 3663
rect 5060 3657 5116 3663
rect 5124 3657 5516 3663
rect 5524 3657 5548 3663
rect 644 3637 764 3643
rect 772 3637 908 3643
rect 1268 3637 1420 3643
rect 1428 3637 1516 3643
rect 212 3617 428 3623
rect 1988 3617 2028 3623
rect 2196 3617 2220 3623
rect 5396 3617 5740 3623
rect 1496 3614 1544 3616
rect 1496 3606 1500 3614
rect 1510 3606 1516 3614
rect 1524 3606 1530 3614
rect 1540 3606 1544 3614
rect 1496 3604 1544 3606
rect 4568 3614 4616 3616
rect 4568 3606 4572 3614
rect 4582 3606 4588 3614
rect 4596 3606 4602 3614
rect 4612 3606 4616 3614
rect 4568 3604 4616 3606
rect 68 3597 92 3603
rect 1924 3597 2108 3603
rect 2356 3597 2412 3603
rect 3684 3597 4380 3603
rect 4804 3597 4828 3603
rect 5332 3597 5548 3603
rect 100 3577 284 3583
rect 1204 3577 1292 3583
rect 1540 3577 1564 3583
rect 2116 3577 2204 3583
rect 2676 3577 2812 3583
rect 420 3557 940 3563
rect 948 3557 2732 3563
rect 5396 3557 5516 3563
rect 564 3537 940 3543
rect 980 3537 1340 3543
rect 1348 3537 1468 3543
rect 1620 3537 3932 3543
rect 4916 3537 5324 3543
rect 5348 3537 5596 3543
rect 436 3517 812 3523
rect 916 3517 1052 3523
rect 1140 3517 1164 3523
rect 1172 3517 1196 3523
rect 1236 3517 1260 3523
rect 2596 3517 2892 3523
rect 3956 3517 4012 3523
rect 4084 3517 4124 3523
rect 4132 3517 4348 3523
rect 4356 3517 4460 3523
rect 5220 3517 5404 3523
rect 5588 3517 5612 3523
rect -19 3497 12 3503
rect 1044 3497 1276 3503
rect 1284 3497 1324 3503
rect 1588 3497 1708 3503
rect 2036 3497 2124 3503
rect 2340 3497 2380 3503
rect 2868 3497 3020 3503
rect 3188 3497 3379 3503
rect 3373 3484 3379 3497
rect 3476 3497 3884 3503
rect 3908 3497 3996 3503
rect 4052 3497 4092 3503
rect 4900 3497 4956 3503
rect 5188 3497 5676 3503
rect 5988 3497 6044 3503
rect 6132 3497 6163 3503
rect 164 3477 236 3483
rect 356 3477 508 3483
rect 564 3477 860 3483
rect 868 3477 924 3483
rect 932 3477 988 3483
rect 1140 3477 1308 3483
rect 2276 3477 2300 3483
rect 2484 3477 2732 3483
rect 2996 3477 3292 3483
rect 3748 3477 4044 3483
rect 4052 3477 4092 3483
rect 4612 3477 5068 3483
rect 5444 3477 5596 3483
rect 5604 3477 5660 3483
rect 5908 3477 6012 3483
rect 6020 3477 6060 3483
rect 180 3457 268 3463
rect 532 3457 2364 3463
rect 2372 3457 3276 3463
rect 3284 3457 3452 3463
rect 3524 3457 3788 3463
rect 4020 3457 4076 3463
rect 4084 3457 4156 3463
rect 4772 3457 5100 3463
rect 5108 3457 5228 3463
rect 1300 3437 1356 3443
rect 1748 3437 1964 3443
rect 3220 3437 3260 3443
rect 3716 3437 4492 3443
rect 100 3417 140 3423
rect 612 3417 812 3423
rect 820 3417 940 3423
rect 1204 3417 1244 3423
rect 1700 3417 1740 3423
rect 1956 3417 2108 3423
rect 2276 3417 2316 3423
rect 2324 3417 2380 3423
rect 3252 3417 3356 3423
rect 4148 3417 4316 3423
rect 5268 3417 5852 3423
rect 3032 3414 3080 3416
rect 3032 3406 3036 3414
rect 3046 3406 3052 3414
rect 3060 3406 3066 3414
rect 3076 3406 3080 3414
rect 3032 3404 3080 3406
rect 84 3397 124 3403
rect 916 3397 1452 3403
rect 1732 3397 1964 3403
rect 2516 3397 2572 3403
rect 2708 3397 2716 3403
rect 2932 3397 2940 3403
rect 3444 3397 3820 3403
rect 4036 3397 4524 3403
rect 4532 3397 4620 3403
rect 5268 3397 5308 3403
rect 5460 3397 6108 3403
rect 2932 3377 3324 3383
rect 3540 3377 4140 3383
rect 4324 3377 4348 3383
rect 5652 3377 5724 3383
rect 5956 3377 6028 3383
rect 516 3357 556 3363
rect 692 3357 764 3363
rect 772 3357 1084 3363
rect 1348 3357 1532 3363
rect 1540 3357 1708 3363
rect 2740 3357 2780 3363
rect 2788 3357 2828 3363
rect 3812 3357 4556 3363
rect 4676 3357 4908 3363
rect 5236 3357 5372 3363
rect 5380 3357 5564 3363
rect 5892 3357 5980 3363
rect 6036 3357 6076 3363
rect 804 3337 972 3343
rect 2548 3337 2684 3343
rect 3268 3337 3564 3343
rect 3764 3337 3916 3343
rect 4020 3337 4396 3343
rect 4516 3337 4652 3343
rect 4692 3337 4892 3343
rect 5380 3337 5388 3343
rect 5716 3337 5900 3343
rect 6084 3337 6092 3343
rect 6116 3337 6163 3343
rect -19 3317 412 3323
rect 548 3317 956 3323
rect 964 3317 1052 3323
rect 1284 3317 1308 3323
rect 1844 3317 1916 3323
rect 2212 3317 2876 3323
rect 2916 3317 2972 3323
rect 2980 3317 3052 3323
rect 3060 3317 3164 3323
rect 3268 3317 3292 3323
rect 3332 3317 3644 3323
rect 3652 3317 3740 3323
rect 3988 3317 4060 3323
rect 4397 3323 4403 3336
rect 4180 3317 4387 3323
rect 4397 3317 4780 3323
rect 1892 3297 2284 3303
rect 2324 3297 2812 3303
rect 2852 3297 2908 3303
rect 2996 3297 3292 3303
rect 3300 3297 3372 3303
rect 3732 3297 3852 3303
rect 3924 3297 4364 3303
rect 4381 3303 4387 3317
rect 4788 3317 4844 3323
rect 4948 3317 4956 3323
rect 5012 3317 5100 3323
rect 5268 3317 5292 3323
rect 5364 3317 5436 3323
rect 5444 3317 5548 3323
rect 5796 3317 5852 3323
rect 5860 3317 5932 3323
rect 5940 3317 5996 3323
rect 4381 3297 4412 3303
rect 4484 3297 4492 3303
rect 4516 3297 4684 3303
rect 4708 3297 4828 3303
rect 4836 3297 5052 3303
rect 2308 3277 2316 3283
rect 2964 3277 3004 3283
rect 3284 3277 3372 3283
rect 3748 3277 3788 3283
rect 4004 3277 4348 3283
rect 4356 3277 4540 3283
rect 4676 3277 4940 3283
rect 2196 3257 2540 3263
rect 3220 3257 3404 3263
rect 3764 3257 3788 3263
rect 4612 3257 4716 3263
rect 4724 3257 4876 3263
rect 132 3237 172 3243
rect 180 3237 316 3243
rect 2084 3237 2588 3243
rect 3380 3237 3772 3243
rect 4436 3237 4492 3243
rect 4500 3237 5468 3243
rect 532 3217 604 3223
rect 1044 3217 1100 3223
rect 2116 3217 2172 3223
rect 3156 3217 3244 3223
rect 3412 3217 3836 3223
rect 4916 3217 5100 3223
rect 5108 3217 5180 3223
rect 5204 3217 5244 3223
rect 5364 3217 5580 3223
rect 1496 3214 1544 3216
rect 1496 3206 1500 3214
rect 1510 3206 1516 3214
rect 1524 3206 1530 3214
rect 1540 3206 1544 3214
rect 1496 3204 1544 3206
rect 20 3197 140 3203
rect 148 3197 380 3203
rect 388 3197 1388 3203
rect 1396 3197 1420 3203
rect 3245 3203 3251 3216
rect 4568 3214 4616 3216
rect 4568 3206 4572 3214
rect 4582 3206 4588 3214
rect 4596 3206 4602 3214
rect 4612 3206 4616 3214
rect 4568 3204 4616 3206
rect 3245 3197 3980 3203
rect 4244 3197 4332 3203
rect 4452 3197 4508 3203
rect 4660 3197 5068 3203
rect 5076 3197 5212 3203
rect 452 3177 476 3183
rect 1028 3177 1100 3183
rect 1300 3177 1612 3183
rect 2068 3177 3468 3183
rect 3604 3177 3756 3183
rect 4004 3177 4044 3183
rect 4372 3177 4604 3183
rect 4621 3177 4812 3183
rect 2388 3157 3884 3163
rect 4036 3157 4188 3163
rect 4548 3157 4572 3163
rect 4621 3163 4627 3177
rect 4820 3177 4899 3183
rect 4596 3157 4627 3163
rect 4660 3157 4876 3163
rect 4893 3163 4899 3177
rect 4916 3177 5020 3183
rect 5028 3177 5132 3183
rect 5140 3177 5228 3183
rect 4893 3157 5004 3163
rect 2660 3137 2700 3143
rect 2900 3137 3116 3143
rect 3348 3137 3580 3143
rect 3588 3137 3724 3143
rect 3764 3137 4652 3143
rect 4788 3137 4812 3143
rect 4852 3137 5020 3143
rect 5044 3137 5084 3143
rect 5284 3137 5324 3143
rect 5844 3137 5868 3143
rect 804 3117 1180 3123
rect 1380 3117 1692 3123
rect 1924 3117 2044 3123
rect 2404 3117 2572 3123
rect 2589 3117 2716 3123
rect 580 3097 876 3103
rect 1044 3097 1292 3103
rect 1476 3097 1564 3103
rect 2340 3097 2380 3103
rect 2589 3103 2595 3117
rect 2740 3117 2748 3123
rect 2852 3117 2924 3123
rect 3492 3117 3708 3123
rect 3860 3117 3964 3123
rect 4020 3117 4076 3123
rect 4116 3117 4124 3123
rect 4756 3117 4796 3123
rect 4868 3117 5068 3123
rect 5124 3117 5212 3123
rect 5220 3117 5228 3123
rect 5300 3117 5388 3123
rect 5764 3117 5852 3123
rect 2484 3097 2595 3103
rect 2628 3097 2844 3103
rect 2852 3097 2972 3103
rect 3716 3097 3756 3103
rect 3796 3097 3836 3103
rect 3924 3097 4044 3103
rect 4084 3097 4172 3103
rect 4244 3097 4380 3103
rect 4676 3097 4684 3103
rect 4724 3097 4764 3103
rect 4964 3097 4988 3103
rect 5060 3097 5116 3103
rect 5268 3097 5340 3103
rect 6132 3097 6163 3103
rect 292 3077 492 3083
rect 724 3077 860 3083
rect 2621 3083 2627 3096
rect 980 3077 2627 3083
rect 2692 3077 2700 3083
rect 2804 3077 2828 3083
rect 2884 3077 2988 3083
rect 2996 3077 3324 3083
rect 3476 3077 3692 3083
rect 3780 3077 3788 3083
rect 3812 3077 3900 3083
rect 3924 3077 3932 3083
rect 3988 3077 4044 3083
rect 4052 3077 4092 3083
rect 4116 3077 4492 3083
rect 4500 3077 4908 3083
rect 5012 3077 5036 3083
rect 5172 3077 5292 3083
rect 5636 3077 5852 3083
rect 5908 3077 5996 3083
rect 324 3057 684 3063
rect 932 3057 2076 3063
rect 2148 3057 2460 3063
rect 2916 3057 3068 3063
rect 3076 3057 3244 3063
rect 3540 3057 3564 3063
rect 3572 3057 3948 3063
rect 3972 3057 4028 3063
rect 4148 3057 4172 3063
rect 4180 3057 4412 3063
rect 4804 3057 4924 3063
rect 4948 3057 5116 3063
rect 5396 3057 5420 3063
rect 5748 3057 5788 3063
rect 5828 3057 5932 3063
rect 5940 3057 6044 3063
rect 1700 3037 1804 3043
rect 1876 3037 2172 3043
rect 2180 3037 2348 3043
rect 2644 3037 2892 3043
rect 3188 3037 3388 3043
rect 4052 3037 4492 3043
rect 4516 3037 4812 3043
rect 5268 3037 5340 3043
rect 5556 3037 5660 3043
rect 5668 3037 5804 3043
rect 5812 3037 5932 3043
rect 1236 3017 1436 3023
rect 1588 3017 2636 3023
rect 2788 3017 2956 3023
rect 3908 3017 4012 3023
rect 4132 3017 4188 3023
rect 4212 3017 4428 3023
rect 4772 3017 4860 3023
rect 4980 3017 5004 3023
rect 5220 3017 5260 3023
rect 5268 3017 5420 3023
rect 5732 3017 5900 3023
rect 3032 3014 3080 3016
rect 3032 3006 3036 3014
rect 3046 3006 3052 3014
rect 3060 3006 3066 3014
rect 3076 3006 3080 3014
rect 3032 3004 3080 3006
rect 4164 2997 4348 3003
rect 4516 2997 4700 3003
rect 4724 2997 4883 3003
rect 2948 2977 2988 2983
rect 3124 2977 3164 2983
rect 3332 2977 3596 2983
rect 3780 2977 3884 2983
rect 3892 2977 4012 2983
rect 4877 2983 4883 2997
rect 4900 2997 5020 3003
rect 5908 2997 5948 3003
rect 4877 2977 4892 2983
rect 4900 2977 4940 2983
rect 5076 2977 5212 2983
rect 292 2957 572 2963
rect 596 2957 860 2963
rect 868 2957 1084 2963
rect 1268 2957 1388 2963
rect 1396 2957 1772 2963
rect 2484 2957 2828 2963
rect 2836 2957 3148 2963
rect 3396 2957 3484 2963
rect 3492 2957 3996 2963
rect 4164 2957 4172 2963
rect 4580 2957 4668 2963
rect 4941 2957 5004 2963
rect 148 2937 172 2943
rect 180 2937 316 2943
rect 324 2937 780 2943
rect 1012 2937 1052 2943
rect 1060 2937 1219 2943
rect 1213 2924 1219 2937
rect 1428 2937 1548 2943
rect 1844 2937 2044 2943
rect 2068 2937 2092 2943
rect 2324 2937 2572 2943
rect 2948 2937 3276 2943
rect 3300 2937 3516 2943
rect 3556 2937 3676 2943
rect 3748 2937 3804 2943
rect 3876 2937 3916 2943
rect 4388 2937 4476 2943
rect 4484 2937 4508 2943
rect 4644 2937 4732 2943
rect 4756 2937 4796 2943
rect 4836 2937 4844 2943
rect 4941 2943 4947 2957
rect 5076 2957 5196 2963
rect 5380 2957 5580 2963
rect 4900 2937 4947 2943
rect 4964 2937 5068 2943
rect 5076 2937 5100 2943
rect 5140 2937 5180 2943
rect 5364 2937 5420 2943
rect 5428 2937 5548 2943
rect 5812 2937 5932 2943
rect 756 2917 1020 2923
rect 1108 2917 1180 2923
rect 1220 2917 1564 2923
rect 1572 2917 1644 2923
rect 2004 2917 2220 2923
rect 2564 2917 2700 2923
rect 2804 2917 3052 2923
rect 3236 2917 3308 2923
rect 3460 2917 3612 2923
rect 3716 2917 4028 2923
rect 4404 2917 4476 2923
rect 4628 2917 4684 2923
rect 4788 2917 4924 2923
rect 4948 2917 4988 2923
rect 5220 2917 5260 2923
rect 5556 2917 5580 2923
rect 548 2897 588 2903
rect 964 2897 1116 2903
rect 1124 2897 1692 2903
rect 1700 2897 1964 2903
rect 2148 2897 2428 2903
rect 2436 2897 2924 2903
rect 2932 2897 3052 2903
rect 3156 2897 3228 2903
rect 3268 2897 3340 2903
rect 3524 2897 3596 2903
rect 3956 2897 4691 2903
rect 1524 2877 1756 2883
rect 2916 2877 3548 2883
rect 3668 2877 3804 2883
rect 3828 2877 4300 2883
rect 4356 2877 4524 2883
rect 4644 2877 4668 2883
rect 4685 2883 4691 2897
rect 4964 2897 5180 2903
rect 5316 2897 5388 2903
rect 5309 2883 5315 2896
rect 4685 2877 5315 2883
rect 1076 2857 1132 2863
rect 1140 2857 2668 2863
rect 3140 2857 3292 2863
rect 3348 2857 3420 2863
rect 3428 2857 3468 2863
rect 3636 2857 3852 2863
rect 3908 2857 3964 2863
rect 4052 2857 4060 2863
rect 4404 2857 4716 2863
rect 5012 2857 5212 2863
rect 404 2837 476 2843
rect 900 2837 940 2843
rect 1444 2837 2060 2843
rect 2084 2837 2364 2843
rect 2372 2837 2444 2843
rect 2932 2837 3148 2843
rect 3204 2837 3276 2843
rect 3700 2837 3836 2843
rect 4004 2837 4636 2843
rect 4660 2837 4812 2843
rect 5140 2837 5452 2843
rect 1876 2817 1916 2823
rect 2292 2817 2492 2823
rect 2676 2817 2764 2823
rect 3220 2817 3244 2823
rect 3364 2817 3644 2823
rect 3652 2817 3788 2823
rect 3796 2817 3852 2823
rect 4788 2817 4796 2823
rect 4884 2817 4972 2823
rect 5076 2817 5132 2823
rect 5140 2817 5308 2823
rect 6036 2817 6060 2823
rect 6068 2817 6092 2823
rect 1496 2814 1544 2816
rect 1496 2806 1500 2814
rect 1510 2806 1516 2814
rect 1524 2806 1530 2814
rect 1540 2806 1544 2814
rect 1496 2804 1544 2806
rect 4568 2814 4616 2816
rect 4568 2806 4572 2814
rect 4582 2806 4588 2814
rect 4596 2806 4602 2814
rect 4612 2806 4616 2814
rect 4568 2804 4616 2806
rect 820 2797 972 2803
rect 1956 2797 1996 2803
rect 2004 2797 2732 2803
rect 2740 2797 2796 2803
rect 2804 2797 2892 2803
rect 2900 2797 3260 2803
rect 3348 2797 3404 2803
rect 3421 2797 4332 2803
rect 2308 2777 2316 2783
rect 3421 2783 3427 2797
rect 4637 2797 4748 2803
rect 2516 2777 3427 2783
rect 3620 2777 3900 2783
rect 4020 2777 4204 2783
rect 4637 2783 4643 2797
rect 4916 2797 5052 2803
rect 5060 2797 5228 2803
rect 5300 2797 5372 2803
rect 4436 2777 4643 2783
rect 4660 2777 4684 2783
rect 4692 2777 5004 2783
rect 5204 2777 5324 2783
rect 1236 2757 1308 2763
rect 1748 2757 1964 2763
rect 1972 2757 3388 2763
rect 3732 2757 3820 2763
rect 4004 2757 4332 2763
rect 4676 2757 4748 2763
rect 4884 2757 5196 2763
rect 5284 2757 5292 2763
rect 5348 2757 5564 2763
rect 5572 2757 5676 2763
rect 5732 2757 5756 2763
rect 5764 2757 5788 2763
rect 852 2737 924 2743
rect 1108 2737 1228 2743
rect 1236 2737 2124 2743
rect 2180 2737 2803 2743
rect 660 2717 684 2723
rect 692 2717 924 2723
rect 1652 2717 1692 2723
rect 2228 2717 2780 2723
rect 2797 2723 2803 2737
rect 2964 2737 2988 2743
rect 3028 2737 3436 2743
rect 3460 2737 3564 2743
rect 3572 2737 3820 2743
rect 3828 2737 3916 2743
rect 4084 2737 4108 2743
rect 4148 2737 4172 2743
rect 4356 2737 4396 2743
rect 4516 2737 4828 2743
rect 4900 2737 5100 2743
rect 5172 2737 5340 2743
rect 5588 2737 5644 2743
rect 5652 2737 5756 2743
rect 2797 2717 3484 2723
rect 3524 2717 3564 2723
rect 3652 2717 3660 2723
rect 3700 2717 3756 2723
rect 3780 2717 4444 2723
rect 4548 2717 4780 2723
rect 4836 2717 5020 2723
rect 5028 2717 5404 2723
rect 5412 2717 5452 2723
rect 5460 2717 5500 2723
rect 260 2697 284 2703
rect 292 2697 460 2703
rect 548 2697 748 2703
rect 756 2697 780 2703
rect 1044 2697 1148 2703
rect 1636 2697 1756 2703
rect 1764 2697 1788 2703
rect 2132 2697 2684 2703
rect 2772 2697 3500 2703
rect 3556 2697 3596 2703
rect 3684 2697 3724 2703
rect 3764 2697 3820 2703
rect 3844 2697 3948 2703
rect 3956 2697 4092 2703
rect 4100 2697 4124 2703
rect 4276 2697 4316 2703
rect 4436 2697 4460 2703
rect 4756 2697 4780 2703
rect 4788 2697 4860 2703
rect 4964 2697 5036 2703
rect 5092 2697 5164 2703
rect 5204 2697 5276 2703
rect 5348 2697 5388 2703
rect 5700 2697 5788 2703
rect 5796 2697 5868 2703
rect 148 2677 748 2683
rect 781 2677 796 2683
rect 804 2677 828 2683
rect 836 2677 876 2683
rect 884 2677 1004 2683
rect 1140 2677 1244 2683
rect 1892 2677 1907 2683
rect 180 2657 540 2663
rect 580 2657 812 2663
rect 916 2657 1180 2663
rect 1684 2657 1884 2663
rect 1901 2663 1907 2677
rect 2084 2677 2124 2683
rect 2452 2677 2700 2683
rect 2996 2677 3004 2683
rect 3092 2677 3228 2683
rect 3284 2677 3404 2683
rect 3444 2677 3948 2683
rect 3972 2677 4044 2683
rect 4164 2677 4323 2683
rect 1901 2657 2204 2663
rect 2644 2657 2780 2663
rect 2852 2657 3004 2663
rect 3156 2657 3244 2663
rect 3252 2657 3260 2663
rect 3876 2657 4012 2663
rect 4020 2657 4076 2663
rect 4084 2657 4204 2663
rect 4317 2663 4323 2677
rect 4340 2677 4412 2683
rect 4749 2677 4764 2683
rect 4749 2663 4755 2677
rect 4868 2677 4972 2683
rect 4980 2677 5100 2683
rect 5108 2677 5420 2683
rect 5428 2677 5484 2683
rect 5556 2677 5644 2683
rect 5780 2677 5980 2683
rect 6036 2677 6044 2683
rect 4317 2657 4755 2663
rect 4772 2657 4796 2663
rect 4804 2657 4844 2663
rect 4852 2657 4956 2663
rect 5012 2657 5148 2663
rect 5172 2657 5244 2663
rect 5268 2657 5436 2663
rect 5444 2657 5484 2663
rect 5876 2657 5948 2663
rect 340 2637 364 2643
rect 372 2637 716 2643
rect 1508 2637 1916 2643
rect 1924 2637 2108 2643
rect 2676 2637 2812 2643
rect 2820 2637 2956 2643
rect 2964 2637 3596 2643
rect 3732 2637 3772 2643
rect 3796 2637 4060 2643
rect 4068 2637 4172 2643
rect 4180 2637 4252 2643
rect 4260 2637 4316 2643
rect 4324 2637 4684 2643
rect 4756 2637 4876 2643
rect 4948 2637 5020 2643
rect 5044 2637 5052 2643
rect 5076 2637 5084 2643
rect 5220 2637 5580 2643
rect 1700 2617 1868 2623
rect 1892 2617 2140 2623
rect 2148 2617 2172 2623
rect 3540 2617 3660 2623
rect 3684 2617 3868 2623
rect 3885 2617 4172 2623
rect 3032 2614 3080 2616
rect 3032 2606 3036 2614
rect 3046 2606 3052 2614
rect 3060 2606 3066 2614
rect 3076 2606 3080 2614
rect 3032 2604 3080 2606
rect 1156 2597 1196 2603
rect 1668 2597 1852 2603
rect 1940 2597 1996 2603
rect 3508 2597 3628 2603
rect 3885 2603 3891 2617
rect 4276 2617 4300 2623
rect 4340 2617 4636 2623
rect 4724 2617 4780 2623
rect 4852 2617 4956 2623
rect 5028 2617 5196 2623
rect 5364 2617 5420 2623
rect 3684 2597 3891 2603
rect 4036 2597 4140 2603
rect 4164 2597 4204 2603
rect 4212 2597 4284 2603
rect 4292 2597 4412 2603
rect 4548 2597 4652 2603
rect 4660 2597 4780 2603
rect 4788 2597 5004 2603
rect 5044 2597 5148 2603
rect 5236 2597 5308 2603
rect 5476 2597 5772 2603
rect 2436 2577 2668 2583
rect 2708 2577 2860 2583
rect 2916 2577 3171 2583
rect 388 2557 748 2563
rect 1012 2557 1116 2563
rect 1124 2557 1260 2563
rect 1268 2557 1612 2563
rect 2484 2557 2604 2563
rect 2612 2557 2668 2563
rect 2852 2557 2876 2563
rect 2884 2557 3132 2563
rect 3165 2563 3171 2577
rect 3188 2577 3900 2583
rect 3924 2577 4668 2583
rect 4724 2577 4924 2583
rect 5028 2577 5068 2583
rect 5124 2577 5180 2583
rect 5188 2577 5292 2583
rect 5300 2577 5468 2583
rect 5620 2577 5708 2583
rect 3165 2557 3276 2563
rect 3284 2557 3372 2563
rect 3396 2557 3500 2563
rect 3508 2557 3756 2563
rect 3988 2557 4060 2563
rect 4196 2557 4236 2563
rect 4308 2557 4364 2563
rect 4420 2557 4508 2563
rect 4804 2557 4828 2563
rect 4845 2557 4892 2563
rect 1652 2537 1820 2543
rect 2084 2537 2332 2543
rect 2372 2537 2396 2543
rect 2740 2537 2908 2543
rect 2964 2537 3036 2543
rect 3092 2537 3148 2543
rect 3428 2537 3468 2543
rect 3476 2537 3660 2543
rect 4148 2537 4268 2543
rect 4404 2537 4476 2543
rect 4532 2537 4556 2543
rect 4580 2537 4700 2543
rect 4845 2543 4851 2557
rect 5060 2557 5100 2563
rect 5108 2557 5292 2563
rect 5300 2557 5340 2563
rect 5364 2557 5420 2563
rect 5428 2557 5452 2563
rect 4708 2537 4851 2543
rect 4884 2537 4892 2543
rect 4900 2537 4972 2543
rect 4980 2537 5260 2543
rect 5332 2537 5372 2543
rect 5652 2537 5900 2543
rect 260 2517 412 2523
rect 644 2517 684 2523
rect 1252 2517 1308 2523
rect 1380 2517 1532 2523
rect 1540 2517 2252 2523
rect 2260 2517 2476 2523
rect 3085 2523 3091 2536
rect 2980 2517 3091 2523
rect 3204 2517 3212 2523
rect 3220 2517 3468 2523
rect 4004 2517 4044 2523
rect 4084 2517 4204 2523
rect 4244 2517 4524 2523
rect 4596 2517 4716 2523
rect 4852 2517 5084 2523
rect 5108 2517 5116 2523
rect 5124 2517 5180 2523
rect 5204 2517 5276 2523
rect 5284 2517 5388 2523
rect 3156 2497 3180 2503
rect 3252 2497 3436 2503
rect 4148 2497 4172 2503
rect 4212 2497 4236 2503
rect 4244 2497 4284 2503
rect 4340 2497 4396 2503
rect 4404 2497 4524 2503
rect 4564 2497 4652 2503
rect 4836 2497 4844 2503
rect 4964 2497 5020 2503
rect 5172 2497 5388 2503
rect 2452 2477 2588 2483
rect 3172 2477 3196 2483
rect 3252 2477 3292 2483
rect 3380 2477 3452 2483
rect 3476 2477 4652 2483
rect 4676 2477 5612 2483
rect 3012 2457 3148 2463
rect 3172 2457 3468 2463
rect 4020 2457 4092 2463
rect 4100 2457 4476 2463
rect 4532 2457 4844 2463
rect 5012 2457 5052 2463
rect 5108 2457 5452 2463
rect 516 2437 956 2443
rect 1364 2437 1452 2443
rect 1460 2437 1788 2443
rect 2420 2437 2508 2443
rect 2516 2437 2924 2443
rect 3108 2437 3212 2443
rect 3252 2437 3260 2443
rect 3460 2437 4060 2443
rect 4116 2437 4220 2443
rect 4244 2437 4652 2443
rect 4916 2437 5036 2443
rect 5044 2437 5356 2443
rect 5396 2437 5516 2443
rect 372 2417 716 2423
rect 724 2417 780 2423
rect 1636 2417 1820 2423
rect 1828 2417 1868 2423
rect 2212 2417 3532 2423
rect 3540 2417 4108 2423
rect 4180 2417 4188 2423
rect 4644 2417 4684 2423
rect 4724 2417 4812 2423
rect 4836 2417 5004 2423
rect 5044 2417 5372 2423
rect 1496 2414 1544 2416
rect 1496 2406 1500 2414
rect 1510 2406 1516 2414
rect 1524 2406 1530 2414
rect 1540 2406 1544 2414
rect 1496 2404 1544 2406
rect 4568 2414 4616 2416
rect 4568 2406 4572 2414
rect 4582 2406 4588 2414
rect 4596 2406 4602 2414
rect 4612 2406 4616 2414
rect 4568 2404 4616 2406
rect 228 2397 524 2403
rect 2788 2397 3619 2403
rect 1828 2377 1932 2383
rect 2276 2377 3468 2383
rect 3524 2377 3596 2383
rect 3613 2383 3619 2397
rect 3844 2397 3884 2403
rect 3892 2397 4236 2403
rect 4372 2397 4540 2403
rect 4756 2397 4908 2403
rect 5156 2397 5228 2403
rect 5236 2397 5411 2403
rect 5405 2384 5411 2397
rect 3613 2377 4636 2383
rect 4964 2377 5068 2383
rect 5412 2377 5548 2383
rect 5668 2377 5740 2383
rect 5876 2377 5884 2383
rect 196 2357 300 2363
rect 308 2357 332 2363
rect 3028 2357 3532 2363
rect 4052 2357 4076 2363
rect 4100 2357 5052 2363
rect 5076 2357 5116 2363
rect 5268 2357 5308 2363
rect 5332 2357 5660 2363
rect -19 2337 12 2343
rect 132 2337 156 2343
rect 836 2337 1244 2343
rect 3220 2337 3356 2343
rect 3364 2337 3420 2343
rect 3428 2337 3484 2343
rect 3492 2337 3516 2343
rect 4004 2337 4044 2343
rect 4052 2337 4764 2343
rect 4884 2337 4924 2343
rect 5092 2337 5196 2343
rect 5204 2337 5308 2343
rect 5316 2337 5436 2343
rect 5972 2337 6044 2343
rect 100 2317 220 2323
rect 260 2317 332 2323
rect 948 2317 988 2323
rect 2724 2317 2732 2323
rect 2996 2317 3020 2323
rect 3044 2317 3132 2323
rect 3156 2317 3404 2323
rect 3476 2317 3516 2323
rect 3556 2317 4076 2323
rect 4292 2317 4508 2323
rect 4516 2317 4700 2323
rect 4708 2317 4716 2323
rect 4756 2317 4780 2323
rect 4820 2317 4844 2323
rect 4852 2317 4876 2323
rect 4964 2317 5244 2323
rect 5316 2317 5324 2323
rect 5460 2317 5484 2323
rect 5508 2317 5628 2323
rect 5876 2317 6044 2323
rect -19 2297 44 2303
rect 164 2297 188 2303
rect 244 2297 268 2303
rect 276 2297 764 2303
rect 772 2297 828 2303
rect 836 2297 1308 2303
rect 1316 2297 1340 2303
rect 2445 2297 2652 2303
rect 2445 2284 2451 2297
rect 2676 2297 2876 2303
rect 2980 2297 3116 2303
rect 3204 2297 3212 2303
rect 3588 2297 3596 2303
rect 3652 2297 4012 2303
rect 4116 2297 4140 2303
rect 4532 2297 4780 2303
rect 4948 2297 4972 2303
rect 5012 2297 5068 2303
rect 5076 2297 5308 2303
rect 5396 2297 5420 2303
rect 5588 2297 5628 2303
rect 6036 2297 6044 2303
rect 36 2277 76 2283
rect 196 2277 332 2283
rect 436 2277 572 2283
rect 852 2277 1020 2283
rect 1860 2277 2275 2283
rect 68 2257 204 2263
rect 228 2257 412 2263
rect 692 2257 2252 2263
rect 2269 2263 2275 2277
rect 2308 2277 2316 2283
rect 2644 2277 2748 2283
rect 2948 2277 3036 2283
rect 3060 2277 3484 2283
rect 3572 2277 3708 2283
rect 3732 2277 3804 2283
rect 3828 2277 4156 2283
rect 4164 2277 4284 2283
rect 4292 2277 4300 2283
rect 4484 2277 4556 2283
rect 4692 2277 4716 2283
rect 4836 2277 5084 2283
rect 5140 2277 5196 2283
rect 5348 2277 5596 2283
rect 5732 2277 6028 2283
rect 2269 2257 2828 2263
rect 2836 2257 3340 2263
rect 3348 2257 3548 2263
rect 3668 2257 4108 2263
rect 4452 2257 4668 2263
rect 5204 2257 5260 2263
rect 5268 2257 5516 2263
rect 5860 2257 6044 2263
rect 884 2237 1324 2243
rect 2180 2237 2204 2243
rect 2452 2237 3500 2243
rect 3508 2237 4348 2243
rect 4356 2237 4460 2243
rect 4468 2237 4588 2243
rect 4660 2237 4684 2243
rect 5316 2237 5484 2243
rect 564 2217 844 2223
rect 2020 2217 2092 2223
rect 2500 2217 2956 2223
rect 3380 2217 3820 2223
rect 4020 2217 5004 2223
rect 5012 2217 5180 2223
rect 5188 2217 5228 2223
rect 5236 2217 5292 2223
rect 5476 2217 5692 2223
rect 3032 2214 3080 2216
rect 3032 2206 3036 2214
rect 3046 2206 3052 2214
rect 3060 2206 3066 2214
rect 3076 2206 3080 2214
rect 3032 2204 3080 2206
rect 612 2197 668 2203
rect 3476 2197 3516 2203
rect 3684 2197 3836 2203
rect 4420 2197 4604 2203
rect 4644 2197 4748 2203
rect 4980 2197 5052 2203
rect 5060 2197 5388 2203
rect 5396 2197 5532 2203
rect 5572 2197 5916 2203
rect 932 2177 956 2183
rect 964 2177 1068 2183
rect 1076 2177 1500 2183
rect 1508 2177 1660 2183
rect 1732 2177 1980 2183
rect 2292 2177 2476 2183
rect 3012 2177 4828 2183
rect 5332 2177 5580 2183
rect 164 2157 316 2163
rect 756 2157 1004 2163
rect 1188 2157 1228 2163
rect 1661 2163 1667 2176
rect 1661 2157 1948 2163
rect 1956 2157 2044 2163
rect 2612 2157 2668 2163
rect 2756 2157 3180 2163
rect 3412 2157 3564 2163
rect 3716 2157 3868 2163
rect 4564 2157 4812 2163
rect 5124 2157 5676 2163
rect 244 2137 332 2143
rect 340 2137 396 2143
rect 404 2137 460 2143
rect 932 2137 1020 2143
rect 1108 2137 1244 2143
rect 1252 2137 1436 2143
rect 1652 2137 1756 2143
rect 2228 2137 2252 2143
rect 2644 2137 2796 2143
rect 2980 2137 3020 2143
rect 3028 2137 3372 2143
rect 3508 2137 3852 2143
rect 4116 2137 4204 2143
rect 4260 2137 4460 2143
rect 5172 2137 5356 2143
rect 5364 2137 5468 2143
rect 5556 2137 5788 2143
rect 52 2117 60 2123
rect 68 2117 92 2123
rect 148 2117 188 2123
rect 836 2117 1084 2123
rect 1140 2117 1164 2123
rect 2052 2117 2124 2123
rect 2132 2117 2156 2123
rect 2324 2117 3900 2123
rect 4852 2117 5196 2123
rect 5684 2117 5772 2123
rect -19 2097 12 2103
rect 100 2097 188 2103
rect 228 2097 268 2103
rect 276 2097 332 2103
rect 1085 2103 1091 2116
rect 1085 2097 1212 2103
rect 1348 2097 1484 2103
rect 3828 2097 3884 2103
rect 4116 2097 4124 2103
rect 4132 2097 4268 2103
rect 4900 2097 5036 2103
rect 5124 2097 5132 2103
rect 5652 2097 5740 2103
rect 260 2077 348 2083
rect 772 2077 796 2083
rect 804 2077 1052 2083
rect 1316 2077 1372 2083
rect 1460 2077 1660 2083
rect 2836 2057 2876 2063
rect 2884 2057 5164 2063
rect 2308 2037 2316 2043
rect 2372 2037 2444 2043
rect 3220 2037 3244 2043
rect 3460 2037 3468 2043
rect 3908 2037 5116 2043
rect 5684 2037 5724 2043
rect 788 2017 844 2023
rect 3108 2017 3116 2023
rect 3748 2017 3788 2023
rect 1496 2014 1544 2016
rect 1496 2006 1500 2014
rect 1510 2006 1516 2014
rect 1524 2006 1530 2014
rect 1540 2006 1544 2014
rect 1496 2004 1544 2006
rect 4568 2014 4616 2016
rect 4568 2006 4572 2014
rect 4582 2006 4588 2014
rect 4596 2006 4602 2014
rect 4612 2006 4616 2014
rect 4568 2004 4616 2006
rect 4340 1997 4428 2003
rect 4436 1997 4508 2003
rect 852 1977 860 1983
rect 996 1977 1068 1983
rect 1076 1977 1116 1983
rect 1124 1977 1356 1983
rect 1364 1977 1420 1983
rect 1428 1977 1612 1983
rect 1620 1977 1644 1983
rect 4116 1977 4172 1983
rect 5780 1977 5900 1983
rect 580 1957 700 1963
rect 2724 1957 2908 1963
rect 2916 1957 3180 1963
rect 3188 1957 3404 1963
rect 3412 1957 3676 1963
rect 3684 1957 3820 1963
rect 4804 1957 5068 1963
rect 388 1937 716 1943
rect 724 1937 732 1943
rect 740 1937 1148 1943
rect 2452 1937 2860 1943
rect 2868 1937 2876 1943
rect 3540 1937 3580 1943
rect 3588 1937 3660 1943
rect 4132 1937 4812 1943
rect 5044 1937 5180 1943
rect 5268 1937 5948 1943
rect 260 1917 476 1923
rect 596 1917 668 1923
rect 708 1917 780 1923
rect 948 1917 1084 1923
rect 1124 1917 1212 1923
rect 2004 1917 2476 1923
rect 4772 1917 4956 1923
rect 4996 1917 5020 1923
rect 5108 1917 5372 1923
rect 5764 1917 5980 1923
rect 484 1897 588 1903
rect 628 1897 716 1903
rect 1028 1897 1084 1903
rect 1284 1897 1356 1903
rect 1364 1897 1452 1903
rect 1524 1897 1596 1903
rect 1604 1897 1708 1903
rect 2068 1897 2076 1903
rect 2100 1897 2348 1903
rect 2500 1897 2588 1903
rect 2868 1897 2956 1903
rect 3124 1897 3132 1903
rect 3140 1897 3180 1903
rect 3188 1897 3468 1903
rect 3476 1897 3612 1903
rect 3620 1897 3660 1903
rect 3668 1897 4028 1903
rect 4676 1897 4684 1903
rect 4772 1897 4796 1903
rect 4948 1897 5132 1903
rect 5140 1897 5292 1903
rect 5604 1897 5660 1903
rect 5956 1897 6028 1903
rect 6132 1897 6163 1903
rect 68 1877 140 1883
rect 340 1877 380 1883
rect 692 1877 892 1883
rect 932 1877 1244 1883
rect 1252 1877 1276 1883
rect 1284 1877 1324 1883
rect 1732 1877 1932 1883
rect 2116 1877 2156 1883
rect 2244 1877 2316 1883
rect 2324 1877 2380 1883
rect 2484 1877 2684 1883
rect 2964 1877 3004 1883
rect 3636 1877 3852 1883
rect 3972 1877 4044 1883
rect 4052 1877 4348 1883
rect 4356 1877 4380 1883
rect 4516 1877 4812 1883
rect 5204 1877 5756 1883
rect 6036 1877 6092 1883
rect 68 1857 172 1863
rect 180 1857 412 1863
rect 500 1857 796 1863
rect 804 1857 1340 1863
rect 1348 1857 1500 1863
rect 1780 1857 1900 1863
rect 2068 1857 2124 1863
rect 2237 1863 2243 1876
rect 2132 1857 2243 1863
rect 2932 1857 3084 1863
rect 3828 1857 4156 1863
rect 4388 1857 5036 1863
rect 5044 1857 5228 1863
rect 5460 1857 5548 1863
rect 5748 1857 5788 1863
rect 372 1837 380 1843
rect 1140 1837 1212 1843
rect 2052 1837 2140 1843
rect 2148 1837 2332 1843
rect 2340 1837 2396 1843
rect 2404 1837 2940 1843
rect 3412 1837 3436 1843
rect 4052 1837 4076 1843
rect 4324 1837 5004 1843
rect 5172 1837 5228 1843
rect 6020 1837 6076 1843
rect 324 1817 380 1823
rect 388 1817 652 1823
rect 676 1817 828 1823
rect 1908 1817 2252 1823
rect 2260 1817 2540 1823
rect 3172 1817 3436 1823
rect 3444 1817 3468 1823
rect 3812 1817 4124 1823
rect 4484 1817 4508 1823
rect 5156 1817 5196 1823
rect 5732 1817 5804 1823
rect 3032 1814 3080 1816
rect 3032 1806 3036 1814
rect 3046 1806 3052 1814
rect 3060 1806 3066 1814
rect 3076 1806 3080 1814
rect 3032 1804 3080 1806
rect 788 1797 1100 1803
rect 1236 1797 1388 1803
rect 2084 1797 2188 1803
rect 2196 1797 2860 1803
rect 3220 1797 3372 1803
rect 3540 1797 3980 1803
rect 4980 1797 5100 1803
rect 5796 1797 5820 1803
rect 308 1777 396 1783
rect 532 1777 732 1783
rect 740 1777 876 1783
rect 884 1777 940 1783
rect 1044 1777 1148 1783
rect 1156 1777 1228 1783
rect 1940 1777 2220 1783
rect 2260 1777 2284 1783
rect 2756 1777 2892 1783
rect 3476 1777 3564 1783
rect 3716 1777 3916 1783
rect 4244 1777 4748 1783
rect 4756 1777 4988 1783
rect 5028 1777 5548 1783
rect 260 1757 300 1763
rect 644 1757 812 1763
rect 836 1757 908 1763
rect 1268 1757 1468 1763
rect 1476 1757 1788 1763
rect 1956 1757 2092 1763
rect 2132 1757 2412 1763
rect 2996 1757 3148 1763
rect 3197 1757 3500 1763
rect 772 1737 828 1743
rect 852 1737 1052 1743
rect 1060 1737 1292 1743
rect 1940 1737 2460 1743
rect 2564 1737 2764 1743
rect 2820 1737 2908 1743
rect 3197 1743 3203 1757
rect 3988 1757 4108 1763
rect 4148 1757 4172 1763
rect 4708 1757 5452 1763
rect 5524 1757 5676 1763
rect 5812 1757 5916 1763
rect 3156 1737 3203 1743
rect 3444 1737 3484 1743
rect 3572 1737 3644 1743
rect 3700 1737 3772 1743
rect 4020 1737 4332 1743
rect 4468 1737 4700 1743
rect 4836 1737 4924 1743
rect 5076 1737 5212 1743
rect 5300 1737 5436 1743
rect 5444 1737 5516 1743
rect 5860 1737 5996 1743
rect 100 1717 204 1723
rect 244 1717 316 1723
rect 804 1717 812 1723
rect 820 1717 1132 1723
rect 1220 1717 1292 1723
rect 1300 1717 1404 1723
rect 1412 1717 1564 1723
rect 1812 1717 1820 1723
rect 1828 1717 1852 1723
rect 2020 1717 2284 1723
rect 3268 1717 3324 1723
rect 3460 1717 3644 1723
rect 3700 1717 4316 1723
rect 4340 1717 4492 1723
rect 4724 1717 4780 1723
rect 5044 1717 5276 1723
rect 5380 1717 5580 1723
rect 5668 1717 5740 1723
rect 212 1697 236 1703
rect 660 1697 828 1703
rect 1380 1697 1964 1703
rect 1972 1697 1996 1703
rect 2020 1697 2092 1703
rect 2100 1697 2156 1703
rect 3348 1697 3404 1703
rect 3412 1697 3420 1703
rect 3556 1697 3628 1703
rect 3636 1697 3740 1703
rect 3812 1697 3820 1703
rect 3860 1697 4092 1703
rect 4100 1697 4172 1703
rect 4452 1697 4524 1703
rect 4660 1697 4748 1703
rect 4772 1697 4892 1703
rect 5124 1697 5196 1703
rect 5252 1697 5340 1703
rect 5348 1697 5452 1703
rect 5572 1697 5628 1703
rect 5652 1697 5996 1703
rect 6132 1697 6163 1703
rect 196 1677 204 1683
rect 212 1677 284 1683
rect 420 1677 1356 1683
rect 1364 1677 1580 1683
rect 1684 1677 1772 1683
rect 1780 1677 2252 1683
rect 3524 1677 3612 1683
rect 4164 1677 4204 1683
rect 4212 1677 4460 1683
rect 4532 1677 4572 1683
rect 4868 1677 4924 1683
rect 5117 1683 5123 1696
rect 4932 1677 5123 1683
rect 5300 1677 5420 1683
rect 5604 1677 5628 1683
rect 5636 1677 5644 1683
rect 5684 1677 5996 1683
rect 6004 1677 6028 1683
rect 788 1657 988 1663
rect 1076 1657 1420 1663
rect 1428 1657 1516 1663
rect 3188 1657 3404 1663
rect 3412 1657 3804 1663
rect 4548 1657 4684 1663
rect 4692 1657 4828 1663
rect 5028 1657 5196 1663
rect 1428 1637 2060 1643
rect 4084 1637 5292 1643
rect 1620 1617 1916 1623
rect 4068 1617 4108 1623
rect 1496 1614 1544 1616
rect 1496 1606 1500 1614
rect 1510 1606 1516 1614
rect 1524 1606 1530 1614
rect 1540 1606 1544 1614
rect 1496 1604 1544 1606
rect 4568 1614 4616 1616
rect 4568 1606 4572 1614
rect 4582 1606 4588 1614
rect 4596 1606 4602 1614
rect 4612 1606 4616 1614
rect 4568 1604 4616 1606
rect 276 1597 428 1603
rect 436 1597 572 1603
rect 580 1597 1404 1603
rect 2420 1597 2588 1603
rect 2596 1597 2812 1603
rect 2820 1597 2844 1603
rect 2980 1597 3196 1603
rect 4708 1597 5068 1603
rect 5140 1597 5388 1603
rect 5396 1597 5516 1603
rect 5828 1597 5852 1603
rect 5972 1597 5980 1603
rect 292 1577 1036 1583
rect 1709 1583 1715 1596
rect 1524 1577 1715 1583
rect 4052 1577 4092 1583
rect 4132 1577 4796 1583
rect 4852 1577 5180 1583
rect 692 1557 732 1563
rect 948 1557 1068 1563
rect 1124 1557 1148 1563
rect 1172 1557 1228 1563
rect 1348 1557 1356 1563
rect 1412 1557 1612 1563
rect 2244 1557 2572 1563
rect 2580 1557 2924 1563
rect 3572 1557 3708 1563
rect 3908 1557 4028 1563
rect 4292 1557 4604 1563
rect 4676 1557 4700 1563
rect 4852 1557 5244 1563
rect 5460 1557 5756 1563
rect 276 1537 380 1543
rect 564 1537 636 1543
rect 644 1537 892 1543
rect 1124 1537 1292 1543
rect 2724 1537 2780 1543
rect 3524 1537 3580 1543
rect 3588 1537 3660 1543
rect 3988 1537 4044 1543
rect 4516 1537 4556 1543
rect 4884 1537 5052 1543
rect 468 1517 508 1523
rect 516 1517 780 1523
rect 964 1517 1020 1523
rect 1092 1517 1164 1523
rect 1316 1517 2140 1523
rect 2148 1517 2604 1523
rect 3716 1517 3772 1523
rect 3789 1517 3852 1523
rect 84 1497 332 1503
rect 404 1497 636 1503
rect 676 1497 764 1503
rect 932 1497 1052 1503
rect 1188 1497 1276 1503
rect 2020 1497 2044 1503
rect 2052 1497 2140 1503
rect 2148 1497 2204 1503
rect 2212 1497 2524 1503
rect 3108 1497 3116 1503
rect 3444 1497 3596 1503
rect 3789 1503 3795 1517
rect 3892 1517 3964 1523
rect 4020 1517 4140 1523
rect 4148 1517 4284 1523
rect 4324 1517 4476 1523
rect 4500 1517 4508 1523
rect 4900 1517 5100 1523
rect 5108 1517 5164 1523
rect 6132 1517 6163 1523
rect 3764 1497 3795 1503
rect 3860 1497 3932 1503
rect 4004 1497 4060 1503
rect 4308 1497 4412 1503
rect 4484 1497 4668 1503
rect 4820 1497 4908 1503
rect 5092 1497 5276 1503
rect 5332 1497 5372 1503
rect 5412 1497 5500 1503
rect 196 1477 316 1483
rect 324 1477 460 1483
rect 548 1477 684 1483
rect 1124 1477 1244 1483
rect 1284 1477 1372 1483
rect 1748 1477 1980 1483
rect 2180 1477 2220 1483
rect 2788 1477 2988 1483
rect 3332 1477 3548 1483
rect 3828 1477 3900 1483
rect 3956 1477 4124 1483
rect 4180 1477 4716 1483
rect 4820 1477 4892 1483
rect 5044 1477 5068 1483
rect 5332 1477 5452 1483
rect 5636 1477 5692 1483
rect 5876 1477 5884 1483
rect 6052 1477 6163 1483
rect 372 1457 396 1463
rect 996 1457 1196 1463
rect 1236 1457 1260 1463
rect 1348 1457 1404 1463
rect 1412 1457 1484 1463
rect 2052 1457 2188 1463
rect 2196 1457 2492 1463
rect 2900 1457 3228 1463
rect 3364 1457 3484 1463
rect 3556 1457 3692 1463
rect 3700 1457 4380 1463
rect 4724 1457 4828 1463
rect 4868 1457 5004 1463
rect 5252 1457 5356 1463
rect 260 1437 380 1443
rect 388 1437 684 1443
rect 1028 1437 1356 1443
rect 2164 1437 2380 1443
rect 3092 1437 3644 1443
rect 3748 1437 4316 1443
rect 4644 1437 4780 1443
rect 5236 1437 5372 1443
rect 5700 1437 5708 1443
rect 388 1417 412 1423
rect 724 1417 828 1423
rect 1780 1417 1804 1423
rect 3812 1417 4972 1423
rect 5364 1417 5788 1423
rect 5860 1417 5868 1423
rect 5876 1417 5916 1423
rect 3032 1414 3080 1416
rect 3032 1406 3036 1414
rect 3046 1406 3052 1414
rect 3060 1406 3066 1414
rect 3076 1406 3080 1414
rect 3032 1404 3080 1406
rect 468 1397 1292 1403
rect 1396 1397 1436 1403
rect 1860 1397 1932 1403
rect 2820 1397 2931 1403
rect 788 1377 860 1383
rect 964 1377 1564 1383
rect 2925 1383 2931 1397
rect 3940 1397 4124 1403
rect 4404 1397 4819 1403
rect 4813 1384 4819 1397
rect 5028 1397 5596 1403
rect 6036 1397 6092 1403
rect 2925 1377 3372 1383
rect 3636 1377 3692 1383
rect 4116 1377 4316 1383
rect 4324 1377 4636 1383
rect 4740 1377 4796 1383
rect 4820 1377 5020 1383
rect 5028 1377 5180 1383
rect 5492 1377 5852 1383
rect 68 1357 188 1363
rect 228 1357 412 1363
rect 692 1357 812 1363
rect 820 1357 892 1363
rect 1396 1357 1580 1363
rect 1908 1357 2076 1363
rect 2084 1357 2540 1363
rect 3604 1357 3820 1363
rect 3956 1357 4140 1363
rect 4420 1357 4732 1363
rect 4740 1357 5036 1363
rect 5076 1357 5132 1363
rect 5156 1357 5452 1363
rect 5460 1357 5564 1363
rect 5572 1357 5580 1363
rect 5588 1357 5628 1363
rect 372 1337 460 1343
rect 468 1337 572 1343
rect 772 1337 1036 1343
rect 1284 1337 1340 1343
rect 1428 1337 1500 1343
rect 1972 1337 2012 1343
rect 2036 1337 2188 1343
rect 2308 1337 2444 1343
rect 2500 1337 2604 1343
rect 2628 1337 2876 1343
rect 2980 1337 3340 1343
rect 3636 1337 3644 1343
rect 3652 1337 3676 1343
rect 3780 1337 3916 1343
rect 4100 1337 4332 1343
rect 4340 1337 4380 1343
rect 4388 1337 4524 1343
rect 4532 1337 4764 1343
rect 4788 1337 4828 1343
rect 4852 1337 4892 1343
rect 5092 1337 5116 1343
rect 5124 1337 5388 1343
rect 5396 1337 5436 1343
rect 5444 1337 5884 1343
rect 5892 1337 6028 1343
rect 340 1317 444 1323
rect 484 1317 556 1323
rect 660 1317 748 1323
rect 980 1317 1004 1323
rect 1108 1317 1244 1323
rect 1252 1317 1356 1323
rect 1364 1317 1420 1323
rect 1428 1317 1452 1323
rect 1837 1323 1843 1336
rect 1572 1317 1843 1323
rect 1940 1317 2028 1323
rect 2068 1317 2092 1323
rect 2532 1317 2620 1323
rect 2852 1317 3068 1323
rect 3348 1317 3532 1323
rect 3540 1317 3660 1323
rect 4068 1317 4444 1323
rect 4452 1317 4492 1323
rect 4516 1317 4940 1323
rect 5108 1317 5404 1323
rect 5524 1317 5644 1323
rect 5684 1317 5836 1323
rect 5860 1317 5948 1323
rect 36 1297 140 1303
rect 148 1297 396 1303
rect 580 1297 1068 1303
rect 1140 1297 1244 1303
rect 1252 1297 1324 1303
rect 1348 1297 1468 1303
rect 1588 1297 2092 1303
rect 2580 1297 2764 1303
rect 4052 1297 4332 1303
rect 4340 1297 4524 1303
rect 4852 1297 4876 1303
rect 4932 1297 5292 1303
rect 5540 1297 5564 1303
rect 5620 1297 5676 1303
rect 5684 1297 5708 1303
rect 5716 1297 6076 1303
rect 436 1277 668 1283
rect 1316 1277 1388 1283
rect 1556 1277 1612 1283
rect 1620 1277 2380 1283
rect 3732 1277 3740 1283
rect 3748 1277 4108 1283
rect 4340 1277 4508 1283
rect 4669 1277 4748 1283
rect 548 1257 1212 1263
rect 1549 1263 1555 1276
rect 1364 1257 1555 1263
rect 4276 1257 4476 1263
rect 4669 1263 4675 1277
rect 4877 1283 4883 1296
rect 4877 1277 5196 1283
rect 5204 1277 5468 1283
rect 4484 1257 4675 1263
rect 4692 1257 5068 1263
rect 420 1237 428 1243
rect 468 1237 620 1243
rect 692 1237 1196 1243
rect 1204 1237 1260 1243
rect 1476 1237 1500 1243
rect 1540 1237 1580 1243
rect 3460 1237 3948 1243
rect 3956 1237 5100 1243
rect 5236 1237 5692 1243
rect 621 1223 627 1236
rect 621 1217 844 1223
rect 852 1217 876 1223
rect 996 1217 1004 1223
rect 1044 1217 1420 1223
rect 2292 1217 2652 1223
rect 3780 1217 4012 1223
rect 4068 1217 4284 1223
rect 4292 1217 4364 1223
rect 4820 1217 5036 1223
rect 5076 1217 5100 1223
rect 1496 1214 1544 1216
rect 1496 1206 1500 1214
rect 1510 1206 1516 1214
rect 1524 1206 1530 1214
rect 1540 1206 1544 1214
rect 1496 1204 1544 1206
rect 4568 1214 4616 1216
rect 4568 1206 4572 1214
rect 4582 1206 4588 1214
rect 4596 1206 4602 1214
rect 4612 1206 4616 1214
rect 4568 1204 4616 1206
rect 1716 1197 1804 1203
rect 2244 1197 2476 1203
rect 2580 1197 2668 1203
rect 3316 1197 3372 1203
rect 4260 1197 4460 1203
rect 4884 1197 5052 1203
rect 5844 1197 5964 1203
rect 1940 1177 2268 1183
rect 2500 1177 2620 1183
rect 2628 1177 2828 1183
rect 4228 1177 4428 1183
rect 4500 1177 4892 1183
rect 4900 1177 4956 1183
rect 4964 1177 5420 1183
rect 5860 1177 5900 1183
rect 5908 1177 6028 1183
rect 244 1157 508 1163
rect 884 1157 1132 1163
rect 1188 1157 1932 1163
rect 1940 1157 1980 1163
rect 2388 1157 2508 1163
rect 3668 1157 3692 1163
rect 4292 1157 4316 1163
rect 4452 1157 4508 1163
rect 5044 1157 5676 1163
rect 196 1137 268 1143
rect 276 1137 540 1143
rect 868 1137 956 1143
rect 1076 1137 1196 1143
rect 1204 1137 1356 1143
rect 2212 1137 2236 1143
rect 2276 1137 2604 1143
rect 2772 1137 2860 1143
rect 2868 1137 2908 1143
rect 4308 1137 4412 1143
rect 4468 1137 4716 1143
rect 5044 1137 5228 1143
rect 5348 1137 5500 1143
rect 308 1117 508 1123
rect 516 1117 588 1123
rect 596 1117 732 1123
rect 836 1117 940 1123
rect 948 1117 1212 1123
rect 1220 1117 1228 1123
rect 1332 1117 1420 1123
rect 1428 1117 1500 1123
rect 1508 1117 1644 1123
rect 2148 1117 2188 1123
rect 2516 1117 2572 1123
rect 4228 1117 4396 1123
rect 4452 1117 4460 1123
rect 4477 1117 5100 1123
rect 100 1097 220 1103
rect 548 1097 684 1103
rect 996 1097 1100 1103
rect 1428 1097 1532 1103
rect 1764 1097 1852 1103
rect 1860 1097 1980 1103
rect 2036 1097 2188 1103
rect 2196 1097 2220 1103
rect 2228 1097 2252 1103
rect 2340 1097 2364 1103
rect 2372 1097 2444 1103
rect 2612 1097 2844 1103
rect 3444 1097 3500 1103
rect 3876 1097 4156 1103
rect 4196 1097 4284 1103
rect 4477 1103 4483 1117
rect 5220 1117 5308 1123
rect 5316 1117 5372 1123
rect 5700 1117 6044 1123
rect 4420 1097 4483 1103
rect 4564 1097 4684 1103
rect 4772 1097 4812 1103
rect 4836 1097 4892 1103
rect 5044 1097 5148 1103
rect 5188 1097 5260 1103
rect 5300 1097 5484 1103
rect 5652 1097 5708 1103
rect 6004 1097 6060 1103
rect 6068 1097 6076 1103
rect 212 1077 268 1083
rect 356 1077 476 1083
rect 484 1077 492 1083
rect 980 1077 1020 1083
rect 1140 1077 1212 1083
rect 1284 1077 1388 1083
rect 1396 1077 1468 1083
rect 1812 1077 1868 1083
rect 1924 1077 2092 1083
rect 2100 1077 2172 1083
rect 2180 1077 2188 1083
rect 2196 1077 2268 1083
rect 2349 1077 2796 1083
rect 2349 1064 2355 1077
rect 2820 1077 2924 1083
rect 2964 1077 3020 1083
rect 3188 1077 3340 1083
rect 3540 1077 3644 1083
rect 3700 1077 3836 1083
rect 4084 1077 4108 1083
rect 4436 1077 4620 1083
rect 4724 1077 4780 1083
rect 4916 1077 4940 1083
rect 4948 1077 5004 1083
rect 5012 1077 5084 1083
rect 5092 1077 5116 1083
rect 5364 1077 5388 1083
rect 5396 1077 5628 1083
rect 5636 1077 5676 1083
rect 5908 1077 6044 1083
rect 260 1057 268 1063
rect 276 1057 604 1063
rect 1076 1057 1084 1063
rect 1252 1057 1564 1063
rect 1572 1057 1836 1063
rect 1844 1057 2108 1063
rect 2116 1057 2348 1063
rect 2372 1057 2412 1063
rect 2420 1057 2572 1063
rect 2900 1057 3084 1063
rect 3533 1063 3539 1076
rect 3092 1057 3539 1063
rect 3828 1057 4444 1063
rect 4484 1057 4492 1063
rect 4500 1057 4684 1063
rect 5076 1057 5212 1063
rect 5540 1057 5868 1063
rect 212 1037 396 1043
rect 452 1037 460 1043
rect 1460 1037 1580 1043
rect 1588 1037 1740 1043
rect 1748 1037 2044 1043
rect 2164 1037 2236 1043
rect 2436 1037 2476 1043
rect 4052 1037 4492 1043
rect 4532 1037 5107 1043
rect 404 1017 892 1023
rect 2557 1017 2716 1023
rect 2557 1004 2563 1017
rect 3636 1017 4012 1023
rect 4020 1017 4028 1023
rect 4116 1017 4348 1023
rect 4356 1017 4636 1023
rect 4644 1017 4860 1023
rect 4868 1017 5084 1023
rect 5101 1023 5107 1037
rect 5156 1037 5660 1043
rect 5716 1037 5724 1043
rect 5101 1017 5212 1023
rect 5220 1017 5564 1023
rect 3032 1014 3080 1016
rect 3032 1006 3036 1014
rect 3046 1006 3052 1014
rect 3060 1006 3066 1014
rect 3076 1006 3080 1014
rect 3032 1004 3080 1006
rect 1380 997 2556 1003
rect 2612 997 2668 1003
rect 3492 997 3820 1003
rect 3828 997 3868 1003
rect 4196 997 4412 1003
rect 4516 997 4828 1003
rect 4964 997 5420 1003
rect 324 977 428 983
rect 612 977 732 983
rect 740 977 796 983
rect 2276 977 2396 983
rect 3332 977 3340 983
rect 4292 977 4844 983
rect 4852 977 4972 983
rect 5076 977 5484 983
rect 5636 977 5692 983
rect 5700 977 5868 983
rect 5892 977 5964 983
rect 6036 977 6076 983
rect 244 957 364 963
rect 596 957 684 963
rect 724 957 796 963
rect 932 957 1052 963
rect 1060 957 1132 963
rect 1140 957 1324 963
rect 2276 957 2316 963
rect 2324 957 2444 963
rect 2452 957 2508 963
rect 3012 957 3308 963
rect 4212 957 4476 963
rect 4532 957 4636 963
rect 4676 957 4755 963
rect 228 937 252 943
rect 260 937 332 943
rect 356 937 636 943
rect 820 937 828 943
rect 1204 937 1276 943
rect 1796 937 1900 943
rect 2228 937 2412 943
rect 2420 937 2956 943
rect 2964 937 3164 943
rect 3524 937 3596 943
rect 4084 937 4140 943
rect 4340 937 4380 943
rect 4388 937 4476 943
rect 4564 937 4732 943
rect 4749 943 4755 957
rect 5108 957 5244 963
rect 5252 957 5276 963
rect 5348 957 5372 963
rect 5620 957 5916 963
rect 4749 937 5036 943
rect 5124 937 5404 943
rect 5412 937 5644 943
rect 292 917 364 923
rect 420 917 748 923
rect 852 917 876 923
rect 1012 917 1180 923
rect 1188 917 1292 923
rect 1300 917 1372 923
rect 2132 917 2156 923
rect 2180 917 2268 923
rect 2404 917 2700 923
rect 2804 917 2876 923
rect 3588 917 3660 923
rect 3668 917 3692 923
rect 4260 917 4300 923
rect 4308 917 4332 923
rect 4420 917 4428 923
rect 4500 917 4556 923
rect 4660 917 4748 923
rect 4804 917 4908 923
rect 4932 917 4988 923
rect 5188 917 5228 923
rect 5332 917 5564 923
rect 5716 917 6012 923
rect 148 897 284 903
rect 404 897 428 903
rect 676 897 764 903
rect 948 897 1068 903
rect 1076 897 1100 903
rect 1124 897 1212 903
rect 1220 897 1308 903
rect 1316 897 1420 903
rect 2052 897 2124 903
rect 2164 897 2348 903
rect 4260 897 4444 903
rect 4500 897 4572 903
rect 4772 897 5196 903
rect 5204 897 5340 903
rect 5348 897 5452 903
rect 5684 897 5740 903
rect 397 883 403 896
rect 20 877 403 883
rect 660 877 684 883
rect 765 883 771 896
rect 765 877 1036 883
rect 1092 877 1148 883
rect 1252 877 1324 883
rect 1412 877 1468 883
rect 4164 877 4284 883
rect 5140 877 5244 883
rect 5252 877 5692 883
rect 740 857 844 863
rect 1325 863 1331 876
rect 1325 857 1436 863
rect 1444 857 1756 863
rect 4596 857 5612 863
rect 628 837 908 843
rect 3988 837 4060 843
rect 4068 837 4252 843
rect 4308 837 4780 843
rect 388 817 524 823
rect 788 817 988 823
rect 1236 817 1388 823
rect 1716 817 1868 823
rect 3796 817 3980 823
rect 4660 817 5004 823
rect 5012 817 5228 823
rect 5636 817 6060 823
rect 1496 814 1544 816
rect 1496 806 1500 814
rect 1510 806 1516 814
rect 1524 806 1530 814
rect 1540 806 1544 814
rect 1496 804 1544 806
rect 4568 814 4616 816
rect 4568 806 4572 814
rect 4582 806 4588 814
rect 4596 806 4602 814
rect 4612 806 4616 814
rect 4568 804 4616 806
rect 1620 797 1900 803
rect 2084 797 2460 803
rect 2468 797 2844 803
rect 3268 797 3372 803
rect 3380 797 3596 803
rect 3604 797 3676 803
rect 4244 797 4460 803
rect 4932 797 5116 803
rect 1588 777 1820 783
rect 3620 777 3644 783
rect 3652 777 4291 783
rect 308 757 412 763
rect 1316 757 1500 763
rect 3188 757 4268 763
rect 4285 763 4291 777
rect 4372 777 4380 783
rect 4388 777 5068 783
rect 5924 777 5948 783
rect 4285 757 4556 763
rect 4580 757 4915 763
rect 84 737 108 743
rect 292 737 380 743
rect 388 737 620 743
rect 644 737 780 743
rect 804 737 1196 743
rect 1460 737 1484 743
rect 1572 737 1884 743
rect 1940 737 1996 743
rect 2532 737 2588 743
rect 3044 737 3548 743
rect 3876 737 3900 743
rect 3956 737 4108 743
rect 4125 737 4444 743
rect 116 717 172 723
rect 276 717 316 723
rect 372 717 492 723
rect 708 717 716 723
rect 836 717 1212 723
rect 1460 717 1964 723
rect 2036 717 2380 723
rect 3716 717 3740 723
rect 3748 717 3820 723
rect 3828 717 3948 723
rect 3956 717 4012 723
rect 4125 723 4131 737
rect 4468 737 4636 743
rect 4724 737 4892 743
rect 4909 743 4915 757
rect 4996 757 5148 763
rect 5444 757 5468 763
rect 5716 757 6028 763
rect 4909 737 5356 743
rect 5428 737 5436 743
rect 5588 737 5724 743
rect 5764 737 5836 743
rect 4020 717 4131 723
rect 4148 717 4172 723
rect 4212 717 4252 723
rect 4452 717 4460 723
rect 4468 717 4524 723
rect 4708 717 4844 723
rect 5060 717 5260 723
rect 5620 717 5644 723
rect 5652 717 5964 723
rect -19 697 12 703
rect 52 697 60 703
rect 260 697 332 703
rect 420 697 460 703
rect 468 697 524 703
rect 532 697 652 703
rect 660 697 716 703
rect 724 697 908 703
rect 996 697 1340 703
rect 1476 697 1628 703
rect 1828 697 1916 703
rect 2020 697 2076 703
rect 3396 697 3580 703
rect 3588 697 3660 703
rect 3668 697 3756 703
rect 4244 697 4268 703
rect 4404 697 4748 703
rect 4804 697 4924 703
rect 5028 697 5052 703
rect 5092 697 5356 703
rect 5556 697 5612 703
rect 5716 697 5756 703
rect 228 677 460 683
rect 756 677 924 683
rect 1012 677 1180 683
rect 1412 677 1644 683
rect 1652 677 1772 683
rect 1876 677 1932 683
rect 2020 677 2172 683
rect 2580 677 2780 683
rect 2900 677 2924 683
rect 3444 677 3532 683
rect 3572 677 3612 683
rect 4084 677 4156 683
rect 4164 677 4220 683
rect 4260 677 4284 683
rect 4484 677 4828 683
rect 4900 677 5004 683
rect 5044 677 5084 683
rect 5172 677 5404 683
rect 5444 677 5484 683
rect 5876 677 5980 683
rect 6020 677 6060 683
rect 180 657 332 663
rect 372 657 428 663
rect 436 657 636 663
rect 644 657 700 663
rect 804 657 860 663
rect 932 657 1020 663
rect 1028 657 1084 663
rect 1972 657 2204 663
rect 2676 657 2748 663
rect 2756 657 3196 663
rect 3236 657 3628 663
rect 3684 657 3724 663
rect 4132 657 4236 663
rect 4244 657 4540 663
rect 4548 657 4668 663
rect 5140 657 5452 663
rect 36 637 140 643
rect 148 637 348 643
rect 452 637 460 643
rect 692 637 988 643
rect 2852 637 3100 643
rect 3396 637 3708 643
rect 3716 637 3932 643
rect 3940 637 4092 643
rect 4100 637 4172 643
rect 4420 637 5132 643
rect 5604 637 5804 643
rect 100 617 140 623
rect 164 617 364 623
rect 756 617 892 623
rect 1748 617 2524 623
rect 3716 617 3772 623
rect 4004 617 4012 623
rect 4196 617 4732 623
rect 4740 617 4844 623
rect 5316 617 5564 623
rect 3032 614 3080 616
rect 3032 606 3036 614
rect 3046 606 3052 614
rect 3060 606 3066 614
rect 3076 606 3080 614
rect 3032 604 3080 606
rect 132 597 172 603
rect 244 597 636 603
rect 644 597 844 603
rect 1636 597 1788 603
rect 3540 597 3900 603
rect 4052 597 4204 603
rect 4228 597 4348 603
rect 4500 597 4796 603
rect 5284 597 5420 603
rect 5428 597 5772 603
rect 5988 597 6028 603
rect 932 577 1052 583
rect 2068 577 2124 583
rect 2228 577 2460 583
rect 3124 577 3196 583
rect 3268 577 3420 583
rect 3428 577 3548 583
rect 3556 577 3628 583
rect 3684 577 3884 583
rect 4356 577 4396 583
rect 5172 577 5388 583
rect 5684 577 5788 583
rect 180 557 492 563
rect 564 557 604 563
rect 612 557 1116 563
rect 1204 557 1404 563
rect 1412 557 1452 563
rect 1476 557 1548 563
rect 1940 557 2204 563
rect 2324 557 2364 563
rect 2420 557 2748 563
rect 3620 557 3692 563
rect 3828 557 3852 563
rect 3892 557 4092 563
rect 4276 557 4364 563
rect 4372 557 4444 563
rect 4468 557 4524 563
rect 4564 557 4652 563
rect 4724 557 4764 563
rect 4772 557 4796 563
rect 5284 557 5356 563
rect 5364 557 5436 563
rect 468 537 748 543
rect 772 537 828 543
rect 868 537 956 543
rect 1124 537 1596 543
rect 1604 537 1660 543
rect 1700 537 1788 543
rect 1796 537 1964 543
rect 2196 537 2236 543
rect 2244 537 2284 543
rect 2292 537 2380 543
rect 2788 537 2892 543
rect 3092 537 3468 543
rect 3572 537 3596 543
rect 3604 537 3788 543
rect 3860 537 3948 543
rect 4148 537 4396 543
rect 4420 537 4508 543
rect 4516 537 4940 543
rect 4948 537 5164 543
rect 5172 537 5308 543
rect 5332 537 5548 543
rect 724 517 940 523
rect 1364 517 1468 523
rect 2052 517 2460 523
rect 2708 517 2796 523
rect 3492 517 3612 523
rect 3620 517 3644 523
rect 3668 517 3756 523
rect 4244 517 4316 523
rect 4404 517 4492 523
rect 4660 517 4732 523
rect 4980 517 5052 523
rect 5060 517 5292 523
rect 5300 517 5548 523
rect 420 497 716 503
rect 884 497 1244 503
rect 1380 497 1628 503
rect 2372 497 2556 503
rect 2836 497 2940 503
rect 3284 497 3452 503
rect 3460 497 3580 503
rect 3636 497 4220 503
rect 4324 497 4348 503
rect 4404 497 4428 503
rect 4452 497 4476 503
rect 4756 497 5116 503
rect 5252 497 5404 503
rect 5876 497 5948 503
rect 1460 477 1484 483
rect 1492 477 1596 483
rect 4452 477 4636 483
rect 5348 477 5372 483
rect 5412 477 5516 483
rect 884 457 908 463
rect 1348 457 1532 463
rect 3412 457 3468 463
rect 3476 457 3548 463
rect 5364 457 5756 463
rect 5764 457 5804 463
rect 2900 437 3132 443
rect 4564 437 4748 443
rect 5268 437 5500 443
rect 6052 417 6092 423
rect 1496 414 1544 416
rect 1496 406 1500 414
rect 1510 406 1516 414
rect 1524 406 1530 414
rect 1540 406 1544 414
rect 1496 404 1544 406
rect 4568 414 4616 416
rect 4568 406 4572 414
rect 4582 406 4588 414
rect 4596 406 4602 414
rect 4612 406 4616 414
rect 4568 404 4616 406
rect 388 397 412 403
rect 2468 397 2796 403
rect 5028 397 5036 403
rect 5092 397 5244 403
rect 5252 397 5532 403
rect 180 377 220 383
rect 1412 377 1452 383
rect 5396 377 5740 383
rect 644 357 892 363
rect 1140 357 1212 363
rect 1220 357 1308 363
rect 4084 357 5356 363
rect 5524 357 5708 363
rect 628 337 828 343
rect 836 337 1148 343
rect 1156 337 1276 343
rect 1284 337 1340 343
rect 4308 337 4428 343
rect 5092 337 5164 343
rect 5444 337 5532 343
rect 564 317 700 323
rect 772 317 844 323
rect 900 317 924 323
rect 1028 317 1164 323
rect 1300 317 1340 323
rect 1684 317 1802 323
rect 1810 317 2220 323
rect 3284 317 3388 323
rect 4276 317 4364 323
rect 4772 317 4844 323
rect 4925 317 5196 323
rect 4925 304 4931 317
rect 5204 317 5324 323
rect 5476 317 5516 323
rect 5572 317 5628 323
rect 6132 317 6163 323
rect -19 297 12 303
rect 68 297 444 303
rect 612 297 652 303
rect 852 297 908 303
rect 932 297 1244 303
rect 1252 297 1372 303
rect 1540 297 1564 303
rect 2180 297 2204 303
rect 2580 297 2732 303
rect 2852 297 3148 303
rect 4244 297 4268 303
rect 4292 297 4316 303
rect 4324 297 4444 303
rect 4660 297 4812 303
rect 4900 297 4924 303
rect 4980 297 5132 303
rect 5220 297 5420 303
rect 5492 297 6060 303
rect 196 277 396 283
rect 900 277 940 283
rect 948 277 1260 283
rect 2004 277 2060 283
rect 2228 277 2284 283
rect 2836 277 2876 283
rect 3044 277 3148 283
rect 3156 277 3180 283
rect 3460 277 3484 283
rect 3796 277 3820 283
rect 4468 277 4700 283
rect 4708 277 5020 283
rect 5028 277 5228 283
rect 5236 277 5260 283
rect 5396 277 5436 283
rect 5524 277 5596 283
rect 5620 277 5900 283
rect 6068 277 6163 283
rect 1300 257 1468 263
rect 3364 257 3468 263
rect 3540 257 3596 263
rect 3604 257 3612 263
rect 3620 257 3628 263
rect 4580 257 4780 263
rect 4788 257 4828 263
rect 4836 257 5100 263
rect 5108 257 5244 263
rect 5588 257 5628 263
rect 5876 257 5900 263
rect 868 237 908 243
rect 1476 237 1628 243
rect 4532 237 4892 243
rect 4900 237 5212 243
rect 5220 237 5388 243
rect 5396 237 5452 243
rect 308 217 1548 223
rect 2324 217 2524 223
rect 3764 217 3804 223
rect 4244 217 4332 223
rect 4340 217 4636 223
rect 3032 214 3080 216
rect 3032 206 3036 214
rect 3046 206 3052 214
rect 3060 206 3066 214
rect 3076 206 3080 214
rect 3032 204 3080 206
rect 180 197 220 203
rect 228 197 540 203
rect 772 197 1004 203
rect 1268 197 1308 203
rect 1316 197 1388 203
rect 1396 197 1644 203
rect 1844 197 1852 203
rect 1860 197 1884 203
rect 2612 197 2748 203
rect 3284 197 3340 203
rect 4340 197 4476 203
rect 4484 197 4652 203
rect 372 177 508 183
rect 516 177 732 183
rect 1108 177 1340 183
rect 2372 177 2492 183
rect 2500 177 2588 183
rect 2596 177 2860 183
rect 2868 177 3116 183
rect 3124 177 3308 183
rect 3316 177 3948 183
rect 3972 177 4044 183
rect 5604 177 5644 183
rect 5652 177 5900 183
rect 340 157 412 163
rect 788 157 828 163
rect 980 157 1340 163
rect 1636 157 1964 163
rect 3508 157 3596 163
rect 3812 157 4092 163
rect 5540 157 5932 163
rect 148 137 428 143
rect 836 137 1020 143
rect 1668 137 1724 143
rect 1940 137 2172 143
rect 2244 137 2332 143
rect 3604 137 3772 143
rect 4116 137 4252 143
rect 4468 137 4524 143
rect 4564 137 4668 143
rect 4788 137 4844 143
rect 4900 137 4940 143
rect 5220 137 5308 143
rect 5316 137 5436 143
rect 5460 137 5660 143
rect 52 117 348 123
rect 356 117 380 123
rect 532 117 780 123
rect 788 117 972 123
rect 1012 117 1164 123
rect 1236 117 1324 123
rect 1780 117 1836 123
rect 2052 117 2236 123
rect 2980 117 3180 123
rect 4308 117 4748 123
rect 4820 117 5180 123
rect 5188 117 5228 123
rect 5300 117 5548 123
rect 5684 117 5836 123
rect 4500 97 4524 103
rect 4804 97 4892 103
rect 4900 97 5036 103
rect 5044 97 5132 103
rect 5188 97 5260 103
rect 5524 97 5708 103
rect 6116 97 6163 103
rect 4228 77 4252 83
rect 4260 77 4348 83
rect 4884 77 5004 83
rect 5668 17 5676 23
rect 1496 14 1544 16
rect 1496 6 1500 14
rect 1510 6 1516 14
rect 1524 6 1530 14
rect 1540 6 1544 14
rect 1496 4 1544 6
rect 4568 14 4616 16
rect 4568 6 4572 14
rect 4582 6 4588 14
rect 4596 6 4602 14
rect 4612 6 4616 14
rect 4568 4 4616 6
<< m4contact >>
rect 1500 5606 1502 5614
rect 1502 5606 1508 5614
rect 1516 5606 1524 5614
rect 1532 5606 1538 5614
rect 1538 5606 1540 5614
rect 4572 5606 4574 5614
rect 4574 5606 4580 5614
rect 4588 5606 4596 5614
rect 4604 5606 4610 5614
rect 4610 5606 4612 5614
rect 6092 5596 6100 5604
rect 1228 5496 1236 5504
rect 332 5456 340 5464
rect 2508 5436 2516 5444
rect 5580 5436 5588 5444
rect 1228 5416 1236 5424
rect 3036 5406 3038 5414
rect 3038 5406 3044 5414
rect 3052 5406 3060 5414
rect 3068 5406 3074 5414
rect 3074 5406 3076 5414
rect 3724 5376 3732 5384
rect 460 5356 468 5364
rect 2444 5356 2452 5364
rect 5260 5356 5268 5364
rect 972 5336 980 5344
rect 5612 5336 5620 5344
rect 524 5316 532 5324
rect 364 5296 372 5304
rect 5196 5316 5204 5324
rect 5900 5296 5908 5304
rect 5996 5256 6004 5264
rect 652 5236 660 5244
rect 4428 5216 4436 5224
rect 1500 5206 1502 5214
rect 1502 5206 1508 5214
rect 1516 5206 1524 5214
rect 1532 5206 1538 5214
rect 1538 5206 1540 5214
rect 4572 5206 4574 5214
rect 4574 5206 4580 5214
rect 4588 5206 4596 5214
rect 4604 5206 4610 5214
rect 4610 5206 4612 5214
rect 4108 5176 4116 5184
rect 5420 5176 5428 5184
rect 460 5136 468 5144
rect 3724 5136 3732 5144
rect 3980 5136 3988 5144
rect 4396 5116 4404 5124
rect 4652 5116 4660 5124
rect 460 5096 468 5104
rect 4140 5096 4148 5104
rect 1900 5076 1908 5084
rect 4876 5076 4884 5084
rect 5260 5076 5268 5084
rect 2956 5036 2964 5044
rect 4876 5036 4884 5044
rect 1708 5016 1716 5024
rect 3036 5006 3038 5014
rect 3038 5006 3044 5014
rect 3052 5006 3060 5014
rect 3068 5006 3074 5014
rect 3074 5006 3076 5014
rect 3916 4996 3924 5004
rect 2252 4976 2260 4984
rect 3308 4976 3316 4984
rect 908 4956 916 4964
rect 2444 4956 2452 4964
rect 5036 4956 5044 4964
rect 972 4936 980 4944
rect 2764 4936 2772 4944
rect 5580 4936 5588 4944
rect 876 4916 884 4924
rect 2828 4916 2836 4924
rect 652 4896 660 4904
rect 1036 4896 1044 4904
rect 2956 4896 2964 4904
rect 4268 4896 4276 4904
rect 1964 4856 1972 4864
rect 4108 4856 4116 4864
rect 4396 4856 4404 4864
rect 172 4836 180 4844
rect 5196 4836 5204 4844
rect 6028 4836 6036 4844
rect 4492 4816 4500 4824
rect 4652 4816 4660 4824
rect 1500 4806 1502 4814
rect 1502 4806 1508 4814
rect 1516 4806 1524 4814
rect 1532 4806 1538 4814
rect 1538 4806 1540 4814
rect 4572 4806 4574 4814
rect 4574 4806 4580 4814
rect 4588 4806 4596 4814
rect 4604 4806 4610 4814
rect 4610 4806 4612 4814
rect 1356 4796 1364 4804
rect 3980 4796 3988 4804
rect 3820 4756 3828 4764
rect 3916 4756 3924 4764
rect 4492 4756 4500 4764
rect 5452 4756 5460 4764
rect 940 4716 948 4724
rect 3308 4716 3316 4724
rect 4684 4716 4692 4724
rect 5036 4716 5044 4724
rect 1356 4696 1364 4704
rect 2412 4696 2420 4704
rect 940 4676 948 4684
rect 1708 4676 1716 4684
rect 4268 4676 4276 4684
rect 4940 4676 4948 4684
rect 5196 4656 5204 4664
rect 3404 4636 3412 4644
rect 4140 4636 4148 4644
rect 3980 4616 3988 4624
rect 3036 4606 3038 4614
rect 3038 4606 3044 4614
rect 3052 4606 3060 4614
rect 3068 4606 3074 4614
rect 3074 4606 3076 4614
rect 1772 4596 1780 4604
rect 5164 4596 5172 4604
rect 5836 4596 5844 4604
rect 460 4576 468 4584
rect 5068 4556 5076 4564
rect 428 4536 436 4544
rect 524 4536 532 4544
rect 1036 4516 1044 4524
rect 4684 4536 4692 4544
rect 4748 4536 4756 4544
rect 5164 4516 5172 4524
rect 5900 4516 5908 4524
rect 5932 4516 5940 4524
rect 1900 4496 1908 4504
rect 2764 4496 2772 4504
rect 1324 4456 1332 4464
rect 2988 4456 2996 4464
rect 1612 4436 1620 4444
rect 876 4416 884 4424
rect 1356 4416 1364 4424
rect 2508 4416 2516 4424
rect 5228 4416 5236 4424
rect 5740 4416 5748 4424
rect 1500 4406 1502 4414
rect 1502 4406 1508 4414
rect 1516 4406 1524 4414
rect 1532 4406 1538 4414
rect 1538 4406 1540 4414
rect 4572 4406 4574 4414
rect 4574 4406 4580 4414
rect 4588 4406 4596 4414
rect 4604 4406 4610 4414
rect 4610 4406 4612 4414
rect 2956 4396 2964 4404
rect 1676 4376 1684 4384
rect 2668 4376 2676 4384
rect 5068 4376 5076 4384
rect 5356 4376 5364 4384
rect 172 4356 180 4364
rect 2220 4316 2228 4324
rect 4940 4316 4948 4324
rect 588 4296 596 4304
rect 1964 4296 1972 4304
rect 140 4276 148 4284
rect 364 4276 372 4284
rect 2028 4276 2036 4284
rect 3980 4276 3988 4284
rect 1356 4236 1364 4244
rect 5612 4236 5620 4244
rect 1292 4216 1300 4224
rect 2316 4216 2324 4224
rect 3372 4216 3380 4224
rect 3036 4206 3038 4214
rect 3038 4206 3044 4214
rect 3052 4206 3060 4214
rect 3068 4206 3074 4214
rect 3074 4206 3076 4214
rect 1900 4196 1908 4204
rect 4204 4196 4212 4204
rect 1164 4156 1172 4164
rect 5100 4156 5108 4164
rect 5900 4136 5908 4144
rect 332 4116 340 4124
rect 1612 4116 1620 4124
rect 1772 4116 1780 4124
rect 5100 4116 5108 4124
rect 1676 4096 1684 4104
rect 3820 4096 3828 4104
rect 3436 4076 3444 4084
rect 4748 4056 4756 4064
rect 4908 4036 4916 4044
rect 2028 4016 2036 4024
rect 1500 4006 1502 4014
rect 1502 4006 1508 4014
rect 1516 4006 1524 4014
rect 1532 4006 1538 4014
rect 1538 4006 1540 4014
rect 4572 4006 4574 4014
rect 4574 4006 4580 4014
rect 4588 4006 4596 4014
rect 4604 4006 4610 4014
rect 4610 4006 4612 4014
rect 460 3976 468 3984
rect 5996 3996 6004 4004
rect 2924 3976 2932 3984
rect 3404 3976 3412 3984
rect 908 3916 916 3924
rect 588 3896 596 3904
rect 2252 3916 2260 3924
rect 2668 3896 2676 3904
rect 428 3876 436 3884
rect 5740 3876 5748 3884
rect 460 3836 468 3844
rect 1068 3816 1076 3824
rect 2828 3816 2836 3824
rect 3036 3806 3038 3814
rect 3038 3806 3044 3814
rect 3052 3806 3060 3814
rect 3068 3806 3074 3814
rect 3074 3806 3076 3814
rect 1292 3776 1300 3784
rect 4748 3796 4756 3804
rect 1068 3756 1076 3764
rect 1324 3756 1332 3764
rect 1900 3756 1908 3764
rect 4428 3756 4436 3764
rect 908 3736 916 3744
rect 2764 3736 2772 3744
rect 4204 3716 4212 3724
rect 5900 3716 5908 3724
rect 2380 3696 2388 3704
rect 3788 3696 3796 3704
rect 2444 3656 2452 3664
rect 2220 3616 2228 3624
rect 5388 3616 5396 3624
rect 1500 3606 1502 3614
rect 1502 3606 1508 3614
rect 1516 3606 1524 3614
rect 1532 3606 1538 3614
rect 1538 3606 1540 3614
rect 4572 3606 4574 3614
rect 4574 3606 4580 3614
rect 4588 3606 4596 3614
rect 4604 3606 4610 3614
rect 4610 3606 4612 3614
rect 2412 3596 2420 3604
rect 1292 3576 1300 3584
rect 5420 3576 5428 3584
rect 940 3556 948 3564
rect 4140 3536 4148 3544
rect 4908 3536 4916 3544
rect 1164 3516 1172 3524
rect 2284 3496 2292 3504
rect 3468 3496 3476 3504
rect 4044 3496 4052 3504
rect 3372 3476 3380 3484
rect 5292 3456 5300 3464
rect 1964 3436 1972 3444
rect 2316 3416 2324 3424
rect 4108 3416 4116 3424
rect 3036 3406 3038 3414
rect 3038 3406 3044 3414
rect 3052 3406 3060 3414
rect 3068 3406 3074 3414
rect 3074 3406 3076 3414
rect 2700 3396 2708 3404
rect 2924 3396 2932 3404
rect 3436 3396 3444 3404
rect 5388 3336 5396 3344
rect 6092 3336 6100 3344
rect 2284 3296 2292 3304
rect 2988 3296 2996 3304
rect 4940 3316 4948 3324
rect 5292 3316 5300 3324
rect 5548 3316 5556 3324
rect 4492 3296 4500 3304
rect 2316 3276 2324 3284
rect 2956 3276 2964 3284
rect 3756 3256 3764 3264
rect 3788 3256 3796 3264
rect 1100 3216 1108 3224
rect 3244 3216 3252 3224
rect 5100 3216 5108 3224
rect 5196 3216 5204 3224
rect 5356 3216 5364 3224
rect 5580 3216 5588 3224
rect 1500 3206 1502 3214
rect 1502 3206 1508 3214
rect 1516 3206 1524 3214
rect 1532 3206 1538 3214
rect 1538 3206 1540 3214
rect 140 3196 148 3204
rect 1388 3196 1396 3204
rect 4572 3206 4574 3214
rect 4574 3206 4580 3214
rect 4588 3206 4596 3214
rect 4604 3206 4610 3214
rect 4610 3206 4612 3214
rect 4652 3196 4660 3204
rect 1292 3176 1300 3184
rect 2060 3176 2068 3184
rect 3468 3176 3476 3184
rect 2380 3156 2388 3164
rect 3116 3136 3124 3144
rect 4652 3136 4660 3144
rect 5036 3136 5044 3144
rect 5836 3136 5844 3144
rect 5868 3136 5876 3144
rect 1964 3096 1972 3104
rect 2732 3116 2740 3124
rect 2924 3116 2932 3124
rect 4108 3116 4116 3124
rect 5068 3116 5076 3124
rect 5228 3116 5236 3124
rect 3756 3096 3764 3104
rect 4044 3096 4052 3104
rect 4684 3096 4692 3104
rect 5004 3096 5012 3104
rect 2700 3076 2708 3084
rect 3788 3076 3796 3084
rect 3916 3076 3924 3084
rect 4492 3076 4500 3084
rect 5036 3076 5044 3084
rect 3532 3056 3540 3064
rect 4172 3056 4180 3064
rect 4940 3056 4948 3064
rect 5388 3056 5396 3064
rect 3148 3036 3156 3044
rect 4044 3036 4052 3044
rect 2956 3016 2964 3024
rect 4012 3016 4020 3024
rect 5004 3016 5012 3024
rect 5420 3016 5428 3024
rect 3036 3006 3038 3014
rect 3038 3006 3044 3014
rect 3052 3006 3060 3014
rect 3068 3006 3074 3014
rect 3074 3006 3076 3014
rect 3116 2976 3124 2984
rect 5068 2976 5076 2984
rect 3148 2956 3156 2964
rect 4172 2956 4180 2964
rect 3916 2936 3924 2944
rect 4844 2936 4852 2944
rect 5196 2956 5204 2964
rect 5068 2936 5076 2944
rect 5100 2936 5108 2944
rect 5804 2936 5812 2944
rect 5932 2936 5940 2944
rect 5548 2916 5556 2924
rect 3948 2896 3956 2904
rect 3660 2876 3668 2884
rect 3820 2876 3828 2884
rect 4300 2876 4308 2884
rect 3628 2856 3636 2864
rect 4044 2856 4052 2864
rect 2060 2836 2068 2844
rect 2444 2836 2452 2844
rect 2508 2836 2516 2844
rect 2924 2836 2932 2844
rect 3276 2836 3284 2844
rect 5132 2836 5140 2844
rect 2284 2816 2292 2824
rect 3212 2816 3220 2824
rect 3244 2816 3252 2824
rect 4780 2816 4788 2824
rect 1500 2806 1502 2814
rect 1502 2806 1508 2814
rect 1516 2806 1524 2814
rect 1532 2806 1538 2814
rect 1538 2806 1540 2814
rect 4572 2806 4574 2814
rect 4574 2806 4580 2814
rect 4588 2806 4596 2814
rect 4604 2806 4610 2814
rect 4610 2806 4612 2814
rect 1996 2796 2004 2804
rect 2732 2796 2740 2804
rect 2316 2776 2324 2784
rect 2508 2776 2516 2784
rect 4332 2796 4340 2804
rect 4012 2776 4020 2784
rect 1964 2756 1972 2764
rect 3596 2756 3604 2764
rect 3820 2756 3828 2764
rect 5196 2756 5204 2764
rect 5292 2756 5300 2764
rect 1100 2736 1108 2744
rect 5580 2736 5588 2744
rect 3660 2716 3668 2724
rect 5196 2696 5204 2704
rect 1388 2676 1396 2684
rect 2860 2676 2868 2684
rect 2988 2676 2996 2684
rect 3276 2676 3284 2684
rect 3948 2676 3956 2684
rect 3148 2656 3156 2664
rect 3244 2656 3252 2664
rect 4204 2656 4212 2664
rect 5100 2676 5108 2684
rect 5420 2676 5428 2684
rect 6028 2676 6036 2684
rect 5260 2656 5268 2664
rect 5484 2656 5492 2664
rect 364 2636 372 2644
rect 3596 2636 3604 2644
rect 3724 2636 3732 2644
rect 3788 2636 3796 2644
rect 4684 2636 4692 2644
rect 4748 2636 4756 2644
rect 4876 2636 4884 2644
rect 5036 2636 5044 2644
rect 5068 2636 5076 2644
rect 3036 2606 3038 2614
rect 3038 2606 3044 2614
rect 3052 2606 3060 2614
rect 3068 2606 3074 2614
rect 3074 2606 3076 2614
rect 1996 2596 2004 2604
rect 3500 2596 3508 2604
rect 3628 2596 3636 2604
rect 4172 2616 4180 2624
rect 4332 2616 4340 2624
rect 4780 2596 4788 2604
rect 2604 2556 2612 2564
rect 4300 2556 4308 2564
rect 2732 2536 2740 2544
rect 2956 2536 2964 2544
rect 3660 2536 3668 2544
rect 5292 2556 5300 2564
rect 4876 2536 4884 2544
rect 5260 2536 5268 2544
rect 5324 2536 5332 2544
rect 3212 2516 3220 2524
rect 5100 2516 5108 2524
rect 2860 2496 2868 2504
rect 4204 2496 4212 2504
rect 4844 2496 4852 2504
rect 3468 2476 3476 2484
rect 3148 2456 3156 2464
rect 2412 2436 2420 2444
rect 3244 2436 3252 2444
rect 4236 2436 4244 2444
rect 4652 2436 4660 2444
rect 5036 2436 5044 2444
rect 5388 2436 5396 2444
rect 5516 2436 5524 2444
rect 3532 2416 3540 2424
rect 4172 2416 4180 2424
rect 4684 2416 4692 2424
rect 4716 2416 4724 2424
rect 1500 2406 1502 2414
rect 1502 2406 1508 2414
rect 1516 2406 1524 2414
rect 1532 2406 1538 2414
rect 1538 2406 1540 2414
rect 4572 2406 4574 2414
rect 4574 2406 4580 2414
rect 4588 2406 4596 2414
rect 4604 2406 4610 2414
rect 4610 2406 4612 2414
rect 3468 2376 3476 2384
rect 4236 2396 4244 2404
rect 5740 2376 5748 2384
rect 5868 2376 5876 2384
rect 4044 2356 4052 2364
rect 4076 2356 4084 2364
rect 5324 2356 5332 2364
rect 940 2316 948 2324
rect 2732 2316 2740 2324
rect 2988 2316 2996 2324
rect 3148 2316 3156 2324
rect 4716 2316 4724 2324
rect 5324 2316 5332 2324
rect 5484 2316 5492 2324
rect 5868 2316 5876 2324
rect 3212 2296 3220 2304
rect 3404 2296 3412 2304
rect 3596 2296 3604 2304
rect 4140 2296 4148 2304
rect 6028 2296 6036 2304
rect 2316 2276 2324 2284
rect 3820 2276 3828 2284
rect 4684 2276 4692 2284
rect 3660 2256 3668 2264
rect 3500 2236 3508 2244
rect 4652 2236 4660 2244
rect 556 2216 564 2224
rect 3116 2216 3124 2224
rect 3820 2216 3828 2224
rect 3036 2206 3038 2214
rect 3038 2206 3044 2214
rect 3052 2206 3060 2214
rect 3068 2206 3074 2214
rect 3074 2206 3076 2214
rect 2604 2156 2612 2164
rect 2220 2136 2228 2144
rect 44 2116 52 2124
rect 2316 2116 2324 2124
rect 3820 2096 3828 2104
rect 5132 2096 5140 2104
rect 5644 2096 5652 2104
rect 2316 2036 2324 2044
rect 3212 2036 3220 2044
rect 3468 2036 3476 2044
rect 5676 2036 5684 2044
rect 3116 2016 3124 2024
rect 1500 2006 1502 2014
rect 1502 2006 1508 2014
rect 1516 2006 1524 2014
rect 1532 2006 1538 2014
rect 1538 2006 1540 2014
rect 4572 2006 4574 2014
rect 4574 2006 4580 2014
rect 4588 2006 4596 2014
rect 4604 2006 4610 2014
rect 4610 2006 4612 2014
rect 844 1976 852 1984
rect 4108 1976 4116 1984
rect 5900 1976 5908 1984
rect 3180 1956 3188 1964
rect 5068 1956 5076 1964
rect 3436 1936 3444 1944
rect 4812 1936 4820 1944
rect 5100 1916 5108 1924
rect 140 1896 148 1904
rect 1452 1896 1460 1904
rect 2060 1896 2068 1904
rect 2092 1896 2100 1904
rect 2860 1896 2868 1904
rect 3116 1896 3124 1904
rect 3468 1896 3476 1904
rect 4684 1896 4692 1904
rect 6092 1876 6100 1884
rect 5740 1856 5748 1864
rect 364 1836 372 1844
rect 4076 1836 4084 1844
rect 5228 1836 5236 1844
rect 3436 1816 3444 1824
rect 5196 1816 5204 1824
rect 5804 1816 5812 1824
rect 3036 1806 3038 1814
rect 3038 1806 3044 1814
rect 3052 1806 3060 1814
rect 3068 1806 3074 1814
rect 3074 1806 3076 1814
rect 1228 1796 1236 1804
rect 2860 1796 2868 1804
rect 2220 1776 2228 1784
rect 2092 1756 2100 1764
rect 2412 1756 2420 1764
rect 3180 1756 3188 1764
rect 5804 1756 5812 1764
rect 812 1716 820 1724
rect 5036 1716 5044 1724
rect 2156 1696 2164 1704
rect 3404 1696 3412 1704
rect 3820 1696 3828 1704
rect 1580 1676 1588 1684
rect 4844 1676 4852 1684
rect 5644 1676 5652 1684
rect 1420 1636 1428 1644
rect 2060 1636 2068 1644
rect 1500 1606 1502 1614
rect 1502 1606 1508 1614
rect 1516 1606 1524 1614
rect 1532 1606 1538 1614
rect 1538 1606 1540 1614
rect 4572 1606 4574 1614
rect 4574 1606 4580 1614
rect 4588 1606 4596 1614
rect 4604 1606 4610 1614
rect 4610 1606 4612 1614
rect 428 1596 436 1604
rect 5964 1596 5972 1604
rect 4844 1576 4852 1584
rect 1356 1556 1364 1564
rect 1612 1556 1620 1564
rect 364 1516 372 1524
rect 3116 1496 3124 1504
rect 4492 1516 4500 1524
rect 4812 1496 4820 1504
rect 5868 1476 5876 1484
rect 5228 1436 5236 1444
rect 5708 1436 5716 1444
rect 3036 1406 3038 1414
rect 3038 1406 3044 1414
rect 3052 1406 3060 1414
rect 3068 1406 3074 1414
rect 3074 1406 3076 1414
rect 1388 1396 1396 1404
rect 3692 1396 3700 1404
rect 5036 1356 5044 1364
rect 5068 1356 5076 1364
rect 6028 1336 6036 1344
rect 940 1316 948 1324
rect 972 1316 980 1324
rect 2060 1316 2068 1324
rect 3340 1316 3348 1324
rect 140 1296 148 1304
rect 1580 1296 1588 1304
rect 4044 1296 4052 1304
rect 3724 1276 3732 1284
rect 5196 1276 5204 1284
rect 4684 1256 4692 1264
rect 428 1236 436 1244
rect 5100 1236 5108 1244
rect 1004 1216 1012 1224
rect 1420 1216 1428 1224
rect 5036 1216 5044 1224
rect 5068 1216 5076 1224
rect 1500 1206 1502 1214
rect 1502 1206 1508 1214
rect 1516 1206 1524 1214
rect 1532 1206 1538 1214
rect 1538 1206 1540 1214
rect 4572 1206 4574 1214
rect 4574 1206 4580 1214
rect 4588 1206 4596 1214
rect 4604 1206 4610 1214
rect 4610 1206 4612 1214
rect 2572 1196 2580 1204
rect 5836 1196 5844 1204
rect 4428 1176 4436 1184
rect 4492 1176 4500 1184
rect 5420 1176 5428 1184
rect 5900 1176 5908 1184
rect 6028 1176 6036 1184
rect 1932 1156 1940 1164
rect 2860 1136 2868 1144
rect 3692 1136 3700 1144
rect 4300 1136 4308 1144
rect 5036 1136 5044 1144
rect 940 1116 948 1124
rect 1228 1116 1236 1124
rect 4460 1116 4468 1124
rect 5708 1096 5716 1104
rect 1388 1076 1396 1084
rect 2956 1076 2964 1084
rect 4076 1076 4084 1084
rect 4108 1076 4116 1084
rect 5676 1076 5684 1084
rect 1068 1056 1076 1064
rect 3820 1056 3828 1064
rect 460 1036 468 1044
rect 4012 1016 4020 1024
rect 4108 1016 4116 1024
rect 5708 1036 5716 1044
rect 3036 1006 3038 1014
rect 3038 1006 3044 1014
rect 3052 1006 3060 1014
rect 3068 1006 3074 1014
rect 3074 1006 3076 1014
rect 3340 976 3348 984
rect 4844 976 4852 984
rect 5068 976 5076 984
rect 5868 976 5876 984
rect 5964 976 5972 984
rect 6028 976 6036 984
rect 364 956 372 964
rect 812 936 820 944
rect 972 936 980 944
rect 2956 936 2964 944
rect 3596 936 3604 944
rect 844 916 852 924
rect 1004 916 1012 924
rect 3660 916 3668 924
rect 4300 916 4308 924
rect 4364 916 4372 924
rect 4428 916 4436 924
rect 4492 916 4500 924
rect 1356 876 1364 884
rect 1068 856 1076 864
rect 524 816 532 824
rect 4652 816 4660 824
rect 1500 806 1502 814
rect 1502 806 1508 814
rect 1516 806 1524 814
rect 1532 806 1538 814
rect 1538 806 1540 814
rect 4572 806 4574 814
rect 4574 806 4580 814
rect 4588 806 4596 814
rect 4604 806 4610 814
rect 4610 806 4612 814
rect 1612 796 1620 804
rect 3180 756 3188 764
rect 4364 776 4372 784
rect 1932 736 1940 744
rect 3948 736 3956 744
rect 716 716 724 724
rect 1452 716 1460 724
rect 5420 736 5428 744
rect 4460 716 4468 724
rect 44 696 52 704
rect 4108 696 4116 704
rect 5548 696 5556 704
rect 716 676 724 684
rect 5164 676 5172 684
rect 5868 676 5876 684
rect 460 636 468 644
rect 4012 616 4020 624
rect 3036 606 3038 614
rect 3038 606 3044 614
rect 3052 606 3060 614
rect 3068 606 3074 614
rect 3074 606 3076 614
rect 2060 576 2068 584
rect 556 556 564 564
rect 1452 556 1460 564
rect 3820 556 3828 564
rect 4652 556 4660 564
rect 2156 536 2164 544
rect 3596 536 3604 544
rect 3948 536 3956 544
rect 3660 516 3668 524
rect 5548 516 5556 524
rect 5804 456 5812 464
rect 6092 416 6100 424
rect 1500 406 1502 414
rect 1502 406 1508 414
rect 1516 406 1524 414
rect 1532 406 1538 414
rect 1538 406 1540 414
rect 4572 406 4574 414
rect 4574 406 4580 414
rect 4588 406 4596 414
rect 4604 406 4610 414
rect 4610 406 4612 414
rect 5036 396 5044 404
rect 4076 356 4084 364
rect 5164 336 5172 344
rect 5708 336 5716 344
rect 2572 296 2580 304
rect 2060 276 2068 284
rect 2828 276 2836 284
rect 3180 276 3188 284
rect 3820 276 3828 284
rect 4076 276 4084 284
rect 3036 206 3038 214
rect 3038 206 3044 214
rect 3052 206 3060 214
rect 3068 206 3074 214
rect 3074 206 3076 214
rect 4044 176 4052 184
rect 972 156 980 164
rect 2828 136 2836 144
rect 5452 136 5460 144
rect 5676 136 5684 144
rect 524 116 532 124
rect 972 116 980 124
rect 5836 116 5844 124
rect 5036 96 5044 104
rect 5516 96 5524 104
rect 5676 16 5684 24
rect 1500 6 1502 14
rect 1502 6 1508 14
rect 1516 6 1524 14
rect 1532 6 1538 14
rect 1538 6 1540 14
rect 4572 6 4574 14
rect 4574 6 4580 14
rect 4588 6 4596 14
rect 4604 6 4610 14
rect 4610 6 4612 14
<< metal4 >>
rect 1496 5614 1544 5640
rect 1496 5606 1500 5614
rect 1508 5606 1516 5614
rect 1524 5606 1532 5614
rect 1540 5606 1544 5614
rect 1226 5504 1238 5506
rect 1226 5496 1228 5504
rect 1236 5496 1238 5504
rect 330 5464 342 5466
rect 330 5456 332 5464
rect 340 5456 342 5464
rect 170 4844 182 4846
rect 170 4836 172 4844
rect 180 4836 182 4844
rect 170 4364 182 4836
rect 170 4356 172 4364
rect 180 4356 182 4364
rect 170 4354 182 4356
rect 138 4284 150 4286
rect 138 4276 140 4284
rect 148 4276 150 4284
rect 138 3204 150 4276
rect 330 4124 342 5456
rect 1226 5424 1238 5496
rect 1226 5416 1228 5424
rect 1236 5416 1238 5424
rect 1226 5414 1238 5416
rect 458 5364 470 5366
rect 458 5356 460 5364
rect 468 5356 470 5364
rect 362 5304 374 5306
rect 362 5296 364 5304
rect 372 5296 374 5304
rect 362 4284 374 5296
rect 458 5144 470 5356
rect 970 5344 982 5346
rect 970 5336 972 5344
rect 980 5336 982 5344
rect 458 5136 460 5144
rect 468 5136 470 5144
rect 458 5134 470 5136
rect 522 5324 534 5326
rect 522 5316 524 5324
rect 532 5316 534 5324
rect 458 5104 470 5106
rect 458 5096 460 5104
rect 468 5096 470 5104
rect 458 4584 470 5096
rect 458 4576 460 4584
rect 468 4576 470 4584
rect 458 4574 470 4576
rect 362 4276 364 4284
rect 372 4276 374 4284
rect 362 4274 374 4276
rect 426 4544 438 4546
rect 426 4536 428 4544
rect 436 4536 438 4544
rect 330 4116 332 4124
rect 340 4116 342 4124
rect 330 4114 342 4116
rect 426 3884 438 4536
rect 522 4544 534 5316
rect 650 5244 662 5246
rect 650 5236 652 5244
rect 660 5236 662 5244
rect 650 4904 662 5236
rect 906 4964 918 4966
rect 906 4956 908 4964
rect 916 4956 918 4964
rect 650 4896 652 4904
rect 660 4896 662 4904
rect 650 4894 662 4896
rect 874 4924 886 4926
rect 874 4916 876 4924
rect 884 4916 886 4924
rect 522 4536 524 4544
rect 532 4536 534 4544
rect 522 4534 534 4536
rect 874 4424 886 4916
rect 874 4416 876 4424
rect 884 4416 886 4424
rect 874 4414 886 4416
rect 586 4304 598 4306
rect 586 4296 588 4304
rect 596 4296 598 4304
rect 426 3876 428 3884
rect 436 3876 438 3884
rect 426 3874 438 3876
rect 458 3984 470 3986
rect 458 3976 460 3984
rect 468 3976 470 3984
rect 458 3844 470 3976
rect 586 3904 598 4296
rect 586 3896 588 3904
rect 596 3896 598 3904
rect 586 3894 598 3896
rect 906 3924 918 4956
rect 970 4944 982 5336
rect 970 4936 972 4944
rect 980 4936 982 4944
rect 970 4934 982 4936
rect 1496 5214 1544 5606
rect 2506 5444 2518 5446
rect 2506 5436 2508 5444
rect 2516 5436 2518 5444
rect 1496 5206 1500 5214
rect 1508 5206 1516 5214
rect 1524 5206 1532 5214
rect 1540 5206 1544 5214
rect 1034 4904 1046 4906
rect 1034 4896 1036 4904
rect 1044 4896 1046 4904
rect 938 4724 950 4726
rect 938 4716 940 4724
rect 948 4716 950 4724
rect 938 4684 950 4716
rect 938 4676 940 4684
rect 948 4676 950 4684
rect 938 4674 950 4676
rect 1034 4524 1046 4896
rect 1496 4814 1544 5206
rect 2442 5364 2454 5366
rect 2442 5356 2444 5364
rect 2452 5356 2454 5364
rect 1898 5084 1910 5086
rect 1898 5076 1900 5084
rect 1908 5076 1910 5084
rect 1496 4806 1500 4814
rect 1508 4806 1516 4814
rect 1524 4806 1532 4814
rect 1540 4806 1544 4814
rect 1354 4804 1366 4806
rect 1354 4796 1356 4804
rect 1364 4796 1366 4804
rect 1354 4704 1366 4796
rect 1354 4696 1356 4704
rect 1364 4696 1366 4704
rect 1354 4694 1366 4696
rect 1034 4516 1036 4524
rect 1044 4516 1046 4524
rect 1034 4514 1046 4516
rect 1322 4464 1334 4466
rect 1322 4456 1324 4464
rect 1332 4456 1334 4464
rect 1290 4224 1302 4226
rect 1290 4216 1292 4224
rect 1300 4216 1302 4224
rect 906 3916 908 3924
rect 916 3916 918 3924
rect 458 3836 460 3844
rect 468 3836 470 3844
rect 458 3834 470 3836
rect 906 3744 918 3916
rect 1162 4164 1174 4166
rect 1162 4156 1164 4164
rect 1172 4156 1174 4164
rect 1066 3824 1078 3826
rect 1066 3816 1068 3824
rect 1076 3816 1078 3824
rect 1066 3764 1078 3816
rect 1066 3756 1068 3764
rect 1076 3756 1078 3764
rect 1066 3754 1078 3756
rect 906 3736 908 3744
rect 916 3736 918 3744
rect 906 3734 918 3736
rect 138 3196 140 3204
rect 148 3196 150 3204
rect 138 3194 150 3196
rect 938 3564 950 3566
rect 938 3556 940 3564
rect 948 3556 950 3564
rect 362 2644 374 2646
rect 362 2636 364 2644
rect 372 2636 374 2644
rect 42 2124 54 2126
rect 42 2116 44 2124
rect 52 2116 54 2124
rect 42 704 54 2116
rect 138 1904 150 1906
rect 138 1896 140 1904
rect 148 1896 150 1904
rect 138 1304 150 1896
rect 362 1844 374 2636
rect 938 2324 950 3556
rect 1162 3524 1174 4156
rect 1290 3784 1302 4216
rect 1290 3776 1292 3784
rect 1300 3776 1302 3784
rect 1290 3774 1302 3776
rect 1322 3764 1334 4456
rect 1354 4424 1366 4426
rect 1354 4416 1356 4424
rect 1364 4416 1366 4424
rect 1354 4244 1366 4416
rect 1354 4236 1356 4244
rect 1364 4236 1366 4244
rect 1354 4234 1366 4236
rect 1496 4414 1544 4806
rect 1706 5024 1718 5026
rect 1706 5016 1708 5024
rect 1716 5016 1718 5024
rect 1706 4684 1718 5016
rect 1706 4676 1708 4684
rect 1716 4676 1718 4684
rect 1706 4674 1718 4676
rect 1770 4604 1782 4606
rect 1770 4596 1772 4604
rect 1780 4596 1782 4604
rect 1496 4406 1500 4414
rect 1508 4406 1516 4414
rect 1524 4406 1532 4414
rect 1540 4406 1544 4414
rect 1322 3756 1324 3764
rect 1332 3756 1334 3764
rect 1322 3754 1334 3756
rect 1496 4014 1544 4406
rect 1610 4444 1622 4446
rect 1610 4436 1612 4444
rect 1620 4436 1622 4444
rect 1610 4124 1622 4436
rect 1610 4116 1612 4124
rect 1620 4116 1622 4124
rect 1610 4114 1622 4116
rect 1674 4384 1686 4386
rect 1674 4376 1676 4384
rect 1684 4376 1686 4384
rect 1674 4104 1686 4376
rect 1770 4124 1782 4596
rect 1898 4504 1910 5076
rect 2250 4984 2262 4986
rect 2250 4976 2252 4984
rect 2260 4976 2262 4984
rect 1898 4496 1900 4504
rect 1908 4496 1910 4504
rect 1898 4494 1910 4496
rect 1962 4864 1974 4866
rect 1962 4856 1964 4864
rect 1972 4856 1974 4864
rect 1962 4304 1974 4856
rect 1962 4296 1964 4304
rect 1972 4296 1974 4304
rect 1962 4294 1974 4296
rect 2218 4324 2230 4326
rect 2218 4316 2220 4324
rect 2228 4316 2230 4324
rect 2026 4284 2038 4286
rect 2026 4276 2028 4284
rect 2036 4276 2038 4284
rect 1770 4116 1772 4124
rect 1780 4116 1782 4124
rect 1770 4114 1782 4116
rect 1898 4204 1910 4206
rect 1898 4196 1900 4204
rect 1908 4196 1910 4204
rect 1674 4096 1676 4104
rect 1684 4096 1686 4104
rect 1674 4094 1686 4096
rect 1496 4006 1500 4014
rect 1508 4006 1516 4014
rect 1524 4006 1532 4014
rect 1540 4006 1544 4014
rect 1496 3614 1544 4006
rect 1898 3764 1910 4196
rect 2026 4024 2038 4276
rect 2026 4016 2028 4024
rect 2036 4016 2038 4024
rect 2026 4014 2038 4016
rect 1898 3756 1900 3764
rect 1908 3756 1910 3764
rect 1898 3754 1910 3756
rect 2218 3624 2230 4316
rect 2250 3924 2262 4976
rect 2442 4964 2454 5356
rect 2442 4956 2444 4964
rect 2452 4956 2454 4964
rect 2442 4954 2454 4956
rect 2410 4704 2422 4706
rect 2410 4696 2412 4704
rect 2420 4696 2422 4704
rect 2250 3916 2252 3924
rect 2260 3916 2262 3924
rect 2250 3914 2262 3916
rect 2314 4224 2326 4226
rect 2314 4216 2316 4224
rect 2324 4216 2326 4224
rect 2218 3616 2220 3624
rect 2228 3616 2230 3624
rect 2218 3614 2230 3616
rect 1496 3606 1500 3614
rect 1508 3606 1516 3614
rect 1524 3606 1532 3614
rect 1540 3606 1544 3614
rect 1162 3516 1164 3524
rect 1172 3516 1174 3524
rect 1162 3514 1174 3516
rect 1290 3584 1302 3586
rect 1290 3576 1292 3584
rect 1300 3576 1302 3584
rect 1098 3224 1110 3226
rect 1098 3216 1100 3224
rect 1108 3216 1110 3224
rect 1098 2744 1110 3216
rect 1290 3184 1302 3576
rect 1496 3214 1544 3606
rect 2282 3504 2294 3506
rect 2282 3496 2284 3504
rect 2292 3496 2294 3504
rect 1496 3206 1500 3214
rect 1508 3206 1516 3214
rect 1524 3206 1532 3214
rect 1540 3206 1544 3214
rect 1290 3176 1292 3184
rect 1300 3176 1302 3184
rect 1290 3174 1302 3176
rect 1386 3204 1398 3206
rect 1386 3196 1388 3204
rect 1396 3196 1398 3204
rect 1098 2736 1100 2744
rect 1108 2736 1110 2744
rect 1098 2734 1110 2736
rect 1386 2684 1398 3196
rect 1386 2676 1388 2684
rect 1396 2676 1398 2684
rect 1386 2674 1398 2676
rect 1496 2814 1544 3206
rect 1496 2806 1500 2814
rect 1508 2806 1516 2814
rect 1524 2806 1532 2814
rect 1540 2806 1544 2814
rect 938 2316 940 2324
rect 948 2316 950 2324
rect 938 2314 950 2316
rect 1496 2414 1544 2806
rect 1962 3444 1974 3446
rect 1962 3436 1964 3444
rect 1972 3436 1974 3444
rect 1962 3104 1974 3436
rect 2282 3304 2294 3496
rect 2314 3424 2326 4216
rect 2314 3416 2316 3424
rect 2324 3416 2326 3424
rect 2314 3414 2326 3416
rect 2378 3704 2390 3706
rect 2378 3696 2380 3704
rect 2388 3696 2390 3704
rect 2282 3296 2284 3304
rect 2292 3296 2294 3304
rect 1962 3096 1964 3104
rect 1972 3096 1974 3104
rect 1962 2764 1974 3096
rect 2058 3184 2070 3186
rect 2058 3176 2060 3184
rect 2068 3176 2070 3184
rect 2058 2844 2070 3176
rect 2058 2836 2060 2844
rect 2068 2836 2070 2844
rect 2058 2834 2070 2836
rect 2282 2824 2294 3296
rect 2282 2816 2284 2824
rect 2292 2816 2294 2824
rect 2282 2814 2294 2816
rect 2314 3284 2326 3286
rect 2314 3276 2316 3284
rect 2324 3276 2326 3284
rect 1962 2756 1964 2764
rect 1972 2756 1974 2764
rect 1962 2754 1974 2756
rect 1994 2804 2006 2806
rect 1994 2796 1996 2804
rect 2004 2796 2006 2804
rect 1994 2604 2006 2796
rect 2314 2784 2326 3276
rect 2378 3164 2390 3696
rect 2410 3604 2422 4696
rect 2506 4424 2518 5436
rect 3032 5414 3080 5640
rect 3032 5406 3036 5414
rect 3044 5406 3052 5414
rect 3060 5406 3068 5414
rect 3076 5406 3080 5414
rect 2954 5044 2966 5046
rect 2954 5036 2956 5044
rect 2964 5036 2966 5044
rect 2506 4416 2508 4424
rect 2516 4416 2518 4424
rect 2506 4414 2518 4416
rect 2762 4944 2774 4946
rect 2762 4936 2764 4944
rect 2772 4936 2774 4944
rect 2762 4504 2774 4936
rect 2762 4496 2764 4504
rect 2772 4496 2774 4504
rect 2666 4384 2678 4386
rect 2666 4376 2668 4384
rect 2676 4376 2678 4384
rect 2666 3904 2678 4376
rect 2666 3896 2668 3904
rect 2676 3896 2678 3904
rect 2666 3894 2678 3896
rect 2762 3744 2774 4496
rect 2826 4924 2838 4926
rect 2826 4916 2828 4924
rect 2836 4916 2838 4924
rect 2826 3824 2838 4916
rect 2954 4904 2966 5036
rect 2954 4896 2956 4904
rect 2964 4896 2966 4904
rect 2954 4894 2966 4896
rect 3032 5014 3080 5406
rect 4568 5614 4616 5640
rect 4568 5606 4572 5614
rect 4580 5606 4588 5614
rect 4596 5606 4604 5614
rect 4612 5606 4616 5614
rect 3722 5384 3734 5386
rect 3722 5376 3724 5384
rect 3732 5376 3734 5384
rect 3722 5144 3734 5376
rect 4426 5224 4438 5226
rect 4426 5216 4428 5224
rect 4436 5216 4438 5224
rect 4106 5184 4118 5186
rect 4106 5176 4108 5184
rect 4116 5176 4118 5184
rect 3722 5136 3724 5144
rect 3732 5136 3734 5144
rect 3722 5134 3734 5136
rect 3978 5144 3990 5146
rect 3978 5136 3980 5144
rect 3988 5136 3990 5144
rect 3032 5006 3036 5014
rect 3044 5006 3052 5014
rect 3060 5006 3068 5014
rect 3076 5006 3080 5014
rect 3032 4614 3080 5006
rect 3914 5004 3926 5006
rect 3914 4996 3916 5004
rect 3924 4996 3926 5004
rect 3306 4984 3318 4986
rect 3306 4976 3308 4984
rect 3316 4976 3318 4984
rect 3306 4724 3318 4976
rect 3306 4716 3308 4724
rect 3316 4716 3318 4724
rect 3306 4714 3318 4716
rect 3818 4764 3830 4766
rect 3818 4756 3820 4764
rect 3828 4756 3830 4764
rect 3032 4606 3036 4614
rect 3044 4606 3052 4614
rect 3060 4606 3068 4614
rect 3076 4606 3080 4614
rect 2986 4464 2998 4466
rect 2986 4456 2988 4464
rect 2996 4456 2998 4464
rect 2954 4404 2966 4406
rect 2954 4396 2956 4404
rect 2964 4396 2966 4404
rect 2826 3816 2828 3824
rect 2836 3816 2838 3824
rect 2826 3814 2838 3816
rect 2922 3984 2934 3986
rect 2922 3976 2924 3984
rect 2932 3976 2934 3984
rect 2762 3736 2764 3744
rect 2772 3736 2774 3744
rect 2762 3734 2774 3736
rect 2410 3596 2412 3604
rect 2420 3596 2422 3604
rect 2410 3594 2422 3596
rect 2442 3664 2454 3666
rect 2442 3656 2444 3664
rect 2452 3656 2454 3664
rect 2378 3156 2380 3164
rect 2388 3156 2390 3164
rect 2378 3154 2390 3156
rect 2442 2844 2454 3656
rect 2698 3404 2710 3406
rect 2698 3396 2700 3404
rect 2708 3396 2710 3404
rect 2698 3084 2710 3396
rect 2922 3404 2934 3976
rect 2922 3396 2924 3404
rect 2932 3396 2934 3404
rect 2922 3394 2934 3396
rect 2954 3284 2966 4396
rect 2986 3304 2998 4456
rect 2986 3296 2988 3304
rect 2996 3296 2998 3304
rect 2986 3294 2998 3296
rect 3032 4214 3080 4606
rect 3402 4644 3414 4646
rect 3402 4636 3404 4644
rect 3412 4636 3414 4644
rect 3032 4206 3036 4214
rect 3044 4206 3052 4214
rect 3060 4206 3068 4214
rect 3076 4206 3080 4214
rect 3032 3814 3080 4206
rect 3032 3806 3036 3814
rect 3044 3806 3052 3814
rect 3060 3806 3068 3814
rect 3076 3806 3080 3814
rect 3032 3414 3080 3806
rect 3370 4224 3382 4226
rect 3370 4216 3372 4224
rect 3380 4216 3382 4224
rect 3370 3484 3382 4216
rect 3402 3984 3414 4636
rect 3818 4104 3830 4756
rect 3914 4764 3926 4996
rect 3978 4804 3990 5136
rect 4106 4864 4118 5176
rect 4394 5124 4406 5126
rect 4394 5116 4396 5124
rect 4404 5116 4406 5124
rect 4106 4856 4108 4864
rect 4116 4856 4118 4864
rect 4106 4854 4118 4856
rect 4138 5104 4150 5106
rect 4138 5096 4140 5104
rect 4148 5096 4150 5104
rect 3978 4796 3980 4804
rect 3988 4796 3990 4804
rect 3978 4794 3990 4796
rect 3914 4756 3916 4764
rect 3924 4756 3926 4764
rect 3914 4754 3926 4756
rect 4138 4644 4150 5096
rect 4266 4904 4278 4906
rect 4266 4896 4268 4904
rect 4276 4896 4278 4904
rect 4266 4684 4278 4896
rect 4394 4864 4406 5116
rect 4394 4856 4396 4864
rect 4404 4856 4406 4864
rect 4394 4854 4406 4856
rect 4266 4676 4268 4684
rect 4276 4676 4278 4684
rect 4266 4674 4278 4676
rect 4138 4636 4140 4644
rect 4148 4636 4150 4644
rect 4138 4634 4150 4636
rect 3978 4624 3990 4626
rect 3978 4616 3980 4624
rect 3988 4616 3990 4624
rect 3978 4284 3990 4616
rect 3978 4276 3980 4284
rect 3988 4276 3990 4284
rect 3978 4274 3990 4276
rect 3818 4096 3820 4104
rect 3828 4096 3830 4104
rect 3818 4094 3830 4096
rect 4202 4204 4214 4206
rect 4202 4196 4204 4204
rect 4212 4196 4214 4204
rect 3402 3976 3404 3984
rect 3412 3976 3414 3984
rect 3402 3974 3414 3976
rect 3434 4084 3446 4086
rect 3434 4076 3436 4084
rect 3444 4076 3446 4084
rect 3370 3476 3372 3484
rect 3380 3476 3382 3484
rect 3370 3474 3382 3476
rect 3032 3406 3036 3414
rect 3044 3406 3052 3414
rect 3060 3406 3068 3414
rect 3076 3406 3080 3414
rect 2954 3276 2956 3284
rect 2964 3276 2966 3284
rect 2954 3274 2966 3276
rect 2698 3076 2700 3084
rect 2708 3076 2710 3084
rect 2698 3074 2710 3076
rect 2730 3124 2742 3126
rect 2730 3116 2732 3124
rect 2740 3116 2742 3124
rect 2442 2836 2444 2844
rect 2452 2836 2454 2844
rect 2442 2834 2454 2836
rect 2506 2844 2518 2846
rect 2506 2836 2508 2844
rect 2516 2836 2518 2844
rect 2314 2776 2316 2784
rect 2324 2776 2326 2784
rect 2314 2774 2326 2776
rect 2506 2784 2518 2836
rect 2730 2804 2742 3116
rect 2922 3124 2934 3126
rect 2922 3116 2924 3124
rect 2932 3116 2934 3124
rect 2922 2844 2934 3116
rect 2922 2836 2924 2844
rect 2932 2836 2934 2844
rect 2922 2834 2934 2836
rect 2954 3024 2966 3026
rect 2954 3016 2956 3024
rect 2964 3016 2966 3024
rect 2730 2796 2732 2804
rect 2740 2796 2742 2804
rect 2730 2794 2742 2796
rect 2506 2776 2508 2784
rect 2516 2776 2518 2784
rect 2506 2774 2518 2776
rect 1994 2596 1996 2604
rect 2004 2596 2006 2604
rect 1994 2594 2006 2596
rect 2858 2684 2870 2686
rect 2858 2676 2860 2684
rect 2868 2676 2870 2684
rect 2602 2564 2614 2566
rect 2602 2556 2604 2564
rect 2612 2556 2614 2564
rect 1496 2406 1500 2414
rect 1508 2406 1516 2414
rect 1524 2406 1532 2414
rect 1540 2406 1544 2414
rect 362 1836 364 1844
rect 372 1836 374 1844
rect 362 1834 374 1836
rect 554 2224 566 2226
rect 554 2216 556 2224
rect 564 2216 566 2224
rect 426 1604 438 1606
rect 426 1596 428 1604
rect 436 1596 438 1604
rect 138 1296 140 1304
rect 148 1296 150 1304
rect 138 1294 150 1296
rect 362 1524 374 1526
rect 362 1516 364 1524
rect 372 1516 374 1524
rect 362 964 374 1516
rect 426 1244 438 1596
rect 426 1236 428 1244
rect 436 1236 438 1244
rect 426 1234 438 1236
rect 362 956 364 964
rect 372 956 374 964
rect 362 954 374 956
rect 458 1044 470 1046
rect 458 1036 460 1044
rect 468 1036 470 1044
rect 42 696 44 704
rect 52 696 54 704
rect 42 694 54 696
rect 458 644 470 1036
rect 458 636 460 644
rect 468 636 470 644
rect 458 634 470 636
rect 522 824 534 826
rect 522 816 524 824
rect 532 816 534 824
rect 522 124 534 816
rect 554 564 566 2216
rect 1496 2014 1544 2406
rect 2410 2444 2422 2446
rect 2410 2436 2412 2444
rect 2420 2436 2422 2444
rect 2314 2284 2326 2286
rect 2314 2276 2316 2284
rect 2324 2276 2326 2284
rect 1496 2006 1500 2014
rect 1508 2006 1516 2014
rect 1524 2006 1532 2014
rect 1540 2006 1544 2014
rect 842 1984 854 1986
rect 842 1976 844 1984
rect 852 1976 854 1984
rect 810 1724 822 1726
rect 810 1716 812 1724
rect 820 1716 822 1724
rect 810 944 822 1716
rect 810 936 812 944
rect 820 936 822 944
rect 810 934 822 936
rect 842 924 854 1976
rect 1450 1904 1462 1906
rect 1450 1896 1452 1904
rect 1460 1896 1462 1904
rect 1226 1804 1238 1806
rect 1226 1796 1228 1804
rect 1236 1796 1238 1804
rect 938 1324 950 1326
rect 938 1316 940 1324
rect 948 1316 950 1324
rect 938 1124 950 1316
rect 938 1116 940 1124
rect 948 1116 950 1124
rect 938 1114 950 1116
rect 970 1324 982 1326
rect 970 1316 972 1324
rect 980 1316 982 1324
rect 970 944 982 1316
rect 970 936 972 944
rect 980 936 982 944
rect 970 934 982 936
rect 1002 1224 1014 1226
rect 1002 1216 1004 1224
rect 1012 1216 1014 1224
rect 842 916 844 924
rect 852 916 854 924
rect 842 914 854 916
rect 1002 924 1014 1216
rect 1226 1124 1238 1796
rect 1418 1644 1430 1646
rect 1418 1636 1420 1644
rect 1428 1636 1430 1644
rect 1226 1116 1228 1124
rect 1236 1116 1238 1124
rect 1226 1114 1238 1116
rect 1354 1564 1366 1566
rect 1354 1556 1356 1564
rect 1364 1556 1366 1564
rect 1002 916 1004 924
rect 1012 916 1014 924
rect 1002 914 1014 916
rect 1066 1064 1078 1066
rect 1066 1056 1068 1064
rect 1076 1056 1078 1064
rect 1066 864 1078 1056
rect 1354 884 1366 1556
rect 1386 1404 1398 1406
rect 1386 1396 1388 1404
rect 1396 1396 1398 1404
rect 1386 1084 1398 1396
rect 1418 1224 1430 1636
rect 1418 1216 1420 1224
rect 1428 1216 1430 1224
rect 1418 1214 1430 1216
rect 1386 1076 1388 1084
rect 1396 1076 1398 1084
rect 1386 1074 1398 1076
rect 1354 876 1356 884
rect 1364 876 1366 884
rect 1354 874 1366 876
rect 1066 856 1068 864
rect 1076 856 1078 864
rect 1066 854 1078 856
rect 714 724 726 726
rect 714 716 716 724
rect 724 716 726 724
rect 714 684 726 716
rect 714 676 716 684
rect 724 676 726 684
rect 714 674 726 676
rect 1450 724 1462 1896
rect 1450 716 1452 724
rect 1460 716 1462 724
rect 554 556 556 564
rect 564 556 566 564
rect 554 554 566 556
rect 1450 564 1462 716
rect 1450 556 1452 564
rect 1460 556 1462 564
rect 1450 554 1462 556
rect 1496 1614 1544 2006
rect 2218 2144 2230 2146
rect 2218 2136 2220 2144
rect 2228 2136 2230 2144
rect 2058 1904 2070 1906
rect 2058 1896 2060 1904
rect 2068 1896 2070 1904
rect 1496 1606 1500 1614
rect 1508 1606 1516 1614
rect 1524 1606 1532 1614
rect 1540 1606 1544 1614
rect 1496 1214 1544 1606
rect 1578 1684 1590 1686
rect 1578 1676 1580 1684
rect 1588 1676 1590 1684
rect 1578 1304 1590 1676
rect 2058 1644 2070 1896
rect 2090 1904 2102 1906
rect 2090 1896 2092 1904
rect 2100 1896 2102 1904
rect 2090 1764 2102 1896
rect 2218 1784 2230 2136
rect 2314 2124 2326 2276
rect 2314 2116 2316 2124
rect 2324 2116 2326 2124
rect 2314 2044 2326 2116
rect 2314 2036 2316 2044
rect 2324 2036 2326 2044
rect 2314 2034 2326 2036
rect 2218 1776 2220 1784
rect 2228 1776 2230 1784
rect 2218 1774 2230 1776
rect 2090 1756 2092 1764
rect 2100 1756 2102 1764
rect 2090 1754 2102 1756
rect 2410 1764 2422 2436
rect 2602 2164 2614 2556
rect 2730 2544 2742 2546
rect 2730 2536 2732 2544
rect 2740 2536 2742 2544
rect 2730 2324 2742 2536
rect 2858 2504 2870 2676
rect 2954 2544 2966 3016
rect 3032 3014 3080 3406
rect 3434 3404 3446 4076
rect 4202 3724 4214 4196
rect 4426 3764 4438 5216
rect 4568 5214 4616 5606
rect 6090 5604 6102 5606
rect 6090 5596 6092 5604
rect 6100 5596 6102 5604
rect 5578 5444 5590 5446
rect 5578 5436 5580 5444
rect 5588 5436 5590 5444
rect 5258 5364 5270 5366
rect 5258 5356 5260 5364
rect 5268 5356 5270 5364
rect 4568 5206 4572 5214
rect 4580 5206 4588 5214
rect 4596 5206 4604 5214
rect 4612 5206 4616 5214
rect 4490 4824 4502 4826
rect 4490 4816 4492 4824
rect 4500 4816 4502 4824
rect 4490 4764 4502 4816
rect 4490 4756 4492 4764
rect 4500 4756 4502 4764
rect 4490 4754 4502 4756
rect 4568 4814 4616 5206
rect 5194 5324 5206 5326
rect 5194 5316 5196 5324
rect 5204 5316 5206 5324
rect 4650 5124 4662 5126
rect 4650 5116 4652 5124
rect 4660 5116 4662 5124
rect 4650 4824 4662 5116
rect 4874 5084 4886 5086
rect 4874 5076 4876 5084
rect 4884 5076 4886 5084
rect 4874 5044 4886 5076
rect 4874 5036 4876 5044
rect 4884 5036 4886 5044
rect 4874 5034 4886 5036
rect 4650 4816 4652 4824
rect 4660 4816 4662 4824
rect 4650 4814 4662 4816
rect 5034 4964 5046 4966
rect 5034 4956 5036 4964
rect 5044 4956 5046 4964
rect 4568 4806 4572 4814
rect 4580 4806 4588 4814
rect 4596 4806 4604 4814
rect 4612 4806 4616 4814
rect 4426 3756 4428 3764
rect 4436 3756 4438 3764
rect 4426 3754 4438 3756
rect 4568 4414 4616 4806
rect 4682 4724 4694 4726
rect 4682 4716 4684 4724
rect 4692 4716 4694 4724
rect 4682 4544 4694 4716
rect 5034 4724 5046 4956
rect 5194 4844 5206 5316
rect 5258 5084 5270 5356
rect 5258 5076 5260 5084
rect 5268 5076 5270 5084
rect 5258 5074 5270 5076
rect 5418 5184 5430 5186
rect 5418 5176 5420 5184
rect 5428 5176 5430 5184
rect 5194 4836 5196 4844
rect 5204 4836 5206 4844
rect 5194 4834 5206 4836
rect 5034 4716 5036 4724
rect 5044 4716 5046 4724
rect 5034 4714 5046 4716
rect 4938 4684 4950 4686
rect 4938 4676 4940 4684
rect 4948 4676 4950 4684
rect 4682 4536 4684 4544
rect 4692 4536 4694 4544
rect 4682 4534 4694 4536
rect 4746 4544 4758 4546
rect 4746 4536 4748 4544
rect 4756 4536 4758 4544
rect 4568 4406 4572 4414
rect 4580 4406 4588 4414
rect 4596 4406 4604 4414
rect 4612 4406 4616 4414
rect 4568 4014 4616 4406
rect 4746 4064 4758 4536
rect 4938 4324 4950 4676
rect 5194 4664 5206 4666
rect 5194 4656 5196 4664
rect 5204 4656 5206 4664
rect 5162 4604 5174 4606
rect 5162 4596 5164 4604
rect 5172 4596 5174 4604
rect 5066 4564 5078 4566
rect 5066 4556 5068 4564
rect 5076 4556 5078 4564
rect 5066 4384 5078 4556
rect 5162 4524 5174 4596
rect 5162 4516 5164 4524
rect 5172 4516 5174 4524
rect 5162 4514 5174 4516
rect 5066 4376 5068 4384
rect 5076 4376 5078 4384
rect 5066 4374 5078 4376
rect 4938 4316 4940 4324
rect 4948 4316 4950 4324
rect 4938 4314 4950 4316
rect 5098 4164 5110 4166
rect 5098 4156 5100 4164
rect 5108 4156 5110 4164
rect 5098 4124 5110 4156
rect 5098 4116 5100 4124
rect 5108 4116 5110 4124
rect 5098 4114 5110 4116
rect 4746 4056 4748 4064
rect 4756 4056 4758 4064
rect 4746 4054 4758 4056
rect 4568 4006 4572 4014
rect 4580 4006 4588 4014
rect 4596 4006 4604 4014
rect 4612 4006 4616 4014
rect 4202 3716 4204 3724
rect 4212 3716 4214 3724
rect 4202 3714 4214 3716
rect 3786 3704 3798 3706
rect 3786 3696 3788 3704
rect 3796 3696 3798 3704
rect 3434 3396 3436 3404
rect 3444 3396 3446 3404
rect 3434 3394 3446 3396
rect 3466 3504 3478 3506
rect 3466 3496 3468 3504
rect 3476 3496 3478 3504
rect 3242 3224 3254 3226
rect 3242 3216 3244 3224
rect 3252 3216 3254 3224
rect 3032 3006 3036 3014
rect 3044 3006 3052 3014
rect 3060 3006 3068 3014
rect 3076 3006 3080 3014
rect 2954 2536 2956 2544
rect 2964 2536 2966 2544
rect 2954 2534 2966 2536
rect 2986 2684 2998 2686
rect 2986 2676 2988 2684
rect 2996 2676 2998 2684
rect 2858 2496 2860 2504
rect 2868 2496 2870 2504
rect 2858 2494 2870 2496
rect 2730 2316 2732 2324
rect 2740 2316 2742 2324
rect 2730 2314 2742 2316
rect 2986 2324 2998 2676
rect 2986 2316 2988 2324
rect 2996 2316 2998 2324
rect 2986 2314 2998 2316
rect 3032 2614 3080 3006
rect 3114 3144 3126 3146
rect 3114 3136 3116 3144
rect 3124 3136 3126 3144
rect 3114 2984 3126 3136
rect 3114 2976 3116 2984
rect 3124 2976 3126 2984
rect 3114 2974 3126 2976
rect 3146 3044 3158 3046
rect 3146 3036 3148 3044
rect 3156 3036 3158 3044
rect 3146 2964 3158 3036
rect 3146 2956 3148 2964
rect 3156 2956 3158 2964
rect 3146 2664 3158 2956
rect 3146 2656 3148 2664
rect 3156 2656 3158 2664
rect 3146 2654 3158 2656
rect 3210 2824 3222 2826
rect 3210 2816 3212 2824
rect 3220 2816 3222 2824
rect 3032 2606 3036 2614
rect 3044 2606 3052 2614
rect 3060 2606 3068 2614
rect 3076 2606 3080 2614
rect 2602 2156 2604 2164
rect 2612 2156 2614 2164
rect 2602 2154 2614 2156
rect 3032 2214 3080 2606
rect 3210 2524 3222 2816
rect 3242 2824 3254 3216
rect 3466 3184 3478 3496
rect 3466 3176 3468 3184
rect 3476 3176 3478 3184
rect 3466 3174 3478 3176
rect 3754 3264 3766 3266
rect 3754 3256 3756 3264
rect 3764 3256 3766 3264
rect 3754 3104 3766 3256
rect 3786 3264 3798 3696
rect 4568 3614 4616 4006
rect 4906 4044 4918 4046
rect 4906 4036 4908 4044
rect 4916 4036 4918 4044
rect 4568 3606 4572 3614
rect 4580 3606 4588 3614
rect 4596 3606 4604 3614
rect 4612 3606 4616 3614
rect 4138 3544 4150 3546
rect 4138 3536 4140 3544
rect 4148 3536 4150 3544
rect 3786 3256 3788 3264
rect 3796 3256 3798 3264
rect 3786 3254 3798 3256
rect 4042 3504 4054 3506
rect 4042 3496 4044 3504
rect 4052 3496 4054 3504
rect 3754 3096 3756 3104
rect 3764 3096 3766 3104
rect 3754 3094 3766 3096
rect 4042 3104 4054 3496
rect 4106 3424 4118 3426
rect 4106 3416 4108 3424
rect 4116 3416 4118 3424
rect 4106 3124 4118 3416
rect 4106 3116 4108 3124
rect 4116 3116 4118 3124
rect 4106 3114 4118 3116
rect 4042 3096 4044 3104
rect 4052 3096 4054 3104
rect 3786 3084 3798 3086
rect 3786 3076 3788 3084
rect 3796 3076 3798 3084
rect 3530 3064 3542 3066
rect 3530 3056 3532 3064
rect 3540 3056 3542 3064
rect 3242 2816 3244 2824
rect 3252 2816 3254 2824
rect 3242 2814 3254 2816
rect 3274 2844 3286 2846
rect 3274 2836 3276 2844
rect 3284 2836 3286 2844
rect 3274 2684 3286 2836
rect 3274 2676 3276 2684
rect 3284 2676 3286 2684
rect 3274 2674 3286 2676
rect 3210 2516 3212 2524
rect 3220 2516 3222 2524
rect 3210 2514 3222 2516
rect 3242 2664 3254 2666
rect 3242 2656 3244 2664
rect 3252 2656 3254 2664
rect 3146 2464 3158 2466
rect 3146 2456 3148 2464
rect 3156 2456 3158 2464
rect 3146 2324 3158 2456
rect 3242 2444 3254 2656
rect 3498 2604 3510 2606
rect 3498 2596 3500 2604
rect 3508 2596 3510 2604
rect 3242 2436 3244 2444
rect 3252 2436 3254 2444
rect 3242 2434 3254 2436
rect 3466 2484 3478 2486
rect 3466 2476 3468 2484
rect 3476 2476 3478 2484
rect 3466 2384 3478 2476
rect 3466 2376 3468 2384
rect 3476 2376 3478 2384
rect 3466 2374 3478 2376
rect 3146 2316 3148 2324
rect 3156 2316 3158 2324
rect 3146 2314 3158 2316
rect 3210 2304 3222 2306
rect 3210 2296 3212 2304
rect 3220 2296 3222 2304
rect 3032 2206 3036 2214
rect 3044 2206 3052 2214
rect 3060 2206 3068 2214
rect 3076 2206 3080 2214
rect 2410 1756 2412 1764
rect 2420 1756 2422 1764
rect 2410 1754 2422 1756
rect 2858 1904 2870 1906
rect 2858 1896 2860 1904
rect 2868 1896 2870 1904
rect 2858 1804 2870 1896
rect 2858 1796 2860 1804
rect 2868 1796 2870 1804
rect 2058 1636 2060 1644
rect 2068 1636 2070 1644
rect 2058 1634 2070 1636
rect 2154 1704 2166 1706
rect 2154 1696 2156 1704
rect 2164 1696 2166 1704
rect 1578 1296 1580 1304
rect 1588 1296 1590 1304
rect 1578 1294 1590 1296
rect 1610 1564 1622 1566
rect 1610 1556 1612 1564
rect 1620 1556 1622 1564
rect 1496 1206 1500 1214
rect 1508 1206 1516 1214
rect 1524 1206 1532 1214
rect 1540 1206 1544 1214
rect 1496 814 1544 1206
rect 1496 806 1500 814
rect 1508 806 1516 814
rect 1524 806 1532 814
rect 1540 806 1544 814
rect 1496 414 1544 806
rect 1610 804 1622 1556
rect 2058 1324 2070 1326
rect 2058 1316 2060 1324
rect 2068 1316 2070 1324
rect 1610 796 1612 804
rect 1620 796 1622 804
rect 1610 794 1622 796
rect 1930 1164 1942 1166
rect 1930 1156 1932 1164
rect 1940 1156 1942 1164
rect 1930 744 1942 1156
rect 1930 736 1932 744
rect 1940 736 1942 744
rect 1930 734 1942 736
rect 1496 406 1500 414
rect 1508 406 1516 414
rect 1524 406 1532 414
rect 1540 406 1544 414
rect 522 116 524 124
rect 532 116 534 124
rect 522 114 534 116
rect 970 164 982 166
rect 970 156 972 164
rect 980 156 982 164
rect 970 124 982 156
rect 970 116 972 124
rect 980 116 982 124
rect 970 114 982 116
rect 1496 14 1544 406
rect 2058 584 2070 1316
rect 2058 576 2060 584
rect 2068 576 2070 584
rect 2058 284 2070 576
rect 2154 544 2166 1696
rect 2154 536 2156 544
rect 2164 536 2166 544
rect 2154 534 2166 536
rect 2570 1204 2582 1206
rect 2570 1196 2572 1204
rect 2580 1196 2582 1204
rect 2570 304 2582 1196
rect 2858 1144 2870 1796
rect 2858 1136 2860 1144
rect 2868 1136 2870 1144
rect 2858 1134 2870 1136
rect 3032 1814 3080 2206
rect 3114 2224 3126 2226
rect 3114 2216 3116 2224
rect 3124 2216 3126 2224
rect 3114 2024 3126 2216
rect 3210 2044 3222 2296
rect 3210 2036 3212 2044
rect 3220 2036 3222 2044
rect 3210 2034 3222 2036
rect 3402 2304 3414 2306
rect 3402 2296 3404 2304
rect 3412 2296 3414 2304
rect 3114 2016 3116 2024
rect 3124 2016 3126 2024
rect 3114 2014 3126 2016
rect 3178 1964 3190 1966
rect 3178 1956 3180 1964
rect 3188 1956 3190 1964
rect 3032 1806 3036 1814
rect 3044 1806 3052 1814
rect 3060 1806 3068 1814
rect 3076 1806 3080 1814
rect 3032 1414 3080 1806
rect 3114 1904 3126 1906
rect 3114 1896 3116 1904
rect 3124 1896 3126 1904
rect 3114 1504 3126 1896
rect 3178 1764 3190 1956
rect 3178 1756 3180 1764
rect 3188 1756 3190 1764
rect 3178 1754 3190 1756
rect 3402 1704 3414 2296
rect 3498 2244 3510 2596
rect 3530 2424 3542 3056
rect 3658 2884 3670 2886
rect 3658 2876 3660 2884
rect 3668 2876 3670 2884
rect 3626 2864 3638 2866
rect 3626 2856 3628 2864
rect 3636 2856 3638 2864
rect 3530 2416 3532 2424
rect 3540 2416 3542 2424
rect 3530 2414 3542 2416
rect 3594 2764 3606 2766
rect 3594 2756 3596 2764
rect 3604 2756 3606 2764
rect 3594 2644 3606 2756
rect 3594 2636 3596 2644
rect 3604 2636 3606 2644
rect 3594 2304 3606 2636
rect 3626 2604 3638 2856
rect 3658 2724 3670 2876
rect 3658 2716 3660 2724
rect 3668 2716 3670 2724
rect 3658 2714 3670 2716
rect 3626 2596 3628 2604
rect 3636 2596 3638 2604
rect 3626 2594 3638 2596
rect 3722 2644 3734 2646
rect 3722 2636 3724 2644
rect 3732 2636 3734 2644
rect 3594 2296 3596 2304
rect 3604 2296 3606 2304
rect 3594 2294 3606 2296
rect 3658 2544 3670 2546
rect 3658 2536 3660 2544
rect 3668 2536 3670 2544
rect 3658 2264 3670 2536
rect 3658 2256 3660 2264
rect 3668 2256 3670 2264
rect 3658 2254 3670 2256
rect 3498 2236 3500 2244
rect 3508 2236 3510 2244
rect 3498 2234 3510 2236
rect 3466 2044 3478 2046
rect 3466 2036 3468 2044
rect 3476 2036 3478 2044
rect 3434 1944 3446 1946
rect 3434 1936 3436 1944
rect 3444 1936 3446 1944
rect 3434 1824 3446 1936
rect 3466 1904 3478 2036
rect 3466 1896 3468 1904
rect 3476 1896 3478 1904
rect 3466 1894 3478 1896
rect 3434 1816 3436 1824
rect 3444 1816 3446 1824
rect 3434 1814 3446 1816
rect 3402 1696 3404 1704
rect 3412 1696 3414 1704
rect 3402 1694 3414 1696
rect 3114 1496 3116 1504
rect 3124 1496 3126 1504
rect 3114 1494 3126 1496
rect 3032 1406 3036 1414
rect 3044 1406 3052 1414
rect 3060 1406 3068 1414
rect 3076 1406 3080 1414
rect 2954 1084 2966 1086
rect 2954 1076 2956 1084
rect 2964 1076 2966 1084
rect 2954 944 2966 1076
rect 2954 936 2956 944
rect 2964 936 2966 944
rect 2954 934 2966 936
rect 3032 1014 3080 1406
rect 3690 1404 3702 1406
rect 3690 1396 3692 1404
rect 3700 1396 3702 1404
rect 3032 1006 3036 1014
rect 3044 1006 3052 1014
rect 3060 1006 3068 1014
rect 3076 1006 3080 1014
rect 2570 296 2572 304
rect 2580 296 2582 304
rect 2570 294 2582 296
rect 3032 614 3080 1006
rect 3338 1324 3350 1326
rect 3338 1316 3340 1324
rect 3348 1316 3350 1324
rect 3338 984 3350 1316
rect 3690 1144 3702 1396
rect 3722 1284 3734 2636
rect 3786 2644 3798 3076
rect 3914 3084 3926 3086
rect 3914 3076 3916 3084
rect 3924 3076 3926 3084
rect 3914 2944 3926 3076
rect 4042 3044 4054 3096
rect 4042 3036 4044 3044
rect 4052 3036 4054 3044
rect 4042 3034 4054 3036
rect 3914 2936 3916 2944
rect 3924 2936 3926 2944
rect 3914 2934 3926 2936
rect 4010 3024 4022 3026
rect 4010 3016 4012 3024
rect 4020 3016 4022 3024
rect 3946 2904 3958 2906
rect 3946 2896 3948 2904
rect 3956 2896 3958 2904
rect 3818 2884 3830 2886
rect 3818 2876 3820 2884
rect 3828 2876 3830 2884
rect 3818 2764 3830 2876
rect 3818 2756 3820 2764
rect 3828 2756 3830 2764
rect 3818 2754 3830 2756
rect 3946 2684 3958 2896
rect 4010 2784 4022 3016
rect 4010 2776 4012 2784
rect 4020 2776 4022 2784
rect 4010 2774 4022 2776
rect 4042 2864 4054 2866
rect 4042 2856 4044 2864
rect 4052 2856 4054 2864
rect 3946 2676 3948 2684
rect 3956 2676 3958 2684
rect 3946 2674 3958 2676
rect 3786 2636 3788 2644
rect 3796 2636 3798 2644
rect 3786 2634 3798 2636
rect 4042 2364 4054 2856
rect 4042 2356 4044 2364
rect 4052 2356 4054 2364
rect 4042 2354 4054 2356
rect 4074 2364 4086 2366
rect 4074 2356 4076 2364
rect 4084 2356 4086 2364
rect 3818 2284 3830 2286
rect 3818 2276 3820 2284
rect 3828 2276 3830 2284
rect 3818 2224 3830 2276
rect 3818 2216 3820 2224
rect 3828 2216 3830 2224
rect 3818 2214 3830 2216
rect 3722 1276 3724 1284
rect 3732 1276 3734 1284
rect 3722 1274 3734 1276
rect 3818 2104 3830 2106
rect 3818 2096 3820 2104
rect 3828 2096 3830 2104
rect 3818 1704 3830 2096
rect 4074 1844 4086 2356
rect 4138 2304 4150 3536
rect 4490 3304 4502 3306
rect 4490 3296 4492 3304
rect 4500 3296 4502 3304
rect 4490 3084 4502 3296
rect 4490 3076 4492 3084
rect 4500 3076 4502 3084
rect 4490 3074 4502 3076
rect 4568 3214 4616 3606
rect 4568 3206 4572 3214
rect 4580 3206 4588 3214
rect 4596 3206 4604 3214
rect 4612 3206 4616 3214
rect 4746 3804 4758 3806
rect 4746 3796 4748 3804
rect 4756 3796 4758 3804
rect 4170 3064 4182 3066
rect 4170 3056 4172 3064
rect 4180 3056 4182 3064
rect 4170 2964 4182 3056
rect 4170 2956 4172 2964
rect 4180 2956 4182 2964
rect 4170 2624 4182 2956
rect 4298 2884 4310 2886
rect 4298 2876 4300 2884
rect 4308 2876 4310 2884
rect 4170 2616 4172 2624
rect 4180 2616 4182 2624
rect 4170 2424 4182 2616
rect 4202 2664 4214 2666
rect 4202 2656 4204 2664
rect 4212 2656 4214 2664
rect 4202 2504 4214 2656
rect 4298 2564 4310 2876
rect 4568 2814 4616 3206
rect 4650 3204 4662 3206
rect 4650 3196 4652 3204
rect 4660 3196 4662 3204
rect 4650 3144 4662 3196
rect 4650 3136 4652 3144
rect 4660 3136 4662 3144
rect 4650 3134 4662 3136
rect 4568 2806 4572 2814
rect 4580 2806 4588 2814
rect 4596 2806 4604 2814
rect 4612 2806 4616 2814
rect 4330 2804 4342 2806
rect 4330 2796 4332 2804
rect 4340 2796 4342 2804
rect 4330 2624 4342 2796
rect 4330 2616 4332 2624
rect 4340 2616 4342 2624
rect 4330 2614 4342 2616
rect 4298 2556 4300 2564
rect 4308 2556 4310 2564
rect 4298 2554 4310 2556
rect 4202 2496 4204 2504
rect 4212 2496 4214 2504
rect 4202 2494 4214 2496
rect 4170 2416 4172 2424
rect 4180 2416 4182 2424
rect 4170 2414 4182 2416
rect 4234 2444 4246 2446
rect 4234 2436 4236 2444
rect 4244 2436 4246 2444
rect 4234 2404 4246 2436
rect 4234 2396 4236 2404
rect 4244 2396 4246 2404
rect 4234 2394 4246 2396
rect 4568 2414 4616 2806
rect 4682 3104 4694 3106
rect 4682 3096 4684 3104
rect 4692 3096 4694 3104
rect 4682 2644 4694 3096
rect 4682 2636 4684 2644
rect 4692 2636 4694 2644
rect 4682 2634 4694 2636
rect 4746 2644 4758 3796
rect 4906 3544 4918 4036
rect 4906 3536 4908 3544
rect 4916 3536 4918 3544
rect 4906 3534 4918 3536
rect 4938 3324 4950 3326
rect 4938 3316 4940 3324
rect 4948 3316 4950 3324
rect 4938 3064 4950 3316
rect 5098 3224 5110 3226
rect 5098 3216 5100 3224
rect 5108 3216 5110 3224
rect 5034 3144 5046 3146
rect 5034 3136 5036 3144
rect 5044 3136 5046 3144
rect 4938 3056 4940 3064
rect 4948 3056 4950 3064
rect 4938 3054 4950 3056
rect 5002 3104 5014 3106
rect 5002 3096 5004 3104
rect 5012 3096 5014 3104
rect 5002 3024 5014 3096
rect 5034 3084 5046 3136
rect 5034 3076 5036 3084
rect 5044 3076 5046 3084
rect 5034 3074 5046 3076
rect 5066 3124 5078 3126
rect 5066 3116 5068 3124
rect 5076 3116 5078 3124
rect 5002 3016 5004 3024
rect 5012 3016 5014 3024
rect 5002 3014 5014 3016
rect 5066 2984 5078 3116
rect 5066 2976 5068 2984
rect 5076 2976 5078 2984
rect 5066 2974 5078 2976
rect 4842 2944 4854 2946
rect 4842 2936 4844 2944
rect 4852 2936 4854 2944
rect 4746 2636 4748 2644
rect 4756 2636 4758 2644
rect 4746 2634 4758 2636
rect 4778 2824 4790 2826
rect 4778 2816 4780 2824
rect 4788 2816 4790 2824
rect 4778 2604 4790 2816
rect 4778 2596 4780 2604
rect 4788 2596 4790 2604
rect 4778 2594 4790 2596
rect 4842 2504 4854 2936
rect 5066 2944 5078 2946
rect 5066 2936 5068 2944
rect 5076 2936 5078 2944
rect 4874 2644 4886 2646
rect 4874 2636 4876 2644
rect 4884 2636 4886 2644
rect 4874 2544 4886 2636
rect 4874 2536 4876 2544
rect 4884 2536 4886 2544
rect 4874 2534 4886 2536
rect 5034 2644 5046 2646
rect 5034 2636 5036 2644
rect 5044 2636 5046 2644
rect 4842 2496 4844 2504
rect 4852 2496 4854 2504
rect 4842 2494 4854 2496
rect 4568 2406 4572 2414
rect 4580 2406 4588 2414
rect 4596 2406 4604 2414
rect 4612 2406 4616 2414
rect 4138 2296 4140 2304
rect 4148 2296 4150 2304
rect 4138 2294 4150 2296
rect 4568 2014 4616 2406
rect 4650 2444 4662 2446
rect 4650 2436 4652 2444
rect 4660 2436 4662 2444
rect 4650 2244 4662 2436
rect 5034 2444 5046 2636
rect 5066 2644 5078 2936
rect 5098 2944 5110 3216
rect 5194 3224 5206 4656
rect 5194 3216 5196 3224
rect 5204 3216 5206 3224
rect 5194 3214 5206 3216
rect 5226 4424 5238 4426
rect 5226 4416 5228 4424
rect 5236 4416 5238 4424
rect 5226 3124 5238 4416
rect 5354 4384 5366 4386
rect 5354 4376 5356 4384
rect 5364 4376 5366 4384
rect 5290 3464 5302 3466
rect 5290 3456 5292 3464
rect 5300 3456 5302 3464
rect 5290 3324 5302 3456
rect 5290 3316 5292 3324
rect 5300 3316 5302 3324
rect 5290 3314 5302 3316
rect 5354 3224 5366 4376
rect 5386 3624 5398 3626
rect 5386 3616 5388 3624
rect 5396 3616 5398 3624
rect 5386 3344 5398 3616
rect 5418 3584 5430 5176
rect 5578 4944 5590 5436
rect 5578 4936 5580 4944
rect 5588 4936 5590 4944
rect 5578 4934 5590 4936
rect 5610 5344 5622 5346
rect 5610 5336 5612 5344
rect 5620 5336 5622 5344
rect 5418 3576 5420 3584
rect 5428 3576 5430 3584
rect 5418 3574 5430 3576
rect 5450 4764 5462 4766
rect 5450 4756 5452 4764
rect 5460 4756 5462 4764
rect 5386 3336 5388 3344
rect 5396 3336 5398 3344
rect 5386 3334 5398 3336
rect 5354 3216 5356 3224
rect 5364 3216 5366 3224
rect 5354 3214 5366 3216
rect 5226 3116 5228 3124
rect 5236 3116 5238 3124
rect 5226 3114 5238 3116
rect 5386 3064 5398 3066
rect 5386 3056 5388 3064
rect 5396 3056 5398 3064
rect 5098 2936 5100 2944
rect 5108 2936 5110 2944
rect 5098 2934 5110 2936
rect 5194 2964 5206 2966
rect 5194 2956 5196 2964
rect 5204 2956 5206 2964
rect 5130 2844 5142 2846
rect 5130 2836 5132 2844
rect 5140 2836 5142 2844
rect 5066 2636 5068 2644
rect 5076 2636 5078 2644
rect 5066 2634 5078 2636
rect 5098 2684 5110 2686
rect 5098 2676 5100 2684
rect 5108 2676 5110 2684
rect 5098 2524 5110 2676
rect 5098 2516 5100 2524
rect 5108 2516 5110 2524
rect 5098 2514 5110 2516
rect 5034 2436 5036 2444
rect 5044 2436 5046 2444
rect 5034 2434 5046 2436
rect 4682 2424 4694 2426
rect 4682 2416 4684 2424
rect 4692 2416 4694 2424
rect 4682 2284 4694 2416
rect 4714 2424 4726 2426
rect 4714 2416 4716 2424
rect 4724 2416 4726 2424
rect 4714 2324 4726 2416
rect 4714 2316 4716 2324
rect 4724 2316 4726 2324
rect 4714 2314 4726 2316
rect 4682 2276 4684 2284
rect 4692 2276 4694 2284
rect 4682 2274 4694 2276
rect 4650 2236 4652 2244
rect 4660 2236 4662 2244
rect 4650 2234 4662 2236
rect 5130 2104 5142 2836
rect 5194 2764 5206 2956
rect 5194 2756 5196 2764
rect 5204 2756 5206 2764
rect 5194 2704 5206 2756
rect 5194 2696 5196 2704
rect 5204 2696 5206 2704
rect 5194 2694 5206 2696
rect 5290 2764 5302 2766
rect 5290 2756 5292 2764
rect 5300 2756 5302 2764
rect 5258 2664 5270 2666
rect 5258 2656 5260 2664
rect 5268 2656 5270 2664
rect 5258 2544 5270 2656
rect 5290 2564 5302 2756
rect 5290 2556 5292 2564
rect 5300 2556 5302 2564
rect 5290 2554 5302 2556
rect 5258 2536 5260 2544
rect 5268 2536 5270 2544
rect 5258 2534 5270 2536
rect 5322 2544 5334 2546
rect 5322 2536 5324 2544
rect 5332 2536 5334 2544
rect 5322 2364 5334 2536
rect 5386 2444 5398 3056
rect 5418 3024 5430 3026
rect 5418 3016 5420 3024
rect 5428 3016 5430 3024
rect 5418 2684 5430 3016
rect 5418 2676 5420 2684
rect 5428 2676 5430 2684
rect 5418 2674 5430 2676
rect 5386 2436 5388 2444
rect 5396 2436 5398 2444
rect 5386 2434 5398 2436
rect 5322 2356 5324 2364
rect 5332 2356 5334 2364
rect 5322 2324 5334 2356
rect 5322 2316 5324 2324
rect 5332 2316 5334 2324
rect 5322 2314 5334 2316
rect 5130 2096 5132 2104
rect 5140 2096 5142 2104
rect 5130 2094 5142 2096
rect 4568 2006 4572 2014
rect 4580 2006 4588 2014
rect 4596 2006 4604 2014
rect 4612 2006 4616 2014
rect 4074 1836 4076 1844
rect 4084 1836 4086 1844
rect 4074 1834 4086 1836
rect 4106 1984 4118 1986
rect 4106 1976 4108 1984
rect 4116 1976 4118 1984
rect 3818 1696 3820 1704
rect 3828 1696 3830 1704
rect 3690 1136 3692 1144
rect 3700 1136 3702 1144
rect 3690 1134 3702 1136
rect 3818 1064 3830 1696
rect 3818 1056 3820 1064
rect 3828 1056 3830 1064
rect 3818 1054 3830 1056
rect 4042 1304 4054 1306
rect 4042 1296 4044 1304
rect 4052 1296 4054 1304
rect 3338 976 3340 984
rect 3348 976 3350 984
rect 3338 974 3350 976
rect 4010 1024 4022 1026
rect 4010 1016 4012 1024
rect 4020 1016 4022 1024
rect 3594 944 3606 946
rect 3594 936 3596 944
rect 3604 936 3606 944
rect 3032 606 3036 614
rect 3044 606 3052 614
rect 3060 606 3068 614
rect 3076 606 3080 614
rect 2058 276 2060 284
rect 2068 276 2070 284
rect 2058 274 2070 276
rect 2826 284 2838 286
rect 2826 276 2828 284
rect 2836 276 2838 284
rect 2826 144 2838 276
rect 2826 136 2828 144
rect 2836 136 2838 144
rect 2826 134 2838 136
rect 3032 214 3080 606
rect 3178 764 3190 766
rect 3178 756 3180 764
rect 3188 756 3190 764
rect 3178 284 3190 756
rect 3594 544 3606 936
rect 3594 536 3596 544
rect 3604 536 3606 544
rect 3594 534 3606 536
rect 3658 924 3670 926
rect 3658 916 3660 924
rect 3668 916 3670 924
rect 3658 524 3670 916
rect 3946 744 3958 746
rect 3946 736 3948 744
rect 3956 736 3958 744
rect 3658 516 3660 524
rect 3668 516 3670 524
rect 3658 514 3670 516
rect 3818 564 3830 566
rect 3818 556 3820 564
rect 3828 556 3830 564
rect 3178 276 3180 284
rect 3188 276 3190 284
rect 3178 274 3190 276
rect 3818 284 3830 556
rect 3946 544 3958 736
rect 4010 624 4022 1016
rect 4010 616 4012 624
rect 4020 616 4022 624
rect 4010 614 4022 616
rect 3946 536 3948 544
rect 3956 536 3958 544
rect 3946 534 3958 536
rect 3818 276 3820 284
rect 3828 276 3830 284
rect 3818 274 3830 276
rect 3032 206 3036 214
rect 3044 206 3052 214
rect 3060 206 3068 214
rect 3076 206 3080 214
rect 1496 6 1500 14
rect 1508 6 1516 14
rect 1524 6 1532 14
rect 1540 6 1544 14
rect 1496 -40 1544 6
rect 3032 -40 3080 206
rect 4042 184 4054 1296
rect 4074 1084 4086 1086
rect 4074 1076 4076 1084
rect 4084 1076 4086 1084
rect 4074 364 4086 1076
rect 4106 1084 4118 1976
rect 4568 1614 4616 2006
rect 5066 1964 5078 1966
rect 5066 1956 5068 1964
rect 5076 1956 5078 1964
rect 4810 1944 4822 1946
rect 4810 1936 4812 1944
rect 4820 1936 4822 1944
rect 4568 1606 4572 1614
rect 4580 1606 4588 1614
rect 4596 1606 4604 1614
rect 4612 1606 4616 1614
rect 4490 1524 4502 1526
rect 4490 1516 4492 1524
rect 4500 1516 4502 1524
rect 4426 1184 4438 1186
rect 4426 1176 4428 1184
rect 4436 1176 4438 1184
rect 4106 1076 4108 1084
rect 4116 1076 4118 1084
rect 4106 1074 4118 1076
rect 4298 1144 4310 1146
rect 4298 1136 4300 1144
rect 4308 1136 4310 1144
rect 4106 1024 4118 1026
rect 4106 1016 4108 1024
rect 4116 1016 4118 1024
rect 4106 704 4118 1016
rect 4298 924 4310 1136
rect 4298 916 4300 924
rect 4308 916 4310 924
rect 4298 914 4310 916
rect 4362 924 4374 926
rect 4362 916 4364 924
rect 4372 916 4374 924
rect 4362 784 4374 916
rect 4426 924 4438 1176
rect 4490 1184 4502 1516
rect 4490 1176 4492 1184
rect 4500 1176 4502 1184
rect 4426 916 4428 924
rect 4436 916 4438 924
rect 4426 914 4438 916
rect 4458 1124 4470 1126
rect 4458 1116 4460 1124
rect 4468 1116 4470 1124
rect 4362 776 4364 784
rect 4372 776 4374 784
rect 4362 774 4374 776
rect 4458 724 4470 1116
rect 4490 924 4502 1176
rect 4490 916 4492 924
rect 4500 916 4502 924
rect 4490 914 4502 916
rect 4568 1214 4616 1606
rect 4682 1904 4694 1906
rect 4682 1896 4684 1904
rect 4692 1896 4694 1904
rect 4682 1264 4694 1896
rect 4810 1504 4822 1936
rect 5034 1724 5046 1726
rect 5034 1716 5036 1724
rect 5044 1716 5046 1724
rect 4810 1496 4812 1504
rect 4820 1496 4822 1504
rect 4810 1494 4822 1496
rect 4842 1684 4854 1686
rect 4842 1676 4844 1684
rect 4852 1676 4854 1684
rect 4842 1584 4854 1676
rect 4842 1576 4844 1584
rect 4852 1576 4854 1584
rect 4682 1256 4684 1264
rect 4692 1256 4694 1264
rect 4682 1254 4694 1256
rect 4568 1206 4572 1214
rect 4580 1206 4588 1214
rect 4596 1206 4604 1214
rect 4612 1206 4616 1214
rect 4458 716 4460 724
rect 4468 716 4470 724
rect 4458 714 4470 716
rect 4568 814 4616 1206
rect 4842 984 4854 1576
rect 5034 1364 5046 1716
rect 5034 1356 5036 1364
rect 5044 1356 5046 1364
rect 5034 1354 5046 1356
rect 5066 1364 5078 1956
rect 5066 1356 5068 1364
rect 5076 1356 5078 1364
rect 5066 1354 5078 1356
rect 5098 1924 5110 1926
rect 5098 1916 5100 1924
rect 5108 1916 5110 1924
rect 5098 1244 5110 1916
rect 5226 1844 5238 1846
rect 5226 1836 5228 1844
rect 5236 1836 5238 1844
rect 5194 1824 5206 1826
rect 5194 1816 5196 1824
rect 5204 1816 5206 1824
rect 5194 1284 5206 1816
rect 5226 1444 5238 1836
rect 5226 1436 5228 1444
rect 5236 1436 5238 1444
rect 5226 1434 5238 1436
rect 5194 1276 5196 1284
rect 5204 1276 5206 1284
rect 5194 1274 5206 1276
rect 5098 1236 5100 1244
rect 5108 1236 5110 1244
rect 5098 1234 5110 1236
rect 5034 1224 5046 1226
rect 5034 1216 5036 1224
rect 5044 1216 5046 1224
rect 5034 1144 5046 1216
rect 5034 1136 5036 1144
rect 5044 1136 5046 1144
rect 5034 1134 5046 1136
rect 5066 1224 5078 1226
rect 5066 1216 5068 1224
rect 5076 1216 5078 1224
rect 4842 976 4844 984
rect 4852 976 4854 984
rect 4842 974 4854 976
rect 5066 984 5078 1216
rect 5066 976 5068 984
rect 5076 976 5078 984
rect 5066 974 5078 976
rect 5418 1184 5430 1186
rect 5418 1176 5420 1184
rect 5428 1176 5430 1184
rect 4568 806 4572 814
rect 4580 806 4588 814
rect 4596 806 4604 814
rect 4612 806 4616 814
rect 4106 696 4108 704
rect 4116 696 4118 704
rect 4106 694 4118 696
rect 4074 356 4076 364
rect 4084 356 4086 364
rect 4074 284 4086 356
rect 4074 276 4076 284
rect 4084 276 4086 284
rect 4074 274 4086 276
rect 4568 414 4616 806
rect 4650 824 4662 826
rect 4650 816 4652 824
rect 4660 816 4662 824
rect 4650 564 4662 816
rect 5418 744 5430 1176
rect 5418 736 5420 744
rect 5428 736 5430 744
rect 5418 734 5430 736
rect 4650 556 4652 564
rect 4660 556 4662 564
rect 4650 554 4662 556
rect 5162 684 5174 686
rect 5162 676 5164 684
rect 5172 676 5174 684
rect 4568 406 4572 414
rect 4580 406 4588 414
rect 4596 406 4604 414
rect 4612 406 4616 414
rect 4042 176 4044 184
rect 4052 176 4054 184
rect 4042 174 4054 176
rect 4568 14 4616 406
rect 5034 404 5046 406
rect 5034 396 5036 404
rect 5044 396 5046 404
rect 5034 104 5046 396
rect 5162 344 5174 676
rect 5162 336 5164 344
rect 5172 336 5174 344
rect 5162 334 5174 336
rect 5450 144 5462 4756
rect 5610 4244 5622 5336
rect 5898 5304 5910 5306
rect 5898 5296 5900 5304
rect 5908 5296 5910 5304
rect 5834 4604 5846 4606
rect 5834 4596 5836 4604
rect 5844 4596 5846 4604
rect 5610 4236 5612 4244
rect 5620 4236 5622 4244
rect 5610 4234 5622 4236
rect 5738 4424 5750 4426
rect 5738 4416 5740 4424
rect 5748 4416 5750 4424
rect 5738 3884 5750 4416
rect 5738 3876 5740 3884
rect 5748 3876 5750 3884
rect 5738 3874 5750 3876
rect 5546 3324 5558 3326
rect 5546 3316 5548 3324
rect 5556 3316 5558 3324
rect 5546 2924 5558 3316
rect 5546 2916 5548 2924
rect 5556 2916 5558 2924
rect 5546 2914 5558 2916
rect 5578 3224 5590 3226
rect 5578 3216 5580 3224
rect 5588 3216 5590 3224
rect 5578 2744 5590 3216
rect 5834 3144 5846 4596
rect 5898 4524 5910 5296
rect 5994 5264 6006 5266
rect 5994 5256 5996 5264
rect 6004 5256 6006 5264
rect 5898 4516 5900 4524
rect 5908 4516 5910 4524
rect 5898 4514 5910 4516
rect 5930 4524 5942 4526
rect 5930 4516 5932 4524
rect 5940 4516 5942 4524
rect 5898 4144 5910 4146
rect 5898 4136 5900 4144
rect 5908 4136 5910 4144
rect 5898 3724 5910 4136
rect 5898 3716 5900 3724
rect 5908 3716 5910 3724
rect 5898 3714 5910 3716
rect 5834 3136 5836 3144
rect 5844 3136 5846 3144
rect 5834 3134 5846 3136
rect 5866 3144 5878 3146
rect 5866 3136 5868 3144
rect 5876 3136 5878 3144
rect 5578 2736 5580 2744
rect 5588 2736 5590 2744
rect 5578 2734 5590 2736
rect 5802 2944 5814 2946
rect 5802 2936 5804 2944
rect 5812 2936 5814 2944
rect 5482 2664 5494 2666
rect 5482 2656 5484 2664
rect 5492 2656 5494 2664
rect 5482 2324 5494 2656
rect 5482 2316 5484 2324
rect 5492 2316 5494 2324
rect 5482 2314 5494 2316
rect 5514 2444 5526 2446
rect 5514 2436 5516 2444
rect 5524 2436 5526 2444
rect 5450 136 5452 144
rect 5460 136 5462 144
rect 5450 134 5462 136
rect 5034 96 5036 104
rect 5044 96 5046 104
rect 5034 94 5046 96
rect 5514 104 5526 2436
rect 5738 2384 5750 2386
rect 5738 2376 5740 2384
rect 5748 2376 5750 2384
rect 5642 2104 5654 2106
rect 5642 2096 5644 2104
rect 5652 2096 5654 2104
rect 5642 1684 5654 2096
rect 5642 1676 5644 1684
rect 5652 1676 5654 1684
rect 5642 1674 5654 1676
rect 5674 2044 5686 2046
rect 5674 2036 5676 2044
rect 5684 2036 5686 2044
rect 5674 1084 5686 2036
rect 5738 1864 5750 2376
rect 5738 1856 5740 1864
rect 5748 1856 5750 1864
rect 5738 1854 5750 1856
rect 5802 1824 5814 2936
rect 5866 2384 5878 3136
rect 5930 2944 5942 4516
rect 5994 4004 6006 5256
rect 5994 3996 5996 4004
rect 6004 3996 6006 4004
rect 5994 3994 6006 3996
rect 6026 4844 6038 4846
rect 6026 4836 6028 4844
rect 6036 4836 6038 4844
rect 5930 2936 5932 2944
rect 5940 2936 5942 2944
rect 5930 2934 5942 2936
rect 6026 2684 6038 4836
rect 6090 3344 6102 5596
rect 6090 3336 6092 3344
rect 6100 3336 6102 3344
rect 6090 3334 6102 3336
rect 6026 2676 6028 2684
rect 6036 2676 6038 2684
rect 6026 2674 6038 2676
rect 5866 2376 5868 2384
rect 5876 2376 5878 2384
rect 5866 2374 5878 2376
rect 5802 1816 5804 1824
rect 5812 1816 5814 1824
rect 5802 1814 5814 1816
rect 5866 2324 5878 2326
rect 5866 2316 5868 2324
rect 5876 2316 5878 2324
rect 5802 1764 5814 1766
rect 5802 1756 5804 1764
rect 5812 1756 5814 1764
rect 5706 1444 5718 1446
rect 5706 1436 5708 1444
rect 5716 1436 5718 1444
rect 5706 1104 5718 1436
rect 5706 1096 5708 1104
rect 5716 1096 5718 1104
rect 5706 1094 5718 1096
rect 5674 1076 5676 1084
rect 5684 1076 5686 1084
rect 5674 1074 5686 1076
rect 5706 1044 5718 1046
rect 5706 1036 5708 1044
rect 5716 1036 5718 1044
rect 5546 704 5558 706
rect 5546 696 5548 704
rect 5556 696 5558 704
rect 5546 524 5558 696
rect 5546 516 5548 524
rect 5556 516 5558 524
rect 5546 514 5558 516
rect 5706 344 5718 1036
rect 5802 464 5814 1756
rect 5866 1484 5878 2316
rect 6026 2304 6038 2306
rect 6026 2296 6028 2304
rect 6036 2296 6038 2304
rect 5866 1476 5868 1484
rect 5876 1476 5878 1484
rect 5866 1474 5878 1476
rect 5898 1984 5910 1986
rect 5898 1976 5900 1984
rect 5908 1976 5910 1984
rect 5802 456 5804 464
rect 5812 456 5814 464
rect 5802 454 5814 456
rect 5834 1204 5846 1206
rect 5834 1196 5836 1204
rect 5844 1196 5846 1204
rect 5706 336 5708 344
rect 5716 336 5718 344
rect 5706 334 5718 336
rect 5514 96 5516 104
rect 5524 96 5526 104
rect 5514 94 5526 96
rect 5674 144 5686 146
rect 5674 136 5676 144
rect 5684 136 5686 144
rect 5674 24 5686 136
rect 5834 124 5846 1196
rect 5898 1184 5910 1976
rect 5898 1176 5900 1184
rect 5908 1176 5910 1184
rect 5898 1174 5910 1176
rect 5962 1604 5974 1606
rect 5962 1596 5964 1604
rect 5972 1596 5974 1604
rect 5866 984 5878 986
rect 5866 976 5868 984
rect 5876 976 5878 984
rect 5866 684 5878 976
rect 5962 984 5974 1596
rect 6026 1344 6038 2296
rect 6026 1336 6028 1344
rect 6036 1336 6038 1344
rect 6026 1334 6038 1336
rect 6090 1884 6102 1886
rect 6090 1876 6092 1884
rect 6100 1876 6102 1884
rect 5962 976 5964 984
rect 5972 976 5974 984
rect 5962 974 5974 976
rect 6026 1184 6038 1186
rect 6026 1176 6028 1184
rect 6036 1176 6038 1184
rect 6026 984 6038 1176
rect 6026 976 6028 984
rect 6036 976 6038 984
rect 6026 974 6038 976
rect 5866 676 5868 684
rect 5876 676 5878 684
rect 5866 674 5878 676
rect 6090 424 6102 1876
rect 6090 416 6092 424
rect 6100 416 6102 424
rect 6090 414 6102 416
rect 5834 116 5836 124
rect 5844 116 5846 124
rect 5834 114 5846 116
rect 5674 16 5676 24
rect 5684 16 5686 24
rect 5674 14 5686 16
rect 4568 6 4572 14
rect 4580 6 4588 14
rect 4596 6 4604 14
rect 4612 6 4616 14
rect 4568 -40 4616 6
use DFFSR  DFFSR_81
timestamp 1743498307
transform 1 0 8 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_362
timestamp 1743498307
transform 1 0 360 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_22
timestamp 1743498307
transform -1 0 56 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_83
timestamp 1743498307
transform 1 0 56 0 1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_363
timestamp 1743498307
transform -1 0 488 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_102
timestamp 1743498307
transform -1 0 520 0 -1 210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1743498307
transform 1 0 520 0 -1 210
box -4 -6 196 206
use BUFX4  BUFX4_72
timestamp 1743498307
transform -1 0 776 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_367
timestamp 1743498307
transform -1 0 472 0 1 210
box -4 -6 68 206
use INVX1  INVX1_104
timestamp 1743498307
transform -1 0 504 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_44
timestamp 1743498307
transform 1 0 504 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_45
timestamp 1743498307
transform -1 0 632 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1743498307
transform -1 0 824 0 1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_35
timestamp 1743498307
transform 1 0 776 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_34
timestamp 1743498307
transform -1 0 904 0 -1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_18
timestamp 1743498307
transform -1 0 1096 0 -1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_41
timestamp 1743498307
transform 1 0 824 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_40
timestamp 1743498307
transform -1 0 952 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1743498307
transform 1 0 952 0 1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_26
timestamp 1743498307
transform -1 0 1272 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_27
timestamp 1743498307
transform 1 0 1144 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_28
timestamp 1743498307
transform -1 0 1400 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_29
timestamp 1743498307
transform 1 0 1272 0 1 210
box -4 -6 68 206
use FILL  FILL_0_0_2
timestamp 1743498307
transform -1 0 1448 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1743498307
transform -1 0 1432 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1743498307
transform -1 0 1416 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_7
timestamp 1743498307
transform -1 0 1400 0 -1 210
box -4 -6 52 206
use BUFX4  BUFX4_75
timestamp 1743498307
transform -1 0 1352 0 -1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1743498307
transform -1 0 1592 0 1 210
box -4 -6 196 206
use DFFSR  DFFSR_78
timestamp 1743498307
transform -1 0 1800 0 -1 210
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1743498307
transform -1 0 1288 0 -1 210
box -4 -6 196 206
use DFFSR  DFFSR_77
timestamp 1743498307
transform 1 0 1800 0 -1 210
box -4 -6 356 206
use FILL  FILL_1_0_0
timestamp 1743498307
transform 1 0 1592 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1743498307
transform 1 0 1608 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1743498307
transform 1 0 1624 0 1 210
box -4 -6 20 206
use INVX1  INVX1_99
timestamp 1743498307
transform 1 0 1640 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_359
timestamp 1743498307
transform 1 0 1672 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_115
timestamp 1743498307
transform -1 0 1784 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_90
timestamp 1743498307
transform -1 0 2136 0 1 210
box -4 -6 356 206
use BUFX2  BUFX2_6
timestamp 1743498307
transform 1 0 2152 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_98
timestamp 1743498307
transform -1 0 2168 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_358
timestamp 1743498307
transform -1 0 2232 0 1 210
box -4 -6 68 206
use DFFSR  DFFSR_80
timestamp 1743498307
transform 1 0 2200 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_361
timestamp 1743498307
transform -1 0 2296 0 1 210
box -4 -6 68 206
use INVX1  INVX1_101
timestamp 1743498307
transform -1 0 2328 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_92
timestamp 1743498307
transform 1 0 2328 0 1 210
box -4 -6 356 206
use BUFX2  BUFX2_9
timestamp 1743498307
transform 1 0 2552 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1743498307
transform 1 0 2600 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_11
timestamp 1743498307
transform 1 0 2648 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_94
timestamp 1743498307
transform 1 0 2696 0 -1 210
box -4 -6 356 206
use INVX1  INVX1_111
timestamp 1743498307
transform 1 0 2680 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_34
timestamp 1743498307
transform 1 0 2712 0 1 210
box -4 -6 356 206
use FILL  FILL_1_1_0
timestamp 1743498307
transform 1 0 3064 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1743498307
transform 1 0 3064 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1743498307
transform 1 0 3048 0 -1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_4
timestamp 1743498307
transform -1 0 3256 0 1 210
box -4 -6 116 206
use INVX1  INVX1_113
timestamp 1743498307
transform 1 0 3112 0 1 210
box -4 -6 36 206
use FILL  FILL_1_1_2
timestamp 1743498307
transform 1 0 3096 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1743498307
transform 1 0 3080 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_13
timestamp 1743498307
transform 1 0 3096 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_2
timestamp 1743498307
transform 1 0 3080 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_37
timestamp 1743498307
transform 1 0 3144 0 -1 210
box -4 -6 356 206
use OR2X2  OR2X2_3
timestamp 1743498307
transform 1 0 3496 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_12
timestamp 1743498307
transform -1 0 3608 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_25
timestamp 1743498307
transform -1 0 3640 0 -1 210
box -4 -6 36 206
use MUX2X1  MUX2X1_33
timestamp 1743498307
transform 1 0 3256 0 1 210
box -4 -6 100 206
use XOR2X1  XOR2X1_4
timestamp 1743498307
transform 1 0 3352 0 1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_8
timestamp 1743498307
transform 1 0 3464 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_11
timestamp 1743498307
transform 1 0 3528 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_38
timestamp 1743498307
transform -1 0 3928 0 1 210
box -4 -6 356 206
use DFFSR  DFFSR_20
timestamp 1743498307
transform 1 0 3640 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_22
timestamp 1743498307
transform -1 0 4072 0 1 210
box -4 -6 148 206
use BUFX2  BUFX2_10
timestamp 1743498307
transform 1 0 3992 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_47
timestamp 1743498307
transform 1 0 4040 0 -1 210
box -4 -6 196 206
use MUX2X1  MUX2X1_31
timestamp 1743498307
transform 1 0 4232 0 -1 210
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_44
timestamp 1743498307
transform -1 0 4520 0 -1 210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_16
timestamp 1743498307
transform 1 0 4072 0 1 210
box -4 -6 148 206
use OAI21X1  OAI21X1_105
timestamp 1743498307
transform 1 0 4216 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_13
timestamp 1743498307
transform -1 0 4344 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_95
timestamp 1743498307
transform -1 0 4536 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1743498307
transform -1 0 4472 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_104
timestamp 1743498307
transform -1 0 4408 0 1 210
box -4 -6 68 206
use FILL  FILL_1_2_2
timestamp 1743498307
transform 1 0 4568 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_1
timestamp 1743498307
transform 1 0 4552 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_0
timestamp 1743498307
transform 1 0 4536 0 1 210
box -4 -6 20 206
use MUX2X1  MUX2X1_28
timestamp 1743498307
transform 1 0 4632 0 -1 210
box -4 -6 100 206
use FILL  FILL_0_2_2
timestamp 1743498307
transform 1 0 4616 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_1
timestamp 1743498307
transform 1 0 4600 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_0
timestamp 1743498307
transform 1 0 4584 0 -1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_96
timestamp 1743498307
transform -1 0 4584 0 -1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_38
timestamp 1743498307
transform 1 0 4584 0 1 210
box -4 -6 196 206
use MUX2X1  MUX2X1_45
timestamp 1743498307
transform -1 0 4824 0 -1 210
box -4 -6 100 206
use OAI21X1  OAI21X1_134
timestamp 1743498307
transform 1 0 4824 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_133
timestamp 1743498307
transform -1 0 4952 0 -1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_35
timestamp 1743498307
transform 1 0 4952 0 -1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_116
timestamp 1743498307
transform 1 0 4776 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_115
timestamp 1743498307
transform -1 0 4904 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_26
timestamp 1743498307
transform 1 0 4904 0 1 210
box -4 -6 196 206
use MUX2X1  MUX2X1_42
timestamp 1743498307
transform -1 0 5240 0 -1 210
box -4 -6 100 206
use OAI21X1  OAI21X1_128
timestamp 1743498307
transform 1 0 5240 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_127
timestamp 1743498307
transform -1 0 5368 0 -1 210
box -4 -6 68 206
use BUFX4  BUFX4_34
timestamp 1743498307
transform -1 0 5432 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_140
timestamp 1743498307
transform 1 0 5096 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_139
timestamp 1743498307
transform -1 0 5224 0 1 210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_1
timestamp 1743498307
transform -1 0 5368 0 1 210
box -4 -6 148 206
use INVX1  INVX1_40
timestamp 1743498307
transform -1 0 5400 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_383
timestamp 1743498307
transform -1 0 5464 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_32
timestamp 1743498307
transform -1 0 5624 0 -1 210
box -4 -6 196 206
use INVX1  INVX1_116
timestamp 1743498307
transform -1 0 5656 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_402
timestamp 1743498307
transform 1 0 5656 0 -1 210
box -4 -6 68 206
use DFFSR  DFFSR_97
timestamp 1743498307
transform -1 0 6072 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_381
timestamp 1743498307
transform 1 0 5464 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_384
timestamp 1743498307
transform -1 0 5592 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_382
timestamp 1743498307
transform -1 0 5656 0 1 210
box -4 -6 68 206
use INVX1  INVX1_115
timestamp 1743498307
transform -1 0 5688 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_96
timestamp 1743498307
transform -1 0 6040 0 1 210
box -4 -6 356 206
use INVX1  INVX1_119
timestamp 1743498307
transform -1 0 6104 0 -1 210
box -4 -6 36 206
use FILL  FILL_1_1
timestamp 1743498307
transform -1 0 6120 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1743498307
transform -1 0 6136 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_117
timestamp 1743498307
transform -1 0 6072 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_23
timestamp 1743498307
transform 1 0 6072 0 1 210
box -4 -6 52 206
use FILL  FILL_2_1
timestamp 1743498307
transform 1 0 6120 0 1 210
box -4 -6 20 206
use DFFSR  DFFSR_85
timestamp 1743498307
transform 1 0 8 0 -1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_366
timestamp 1743498307
transform 1 0 360 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1743498307
transform -1 0 472 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_18
timestamp 1743498307
transform -1 0 616 0 -1 610
box -4 -6 148 206
use MUX2X1  MUX2X1_19
timestamp 1743498307
transform -1 0 712 0 -1 610
box -4 -6 100 206
use NAND2X1  NAND2X1_3
timestamp 1743498307
transform -1 0 760 0 -1 610
box -4 -6 52 206
use MUX2X1  MUX2X1_14
timestamp 1743498307
transform 1 0 760 0 -1 610
box -4 -6 100 206
use MUX2X1  MUX2X1_17
timestamp 1743498307
transform -1 0 952 0 -1 610
box -4 -6 100 206
use INVX1  INVX1_23
timestamp 1743498307
transform 1 0 952 0 -1 610
box -4 -6 36 206
use CLKBUF1  CLKBUF1_21
timestamp 1743498307
transform -1 0 1128 0 -1 610
box -4 -6 148 206
use MUX2X1  MUX2X1_10
timestamp 1743498307
transform -1 0 1224 0 -1 610
box -4 -6 100 206
use MUX2X1  MUX2X1_11
timestamp 1743498307
transform 1 0 1224 0 -1 610
box -4 -6 100 206
use BUFX4  BUFX4_10
timestamp 1743498307
transform -1 0 1384 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_22
timestamp 1743498307
transform -1 0 1480 0 -1 610
box -4 -6 100 206
use FILL  FILL_2_0_0
timestamp 1743498307
transform 1 0 1480 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1743498307
transform 1 0 1496 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1743498307
transform 1 0 1512 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_51
timestamp 1743498307
transform 1 0 1528 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_50
timestamp 1743498307
transform -1 0 1656 0 -1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_35
timestamp 1743498307
transform 1 0 1656 0 -1 610
box -4 -6 148 206
use DFFSR  DFFSR_88
timestamp 1743498307
transform 1 0 1800 0 -1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_114
timestamp 1743498307
transform 1 0 2152 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_108
timestamp 1743498307
transform -1 0 2232 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_117
timestamp 1743498307
transform 1 0 2232 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_116
timestamp 1743498307
transform 1 0 2280 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_360
timestamp 1743498307
transform -1 0 2392 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_100
timestamp 1743498307
transform -1 0 2424 0 -1 610
box -4 -6 36 206
use DFFSR  DFFSR_79
timestamp 1743498307
transform 1 0 2424 0 -1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_376
timestamp 1743498307
transform 1 0 2776 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_378
timestamp 1743498307
transform -1 0 2904 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_1_0
timestamp 1743498307
transform 1 0 2904 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1743498307
transform 1 0 2920 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1743498307
transform 1 0 2936 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_36
timestamp 1743498307
transform 1 0 2952 0 -1 610
box -4 -6 356 206
use MUX2X1  MUX2X1_34
timestamp 1743498307
transform -1 0 3400 0 -1 610
box -4 -6 100 206
use NAND2X1  NAND2X1_35
timestamp 1743498307
transform 1 0 3400 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_36
timestamp 1743498307
transform -1 0 3496 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_2
timestamp 1743498307
transform 1 0 3496 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_111
timestamp 1743498307
transform 1 0 3560 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_2
timestamp 1743498307
transform 1 0 3624 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_35
timestamp 1743498307
transform 1 0 3688 0 -1 610
box -4 -6 36 206
use DFFSR  DFFSR_33
timestamp 1743498307
transform 1 0 3720 0 -1 610
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_41
timestamp 1743498307
transform 1 0 4072 0 -1 610
box -4 -6 196 206
use INVX1  INVX1_45
timestamp 1743498307
transform 1 0 4264 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_166
timestamp 1743498307
transform 1 0 4296 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_121
timestamp 1743498307
transform -1 0 4424 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_122
timestamp 1743498307
transform -1 0 4488 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_39
timestamp 1743498307
transform -1 0 4584 0 -1 610
box -4 -6 100 206
use FILL  FILL_2_2_0
timestamp 1743498307
transform -1 0 4600 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_1
timestamp 1743498307
transform -1 0 4616 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_2
timestamp 1743498307
transform -1 0 4632 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_154
timestamp 1743498307
transform -1 0 4696 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_39
timestamp 1743498307
transform -1 0 4728 0 -1 610
box -4 -6 36 206
use MUX2X1  MUX2X1_36
timestamp 1743498307
transform 1 0 4728 0 -1 610
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_39
timestamp 1743498307
transform 1 0 4824 0 -1 610
box -4 -6 196 206
use INVX1  INVX1_46
timestamp 1743498307
transform 1 0 5016 0 -1 610
box -4 -6 36 206
use MUX2X1  MUX2X1_48
timestamp 1743498307
transform 1 0 5048 0 -1 610
box -4 -6 100 206
use BUFX4  BUFX4_31
timestamp 1743498307
transform -1 0 5208 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_51
timestamp 1743498307
transform -1 0 5304 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_145
timestamp 1743498307
transform 1 0 5304 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_146
timestamp 1743498307
transform -1 0 5432 0 -1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_29
timestamp 1743498307
transform -1 0 5624 0 -1 610
box -4 -6 196 206
use CLKBUF1  CLKBUF1_42
timestamp 1743498307
transform -1 0 5768 0 -1 610
box -4 -6 148 206
use DFFSR  DFFSR_100
timestamp 1743498307
transform -1 0 6120 0 -1 610
box -4 -6 356 206
use FILL  FILL_3_1
timestamp 1743498307
transform -1 0 6136 0 -1 610
box -4 -6 20 206
use INVX1  INVX1_106
timestamp 1743498307
transform 1 0 8 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_371
timestamp 1743498307
transform 1 0 40 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_370
timestamp 1743498307
transform -1 0 168 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_5
timestamp 1743498307
transform -1 0 216 0 1 610
box -4 -6 52 206
use MUX2X1  MUX2X1_5
timestamp 1743498307
transform -1 0 312 0 1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_16
timestamp 1743498307
transform 1 0 312 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_15
timestamp 1743498307
transform -1 0 440 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_23
timestamp 1743498307
transform 1 0 440 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_9
timestamp 1743498307
transform 1 0 632 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_32
timestamp 1743498307
transform 1 0 696 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_33
timestamp 1743498307
transform -1 0 824 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_13
timestamp 1743498307
transform 1 0 824 0 1 610
box -4 -6 100 206
use BUFX4  BUFX4_41
timestamp 1743498307
transform -1 0 984 0 1 610
box -4 -6 68 206
use INVX1  INVX1_22
timestamp 1743498307
transform 1 0 984 0 1 610
box -4 -6 36 206
use INVX1  INVX1_21
timestamp 1743498307
transform 1 0 1016 0 1 610
box -4 -6 36 206
use INVX1  INVX1_18
timestamp 1743498307
transform 1 0 1048 0 1 610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_17
timestamp 1743498307
transform -1 0 1272 0 1 610
box -4 -6 196 206
use INVX1  INVX1_17
timestamp 1743498307
transform -1 0 1304 0 1 610
box -4 -6 36 206
use INVX1  INVX1_15
timestamp 1743498307
transform 1 0 1304 0 1 610
box -4 -6 36 206
use BUFX4  BUFX4_42
timestamp 1743498307
transform 1 0 1336 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_52
timestamp 1743498307
transform 1 0 1400 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_53
timestamp 1743498307
transform -1 0 1528 0 1 610
box -4 -6 68 206
use FILL  FILL_3_0_0
timestamp 1743498307
transform 1 0 1528 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1743498307
transform 1 0 1544 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1743498307
transform 1 0 1560 0 1 610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1743498307
transform 1 0 1576 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_6
timestamp 1743498307
transform 1 0 1768 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_7
timestamp 1743498307
transform -1 0 1896 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_2
timestamp 1743498307
transform 1 0 1896 0 1 610
box -4 -6 100 206
use NAND2X1  NAND2X1_27
timestamp 1743498307
transform -1 0 2040 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_5
timestamp 1743498307
transform 1 0 2040 0 1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_88
timestamp 1743498307
transform -1 0 2456 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_87
timestamp 1743498307
transform 1 0 2456 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1743498307
transform 1 0 2520 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_4
timestamp 1743498307
transform -1 0 2920 0 1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_120
timestamp 1743498307
transform 1 0 2920 0 1 610
box -4 -6 52 206
use FILL  FILL_3_1_0
timestamp 1743498307
transform -1 0 2984 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1743498307
transform -1 0 3000 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1743498307
transform -1 0 3016 0 1 610
box -4 -6 20 206
use DFFSR  DFFSR_23
timestamp 1743498307
transform -1 0 3368 0 1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_109
timestamp 1743498307
transform 1 0 3368 0 1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_3
timestamp 1743498307
transform 1 0 3432 0 1 610
box -4 -6 116 206
use OAI21X1  OAI21X1_176
timestamp 1743498307
transform -1 0 3608 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_54
timestamp 1743498307
transform 1 0 3608 0 1 610
box -4 -6 52 206
use OR2X2  OR2X2_4
timestamp 1743498307
transform 1 0 3656 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1743498307
transform 1 0 3720 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_112
timestamp 1743498307
transform 1 0 3768 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_37
timestamp 1743498307
transform 1 0 3832 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_110
timestamp 1743498307
transform 1 0 3880 0 1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_6
timestamp 1743498307
transform 1 0 3944 0 1 610
box -4 -6 116 206
use INVX2  INVX2_2
timestamp 1743498307
transform 1 0 4056 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_174
timestamp 1743498307
transform 1 0 4088 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_173
timestamp 1743498307
transform 1 0 4152 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_39
timestamp 1743498307
transform -1 0 4264 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1743498307
transform 1 0 4264 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_37
timestamp 1743498307
transform -1 0 4392 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_168
timestamp 1743498307
transform 1 0 4392 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_107
timestamp 1743498307
transform -1 0 4520 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_156
timestamp 1743498307
transform -1 0 4584 0 1 610
box -4 -6 68 206
use FILL  FILL_3_2_0
timestamp 1743498307
transform -1 0 4600 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_1
timestamp 1743498307
transform -1 0 4616 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_2
timestamp 1743498307
transform -1 0 4632 0 1 610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_48
timestamp 1743498307
transform -1 0 4824 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_118
timestamp 1743498307
transform 1 0 4824 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_117
timestamp 1743498307
transform -1 0 4952 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_141
timestamp 1743498307
transform 1 0 4952 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_142
timestamp 1743498307
transform -1 0 5080 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_167
timestamp 1743498307
transform 1 0 5080 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_27
timestamp 1743498307
transform -1 0 5336 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_155
timestamp 1743498307
transform 1 0 5336 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_43
timestamp 1743498307
transform 1 0 5400 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_49
timestamp 1743498307
transform -1 0 5496 0 1 610
box -4 -6 52 206
use BUFX4  BUFX4_38
timestamp 1743498307
transform 1 0 5496 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_147
timestamp 1743498307
transform 1 0 5560 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_52
timestamp 1743498307
transform 1 0 5624 0 1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_148
timestamp 1743498307
transform -1 0 5784 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_30
timestamp 1743498307
transform 1 0 5784 0 1 610
box -4 -6 196 206
use NAND2X1  NAND2X1_118
timestamp 1743498307
transform 1 0 5976 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_390
timestamp 1743498307
transform -1 0 6088 0 1 610
box -4 -6 68 206
use FILL  FILL_4_1
timestamp 1743498307
transform 1 0 6088 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1743498307
transform 1 0 6104 0 1 610
box -4 -6 20 206
use FILL  FILL_4_3
timestamp 1743498307
transform 1 0 6120 0 1 610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_24
timestamp 1743498307
transform -1 0 200 0 -1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_14
timestamp 1743498307
transform -1 0 264 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_19
timestamp 1743498307
transform 1 0 264 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_6
timestamp 1743498307
transform -1 0 424 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_18
timestamp 1743498307
transform -1 0 488 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_21
timestamp 1743498307
transform 1 0 488 0 -1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_10
timestamp 1743498307
transform -1 0 744 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_3
timestamp 1743498307
transform 1 0 744 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_8
timestamp 1743498307
transform -1 0 904 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_6
timestamp 1743498307
transform 1 0 904 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_77
timestamp 1743498307
transform -1 0 1032 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_4
timestamp 1743498307
transform 1 0 1032 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_9
timestamp 1743498307
transform -1 0 1144 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_69
timestamp 1743498307
transform -1 0 1208 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_17
timestamp 1743498307
transform -1 0 1256 0 -1 1010
box -4 -6 52 206
use MUX2X1  MUX2X1_23
timestamp 1743498307
transform -1 0 1352 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_65
timestamp 1743498307
transform 1 0 1352 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_15
timestamp 1743498307
transform -1 0 1464 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_3
timestamp 1743498307
transform -1 0 1528 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1743498307
transform -1 0 1544 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1743498307
transform -1 0 1560 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1743498307
transform -1 0 1576 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_20
timestamp 1743498307
transform -1 0 1768 0 -1 1010
box -4 -6 196 206
use DFFSR  DFFSR_18
timestamp 1743498307
transform 1 0 1768 0 -1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_21
timestamp 1743498307
transform -1 0 2184 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_7
timestamp 1743498307
transform 1 0 2184 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_8
timestamp 1743498307
transform -1 0 2280 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1743498307
transform -1 0 2344 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1743498307
transform -1 0 2392 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_22
timestamp 1743498307
transform 1 0 2392 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_11
timestamp 1743498307
transform 1 0 2456 0 -1 1010
box -4 -6 36 206
use DFFSR  DFFSR_19
timestamp 1743498307
transform -1 0 2840 0 -1 1010
box -4 -6 356 206
use DFFSR  DFFSR_17
timestamp 1743498307
transform 1 0 2840 0 -1 1010
box -4 -6 356 206
use FILL  FILL_4_1_0
timestamp 1743498307
transform -1 0 3208 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1743498307
transform -1 0 3224 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1743498307
transform -1 0 3240 0 -1 1010
box -4 -6 20 206
use BUFX4  BUFX4_60
timestamp 1743498307
transform -1 0 3304 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_21
timestamp 1743498307
transform -1 0 3656 0 -1 1010
box -4 -6 356 206
use DFFSR  DFFSR_32
timestamp 1743498307
transform 1 0 3656 0 -1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_172
timestamp 1743498307
transform -1 0 4072 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_47
timestamp 1743498307
transform 1 0 4072 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_170
timestamp 1743498307
transform 1 0 4104 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_32
timestamp 1743498307
transform -1 0 4264 0 -1 1010
box -4 -6 100 206
use NOR2X1  NOR2X1_18
timestamp 1743498307
transform -1 0 4312 0 -1 1010
box -4 -6 52 206
use BUFX4  BUFX4_39
timestamp 1743498307
transform -1 0 4376 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_108
timestamp 1743498307
transform 1 0 4376 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_19
timestamp 1743498307
transform -1 0 4488 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_171
timestamp 1743498307
transform -1 0 4552 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_51
timestamp 1743498307
transform -1 0 4600 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_2_0
timestamp 1743498307
transform 1 0 4600 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_1
timestamp 1743498307
transform 1 0 4616 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_2
timestamp 1743498307
transform 1 0 4632 0 -1 1010
box -4 -6 20 206
use MUX2X1  MUX2X1_37
timestamp 1743498307
transform 1 0 4648 0 -1 1010
box -4 -6 100 206
use INVX1  INVX1_48
timestamp 1743498307
transform -1 0 4776 0 -1 1010
box -4 -6 36 206
use BUFX4  BUFX4_54
timestamp 1743498307
transform -1 0 4840 0 -1 1010
box -4 -6 68 206
use BUFX4  BUFX4_55
timestamp 1743498307
transform 1 0 4840 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_94
timestamp 1743498307
transform 1 0 4904 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_49
timestamp 1743498307
transform 1 0 4968 0 -1 1010
box -4 -6 100 206
use BUFX4  BUFX4_36
timestamp 1743498307
transform 1 0 5064 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_31
timestamp 1743498307
transform 1 0 5128 0 -1 1010
box -4 -6 52 206
use MUX2X1  MUX2X1_46
timestamp 1743498307
transform 1 0 5176 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_136
timestamp 1743498307
transform 1 0 5272 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_135
timestamp 1743498307
transform -1 0 5400 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1743498307
transform 1 0 5400 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_36
timestamp 1743498307
transform -1 0 5640 0 -1 1010
box -4 -6 196 206
use NAND2X1  NAND2X1_34
timestamp 1743498307
transform 1 0 5640 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_389
timestamp 1743498307
transform 1 0 5688 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_98
timestamp 1743498307
transform 1 0 5752 0 -1 1010
box -4 -6 356 206
use FILL  FILL_5_1
timestamp 1743498307
transform -1 0 6120 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1743498307
transform -1 0 6136 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1743498307
transform 1 0 8 0 1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_49
timestamp 1743498307
transform -1 0 264 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_48
timestamp 1743498307
transform -1 0 328 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_73
timestamp 1743498307
transform -1 0 392 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_25
timestamp 1743498307
transform -1 0 488 0 1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_46
timestamp 1743498307
transform 1 0 488 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_47
timestamp 1743498307
transform -1 0 616 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_20
timestamp 1743498307
transform -1 0 712 0 1 1010
box -4 -6 100 206
use BUFX4  BUFX4_43
timestamp 1743498307
transform -1 0 776 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_14
timestamp 1743498307
transform -1 0 840 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1743498307
transform 1 0 840 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_7
timestamp 1743498307
transform 1 0 888 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_78
timestamp 1743498307
transform -1 0 1016 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_79
timestamp 1743498307
transform 1 0 1016 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_70
timestamp 1743498307
transform 1 0 1080 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_71
timestamp 1743498307
transform 1 0 1144 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_11
timestamp 1743498307
transform 1 0 1208 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1743498307
transform -1 0 1320 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_14
timestamp 1743498307
transform 1 0 1320 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_67
timestamp 1743498307
transform -1 0 1416 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_84
timestamp 1743498307
transform -1 0 1480 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1743498307
transform -1 0 1496 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1743498307
transform -1 0 1512 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1743498307
transform -1 0 1528 0 1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_85
timestamp 1743498307
transform -1 0 1592 0 1 1010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_14
timestamp 1743498307
transform 1 0 1592 0 1 1010
box -4 -6 148 206
use MUX2X1  MUX2X1_8
timestamp 1743498307
transform 1 0 1736 0 1 1010
box -4 -6 100 206
use MUX2X1  MUX2X1_7
timestamp 1743498307
transform 1 0 1832 0 1 1010
box -4 -6 100 206
use XOR2X1  XOR2X1_2
timestamp 1743498307
transform 1 0 1928 0 1 1010
box -4 -6 116 206
use OR2X2  OR2X2_2
timestamp 1743498307
transform -1 0 2104 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_1
timestamp 1743498307
transform -1 0 2168 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_1
timestamp 1743498307
transform 1 0 2168 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_1
timestamp 1743498307
transform -1 0 2264 0 1 1010
box -4 -6 36 206
use OR2X2  OR2X2_1
timestamp 1743498307
transform 1 0 2264 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_1
timestamp 1743498307
transform 1 0 2328 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_23
timestamp 1743498307
transform -1 0 2440 0 1 1010
box -4 -6 68 206
use DFFSR  DFFSR_2
timestamp 1743498307
transform 1 0 2440 0 1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_20
timestamp 1743498307
transform -1 0 2856 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_97
timestamp 1743498307
transform -1 0 2920 0 1 1010
box -4 -6 68 206
use XOR2X1  XOR2X1_1
timestamp 1743498307
transform 1 0 2920 0 1 1010
box -4 -6 116 206
use FILL  FILL_5_1_0
timestamp 1743498307
transform 1 0 3032 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1743498307
transform 1 0 3048 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1743498307
transform 1 0 3064 0 1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_122
timestamp 1743498307
transform 1 0 3080 0 1 1010
box -4 -6 52 206
use DFFSR  DFFSR_25
timestamp 1743498307
transform -1 0 3480 0 1 1010
box -4 -6 356 206
use BUFX4  BUFX4_78
timestamp 1743498307
transform -1 0 3544 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_79
timestamp 1743498307
transform 1 0 3544 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_110
timestamp 1743498307
transform -1 0 3640 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_375
timestamp 1743498307
transform 1 0 3640 0 1 1010
box -4 -6 68 206
use DFFSR  DFFSR_91
timestamp 1743498307
transform 1 0 3704 0 1 1010
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_42
timestamp 1743498307
transform -1 0 4248 0 1 1010
box -4 -6 196 206
use INVX1  INVX1_29
timestamp 1743498307
transform 1 0 4248 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_124
timestamp 1743498307
transform -1 0 4344 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_40
timestamp 1743498307
transform -1 0 4440 0 1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_160
timestamp 1743498307
transform -1 0 4504 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_158
timestamp 1743498307
transform -1 0 4568 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_2_0
timestamp 1743498307
transform 1 0 4568 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_1
timestamp 1743498307
transform 1 0 4584 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_2
timestamp 1743498307
transform 1 0 4600 0 1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_41
timestamp 1743498307
transform 1 0 4616 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_38
timestamp 1743498307
transform -1 0 4696 0 1 1010
box -4 -6 36 206
use INVX1  INVX1_41
timestamp 1743498307
transform -1 0 4728 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_38
timestamp 1743498307
transform 1 0 4728 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1743498307
transform 1 0 4776 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_159
timestamp 1743498307
transform -1 0 4888 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_45
timestamp 1743498307
transform -1 0 4936 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_103
timestamp 1743498307
transform 1 0 4936 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_33
timestamp 1743498307
transform 1 0 5000 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_42
timestamp 1743498307
transform -1 0 5080 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_106
timestamp 1743498307
transform 1 0 5080 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_43
timestamp 1743498307
transform -1 0 5240 0 1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_130
timestamp 1743498307
transform 1 0 5240 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_129
timestamp 1743498307
transform -1 0 5368 0 1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_33
timestamp 1743498307
transform -1 0 5560 0 1 1010
box -4 -6 196 206
use BUFX4  BUFX4_32
timestamp 1743498307
transform 1 0 5560 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_387
timestamp 1743498307
transform 1 0 5624 0 1 1010
box -4 -6 68 206
use DFFSR  DFFSR_99
timestamp 1743498307
transform -1 0 6040 0 1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_388
timestamp 1743498307
transform -1 0 6104 0 1 1010
box -4 -6 68 206
use FILL  FILL_6_1
timestamp 1743498307
transform 1 0 6104 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1743498307
transform 1 0 6120 0 1 1010
box -4 -6 20 206
use DFFSR  DFFSR_89
timestamp 1743498307
transform -1 0 360 0 -1 1410
box -4 -6 356 206
use NAND2X1  NAND2X1_113
timestamp 1743498307
transform 1 0 360 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_357
timestamp 1743498307
transform -1 0 472 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_21
timestamp 1743498307
transform -1 0 568 0 -1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_56
timestamp 1743498307
transform 1 0 568 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_57
timestamp 1743498307
transform -1 0 696 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1743498307
transform 1 0 696 0 -1 1410
box -4 -6 196 206
use BUFX4  BUFX4_13
timestamp 1743498307
transform -1 0 952 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_81
timestamp 1743498307
transform -1 0 1016 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1743498307
transform 1 0 1016 0 -1 1410
box -4 -6 196 206
use NAND2X1  NAND2X1_12
timestamp 1743498307
transform 1 0 1208 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_24
timestamp 1743498307
transform 1 0 1256 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_23
timestamp 1743498307
transform 1 0 1288 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_82
timestamp 1743498307
transform 1 0 1336 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_66
timestamp 1743498307
transform 1 0 1400 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1743498307
transform -1 0 1512 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_0_0
timestamp 1743498307
transform 1 0 1512 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1743498307
transform 1 0 1528 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1743498307
transform 1 0 1544 0 -1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_83
timestamp 1743498307
transform 1 0 1560 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_14
timestamp 1743498307
transform -1 0 1976 0 -1 1410
box -4 -6 356 206
use NAND2X1  NAND2X1_18
timestamp 1743498307
transform -1 0 2024 0 -1 1410
box -4 -6 52 206
use BUFX4  BUFX4_52
timestamp 1743498307
transform -1 0 2088 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_1
timestamp 1743498307
transform -1 0 2440 0 -1 1410
box -4 -6 356 206
use NOR2X1  NOR2X1_2
timestamp 1743498307
transform -1 0 2488 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_6
timestamp 1743498307
transform 1 0 2488 0 -1 1410
box -4 -6 52 206
use BUFX4  BUFX4_50
timestamp 1743498307
transform 1 0 2536 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_89
timestamp 1743498307
transform 1 0 2600 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_6
timestamp 1743498307
transform -1 0 3016 0 -1 1410
box -4 -6 356 206
use FILL  FILL_6_1_0
timestamp 1743498307
transform -1 0 3032 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1743498307
transform -1 0 3048 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1743498307
transform -1 0 3064 0 -1 1410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_15
timestamp 1743498307
transform -1 0 3208 0 -1 1410
box -4 -6 148 206
use DFFSR  DFFSR_104
timestamp 1743498307
transform 1 0 3208 0 -1 1410
box -4 -6 356 206
use BUFX4  BUFX4_80
timestamp 1743498307
transform 1 0 3560 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_3
timestamp 1743498307
transform -1 0 3672 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_169
timestamp 1743498307
transform 1 0 3672 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_52
timestamp 1743498307
transform 1 0 3736 0 -1 1410
box -4 -6 52 206
use DFFSR  DFFSR_31
timestamp 1743498307
transform 1 0 3784 0 -1 1410
box -4 -6 356 206
use CLKBUF1  CLKBUF1_32
timestamp 1743498307
transform -1 0 4280 0 -1 1410
box -4 -6 148 206
use OAI21X1  OAI21X1_123
timestamp 1743498307
transform -1 0 4344 0 -1 1410
box -4 -6 68 206
use BUFX4  BUFX4_33
timestamp 1743498307
transform 1 0 4344 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_11
timestamp 1743498307
transform -1 0 4472 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1743498307
transform 1 0 4472 0 -1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_5
timestamp 1743498307
transform 1 0 4520 0 -1 1410
box -4 -6 116 206
use FILL  FILL_6_2_0
timestamp 1743498307
transform -1 0 4648 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_1
timestamp 1743498307
transform -1 0 4664 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_2
timestamp 1743498307
transform -1 0 4680 0 -1 1410
box -4 -6 20 206
use INVX1  INVX1_28
timestamp 1743498307
transform -1 0 4712 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_13
timestamp 1743498307
transform 1 0 4712 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_125
timestamp 1743498307
transform 1 0 4760 0 -1 1410
box -4 -6 68 206
use BUFX4  BUFX4_57
timestamp 1743498307
transform -1 0 4888 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_126
timestamp 1743498307
transform -1 0 4952 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_41
timestamp 1743498307
transform -1 0 5048 0 -1 1410
box -4 -6 100 206
use BUFX4  BUFX4_40
timestamp 1743498307
transform -1 0 5112 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_97
timestamp 1743498307
transform 1 0 5112 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_31
timestamp 1743498307
transform -1 0 5368 0 -1 1410
box -4 -6 196 206
use OAI21X1  OAI21X1_90
timestamp 1743498307
transform 1 0 5368 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_26
timestamp 1743498307
transform -1 0 5464 0 -1 1410
box -4 -6 36 206
use BUFX4  BUFX4_56
timestamp 1743498307
transform 1 0 5464 0 -1 1410
box -4 -6 68 206
use BUFX4  BUFX4_35
timestamp 1743498307
transform 1 0 5528 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_44
timestamp 1743498307
transform -1 0 5624 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_131
timestamp 1743498307
transform 1 0 5624 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_44
timestamp 1743498307
transform 1 0 5688 0 -1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_132
timestamp 1743498307
transform 1 0 5784 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_32
timestamp 1743498307
transform -1 0 5896 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_34
timestamp 1743498307
transform 1 0 5896 0 -1 1410
box -4 -6 196 206
use FILL  FILL_7_1
timestamp 1743498307
transform -1 0 6104 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1743498307
transform -1 0 6120 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_3
timestamp 1743498307
transform -1 0 6136 0 -1 1410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1743498307
transform 1 0 8 0 1 1410
box -4 -6 196 206
use OAI21X1  OAI21X1_12
timestamp 1743498307
transform -1 0 264 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_58
timestamp 1743498307
transform 1 0 264 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_59
timestamp 1743498307
transform -1 0 392 0 1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_26
timestamp 1743498307
transform -1 0 488 0 1 1410
box -4 -6 100 206
use MUX2X1  MUX2X1_1
timestamp 1743498307
transform -1 0 584 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_3
timestamp 1743498307
transform 1 0 584 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_4
timestamp 1743498307
transform -1 0 712 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_19
timestamp 1743498307
transform 1 0 712 0 1 1410
box -4 -6 196 206
use NAND3X1  NAND3X1_2
timestamp 1743498307
transform 1 0 904 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_61
timestamp 1743498307
transform 1 0 968 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_5
timestamp 1743498307
transform 1 0 1032 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_74
timestamp 1743498307
transform 1 0 1096 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_73
timestamp 1743498307
transform -1 0 1224 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_62
timestamp 1743498307
transform 1 0 1224 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_75
timestamp 1743498307
transform 1 0 1288 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_63
timestamp 1743498307
transform 1 0 1352 0 1 1410
box -4 -6 68 206
use INVX2  INVX2_1
timestamp 1743498307
transform 1 0 1416 0 1 1410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_3
timestamp 1743498307
transform -1 0 1560 0 1 1410
box -4 -6 116 206
use FILL  FILL_7_0_0
timestamp 1743498307
transform 1 0 1560 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1743498307
transform 1 0 1576 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1743498307
transform 1 0 1592 0 1 1410
box -4 -6 20 206
use DFFSR  DFFSR_9
timestamp 1743498307
transform 1 0 1608 0 1 1410
box -4 -6 356 206
use OAI21X1  OAI21X1_68
timestamp 1743498307
transform -1 0 2024 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_99
timestamp 1743498307
transform -1 0 2088 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_5
timestamp 1743498307
transform -1 0 2136 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_20
timestamp 1743498307
transform -1 0 2184 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_72
timestamp 1743498307
transform 1 0 2184 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_10
timestamp 1743498307
transform 1 0 2248 0 1 1410
box -4 -6 356 206
use NAND2X1  NAND2X1_28
timestamp 1743498307
transform -1 0 2648 0 1 1410
box -4 -6 52 206
use DFFSR  DFFSR_102
timestamp 1743498307
transform 1 0 2648 0 1 1410
box -4 -6 356 206
use INVX1  INVX1_120
timestamp 1743498307
transform -1 0 3032 0 1 1410
box -4 -6 36 206
use FILL  FILL_7_1_0
timestamp 1743498307
transform 1 0 3032 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1743498307
transform 1 0 3048 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1743498307
transform 1 0 3064 0 1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_178
timestamp 1743498307
transform 1 0 3080 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_56
timestamp 1743498307
transform 1 0 3144 0 1 1410
box -4 -6 52 206
use DFFSR  DFFSR_22
timestamp 1743498307
transform 1 0 3192 0 1 1410
box -4 -6 356 206
use NAND2X1  NAND2X1_53
timestamp 1743498307
transform -1 0 3592 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_175
timestamp 1743498307
transform -1 0 3656 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_119
timestamp 1743498307
transform 1 0 3656 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_152
timestamp 1743498307
transform -1 0 3768 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_164
timestamp 1743498307
transform -1 0 3832 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_150
timestamp 1743498307
transform 1 0 3832 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_162
timestamp 1743498307
transform -1 0 3960 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_9
timestamp 1743498307
transform -1 0 4024 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_12
timestamp 1743498307
transform -1 0 4088 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_92
timestamp 1743498307
transform 1 0 4088 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_93
timestamp 1743498307
transform -1 0 4216 0 1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_27
timestamp 1743498307
transform -1 0 4312 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_151
timestamp 1743498307
transform -1 0 4376 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_37
timestamp 1743498307
transform -1 0 4408 0 1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_29
timestamp 1743498307
transform 1 0 4408 0 1 1410
box -4 -6 100 206
use NAND2X1  NAND2X1_40
timestamp 1743498307
transform -1 0 4552 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_2_0
timestamp 1743498307
transform -1 0 4568 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_1
timestamp 1743498307
transform -1 0 4584 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_2
timestamp 1743498307
transform -1 0 4600 0 1 1410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_43
timestamp 1743498307
transform -1 0 4792 0 1 1410
box -4 -6 196 206
use INVX1  INVX1_43
timestamp 1743498307
transform -1 0 4824 0 1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_38
timestamp 1743498307
transform 1 0 4824 0 1 1410
box -4 -6 100 206
use NAND2X1  NAND2X1_47
timestamp 1743498307
transform 1 0 4920 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_163
timestamp 1743498307
transform -1 0 5032 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_120
timestamp 1743498307
transform 1 0 5032 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_119
timestamp 1743498307
transform -1 0 5160 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_40
timestamp 1743498307
transform -1 0 5352 0 1 1410
box -4 -6 196 206
use OAI21X1  OAI21X1_102
timestamp 1743498307
transform 1 0 5352 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_46
timestamp 1743498307
transform -1 0 5608 0 1 1410
box -4 -6 196 206
use OR2X2  OR2X2_10
timestamp 1743498307
transform 1 0 5608 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_103
timestamp 1743498307
transform -1 0 6024 0 1 1410
box -4 -6 356 206
use INVX1  INVX1_118
timestamp 1743498307
transform -1 0 6056 0 1 1410
box -4 -6 36 206
use BUFX2  BUFX2_14
timestamp 1743498307
transform 1 0 6056 0 1 1410
box -4 -6 52 206
use FILL  FILL_8_1
timestamp 1743498307
transform 1 0 6104 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1743498307
transform 1 0 6120 0 1 1410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_22
timestamp 1743498307
transform 1 0 8 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_13
timestamp 1743498307
transform -1 0 264 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_4
timestamp 1743498307
transform 1 0 264 0 -1 1810
box -4 -6 100 206
use BUFX4  BUFX4_74
timestamp 1743498307
transform -1 0 424 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_2
timestamp 1743498307
transform -1 0 488 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_3
timestamp 1743498307
transform -1 0 520 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1743498307
transform -1 0 712 0 -1 1810
box -4 -6 196 206
use MUX2X1  MUX2X1_9
timestamp 1743498307
transform -1 0 808 0 -1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_25
timestamp 1743498307
transform 1 0 808 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_24
timestamp 1743498307
transform -1 0 936 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_12
timestamp 1743498307
transform 1 0 936 0 -1 1810
box -4 -6 36 206
use MUX2X1  MUX2X1_15
timestamp 1743498307
transform -1 0 1064 0 -1 1810
box -4 -6 100 206
use INVX1  INVX1_20
timestamp 1743498307
transform 1 0 1064 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_19
timestamp 1743498307
transform 1 0 1096 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_13
timestamp 1743498307
transform 1 0 1144 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_19
timestamp 1743498307
transform 1 0 1176 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_10
timestamp 1743498307
transform -1 0 1256 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1743498307
transform 1 0 1256 0 -1 1810
box -4 -6 52 206
use BUFX4  BUFX4_76
timestamp 1743498307
transform -1 0 1368 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_16
timestamp 1743498307
transform 1 0 1368 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_3
timestamp 1743498307
transform -1 0 1448 0 -1 1810
box -4 -6 52 206
use FILL  FILL_8_0_0
timestamp 1743498307
transform -1 0 1464 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1743498307
transform -1 0 1480 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1743498307
transform -1 0 1496 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_13
timestamp 1743498307
transform -1 0 1848 0 -1 1810
box -4 -6 356 206
use BUFX4  BUFX4_51
timestamp 1743498307
transform -1 0 1912 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_24
timestamp 1743498307
transform -1 0 1960 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_25
timestamp 1743498307
transform -1 0 2008 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_86
timestamp 1743498307
transform -1 0 2072 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_3
timestamp 1743498307
transform -1 0 2424 0 -1 1810
box -4 -6 356 206
use DFFSR  DFFSR_8
timestamp 1743498307
transform 1 0 2424 0 -1 1810
box -4 -6 356 206
use NAND2X1  NAND2X1_16
timestamp 1743498307
transform -1 0 2824 0 -1 1810
box -4 -6 52 206
use CLKBUF1  CLKBUF1_38
timestamp 1743498307
transform -1 0 2968 0 -1 1810
box -4 -6 148 206
use FILL  FILL_8_1_0
timestamp 1743498307
transform 1 0 2968 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1743498307
transform 1 0 2984 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1743498307
transform 1 0 3000 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_27
timestamp 1743498307
transform 1 0 3016 0 -1 1810
box -4 -6 356 206
use NAND2X1  NAND2X1_48
timestamp 1743498307
transform 1 0 3368 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_153
timestamp 1743498307
transform -1 0 3480 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_44
timestamp 1743498307
transform 1 0 3480 0 -1 1810
box -4 -6 52 206
use BUFX4  BUFX4_59
timestamp 1743498307
transform 1 0 3528 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_42
timestamp 1743498307
transform 1 0 3592 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_177
timestamp 1743498307
transform 1 0 3640 0 -1 1810
box -4 -6 68 206
use BUFX4  BUFX4_77
timestamp 1743498307
transform 1 0 3704 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_55
timestamp 1743498307
transform 1 0 3768 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_36
timestamp 1743498307
transform -1 0 3848 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_37
timestamp 1743498307
transform -1 0 4040 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_113
timestamp 1743498307
transform 1 0 4040 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_114
timestamp 1743498307
transform -1 0 4168 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_35
timestamp 1743498307
transform -1 0 4264 0 -1 1810
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_45
timestamp 1743498307
transform 1 0 4264 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_99
timestamp 1743498307
transform 1 0 4456 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_98
timestamp 1743498307
transform -1 0 4584 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_2_0
timestamp 1743498307
transform 1 0 4584 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_1
timestamp 1743498307
transform 1 0 4600 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_2
timestamp 1743498307
transform 1 0 4616 0 -1 1810
box -4 -6 20 206
use OAI21X1  OAI21X1_137
timestamp 1743498307
transform 1 0 4632 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_138
timestamp 1743498307
transform 1 0 4696 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_47
timestamp 1743498307
transform -1 0 4856 0 -1 1810
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_28
timestamp 1743498307
transform -1 0 5048 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_144
timestamp 1743498307
transform 1 0 5048 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_143
timestamp 1743498307
transform -1 0 5176 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_50
timestamp 1743498307
transform 1 0 5176 0 -1 1810
box -4 -6 100 206
use MUX2X1  MUX2X1_30
timestamp 1743498307
transform 1 0 5272 0 -1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_101
timestamp 1743498307
transform 1 0 5368 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_100
timestamp 1743498307
transform 1 0 5432 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_109
timestamp 1743498307
transform -1 0 5528 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_29
timestamp 1743498307
transform 1 0 5528 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_379
timestamp 1743498307
transform 1 0 5576 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_95
timestamp 1743498307
transform -1 0 5992 0 -1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_380
timestamp 1743498307
transform -1 0 6056 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_114
timestamp 1743498307
transform -1 0 6088 0 -1 1810
box -4 -6 36 206
use FILL  FILL_9_1
timestamp 1743498307
transform -1 0 6104 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1743498307
transform -1 0 6120 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_3
timestamp 1743498307
transform -1 0 6136 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_84
timestamp 1743498307
transform 1 0 8 0 1 1810
box -4 -6 356 206
use INVX1  INVX1_9
timestamp 1743498307
transform -1 0 392 0 1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1743498307
transform 1 0 392 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_55
timestamp 1743498307
transform -1 0 648 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_54
timestamp 1743498307
transform 1 0 648 0 1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_24
timestamp 1743498307
transform -1 0 808 0 1 1810
box -4 -6 100 206
use BUFX4  BUFX4_44
timestamp 1743498307
transform -1 0 872 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1743498307
transform 1 0 872 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_37
timestamp 1743498307
transform 1 0 1064 0 1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_12
timestamp 1743498307
transform 1 0 1128 0 1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_36
timestamp 1743498307
transform -1 0 1288 0 1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_16
timestamp 1743498307
transform 1 0 1288 0 1 1810
box -4 -6 100 206
use BUFX4  BUFX4_12
timestamp 1743498307
transform 1 0 1384 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_4
timestamp 1743498307
transform -1 0 1480 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_8
timestamp 1743498307
transform 1 0 1480 0 1 1810
box -4 -6 52 206
use FILL  FILL_9_0_0
timestamp 1743498307
transform -1 0 1544 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1743498307
transform -1 0 1560 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1743498307
transform -1 0 1576 0 1 1810
box -4 -6 20 206
use INVX1  INVX1_5
timestamp 1743498307
transform -1 0 1608 0 1 1810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_1
timestamp 1743498307
transform 1 0 1608 0 1 1810
box -4 -6 116 206
use DFFSR  DFFSR_15
timestamp 1743498307
transform -1 0 2072 0 1 1810
box -4 -6 356 206
use NAND2X1  NAND2X1_22
timestamp 1743498307
transform -1 0 2120 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_76
timestamp 1743498307
transform 1 0 2120 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_5
timestamp 1743498307
transform 1 0 2184 0 1 1810
box -4 -6 52 206
use INVX8  INVX8_1
timestamp 1743498307
transform -1 0 2312 0 1 1810
box -4 -6 84 206
use OAI21X1  OAI21X1_80
timestamp 1743498307
transform 1 0 2312 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_60
timestamp 1743498307
transform 1 0 2376 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1743498307
transform 1 0 2440 0 1 1810
box -4 -6 52 206
use BUFX4  BUFX4_53
timestamp 1743498307
transform -1 0 2552 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_7
timestamp 1743498307
transform 1 0 2552 0 1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_64
timestamp 1743498307
transform -1 0 2968 0 1 1810
box -4 -6 68 206
use BUFX4  BUFX4_98
timestamp 1743498307
transform 1 0 2968 0 1 1810
box -4 -6 68 206
use FILL  FILL_9_1_0
timestamp 1743498307
transform 1 0 3032 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1743498307
transform 1 0 3048 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1743498307
transform 1 0 3064 0 1 1810
box -4 -6 20 206
use INVX1  INVX1_183
timestamp 1743498307
transform 1 0 3080 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_15
timestamp 1743498307
transform 1 0 3112 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_161
timestamp 1743498307
transform 1 0 3160 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_29
timestamp 1743498307
transform -1 0 3576 0 1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_149
timestamp 1743498307
transform -1 0 3640 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_26
timestamp 1743498307
transform -1 0 3992 0 1 1810
box -4 -6 356 206
use DFFSR  DFFSR_24
timestamp 1743498307
transform 1 0 3992 0 1 1810
box -4 -6 356 206
use DFFSR  DFFSR_35
timestamp 1743498307
transform 1 0 4344 0 1 1810
box -4 -6 356 206
use FILL  FILL_9_2_0
timestamp 1743498307
transform 1 0 4696 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_1
timestamp 1743498307
transform 1 0 4712 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_2
timestamp 1743498307
transform 1 0 4728 0 1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_25
timestamp 1743498307
transform 1 0 4744 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_91
timestamp 1743498307
transform 1 0 4936 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_121
timestamp 1743498307
transform -1 0 5048 0 1 1810
box -4 -6 52 206
use INVX8  INVX8_6
timestamp 1743498307
transform -1 0 5128 0 1 1810
box -4 -6 84 206
use NOR2X1  NOR2X1_14
timestamp 1743498307
transform -1 0 5176 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_377
timestamp 1743498307
transform -1 0 5240 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_112
timestamp 1743498307
transform -1 0 5272 0 1 1810
box -4 -6 36 206
use DFFSR  DFFSR_101
timestamp 1743498307
transform -1 0 5624 0 1 1810
box -4 -6 356 206
use DFFSR  DFFSR_93
timestamp 1743498307
transform 1 0 5624 0 1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_386
timestamp 1743498307
transform -1 0 6040 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_12
timestamp 1743498307
transform 1 0 6040 0 1 1810
box -4 -6 52 206
use FILL  FILL_10_1
timestamp 1743498307
transform 1 0 6088 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_2
timestamp 1743498307
transform 1 0 6104 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_3
timestamp 1743498307
transform 1 0 6120 0 1 1810
box -4 -6 20 206
use INVX1  INVX1_105
timestamp 1743498307
transform 1 0 8 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_369
timestamp 1743498307
transform 1 0 40 0 -1 2210
box -4 -6 68 206
use OR2X2  OR2X2_9
timestamp 1743498307
transform -1 0 168 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_368
timestamp 1743498307
transform 1 0 168 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1743498307
transform 1 0 232 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_17
timestamp 1743498307
transform -1 0 344 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_11
timestamp 1743498307
transform -1 0 408 0 -1 2210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_25
timestamp 1743498307
transform -1 0 552 0 -1 2210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_24
timestamp 1743498307
transform 1 0 552 0 -1 2210
box -4 -6 148 206
use MUX2X1  MUX2X1_18
timestamp 1743498307
transform -1 0 792 0 -1 2210
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1743498307
transform -1 0 984 0 -1 2210
box -4 -6 196 206
use OAI21X1  OAI21X1_43
timestamp 1743498307
transform 1 0 984 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_42
timestamp 1743498307
transform -1 0 1112 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_31
timestamp 1743498307
transform 1 0 1112 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_30
timestamp 1743498307
transform -1 0 1240 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_38
timestamp 1743498307
transform 1 0 1240 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_39
timestamp 1743498307
transform -1 0 1368 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1743498307
transform -1 0 1560 0 -1 2210
box -4 -6 196 206
use FILL  FILL_10_0_0
timestamp 1743498307
transform 1 0 1560 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_1
timestamp 1743498307
transform 1 0 1576 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_2
timestamp 1743498307
transform 1 0 1592 0 -1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_10
timestamp 1743498307
transform 1 0 1608 0 -1 2210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_2
timestamp 1743498307
transform -1 0 1768 0 -1 2210
box -4 -6 116 206
use DFFSR  DFFSR_16
timestamp 1743498307
transform -1 0 2120 0 -1 2210
box -4 -6 356 206
use DFFSR  DFFSR_12
timestamp 1743498307
transform 1 0 2120 0 -1 2210
box -4 -6 356 206
use INVX1  INVX1_182
timestamp 1743498307
transform 1 0 2472 0 -1 2210
box -4 -6 36 206
use DFFSR  DFFSR_171
timestamp 1743498307
transform 1 0 2504 0 -1 2210
box -4 -6 356 206
use INVX1  INVX1_159
timestamp 1743498307
transform -1 0 2888 0 -1 2210
box -4 -6 36 206
use CLKBUF1  CLKBUF1_3
timestamp 1743498307
transform -1 0 3032 0 -1 2210
box -4 -6 148 206
use FILL  FILL_10_1_0
timestamp 1743498307
transform -1 0 3048 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_1
timestamp 1743498307
transform -1 0 3064 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_2
timestamp 1743498307
transform -1 0 3080 0 -1 2210
box -4 -6 20 206
use DFFSR  DFFSR_167
timestamp 1743498307
transform -1 0 3432 0 -1 2210
box -4 -6 356 206
use OAI21X1  OAI21X1_157
timestamp 1743498307
transform 1 0 3432 0 -1 2210
box -4 -6 68 206
use DFFSR  DFFSR_28
timestamp 1743498307
transform -1 0 3848 0 -1 2210
box -4 -6 356 206
use NAND2X1  NAND2X1_46
timestamp 1743498307
transform 1 0 3848 0 -1 2210
box -4 -6 52 206
use INVX8  INVX8_2
timestamp 1743498307
transform 1 0 3896 0 -1 2210
box -4 -6 84 206
use BUFX4  BUFX4_58
timestamp 1743498307
transform 1 0 3976 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_165
timestamp 1743498307
transform 1 0 4040 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_33
timestamp 1743498307
transform 1 0 4104 0 -1 2210
box -4 -6 36 206
use BUFX4  BUFX4_1
timestamp 1743498307
transform 1 0 4136 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_50
timestamp 1743498307
transform 1 0 4200 0 -1 2210
box -4 -6 52 206
use DFFSR  DFFSR_30
timestamp 1743498307
transform -1 0 4600 0 -1 2210
box -4 -6 356 206
use FILL  FILL_10_2_0
timestamp 1743498307
transform 1 0 4600 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_1
timestamp 1743498307
transform 1 0 4616 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_2
timestamp 1743498307
transform 1 0 4632 0 -1 2210
box -4 -6 20 206
use INVX1  INVX1_34
timestamp 1743498307
transform 1 0 4648 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_32
timestamp 1743498307
transform 1 0 4680 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_30
timestamp 1743498307
transform 1 0 4712 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_27
timestamp 1743498307
transform 1 0 4744 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_31
timestamp 1743498307
transform 1 0 4776 0 -1 2210
box -4 -6 36 206
use AND2X2  AND2X2_5
timestamp 1743498307
transform -1 0 4872 0 -1 2210
box -4 -6 68 206
use DFFSR  DFFSR_139
timestamp 1743498307
transform 1 0 4872 0 -1 2210
box -4 -6 356 206
use INVX1  INVX1_146
timestamp 1743498307
transform 1 0 5224 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_426
timestamp 1743498307
transform 1 0 5256 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_139
timestamp 1743498307
transform -1 0 5368 0 -1 2210
box -4 -6 52 206
use DFFSR  DFFSR_136
timestamp 1743498307
transform -1 0 5720 0 -1 2210
box -4 -6 356 206
use OAI21X1  OAI21X1_385
timestamp 1743498307
transform 1 0 5720 0 -1 2210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_13
timestamp 1743498307
transform -1 0 5928 0 -1 2210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_2
timestamp 1743498307
transform 1 0 5928 0 -1 2210
box -4 -6 148 206
use FILL  FILL_11_1
timestamp 1743498307
transform -1 0 6088 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_2
timestamp 1743498307
transform -1 0 6104 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_3
timestamp 1743498307
transform -1 0 6120 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_4
timestamp 1743498307
transform -1 0 6136 0 -1 2210
box -4 -6 20 206
use INVX1  INVX1_107
timestamp 1743498307
transform 1 0 8 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_103
timestamp 1743498307
transform 1 0 40 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_373
timestamp 1743498307
transform 1 0 72 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_372
timestamp 1743498307
transform 1 0 136 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_365
timestamp 1743498307
transform 1 0 200 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_6
timestamp 1743498307
transform 1 0 264 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_364
timestamp 1743498307
transform 1 0 312 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1743498307
transform -1 0 408 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_97
timestamp 1743498307
transform 1 0 408 0 1 2210
box -4 -6 36 206
use DFFSR  DFFSR_87
timestamp 1743498307
transform 1 0 440 0 1 2210
box -4 -6 356 206
use NAND2X1  NAND2X1_2
timestamp 1743498307
transform -1 0 840 0 1 2210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_36
timestamp 1743498307
transform 1 0 840 0 1 2210
box -4 -6 148 206
use BUFX4  BUFX4_4
timestamp 1743498307
transform 1 0 984 0 1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1743498307
transform 1 0 1048 0 1 2210
box -4 -6 196 206
use OAI21X1  OAI21X1_5
timestamp 1743498307
transform -1 0 1304 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_4
timestamp 1743498307
transform -1 0 1352 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1743498307
transform 1 0 1352 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_2
timestamp 1743498307
transform -1 0 1448 0 1 2210
box -4 -6 36 206
use FILL  FILL_11_0_0
timestamp 1743498307
transform 1 0 1448 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_1
timestamp 1743498307
transform 1 0 1464 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_2
timestamp 1743498307
transform 1 0 1480 0 1 2210
box -4 -6 20 206
use DFFSR  DFFSR_159
timestamp 1743498307
transform 1 0 1496 0 1 2210
box -4 -6 356 206
use INVX1  INVX1_157
timestamp 1743498307
transform 1 0 1848 0 1 2210
box -4 -6 36 206
use DFFSR  DFFSR_11
timestamp 1743498307
transform 1 0 1880 0 1 2210
box -4 -6 356 206
use INVX8  INVX8_5
timestamp 1743498307
transform -1 0 2312 0 1 2210
box -4 -6 84 206
use DFFSR  DFFSR_162
timestamp 1743498307
transform 1 0 2312 0 1 2210
box -4 -6 356 206
use NAND2X1  NAND2X1_174
timestamp 1743498307
transform -1 0 2712 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_173
timestamp 1743498307
transform -1 0 2760 0 1 2210
box -4 -6 52 206
use INVX2  INVX2_10
timestamp 1743498307
transform 1 0 2760 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_445
timestamp 1743498307
transform -1 0 2856 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_180
timestamp 1743498307
transform -1 0 2888 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_457
timestamp 1743498307
transform -1 0 2952 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_456
timestamp 1743498307
transform 1 0 2952 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_172
timestamp 1743498307
transform 1 0 3016 0 1 2210
box -4 -6 52 206
use FILL  FILL_11_1_0
timestamp 1743498307
transform 1 0 3064 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_1
timestamp 1743498307
transform 1 0 3080 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_2
timestamp 1743498307
transform 1 0 3096 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_458
timestamp 1743498307
transform 1 0 3112 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_64
timestamp 1743498307
transform 1 0 3176 0 1 2210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_4
timestamp 1743498307
transform -1 0 3384 0 1 2210
box -4 -6 148 206
use NAND3X1  NAND3X1_58
timestamp 1743498307
transform 1 0 3384 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_61
timestamp 1743498307
transform 1 0 3448 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_55
timestamp 1743498307
transform 1 0 3512 0 1 2210
box -4 -6 68 206
use MUX2X1  MUX2X1_121
timestamp 1743498307
transform 1 0 3576 0 1 2210
box -4 -6 100 206
use DFFSR  DFFSR_143
timestamp 1743498307
transform 1 0 3672 0 1 2210
box -4 -6 356 206
use INVX1  INVX1_176
timestamp 1743498307
transform -1 0 4056 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_160
timestamp 1743498307
transform -1 0 4104 0 1 2210
box -4 -6 52 206
use BUFX4  BUFX4_3
timestamp 1743498307
transform 1 0 4104 0 1 2210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_12
timestamp 1743498307
transform -1 0 4312 0 1 2210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_41
timestamp 1743498307
transform 1 0 4312 0 1 2210
box -4 -6 148 206
use AOI22X1  AOI22X1_12
timestamp 1743498307
transform 1 0 4456 0 1 2210
box -4 -6 84 206
use AOI22X1  AOI22X1_11
timestamp 1743498307
transform -1 0 4616 0 1 2210
box -4 -6 84 206
use FILL  FILL_11_2_0
timestamp 1743498307
transform 1 0 4616 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_1
timestamp 1743498307
transform 1 0 4632 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_2
timestamp 1743498307
transform 1 0 4648 0 1 2210
box -4 -6 20 206
use NAND2X1  NAND2X1_153
timestamp 1743498307
transform 1 0 4664 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_45
timestamp 1743498307
transform 1 0 4712 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_154
timestamp 1743498307
transform 1 0 4776 0 1 2210
box -4 -6 52 206
use AOI22X1  AOI22X1_1
timestamp 1743498307
transform 1 0 4824 0 1 2210
box -4 -6 84 206
use NAND3X1  NAND3X1_39
timestamp 1743498307
transform -1 0 4968 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_9
timestamp 1743498307
transform -1 0 5032 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_37
timestamp 1743498307
transform -1 0 5096 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_38
timestamp 1743498307
transform -1 0 5160 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_36
timestamp 1743498307
transform 1 0 5160 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_33
timestamp 1743498307
transform 1 0 5224 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_32
timestamp 1743498307
transform 1 0 5288 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_30
timestamp 1743498307
transform -1 0 5416 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_29
timestamp 1743498307
transform -1 0 5480 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_138
timestamp 1743498307
transform -1 0 5528 0 1 2210
box -4 -6 52 206
use INVX2  INVX2_7
timestamp 1743498307
transform 1 0 5528 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_34
timestamp 1743498307
transform 1 0 5560 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_137
timestamp 1743498307
transform -1 0 5672 0 1 2210
box -4 -6 52 206
use DFFSR  DFFSR_138
timestamp 1743498307
transform -1 0 6024 0 1 2210
box -4 -6 356 206
use OAI21X1  OAI21X1_374
timestamp 1743498307
transform 1 0 6024 0 1 2210
box -4 -6 68 206
use FILL  FILL_12_1
timestamp 1743498307
transform 1 0 6088 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1743498307
transform 1 0 6104 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_3
timestamp 1743498307
transform 1 0 6120 0 1 2210
box -4 -6 20 206
use DFFSR  DFFSR_86
timestamp 1743498307
transform 1 0 8 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_10
timestamp 1743498307
transform -1 0 392 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_82
timestamp 1743498307
transform 1 0 392 0 -1 2610
box -4 -6 356 206
use NOR2X1  NOR2X1_61
timestamp 1743498307
transform 1 0 744 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_17
timestamp 1743498307
transform -1 0 856 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_7
timestamp 1743498307
transform -1 0 888 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_56
timestamp 1743498307
transform -1 0 936 0 -1 2610
box -4 -6 52 206
use DFFSR  DFFSR_174
timestamp 1743498307
transform -1 0 1288 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_6
timestamp 1743498307
transform -1 0 1320 0 -1 2610
box -4 -6 36 206
use BUFX4  BUFX4_67
timestamp 1743498307
transform -1 0 1384 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_0_0
timestamp 1743498307
transform -1 0 1400 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_1
timestamp 1743498307
transform -1 0 1416 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_2
timestamp 1743498307
transform -1 0 1432 0 -1 2610
box -4 -6 20 206
use DFFSR  DFFSR_170
timestamp 1743498307
transform -1 0 1784 0 -1 2610
box -4 -6 356 206
use NAND2X1  NAND2X1_161
timestamp 1743498307
transform 1 0 1784 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_446
timestamp 1743498307
transform -1 0 1896 0 -1 2610
box -4 -6 68 206
use INVX4  INVX4_3
timestamp 1743498307
transform -1 0 1944 0 -1 2610
box -4 -6 52 206
use DFFSR  DFFSR_146
timestamp 1743498307
transform 1 0 1944 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_179
timestamp 1743498307
transform 1 0 2296 0 -1 2610
box -4 -6 36 206
use MUX2X1  MUX2X1_124
timestamp 1743498307
transform -1 0 2424 0 -1 2610
box -4 -6 100 206
use BUFX4  BUFX4_71
timestamp 1743498307
transform -1 0 2488 0 -1 2610
box -4 -6 68 206
use DFFSR  DFFSR_166
timestamp 1743498307
transform -1 0 2840 0 -1 2610
box -4 -6 356 206
use OAI22X1  OAI22X1_8
timestamp 1743498307
transform -1 0 2920 0 -1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_449
timestamp 1743498307
transform -1 0 2984 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_166
timestamp 1743498307
transform 1 0 2984 0 -1 2610
box -4 -6 52 206
use FILL  FILL_12_1_0
timestamp 1743498307
transform 1 0 3032 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_1
timestamp 1743498307
transform 1 0 3048 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_2
timestamp 1743498307
transform 1 0 3064 0 -1 2610
box -4 -6 20 206
use OR2X2  OR2X2_14
timestamp 1743498307
transform 1 0 3080 0 -1 2610
box -4 -6 68 206
use BUFX4  BUFX4_9
timestamp 1743498307
transform -1 0 3208 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_448
timestamp 1743498307
transform -1 0 3272 0 -1 2610
box -4 -6 68 206
use OAI22X1  OAI22X1_7
timestamp 1743498307
transform -1 0 3352 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_163
timestamp 1743498307
transform -1 0 3400 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_60
timestamp 1743498307
transform 1 0 3400 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_1
timestamp 1743498307
transform 1 0 3464 0 -1 2610
box -4 -6 52 206
use DFFSR  DFFSR_144
timestamp 1743498307
transform 1 0 3512 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_177
timestamp 1743498307
transform -1 0 3896 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_63
timestamp 1743498307
transform 1 0 3896 0 -1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_10
timestamp 1743498307
transform -1 0 4040 0 -1 2610
box -4 -6 84 206
use AOI22X1  AOI22X1_4
timestamp 1743498307
transform -1 0 4120 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_149
timestamp 1743498307
transform 1 0 4120 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_42
timestamp 1743498307
transform 1 0 4168 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_150
timestamp 1743498307
transform -1 0 4280 0 -1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_15
timestamp 1743498307
transform 1 0 4280 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_156
timestamp 1743498307
transform 1 0 4360 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_155
timestamp 1743498307
transform -1 0 4456 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_48
timestamp 1743498307
transform 1 0 4456 0 -1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_5
timestamp 1743498307
transform -1 0 4600 0 -1 2610
box -4 -6 84 206
use FILL  FILL_12_2_0
timestamp 1743498307
transform -1 0 4616 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_1
timestamp 1743498307
transform -1 0 4632 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_2
timestamp 1743498307
transform -1 0 4648 0 -1 2610
box -4 -6 20 206
use AOI22X1  AOI22X1_13
timestamp 1743498307
transform -1 0 4728 0 -1 2610
box -4 -6 84 206
use NAND3X1  NAND3X1_46
timestamp 1743498307
transform 1 0 4728 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_48
timestamp 1743498307
transform 1 0 4792 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_49
timestamp 1743498307
transform -1 0 4888 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_154
timestamp 1743498307
transform -1 0 4920 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_153
timestamp 1743498307
transform -1 0 4952 0 -1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_5
timestamp 1743498307
transform 1 0 4952 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_135
timestamp 1743498307
transform -1 0 5064 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_31
timestamp 1743498307
transform -1 0 5128 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_47
timestamp 1743498307
transform -1 0 5176 0 -1 2610
box -4 -6 52 206
use OAI22X1  OAI22X1_1
timestamp 1743498307
transform -1 0 5256 0 -1 2610
box -4 -6 84 206
use OAI22X1  OAI22X1_3
timestamp 1743498307
transform -1 0 5336 0 -1 2610
box -4 -6 84 206
use INVX1  INVX1_149
timestamp 1743498307
transform 1 0 5336 0 -1 2610
box -4 -6 36 206
use OAI22X1  OAI22X1_4
timestamp 1743498307
transform -1 0 5448 0 -1 2610
box -4 -6 84 206
use INVX2  INVX2_5
timestamp 1743498307
transform 1 0 5448 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_425
timestamp 1743498307
transform 1 0 5480 0 -1 2610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_37
timestamp 1743498307
transform 1 0 5544 0 -1 2610
box -4 -6 148 206
use DFFSR  DFFSR_48
timestamp 1743498307
transform -1 0 6040 0 -1 2610
box -4 -6 356 206
use BUFX2  BUFX2_24
timestamp 1743498307
transform 1 0 6040 0 -1 2610
box -4 -6 52 206
use FILL  FILL_13_1
timestamp 1743498307
transform -1 0 6104 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_2
timestamp 1743498307
transform -1 0 6120 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_3
timestamp 1743498307
transform -1 0 6136 0 -1 2610
box -4 -6 20 206
use DFFSR  DFFSR_178
timestamp 1743498307
transform 1 0 8 0 1 2610
box -4 -6 356 206
use DFFSR  DFFSR_140
timestamp 1743498307
transform -1 0 712 0 1 2610
box -4 -6 356 206
use NOR2X1  NOR2X1_60
timestamp 1743498307
transform 1 0 712 0 1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_16
timestamp 1743498307
transform -1 0 824 0 1 2610
box -4 -6 68 206
use DFFSR  DFFSR_155
timestamp 1743498307
transform -1 0 1176 0 1 2610
box -4 -6 356 206
use AOI21X1  AOI21X1_12
timestamp 1743498307
transform -1 0 1240 0 1 2610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_31
timestamp 1743498307
transform -1 0 1384 0 1 2610
box -4 -6 148 206
use CLKBUF1  CLKBUF1_17
timestamp 1743498307
transform 1 0 1384 0 1 2610
box -4 -6 148 206
use FILL  FILL_13_0_0
timestamp 1743498307
transform 1 0 1528 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_1
timestamp 1743498307
transform 1 0 1544 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_2
timestamp 1743498307
transform 1 0 1560 0 1 2610
box -4 -6 20 206
use BUFX4  BUFX4_66
timestamp 1743498307
transform 1 0 1576 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_55
timestamp 1743498307
transform -1 0 1688 0 1 2610
box -4 -6 52 206
use OR2X2  OR2X2_13
timestamp 1743498307
transform -1 0 1752 0 1 2610
box -4 -6 68 206
use DFFSR  DFFSR_160
timestamp 1743498307
transform 1 0 1752 0 1 2610
box -4 -6 356 206
use INVX2  INVX2_8
timestamp 1743498307
transform -1 0 2136 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_167
timestamp 1743498307
transform 1 0 2136 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_168
timestamp 1743498307
transform 1 0 2184 0 1 2610
box -4 -6 52 206
use INVX8  INVX8_9
timestamp 1743498307
transform -1 0 2312 0 1 2610
box -4 -6 84 206
use DFFSR  DFFSR_141
timestamp 1743498307
transform 1 0 2312 0 1 2610
box -4 -6 356 206
use MUX2X1  MUX2X1_119
timestamp 1743498307
transform 1 0 2664 0 1 2610
box -4 -6 100 206
use INVX1  INVX1_174
timestamp 1743498307
transform -1 0 2792 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_453
timestamp 1743498307
transform -1 0 2856 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_452
timestamp 1743498307
transform 1 0 2856 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_181
timestamp 1743498307
transform 1 0 2920 0 1 2610
box -4 -6 36 206
use MUX2X1  MUX2X1_123
timestamp 1743498307
transform 1 0 2952 0 1 2610
box -4 -6 100 206
use FILL  FILL_13_1_0
timestamp 1743498307
transform 1 0 3048 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_1
timestamp 1743498307
transform 1 0 3064 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_2
timestamp 1743498307
transform 1 0 3080 0 1 2610
box -4 -6 20 206
use DFFSR  DFFSR_145
timestamp 1743498307
transform 1 0 3096 0 1 2610
box -4 -6 356 206
use INVX1  INVX1_178
timestamp 1743498307
transform -1 0 3480 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_463
timestamp 1743498307
transform -1 0 3544 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_462
timestamp 1743498307
transform 1 0 3544 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_185
timestamp 1743498307
transform -1 0 3640 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_181
timestamp 1743498307
transform -1 0 3688 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_71
timestamp 1743498307
transform 1 0 3688 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_70
timestamp 1743498307
transform 1 0 3752 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_67
timestamp 1743498307
transform 1 0 3816 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_69
timestamp 1743498307
transform 1 0 3880 0 1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_7
timestamp 1743498307
transform 1 0 3944 0 1 2610
box -4 -6 84 206
use AOI22X1  AOI22X1_2
timestamp 1743498307
transform 1 0 4024 0 1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_148
timestamp 1743498307
transform 1 0 4104 0 1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_3
timestamp 1743498307
transform -1 0 4232 0 1 2610
box -4 -6 84 206
use AOI22X1  AOI22X1_6
timestamp 1743498307
transform -1 0 4312 0 1 2610
box -4 -6 84 206
use NAND3X1  NAND3X1_44
timestamp 1743498307
transform 1 0 4312 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_50
timestamp 1743498307
transform -1 0 4440 0 1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_14
timestamp 1743498307
transform -1 0 4520 0 1 2610
box -4 -6 84 206
use NAND3X1  NAND3X1_43
timestamp 1743498307
transform -1 0 4584 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_2_0
timestamp 1743498307
transform 1 0 4584 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_1
timestamp 1743498307
transform 1 0 4600 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_2
timestamp 1743498307
transform 1 0 4616 0 1 2610
box -4 -6 20 206
use NAND3X1  NAND3X1_41
timestamp 1743498307
transform 1 0 4632 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_49
timestamp 1743498307
transform 1 0 4696 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_40
timestamp 1743498307
transform 1 0 4760 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_41
timestamp 1743498307
transform -1 0 4872 0 1 2610
box -4 -6 52 206
use OAI22X1  OAI22X1_5
timestamp 1743498307
transform -1 0 4952 0 1 2610
box -4 -6 84 206
use AOI21X1  AOI21X1_7
timestamp 1743498307
transform 1 0 4952 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_42
timestamp 1743498307
transform 1 0 5016 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_427
timestamp 1743498307
transform -1 0 5128 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_43
timestamp 1743498307
transform 1 0 5128 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_44
timestamp 1743498307
transform -1 0 5224 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_428
timestamp 1743498307
transform 1 0 5224 0 1 2610
box -4 -6 68 206
use OAI22X1  OAI22X1_2
timestamp 1743498307
transform 1 0 5288 0 1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_133
timestamp 1743498307
transform -1 0 5416 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_147
timestamp 1743498307
transform -1 0 5448 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_134
timestamp 1743498307
transform -1 0 5496 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_136
timestamp 1743498307
transform -1 0 5544 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_250
timestamp 1743498307
transform 1 0 5544 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_76
timestamp 1743498307
transform 1 0 5608 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_267
timestamp 1743498307
transform 1 0 5656 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_84
timestamp 1743498307
transform 1 0 5720 0 1 2610
box -4 -6 52 206
use DFFSR  DFFSR_44
timestamp 1743498307
transform -1 0 6120 0 1 2610
box -4 -6 356 206
use FILL  FILL_14_1
timestamp 1743498307
transform 1 0 6120 0 1 2610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_28
timestamp 1743498307
transform 1 0 8 0 -1 3010
box -4 -6 148 206
use DFFSR  DFFSR_177
timestamp 1743498307
transform 1 0 152 0 -1 3010
box -4 -6 356 206
use NOR2X1  NOR2X1_59
timestamp 1743498307
transform 1 0 504 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_15
timestamp 1743498307
transform -1 0 616 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_176
timestamp 1743498307
transform 1 0 616 0 -1 3010
box -4 -6 356 206
use NOR2X1  NOR2X1_58
timestamp 1743498307
transform 1 0 968 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_14
timestamp 1743498307
transform -1 0 1080 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_164
timestamp 1743498307
transform 1 0 1080 0 -1 3010
box -4 -6 36 206
use MUX2X1  MUX2X1_109
timestamp 1743498307
transform 1 0 1112 0 -1 3010
box -4 -6 100 206
use DFFSR  DFFSR_175
timestamp 1743498307
transform -1 0 1560 0 -1 3010
box -4 -6 356 206
use FILL  FILL_14_0_0
timestamp 1743498307
transform 1 0 1560 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_1
timestamp 1743498307
transform 1 0 1576 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_2
timestamp 1743498307
transform 1 0 1592 0 -1 3010
box -4 -6 20 206
use INVX1  INVX1_158
timestamp 1743498307
transform 1 0 1608 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_444
timestamp 1743498307
transform 1 0 1640 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_165
timestamp 1743498307
transform 1 0 1704 0 -1 3010
box -4 -6 356 206
use INVX2  INVX2_13
timestamp 1743498307
transform 1 0 2056 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_182
timestamp 1743498307
transform 1 0 2088 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_183
timestamp 1743498307
transform 1 0 2136 0 -1 3010
box -4 -6 52 206
use DFFSR  DFFSR_142
timestamp 1743498307
transform 1 0 2184 0 -1 3010
box -4 -6 356 206
use INVX1  INVX1_175
timestamp 1743498307
transform 1 0 2536 0 -1 3010
box -4 -6 36 206
use MUX2X1  MUX2X1_120
timestamp 1743498307
transform -1 0 2664 0 -1 3010
box -4 -6 100 206
use DFFSR  DFFSR_161
timestamp 1743498307
transform 1 0 2664 0 -1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_170
timestamp 1743498307
transform 1 0 3016 0 -1 3010
box -4 -6 52 206
use FILL  FILL_14_1_0
timestamp 1743498307
transform 1 0 3064 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_1
timestamp 1743498307
transform 1 0 3080 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_2
timestamp 1743498307
transform 1 0 3096 0 -1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_171
timestamp 1743498307
transform 1 0 3112 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_169
timestamp 1743498307
transform 1 0 3160 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_455
timestamp 1743498307
transform 1 0 3208 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_454
timestamp 1743498307
transform 1 0 3272 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_164
timestamp 1743498307
transform 1 0 3336 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_54
timestamp 1743498307
transform 1 0 3384 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_160
timestamp 1743498307
transform -1 0 3464 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_53
timestamp 1743498307
transform 1 0 3464 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_54
timestamp 1743498307
transform 1 0 3528 0 -1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_122
timestamp 1743498307
transform 1 0 3592 0 -1 3010
box -4 -6 100 206
use NAND2X1  NAND2X1_178
timestamp 1743498307
transform -1 0 3736 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_68
timestamp 1743498307
transform 1 0 3736 0 -1 3010
box -4 -6 68 206
use INVX4  INVX4_4
timestamp 1743498307
transform 1 0 3800 0 -1 3010
box -4 -6 52 206
use AOI22X1  AOI22X1_18
timestamp 1743498307
transform -1 0 3928 0 -1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_151
timestamp 1743498307
transform 1 0 3928 0 -1 3010
box -4 -6 52 206
use DFFSR  DFFSR_134
timestamp 1743498307
transform -1 0 4328 0 -1 3010
box -4 -6 356 206
use AOI22X1  AOI22X1_8
timestamp 1743498307
transform -1 0 4408 0 -1 3010
box -4 -6 84 206
use AOI22X1  AOI22X1_16
timestamp 1743498307
transform -1 0 4488 0 -1 3010
box -4 -6 84 206
use INVX1  INVX1_151
timestamp 1743498307
transform -1 0 4520 0 -1 3010
box -4 -6 36 206
use INVX1  INVX1_152
timestamp 1743498307
transform -1 0 4552 0 -1 3010
box -4 -6 36 206
use FILL  FILL_14_2_0
timestamp 1743498307
transform 1 0 4552 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_1
timestamp 1743498307
transform 1 0 4568 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_2
timestamp 1743498307
transform 1 0 4584 0 -1 3010
box -4 -6 20 206
use NAND3X1  NAND3X1_51
timestamp 1743498307
transform 1 0 4600 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_47
timestamp 1743498307
transform 1 0 4664 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_10
timestamp 1743498307
transform 1 0 4728 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_158
timestamp 1743498307
transform -1 0 4840 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_11
timestamp 1743498307
transform 1 0 4840 0 -1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_52
timestamp 1743498307
transform 1 0 4904 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_146
timestamp 1743498307
transform 1 0 4952 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_430
timestamp 1743498307
transform -1 0 5064 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_429
timestamp 1743498307
transform 1 0 5064 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_145
timestamp 1743498307
transform 1 0 5128 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_53
timestamp 1743498307
transform -1 0 5224 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_46
timestamp 1743498307
transform 1 0 5224 0 -1 3010
box -4 -6 52 206
use INVX2  INVX2_6
timestamp 1743498307
transform 1 0 5272 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_246
timestamp 1743498307
transform -1 0 5368 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_47
timestamp 1743498307
transform -1 0 5720 0 -1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_127
timestamp 1743498307
transform 1 0 5720 0 -1 3010
box -4 -6 52 206
use DFFSR  DFFSR_105
timestamp 1743498307
transform 1 0 5768 0 -1 3010
box -4 -6 356 206
use FILL  FILL_15_1
timestamp 1743498307
transform -1 0 6136 0 -1 3010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_20
timestamp 1743498307
transform 1 0 8 0 1 3010
box -4 -6 148 206
use DFFSR  DFFSR_156
timestamp 1743498307
transform 1 0 152 0 1 3010
box -4 -6 356 206
use DFFSR  DFFSR_158
timestamp 1743498307
transform -1 0 856 0 1 3010
box -4 -6 356 206
use MUX2X1  MUX2X1_112
timestamp 1743498307
transform -1 0 952 0 1 3010
box -4 -6 100 206
use MUX2X1  MUX2X1_111
timestamp 1743498307
transform 1 0 952 0 1 3010
box -4 -6 100 206
use INVX1  INVX1_166
timestamp 1743498307
transform -1 0 1080 0 1 3010
box -4 -6 36 206
use DFFSR  DFFSR_157
timestamp 1743498307
transform -1 0 1432 0 1 3010
box -4 -6 356 206
use NOR2X1  NOR2X1_57
timestamp 1743498307
transform 1 0 1432 0 1 3010
box -4 -6 52 206
use FILL  FILL_15_0_0
timestamp 1743498307
transform -1 0 1496 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_1
timestamp 1743498307
transform -1 0 1512 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_2
timestamp 1743498307
transform -1 0 1528 0 1 3010
box -4 -6 20 206
use AOI21X1  AOI21X1_13
timestamp 1743498307
transform -1 0 1592 0 1 3010
box -4 -6 68 206
use DFFSR  DFFSR_173
timestamp 1743498307
transform -1 0 1944 0 1 3010
box -4 -6 356 206
use NAND3X1  NAND3X1_52
timestamp 1743498307
transform 1 0 1944 0 1 3010
box -4 -6 68 206
use DFFSR  DFFSR_163
timestamp 1743498307
transform 1 0 2008 0 1 3010
box -4 -6 356 206
use INVX2  INVX2_11
timestamp 1743498307
transform -1 0 2392 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_176
timestamp 1743498307
transform 1 0 2392 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_177
timestamp 1743498307
transform 1 0 2440 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_69
timestamp 1743498307
transform 1 0 2488 0 1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_117
timestamp 1743498307
transform -1 0 2648 0 1 3010
box -4 -6 100 206
use MUX2X1  MUX2X1_115
timestamp 1743498307
transform 1 0 2648 0 1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_459
timestamp 1743498307
transform -1 0 2808 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_175
timestamp 1743498307
transform 1 0 2808 0 1 3010
box -4 -6 52 206
use INVX2  INVX2_12
timestamp 1743498307
transform -1 0 2888 0 1 3010
box -4 -6 36 206
use INVX2  INVX2_9
timestamp 1743498307
transform -1 0 2920 0 1 3010
box -4 -6 36 206
use FILL  FILL_15_1_0
timestamp 1743498307
transform -1 0 2936 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_1
timestamp 1743498307
transform -1 0 2952 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_2
timestamp 1743498307
transform -1 0 2968 0 1 3010
box -4 -6 20 206
use DFFSR  DFFSR_164
timestamp 1743498307
transform -1 0 3320 0 1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_179
timestamp 1743498307
transform 1 0 3320 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_180
timestamp 1743498307
transform 1 0 3368 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_461
timestamp 1743498307
transform -1 0 3480 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_460
timestamp 1743498307
transform -1 0 3544 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_184
timestamp 1743498307
transform -1 0 3576 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_57
timestamp 1743498307
transform 1 0 3576 0 1 3010
box -4 -6 68 206
use INVX4  INVX4_5
timestamp 1743498307
transform -1 0 3688 0 1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_66
timestamp 1743498307
transform 1 0 3688 0 1 3010
box -4 -6 68 206
use AOI22X1  AOI22X1_17
timestamp 1743498307
transform -1 0 3832 0 1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_157
timestamp 1743498307
transform 1 0 3832 0 1 3010
box -4 -6 52 206
use AOI22X1  AOI22X1_9
timestamp 1743498307
transform 1 0 3880 0 1 3010
box -4 -6 84 206
use OAI21X1  OAI21X1_438
timestamp 1743498307
transform 1 0 3960 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_436
timestamp 1743498307
transform 1 0 4024 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_155
timestamp 1743498307
transform -1 0 4120 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_437
timestamp 1743498307
transform -1 0 4184 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_439
timestamp 1743498307
transform 1 0 4184 0 1 3010
box -4 -6 68 206
use DFFSR  DFFSR_135
timestamp 1743498307
transform 1 0 4248 0 1 3010
box -4 -6 356 206
use FILL  FILL_15_2_0
timestamp 1743498307
transform 1 0 4600 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_1
timestamp 1743498307
transform 1 0 4616 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_2
timestamp 1743498307
transform 1 0 4632 0 1 3010
box -4 -6 20 206
use OAI21X1  OAI21X1_431
timestamp 1743498307
transform 1 0 4648 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_150
timestamp 1743498307
transform 1 0 4712 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_433
timestamp 1743498307
transform 1 0 4744 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_442
timestamp 1743498307
transform -1 0 4872 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_435
timestamp 1743498307
transform -1 0 4936 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_8
timestamp 1743498307
transform -1 0 5000 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_441
timestamp 1743498307
transform 1 0 5000 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_440
timestamp 1743498307
transform 1 0 5064 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_159
timestamp 1743498307
transform -1 0 5176 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_144
timestamp 1743498307
transform -1 0 5224 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_242
timestamp 1743498307
transform -1 0 5288 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_2
timestamp 1743498307
transform 1 0 5288 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_74
timestamp 1743498307
transform 1 0 5336 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_26
timestamp 1743498307
transform 1 0 5384 0 1 3010
box -4 -6 68 206
use INVX4  INVX4_2
timestamp 1743498307
transform 1 0 5448 0 1 3010
box -4 -6 52 206
use DFFSR  DFFSR_108
timestamp 1743498307
transform 1 0 5496 0 1 3010
box -4 -6 356 206
use OAI21X1  OAI21X1_395
timestamp 1743498307
transform -1 0 5912 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_125
timestamp 1743498307
transform -1 0 5944 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_392
timestamp 1743498307
transform -1 0 6008 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_122
timestamp 1743498307
transform -1 0 6040 0 1 3010
box -4 -6 36 206
use BUFX2  BUFX2_17
timestamp 1743498307
transform 1 0 6040 0 1 3010
box -4 -6 52 206
use FILL  FILL_16_1
timestamp 1743498307
transform 1 0 6088 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_2
timestamp 1743498307
transform 1 0 6104 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_3
timestamp 1743498307
transform 1 0 6120 0 1 3010
box -4 -6 20 206
use DFFSR  DFFSR_127
timestamp 1743498307
transform 1 0 8 0 -1 3410
box -4 -6 356 206
use BUFX4  BUFX4_2
timestamp 1743498307
transform -1 0 424 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_165
timestamp 1743498307
transform -1 0 456 0 -1 3410
box -4 -6 36 206
use MUX2X1  MUX2X1_110
timestamp 1743498307
transform -1 0 552 0 -1 3410
box -4 -6 100 206
use INVX1  INVX1_167
timestamp 1743498307
transform 1 0 552 0 -1 3410
box -4 -6 36 206
use DFFSR  DFFSR_153
timestamp 1743498307
transform -1 0 936 0 -1 3410
box -4 -6 356 206
use INVX1  INVX1_162
timestamp 1743498307
transform 1 0 936 0 -1 3410
box -4 -6 36 206
use MUX2X1  MUX2X1_107
timestamp 1743498307
transform -1 0 1064 0 -1 3410
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_86
timestamp 1743498307
transform 1 0 1064 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_89
timestamp 1743498307
transform 1 0 1256 0 -1 3410
box -4 -6 196 206
use INVX1  INVX1_78
timestamp 1743498307
transform -1 0 1480 0 -1 3410
box -4 -6 36 206
use FILL  FILL_16_0_0
timestamp 1743498307
transform -1 0 1496 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_1
timestamp 1743498307
transform -1 0 1512 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_2
timestamp 1743498307
transform -1 0 1528 0 -1 3410
box -4 -6 20 206
use DFFSR  DFFSR_154
timestamp 1743498307
transform -1 0 1880 0 -1 3410
box -4 -6 356 206
use BUFX4  BUFX4_70
timestamp 1743498307
transform 1 0 1880 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_151
timestamp 1743498307
transform 1 0 1944 0 -1 3410
box -4 -6 356 206
use INVX8  INVX8_8
timestamp 1743498307
transform 1 0 2296 0 -1 3410
box -4 -6 84 206
use INVX1  INVX1_172
timestamp 1743498307
transform 1 0 2376 0 -1 3410
box -4 -6 36 206
use DFFSR  DFFSR_149
timestamp 1743498307
transform 1 0 2408 0 -1 3410
box -4 -6 356 206
use INVX1  INVX1_170
timestamp 1743498307
transform -1 0 2792 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_65
timestamp 1743498307
transform -1 0 2856 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_59
timestamp 1743498307
transform -1 0 2920 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_56
timestamp 1743498307
transform -1 0 2984 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_62
timestamp 1743498307
transform -1 0 3048 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_1_0
timestamp 1743498307
transform -1 0 3064 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_1
timestamp 1743498307
transform -1 0 3080 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_2
timestamp 1743498307
transform -1 0 3096 0 -1 3410
box -4 -6 20 206
use BUFX4  BUFX4_7
timestamp 1743498307
transform -1 0 3160 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_162
timestamp 1743498307
transform 1 0 3160 0 -1 3410
box -4 -6 52 206
use OAI22X1  OAI22X1_6
timestamp 1743498307
transform 1 0 3208 0 -1 3410
box -4 -6 84 206
use OAI21X1  OAI21X1_447
timestamp 1743498307
transform -1 0 3352 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_169
timestamp 1743498307
transform -1 0 3704 0 -1 3410
box -4 -6 356 206
use OAI21X1  OAI21X1_451
timestamp 1743498307
transform -1 0 3768 0 -1 3410
box -4 -6 68 206
use OAI22X1  OAI22X1_9
timestamp 1743498307
transform -1 0 3848 0 -1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_165
timestamp 1743498307
transform -1 0 3896 0 -1 3410
box -4 -6 52 206
use BUFX4  BUFX4_8
timestamp 1743498307
transform -1 0 3960 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_133
timestamp 1743498307
transform -1 0 4312 0 -1 3410
box -4 -6 356 206
use NAND2X1  NAND2X1_152
timestamp 1743498307
transform -1 0 4360 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_156
timestamp 1743498307
transform 1 0 4360 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_443
timestamp 1743498307
transform 1 0 4392 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_434
timestamp 1743498307
transform 1 0 4456 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_142
timestamp 1743498307
transform 1 0 4520 0 -1 3410
box -4 -6 52 206
use FILL  FILL_16_2_0
timestamp 1743498307
transform 1 0 4568 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_1
timestamp 1743498307
transform 1 0 4584 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_2
timestamp 1743498307
transform 1 0 4600 0 -1 3410
box -4 -6 20 206
use AOI21X1  AOI21X1_6
timestamp 1743498307
transform 1 0 4616 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_50
timestamp 1743498307
transform 1 0 4680 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_51
timestamp 1743498307
transform -1 0 4776 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_432
timestamp 1743498307
transform -1 0 4840 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_143
timestamp 1743498307
transform 1 0 4840 0 -1 3410
box -4 -6 52 206
use INVX4  INVX4_1
timestamp 1743498307
transform 1 0 4888 0 -1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_35
timestamp 1743498307
transform 1 0 4936 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_45
timestamp 1743498307
transform -1 0 5048 0 -1 3410
box -4 -6 52 206
use DFFSR  DFFSR_46
timestamp 1743498307
transform -1 0 5400 0 -1 3410
box -4 -6 356 206
use DFFSR  DFFSR_42
timestamp 1743498307
transform 1 0 5400 0 -1 3410
box -4 -6 356 206
use NAND2X1  NAND2X1_125
timestamp 1743498307
transform -1 0 5800 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_393
timestamp 1743498307
transform -1 0 5864 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_123
timestamp 1743498307
transform -1 0 5896 0 -1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_124
timestamp 1743498307
transform 1 0 5896 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_394
timestamp 1743498307
transform -1 0 6008 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_124
timestamp 1743498307
transform -1 0 6040 0 -1 3410
box -4 -6 36 206
use INVX8  INVX8_7
timestamp 1743498307
transform -1 0 6120 0 -1 3410
box -4 -6 84 206
use FILL  FILL_17_1
timestamp 1743498307
transform -1 0 6136 0 -1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_416
timestamp 1743498307
transform 1 0 136 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_418
timestamp 1743498307
transform 1 0 72 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_139
timestamp 1743498307
transform 1 0 40 0 -1 3810
box -4 -6 36 206
use INVX1  INVX1_140
timestamp 1743498307
transform 1 0 8 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_422
timestamp 1743498307
transform 1 0 40 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_142
timestamp 1743498307
transform 1 0 8 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_417
timestamp 1743498307
transform -1 0 392 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_421
timestamp 1743498307
transform 1 0 264 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_415
timestamp 1743498307
transform -1 0 264 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_124
timestamp 1743498307
transform 1 0 104 0 1 3410
box -4 -6 356 206
use OAI21X1  OAI21X1_275
timestamp 1743498307
transform -1 0 568 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_87
timestamp 1743498307
transform -1 0 504 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_284
timestamp 1743498307
transform -1 0 456 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_89
timestamp 1743498307
transform -1 0 568 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_82
timestamp 1743498307
transform -1 0 520 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_80
timestamp 1743498307
transform 1 0 456 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_305
timestamp 1743498307
transform -1 0 792 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_306
timestamp 1743498307
transform 1 0 664 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_94
timestamp 1743498307
transform 1 0 568 0 -1 3810
box -4 -6 100 206
use INVX1  INVX1_79
timestamp 1743498307
transform -1 0 600 0 1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_80
timestamp 1743498307
transform 1 0 600 0 1 3410
box -4 -6 196 206
use INVX1  INVX1_75
timestamp 1743498307
transform -1 0 824 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_86
timestamp 1743498307
transform -1 0 872 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_272
timestamp 1743498307
transform -1 0 936 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_281
timestamp 1743498307
transform -1 0 1000 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_81
timestamp 1743498307
transform -1 0 1032 0 1 3410
box -4 -6 36 206
use MUX2X1  MUX2X1_88
timestamp 1743498307
transform 1 0 1032 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_291
timestamp 1743498307
transform 1 0 792 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_292
timestamp 1743498307
transform -1 0 920 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_85
timestamp 1743498307
transform -1 0 1112 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_299
timestamp 1743498307
transform 1 0 1208 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_268
timestamp 1743498307
transform -1 0 1208 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_74
timestamp 1743498307
transform 1 0 1112 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_293
timestamp 1743498307
transform -1 0 1256 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_294
timestamp 1743498307
transform 1 0 1128 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_301
timestamp 1743498307
transform 1 0 1368 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_92
timestamp 1743498307
transform 1 0 1272 0 -1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_91
timestamp 1743498307
transform 1 0 1320 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_300
timestamp 1743498307
transform -1 0 1320 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_302
timestamp 1743498307
transform 1 0 1432 0 -1 3810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_26
timestamp 1743498307
transform 1 0 1416 0 1 3410
box -4 -6 148 206
use FILL  FILL_18_0_2
timestamp 1743498307
transform 1 0 1528 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_1
timestamp 1743498307
transform 1 0 1512 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_0
timestamp 1743498307
transform 1 0 1496 0 -1 3810
box -4 -6 20 206
use INVX1  INVX1_163
timestamp 1743498307
transform 1 0 1608 0 1 3410
box -4 -6 36 206
use FILL  FILL_17_0_2
timestamp 1743498307
transform 1 0 1592 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_1
timestamp 1743498307
transform 1 0 1576 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_0
timestamp 1743498307
transform 1 0 1560 0 1 3410
box -4 -6 20 206
use BUFX2  BUFX2_26
timestamp 1743498307
transform 1 0 1736 0 1 3410
box -4 -6 52 206
use MUX2X1  MUX2X1_108
timestamp 1743498307
transform -1 0 1736 0 1 3410
box -4 -6 100 206
use DFFSR  DFFSR_68
timestamp 1743498307
transform 1 0 1736 0 -1 3810
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_90
timestamp 1743498307
transform 1 0 1544 0 -1 3810
box -4 -6 196 206
use DFFSR  DFFSR_65
timestamp 1743498307
transform 1 0 1784 0 1 3410
box -4 -6 356 206
use BUFX4  BUFX4_87
timestamp 1743498307
transform -1 0 2200 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_100
timestamp 1743498307
transform -1 0 2136 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_343
timestamp 1743498307
transform -1 0 2200 0 -1 3810
box -4 -6 68 206
use INVX8  INVX8_4
timestamp 1743498307
transform -1 0 2280 0 1 3410
box -4 -6 84 206
use BUFX4  BUFX4_68
timestamp 1743498307
transform 1 0 2280 0 1 3410
box -4 -6 68 206
use DFFSR  DFFSR_147
timestamp 1743498307
transform 1 0 2344 0 1 3410
box -4 -6 356 206
use OAI21X1  OAI21X1_331
timestamp 1743498307
transform -1 0 2264 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_339
timestamp 1743498307
transform 1 0 2264 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_67
timestamp 1743498307
transform -1 0 2680 0 -1 3810
box -4 -6 356 206
use MUX2X1  MUX2X1_113
timestamp 1743498307
transform 1 0 2696 0 1 3410
box -4 -6 100 206
use INVX1  INVX1_168
timestamp 1743498307
transform -1 0 2824 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_55
timestamp 1743498307
transform 1 0 2824 0 1 3410
box -4 -6 36 206
use DFFSR  DFFSR_150
timestamp 1743498307
transform 1 0 2856 0 1 3410
box -4 -6 356 206
use BUFX4  BUFX4_6
timestamp 1743498307
transform -1 0 2744 0 -1 3810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_33
timestamp 1743498307
transform 1 0 2744 0 -1 3810
box -4 -6 148 206
use CLKBUF1  CLKBUF1_7
timestamp 1743498307
transform 1 0 2888 0 -1 3810
box -4 -6 148 206
use FILL  FILL_17_1_0
timestamp 1743498307
transform 1 0 3208 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_1
timestamp 1743498307
transform 1 0 3224 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_2
timestamp 1743498307
transform 1 0 3240 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_1_0
timestamp 1743498307
transform 1 0 3032 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_1
timestamp 1743498307
transform 1 0 3048 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_2
timestamp 1743498307
transform 1 0 3064 0 -1 3810
box -4 -6 20 206
use MUX2X1  MUX2X1_118
timestamp 1743498307
transform 1 0 3080 0 -1 3810
box -4 -6 100 206
use INVX1  INVX1_173
timestamp 1743498307
transform -1 0 3208 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_450
timestamp 1743498307
transform -1 0 3272 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_116
timestamp 1743498307
transform 1 0 3256 0 1 3410
box -4 -6 100 206
use INVX1  INVX1_171
timestamp 1743498307
transform -1 0 3384 0 1 3410
box -4 -6 36 206
use DFFSR  DFFSR_168
timestamp 1743498307
transform 1 0 3384 0 1 3410
box -4 -6 356 206
use INVX1  INVX1_161
timestamp 1743498307
transform -1 0 3304 0 -1 3810
box -4 -6 36 206
use MUX2X1  MUX2X1_114
timestamp 1743498307
transform 1 0 3304 0 -1 3810
box -4 -6 100 206
use INVX1  INVX1_169
timestamp 1743498307
transform -1 0 3432 0 -1 3810
box -4 -6 36 206
use DFFSR  DFFSR_148
timestamp 1743498307
transform 1 0 3432 0 -1 3810
box -4 -6 356 206
use INVX1  INVX1_148
timestamp 1743498307
transform 1 0 3736 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_141
timestamp 1743498307
transform 1 0 3768 0 1 3410
box -4 -6 52 206
use MUX2X1  MUX2X1_106
timestamp 1743498307
transform -1 0 3912 0 1 3410
box -4 -6 100 206
use MUX2X1  MUX2X1_105
timestamp 1743498307
transform -1 0 4008 0 1 3410
box -4 -6 100 206
use DFFSR  DFFSR_49
timestamp 1743498307
transform -1 0 4136 0 -1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_140
timestamp 1743498307
transform -1 0 4056 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_145
timestamp 1743498307
transform -1 0 4088 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_147
timestamp 1743498307
transform 1 0 4088 0 1 3410
box -4 -6 52 206
use DFFSR  DFFSR_137
timestamp 1743498307
transform -1 0 4488 0 1 3410
box -4 -6 356 206
use BUFX4  BUFX4_5
timestamp 1743498307
transform 1 0 4136 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_78
timestamp 1743498307
transform -1 0 4248 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_254
timestamp 1743498307
transform -1 0 4312 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_238
timestamp 1743498307
transform 1 0 4312 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_2_2
timestamp 1743498307
transform -1 0 4472 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_1
timestamp 1743498307
transform -1 0 4456 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_0
timestamp 1743498307
transform -1 0 4440 0 -1 3810
box -4 -6 20 206
use NAND2X1  NAND2X1_70
timestamp 1743498307
transform 1 0 4376 0 -1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_25
timestamp 1743498307
transform 1 0 4488 0 1 3410
box -4 -6 52 206
use FILL  FILL_17_2_2
timestamp 1743498307
transform -1 0 4584 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_1
timestamp 1743498307
transform -1 0 4568 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_0
timestamp 1743498307
transform -1 0 4552 0 1 3410
box -4 -6 20 206
use DFFSR  DFFSR_45
timestamp 1743498307
transform -1 0 4824 0 -1 3810
box -4 -6 356 206
use DFFSR  DFFSR_116
timestamp 1743498307
transform -1 0 4936 0 1 3410
box -4 -6 356 206
use DFFSR  DFFSR_118
timestamp 1743498307
transform 1 0 4936 0 1 3410
box -4 -6 356 206
use INVX1  INVX1_132
timestamp 1743498307
transform -1 0 4856 0 -1 3810
box -4 -6 36 206
use CLKBUF1  CLKBUF1_9
timestamp 1743498307
transform -1 0 5000 0 -1 3810
box -4 -6 148 206
use BUFX4  BUFX4_30
timestamp 1743498307
transform -1 0 5064 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_72
timestamp 1743498307
transform 1 0 5288 0 1 3410
box -4 -6 52 206
use BUFX4  BUFX4_29
timestamp 1743498307
transform -1 0 5400 0 1 3410
box -4 -6 68 206
use BUFX4  BUFX4_25
timestamp 1743498307
transform 1 0 5400 0 1 3410
box -4 -6 68 206
use BUFX4  BUFX4_28
timestamp 1743498307
transform -1 0 5128 0 -1 3810
box -4 -6 68 206
use BUFX4  BUFX4_24
timestamp 1743498307
transform -1 0 5192 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_40
timestamp 1743498307
transform -1 0 5544 0 -1 3810
box -4 -6 356 206
use INVX8  INVX8_3
timestamp 1743498307
transform 1 0 5464 0 1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_82
timestamp 1743498307
transform -1 0 5592 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_265
timestamp 1743498307
transform 1 0 5592 0 1 3410
box -4 -6 68 206
use DFFSR  DFFSR_106
timestamp 1743498307
transform 1 0 5656 0 1 3410
box -4 -6 356 206
use BUFX4  BUFX4_27
timestamp 1743498307
transform 1 0 5544 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_81
timestamp 1743498307
transform -1 0 5656 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_264
timestamp 1743498307
transform 1 0 5656 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_41
timestamp 1743498307
transform -1 0 6072 0 -1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_126
timestamp 1743498307
transform 1 0 6008 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_15
timestamp 1743498307
transform 1 0 6056 0 1 3410
box -4 -6 52 206
use FILL  FILL_18_1
timestamp 1743498307
transform 1 0 6104 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2
timestamp 1743498307
transform 1 0 6120 0 1 3410
box -4 -6 20 206
use BUFX2  BUFX2_16
timestamp 1743498307
transform 1 0 6072 0 -1 3810
box -4 -6 52 206
use FILL  FILL_19_1
timestamp 1743498307
transform -1 0 6136 0 -1 3810
box -4 -6 20 206
use DFFSR  DFFSR_125
timestamp 1743498307
transform 1 0 8 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_90
timestamp 1743498307
transform -1 0 408 0 1 3810
box -4 -6 52 206
use BUFX4  BUFX4_22
timestamp 1743498307
transform -1 0 472 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_83
timestamp 1743498307
transform 1 0 472 0 1 3810
box -4 -6 196 206
use BUFX4  BUFX4_19
timestamp 1743498307
transform 1 0 664 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_269
timestamp 1743498307
transform -1 0 792 0 1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_87
timestamp 1743498307
transform -1 0 888 0 1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_97
timestamp 1743498307
transform -1 0 984 0 1 3810
box -4 -6 100 206
use INVX1  INVX1_88
timestamp 1743498307
transform -1 0 1016 0 1 3810
box -4 -6 36 206
use BUFX4  BUFX4_83
timestamp 1743498307
transform -1 0 1080 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_34
timestamp 1743498307
transform -1 0 1128 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_77
timestamp 1743498307
transform 1 0 1128 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_323
timestamp 1743498307
transform 1 0 1320 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_324
timestamp 1743498307
transform -1 0 1448 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_45
timestamp 1743498307
transform -1 0 1512 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_0_0
timestamp 1743498307
transform 1 0 1512 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_1
timestamp 1743498307
transform 1 0 1528 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_2
timestamp 1743498307
transform 1 0 1544 0 1 3810
box -4 -6 20 206
use INVX1  INVX1_93
timestamp 1743498307
transform 1 0 1560 0 1 3810
box -4 -6 36 206
use BUFX4  BUFX4_20
timestamp 1743498307
transform -1 0 1656 0 1 3810
box -4 -6 68 206
use DFFSR  DFFSR_58
timestamp 1743498307
transform -1 0 2008 0 1 3810
box -4 -6 356 206
use INVX1  INVX1_95
timestamp 1743498307
transform 1 0 2008 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_106
timestamp 1743498307
transform -1 0 2088 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_110
timestamp 1743498307
transform -1 0 2136 0 1 3810
box -4 -6 52 206
use DFFSR  DFFSR_61
timestamp 1743498307
transform 1 0 2136 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_104
timestamp 1743498307
transform 1 0 2488 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_354
timestamp 1743498307
transform -1 0 2600 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_4
timestamp 1743498307
transform -1 0 2648 0 1 3810
box -4 -6 52 206
use DFFSR  DFFSR_64
timestamp 1743498307
transform 1 0 2648 0 1 3810
box -4 -6 356 206
use FILL  FILL_19_1_0
timestamp 1743498307
transform 1 0 3000 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_1
timestamp 1743498307
transform 1 0 3016 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_2
timestamp 1743498307
transform 1 0 3032 0 1 3810
box -4 -6 20 206
use DFFSR  DFFSR_152
timestamp 1743498307
transform 1 0 3048 0 1 3810
box -4 -6 356 206
use DFFSR  DFFSR_172
timestamp 1743498307
transform -1 0 3752 0 1 3810
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_62
timestamp 1743498307
transform 1 0 3752 0 1 3810
box -4 -6 196 206
use INVX1  INVX1_54
timestamp 1743498307
transform 1 0 3944 0 1 3810
box -4 -6 36 206
use INVX1  INVX1_51
timestamp 1743498307
transform 1 0 3976 0 1 3810
box -4 -6 36 206
use BUFX4  BUFX4_90
timestamp 1743498307
transform 1 0 4008 0 1 3810
box -4 -6 68 206
use DFFSR  DFFSR_50
timestamp 1743498307
transform -1 0 4424 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_80
timestamp 1743498307
transform -1 0 4472 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_258
timestamp 1743498307
transform -1 0 4536 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_2_0
timestamp 1743498307
transform 1 0 4536 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_1
timestamp 1743498307
transform 1 0 4552 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_2
timestamp 1743498307
transform 1 0 4568 0 1 3810
box -4 -6 20 206
use DFFSR  DFFSR_52
timestamp 1743498307
transform 1 0 4584 0 1 3810
box -4 -6 356 206
use CLKBUF1  CLKBUF1_19
timestamp 1743498307
transform -1 0 5080 0 1 3810
box -4 -6 148 206
use NOR2X1  NOR2X1_26
timestamp 1743498307
transform -1 0 5128 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_65
timestamp 1743498307
transform -1 0 5176 0 1 3810
box -4 -6 52 206
use DFFSR  DFFSR_57
timestamp 1743498307
transform 1 0 5176 0 1 3810
box -4 -6 356 206
use NOR2X1  NOR2X1_21
timestamp 1743498307
transform -1 0 5576 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_201
timestamp 1743498307
transform -1 0 5640 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_59
timestamp 1743498307
transform -1 0 5672 0 1 3810
box -4 -6 36 206
use OR2X2  OR2X2_6
timestamp 1743498307
transform -1 0 5736 0 1 3810
box -4 -6 68 206
use DFFSR  DFFSR_43
timestamp 1743498307
transform 1 0 5736 0 1 3810
box -4 -6 356 206
use FILL  FILL_20_1
timestamp 1743498307
transform 1 0 6088 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_2
timestamp 1743498307
transform 1 0 6104 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_3
timestamp 1743498307
transform 1 0 6120 0 1 3810
box -4 -6 20 206
use DFFSR  DFFSR_128
timestamp 1743498307
transform 1 0 8 0 -1 4210
box -4 -6 356 206
use OAI21X1  OAI21X1_423
timestamp 1743498307
transform -1 0 424 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_315
timestamp 1743498307
transform 1 0 424 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_99
timestamp 1743498307
transform 1 0 488 0 -1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_316
timestamp 1743498307
transform -1 0 648 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_73
timestamp 1743498307
transform 1 0 648 0 -1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_312
timestamp 1743498307
transform 1 0 840 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_311
timestamp 1743498307
transform -1 0 968 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_96
timestamp 1743498307
transform 1 0 968 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_333
timestamp 1743498307
transform 1 0 1016 0 -1 4210
box -4 -6 68 206
use BUFX4  BUFX4_84
timestamp 1743498307
transform -1 0 1144 0 -1 4210
box -4 -6 68 206
use BUFX4  BUFX4_82
timestamp 1743498307
transform -1 0 1208 0 -1 4210
box -4 -6 68 206
use BUFX4  BUFX4_81
timestamp 1743498307
transform 1 0 1208 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_94
timestamp 1743498307
transform 1 0 1272 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_334
timestamp 1743498307
transform 1 0 1304 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_103
timestamp 1743498307
transform 1 0 1368 0 -1 4210
box -4 -6 100 206
use NAND2X1  NAND2X1_105
timestamp 1743498307
transform 1 0 1464 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_0_0
timestamp 1743498307
transform 1 0 1512 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_1
timestamp 1743498307
transform 1 0 1528 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_2
timestamp 1743498307
transform 1 0 1544 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_345
timestamp 1743498307
transform 1 0 1560 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_344
timestamp 1743498307
transform 1 0 1624 0 -1 4210
box -4 -6 68 206
use BUFX4  BUFX4_47
timestamp 1743498307
transform 1 0 1688 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_346
timestamp 1743498307
transform 1 0 1752 0 -1 4210
box -4 -6 68 206
use DFFSR  DFFSR_76
timestamp 1743498307
transform 1 0 1816 0 -1 4210
box -4 -6 356 206
use INVX1  INVX1_73
timestamp 1743498307
transform 1 0 2168 0 -1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_32
timestamp 1743498307
transform 1 0 2200 0 -1 4210
box -4 -6 52 206
use AOI21X1  AOI21X1_4
timestamp 1743498307
transform -1 0 2312 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_22
timestamp 1743498307
transform -1 0 2376 0 -1 4210
box -4 -6 68 206
use OR2X2  OR2X2_7
timestamp 1743498307
transform 1 0 2376 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_31
timestamp 1743498307
transform -1 0 2488 0 -1 4210
box -4 -6 52 206
use XOR2X1  XOR2X1_8
timestamp 1743498307
transform 1 0 2488 0 -1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_287
timestamp 1743498307
transform -1 0 2664 0 -1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_7
timestamp 1743498307
transform 1 0 2664 0 -1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_327
timestamp 1743498307
transform 1 0 2776 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_347
timestamp 1743498307
transform 1 0 2840 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_108
timestamp 1743498307
transform 1 0 2904 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_1_0
timestamp 1743498307
transform 1 0 2952 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_1
timestamp 1743498307
transform 1 0 2968 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_2
timestamp 1743498307
transform 1 0 2984 0 -1 4210
box -4 -6 20 206
use DFFSR  DFFSR_69
timestamp 1743498307
transform 1 0 3000 0 -1 4210
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_72
timestamp 1743498307
transform 1 0 3352 0 -1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_196
timestamp 1743498307
transform 1 0 3544 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_197
timestamp 1743498307
transform -1 0 3672 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_71
timestamp 1743498307
transform 1 0 3672 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_204
timestamp 1743498307
transform 1 0 3704 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_205
timestamp 1743498307
transform -1 0 3832 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_63
timestamp 1743498307
transform 1 0 3832 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_243
timestamp 1743498307
transform 1 0 3864 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_17
timestamp 1743498307
transform 1 0 3928 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1743498307
transform 1 0 3992 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_259
timestamp 1743498307
transform 1 0 4056 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_64
timestamp 1743498307
transform 1 0 4120 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_244
timestamp 1743498307
transform 1 0 4152 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_245
timestamp 1743498307
transform 1 0 4216 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_261
timestamp 1743498307
transform 1 0 4280 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_62
timestamp 1743498307
transform -1 0 4424 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_69
timestamp 1743498307
transform 1 0 4344 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_241
timestamp 1743498307
transform 1 0 4424 0 -1 4210
box -4 -6 68 206
use INVX2  INVX2_3
timestamp 1743498307
transform 1 0 4536 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_67
timestamp 1743498307
transform 1 0 4488 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_262
timestamp 1743498307
transform -1 0 4680 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_2_2
timestamp 1743498307
transform -1 0 4616 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_1
timestamp 1743498307
transform -1 0 4600 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_0
timestamp 1743498307
transform -1 0 4584 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_263
timestamp 1743498307
transform -1 0 4744 0 -1 4210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_9
timestamp 1743498307
transform -1 0 4856 0 -1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_199
timestamp 1743498307
transform -1 0 4920 0 -1 4210
box -4 -6 68 206
use AND2X2  AND2X2_3
timestamp 1743498307
transform -1 0 4984 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_3
timestamp 1743498307
transform -1 0 5048 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_64
timestamp 1743498307
transform 1 0 5048 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_63
timestamp 1743498307
transform 1 0 5096 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_15
timestamp 1743498307
transform 1 0 5144 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_49
timestamp 1743498307
transform 1 0 5208 0 -1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_22
timestamp 1743498307
transform 1 0 5240 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_5
timestamp 1743498307
transform -1 0 5352 0 -1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_6
timestamp 1743498307
transform 1 0 5352 0 -1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_200
timestamp 1743498307
transform 1 0 5464 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_198
timestamp 1743498307
transform 1 0 5528 0 -1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_5
timestamp 1743498307
transform 1 0 5592 0 -1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_83
timestamp 1743498307
transform 1 0 5704 0 -1 4210
box -4 -6 52 206
use DFFSR  DFFSR_107
timestamp 1743498307
transform 1 0 5752 0 -1 4210
box -4 -6 356 206
use FILL  FILL_21_1
timestamp 1743498307
transform -1 0 6120 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_2
timestamp 1743498307
transform -1 0 6136 0 -1 4210
box -4 -6 20 206
use INVX1  INVX1_143
timestamp 1743498307
transform 1 0 8 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_424
timestamp 1743498307
transform 1 0 40 0 1 4210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_11
timestamp 1743498307
transform 1 0 104 0 1 4210
box -4 -6 148 206
use OAI21X1  OAI21X1_303
timestamp 1743498307
transform -1 0 312 0 1 4210
box -4 -6 68 206
use OR2X2  OR2X2_12
timestamp 1743498307
transform 1 0 312 0 1 4210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_8
timestamp 1743498307
transform 1 0 376 0 1 4210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_74
timestamp 1743498307
transform 1 0 520 0 1 4210
box -4 -6 196 206
use MUX2X1  MUX2X1_100
timestamp 1743498307
transform 1 0 712 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_318
timestamp 1743498307
transform 1 0 808 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_317
timestamp 1743498307
transform -1 0 936 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_99
timestamp 1743498307
transform 1 0 936 0 1 4210
box -4 -6 52 206
use MUX2X1  MUX2X1_89
timestamp 1743498307
transform 1 0 984 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_296
timestamp 1743498307
transform 1 0 1080 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_295
timestamp 1743498307
transform -1 0 1208 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_87
timestamp 1743498307
transform 1 0 1208 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_332
timestamp 1743498307
transform 1 0 1240 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_84
timestamp 1743498307
transform 1 0 1304 0 1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_87
timestamp 1743498307
transform -1 0 1528 0 1 4210
box -4 -6 196 206
use FILL  FILL_21_0_0
timestamp 1743498307
transform 1 0 1528 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_1
timestamp 1743498307
transform 1 0 1544 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_2
timestamp 1743498307
transform 1 0 1560 0 1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_282
timestamp 1743498307
transform 1 0 1576 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_283
timestamp 1743498307
transform -1 0 1704 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_321
timestamp 1743498307
transform 1 0 1704 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_322
timestamp 1743498307
transform -1 0 1832 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_95
timestamp 1743498307
transform -1 0 2024 0 1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_348
timestamp 1743498307
transform 1 0 2024 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_350
timestamp 1743498307
transform 1 0 2088 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_93
timestamp 1743498307
transform -1 0 2200 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_288
timestamp 1743498307
transform -1 0 2264 0 1 4210
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1743498307
transform -1 0 2328 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_92
timestamp 1743498307
transform 1 0 2328 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_91
timestamp 1743498307
transform 1 0 2376 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_290
timestamp 1743498307
transform -1 0 2488 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_83
timestamp 1743498307
transform -1 0 2520 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_289
timestamp 1743498307
transform -1 0 2584 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_85
timestamp 1743498307
transform 1 0 2584 0 1 4210
box -4 -6 100 206
use MUX2X1  MUX2X1_86
timestamp 1743498307
transform 1 0 2680 0 1 4210
box -4 -6 100 206
use NAND2X1  NAND2X1_98
timestamp 1743498307
transform -1 0 2824 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_57
timestamp 1743498307
transform 1 0 2824 0 1 4210
box -4 -6 36 206
use DFFSR  DFFSR_74
timestamp 1743498307
transform -1 0 3208 0 1 4210
box -4 -6 356 206
use FILL  FILL_21_1_0
timestamp 1743498307
transform 1 0 3208 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_1
timestamp 1743498307
transform 1 0 3224 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_2
timestamp 1743498307
transform 1 0 3240 0 1 4210
box -4 -6 20 206
use INVX1  INVX1_58
timestamp 1743498307
transform 1 0 3256 0 1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_66
timestamp 1743498307
transform 1 0 3288 0 1 4210
box -4 -6 196 206
use MUX2X1  MUX2X1_66
timestamp 1743498307
transform 1 0 3480 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_213
timestamp 1743498307
transform 1 0 3576 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_212
timestamp 1743498307
transform -1 0 3704 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_58
timestamp 1743498307
transform -1 0 3800 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_202
timestamp 1743498307
transform 1 0 3800 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_62
timestamp 1743498307
transform -1 0 3960 0 1 4210
box -4 -6 100 206
use INVX1  INVX1_56
timestamp 1743498307
transform 1 0 3960 0 1 4210
box -4 -6 36 206
use MUX2X1  MUX2X1_68
timestamp 1743498307
transform -1 0 4088 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_217
timestamp 1743498307
transform 1 0 4088 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_56
timestamp 1743498307
transform -1 0 4344 0 1 4210
box -4 -6 196 206
use INVX1  INVX1_60
timestamp 1743498307
transform 1 0 4344 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_239
timestamp 1743498307
transform 1 0 4376 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_69
timestamp 1743498307
transform 1 0 4440 0 1 4210
box -4 -6 196 206
use FILL  FILL_21_2_0
timestamp 1743498307
transform -1 0 4648 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_1
timestamp 1743498307
transform -1 0 4664 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_2
timestamp 1743498307
transform -1 0 4680 0 1 4210
box -4 -6 20 206
use NAND3X1  NAND3X1_18
timestamp 1743498307
transform -1 0 4744 0 1 4210
box -4 -6 68 206
use DFFSR  DFFSR_51
timestamp 1743498307
transform -1 0 5096 0 1 4210
box -4 -6 356 206
use DFFSR  DFFSR_39
timestamp 1743498307
transform -1 0 5448 0 1 4210
box -4 -6 356 206
use MUX2X1  MUX2X1_59
timestamp 1743498307
transform 1 0 5448 0 1 4210
box -4 -6 100 206
use MUX2X1  MUX2X1_60
timestamp 1743498307
transform 1 0 5544 0 1 4210
box -4 -6 100 206
use DFFSR  DFFSR_55
timestamp 1743498307
transform -1 0 5992 0 1 4210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_34
timestamp 1743498307
transform -1 0 6136 0 1 4210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_79
timestamp 1743498307
transform -1 0 200 0 -1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_304
timestamp 1743498307
transform 1 0 200 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_93
timestamp 1743498307
transform -1 0 360 0 -1 4610
box -4 -6 100 206
use INVX1  INVX1_85
timestamp 1743498307
transform 1 0 360 0 -1 4610
box -4 -6 36 206
use BUFX4  BUFX4_23
timestamp 1743498307
transform -1 0 456 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_278
timestamp 1743498307
transform -1 0 520 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_91
timestamp 1743498307
transform 1 0 520 0 -1 4610
box -4 -6 196 206
use MUX2X1  MUX2X1_79
timestamp 1743498307
transform 1 0 712 0 -1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_271
timestamp 1743498307
transform 1 0 808 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_270
timestamp 1743498307
transform -1 0 936 0 -1 4610
box -4 -6 68 206
use BUFX4  BUFX4_21
timestamp 1743498307
transform -1 0 1000 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_329
timestamp 1743498307
transform 1 0 1000 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_23
timestamp 1743498307
transform 1 0 1064 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_24
timestamp 1743498307
transform 1 0 1128 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_102
timestamp 1743498307
transform -1 0 1288 0 -1 4610
box -4 -6 100 206
use INVX1  INVX1_89
timestamp 1743498307
transform 1 0 1288 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_328
timestamp 1743498307
transform 1 0 1320 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_330
timestamp 1743498307
transform 1 0 1384 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_103
timestamp 1743498307
transform 1 0 1448 0 -1 4610
box -4 -6 52 206
use FILL  FILL_22_0_0
timestamp 1743498307
transform -1 0 1512 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_1
timestamp 1743498307
transform -1 0 1528 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_2
timestamp 1743498307
transform -1 0 1544 0 -1 4610
box -4 -6 20 206
use MUX2X1  MUX2X1_83
timestamp 1743498307
transform -1 0 1640 0 -1 4610
box -4 -6 100 206
use NAND3X1  NAND3X1_27
timestamp 1743498307
transform -1 0 1704 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_285
timestamp 1743498307
transform 1 0 1704 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_76
timestamp 1743498307
transform -1 0 1960 0 -1 4610
box -4 -6 196 206
use NAND3X1  NAND3X1_28
timestamp 1743498307
transform 1 0 1960 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_86
timestamp 1743498307
transform 1 0 2024 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_97
timestamp 1743498307
transform -1 0 2104 0 -1 4610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_39
timestamp 1743498307
transform 1 0 2104 0 -1 4610
box -4 -6 148 206
use NAND2X1  NAND2X1_109
timestamp 1743498307
transform -1 0 2296 0 -1 4610
box -4 -6 52 206
use BUFX4  BUFX4_85
timestamp 1743498307
transform 1 0 2296 0 -1 4610
box -4 -6 68 206
use DFFSR  DFFSR_75
timestamp 1743498307
transform -1 0 2712 0 -1 4610
box -4 -6 356 206
use OR2X2  OR2X2_8
timestamp 1743498307
transform -1 0 2776 0 -1 4610
box -4 -6 68 206
use BUFX4  BUFX4_89
timestamp 1743498307
transform 1 0 2776 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_335
timestamp 1743498307
transform 1 0 2840 0 -1 4610
box -4 -6 68 206
use FILL  FILL_22_1_0
timestamp 1743498307
transform -1 0 2920 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_1
timestamp 1743498307
transform -1 0 2936 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_2
timestamp 1743498307
transform -1 0 2952 0 -1 4610
box -4 -6 20 206
use DFFSR  DFFSR_66
timestamp 1743498307
transform -1 0 3304 0 -1 4610
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_55
timestamp 1743498307
transform -1 0 3496 0 -1 4610
box -4 -6 196 206
use INVX1  INVX1_69
timestamp 1743498307
transform 1 0 3496 0 -1 4610
box -4 -6 36 206
use BUFX4  BUFX4_92
timestamp 1743498307
transform 1 0 3528 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_215
timestamp 1743498307
transform 1 0 3592 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_67
timestamp 1743498307
transform 1 0 3656 0 -1 4610
box -4 -6 100 206
use MUX2X1  MUX2X1_61
timestamp 1743498307
transform 1 0 3752 0 -1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_203
timestamp 1743498307
transform 1 0 3848 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_61
timestamp 1743498307
transform 1 0 3912 0 -1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_214
timestamp 1743498307
transform -1 0 4168 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_216
timestamp 1743498307
transform -1 0 4232 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_257
timestamp 1743498307
transform -1 0 4296 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_260
timestamp 1743498307
transform 1 0 4296 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_255
timestamp 1743498307
transform 1 0 4360 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_16
timestamp 1743498307
transform 1 0 4424 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_20
timestamp 1743498307
transform 1 0 4488 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_61
timestamp 1743498307
transform 1 0 4552 0 -1 4610
box -4 -6 36 206
use FILL  FILL_22_2_0
timestamp 1743498307
transform 1 0 4584 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_1
timestamp 1743498307
transform 1 0 4600 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_2
timestamp 1743498307
transform 1 0 4616 0 -1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_240
timestamp 1743498307
transform 1 0 4632 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_187
timestamp 1743498307
transform 1 0 4696 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_188
timestamp 1743498307
transform -1 0 4824 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_55
timestamp 1743498307
transform 1 0 4824 0 -1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_247
timestamp 1743498307
transform -1 0 4984 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_249
timestamp 1743498307
transform 1 0 4984 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_29
timestamp 1743498307
transform -1 0 5096 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_19
timestamp 1743498307
transform -1 0 5160 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_251
timestamp 1743498307
transform -1 0 5224 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_67
timestamp 1743498307
transform 1 0 5224 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_253
timestamp 1743498307
transform -1 0 5320 0 -1 4610
box -4 -6 68 206
use BUFX4  BUFX4_95
timestamp 1743498307
transform 1 0 5320 0 -1 4610
box -4 -6 68 206
use DFFSR  DFFSR_54
timestamp 1743498307
transform -1 0 5736 0 -1 4610
box -4 -6 356 206
use DFFSR  DFFSR_56
timestamp 1743498307
transform -1 0 6088 0 -1 4610
box -4 -6 356 206
use FILL  FILL_23_1
timestamp 1743498307
transform -1 0 6104 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_2
timestamp 1743498307
transform -1 0 6120 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_3
timestamp 1743498307
transform -1 0 6136 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_93
timestamp 1743498307
transform 1 0 8 0 1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_277
timestamp 1743498307
transform 1 0 200 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_276
timestamp 1743498307
transform -1 0 328 0 1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_88
timestamp 1743498307
transform 1 0 328 0 1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_297
timestamp 1743498307
transform 1 0 520 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_298
timestamp 1743498307
transform -1 0 648 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_81
timestamp 1743498307
transform -1 0 744 0 1 4610
box -4 -6 100 206
use NAND2X1  NAND2X1_85
timestamp 1743498307
transform -1 0 792 0 1 4610
box -4 -6 52 206
use MUX2X1  MUX2X1_90
timestamp 1743498307
transform -1 0 888 0 1 4610
box -4 -6 100 206
use BUFX4  BUFX4_49
timestamp 1743498307
transform -1 0 952 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_80
timestamp 1743498307
transform -1 0 1048 0 1 4610
box -4 -6 100 206
use BUFX4  BUFX4_48
timestamp 1743498307
transform -1 0 1112 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_91
timestamp 1743498307
transform 1 0 1112 0 1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_25
timestamp 1743498307
transform 1 0 1144 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_340
timestamp 1743498307
transform -1 0 1272 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_336
timestamp 1743498307
transform -1 0 1336 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_338
timestamp 1743498307
transform 1 0 1336 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_39
timestamp 1743498307
transform 1 0 1400 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_341
timestamp 1743498307
transform 1 0 1448 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_0_0
timestamp 1743498307
transform 1 0 1512 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_1
timestamp 1743498307
transform 1 0 1528 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_2
timestamp 1743498307
transform 1 0 1544 0 1 4610
box -4 -6 20 206
use BUFX4  BUFX4_46
timestamp 1743498307
transform 1 0 1560 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_84
timestamp 1743498307
transform -1 0 1720 0 1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_286
timestamp 1743498307
transform 1 0 1720 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_342
timestamp 1743498307
transform 1 0 1784 0 1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_96
timestamp 1743498307
transform -1 0 2040 0 1 4610
box -4 -6 196 206
use NAND2X1  NAND2X1_95
timestamp 1743498307
transform 1 0 2040 0 1 4610
box -4 -6 52 206
use INVX2  INVX2_4
timestamp 1743498307
transform 1 0 2088 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_352
timestamp 1743498307
transform 1 0 2120 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_351
timestamp 1743498307
transform -1 0 2248 0 1 4610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_12
timestamp 1743498307
transform -1 0 2360 0 1 4610
box -4 -6 116 206
use OAI21X1  OAI21X1_353
timestamp 1743498307
transform -1 0 2424 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_36
timestamp 1743498307
transform -1 0 2472 0 1 4610
box -4 -6 52 206
use BUFX4  BUFX4_88
timestamp 1743498307
transform 1 0 2472 0 1 4610
box -4 -6 68 206
use DFFSR  DFFSR_59
timestamp 1743498307
transform 1 0 2536 0 1 4610
box -4 -6 356 206
use NAND2X1  NAND2X1_102
timestamp 1743498307
transform 1 0 2888 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_35
timestamp 1743498307
transform -1 0 2984 0 1 4610
box -4 -6 52 206
use BUFX4  BUFX4_91
timestamp 1743498307
transform -1 0 3048 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_1_0
timestamp 1743498307
transform 1 0 3048 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_1
timestamp 1743498307
transform 1 0 3064 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_2
timestamp 1743498307
transform 1 0 3080 0 1 4610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_60
timestamp 1743498307
transform 1 0 3096 0 1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_195
timestamp 1743498307
transform -1 0 3352 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_179
timestamp 1743498307
transform 1 0 3352 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_50
timestamp 1743498307
transform -1 0 3448 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_224
timestamp 1743498307
transform 1 0 3448 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_225
timestamp 1743498307
transform -1 0 3576 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_72
timestamp 1743498307
transform -1 0 3672 0 1 4610
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_68
timestamp 1743498307
transform 1 0 3672 0 1 4610
box -4 -6 196 206
use BUFX4  BUFX4_62
timestamp 1743498307
transform -1 0 3928 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_183
timestamp 1743498307
transform -1 0 3992 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_72
timestamp 1743498307
transform 1 0 3992 0 1 4610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_67
timestamp 1743498307
transform 1 0 4024 0 1 4610
box -4 -6 196 206
use NAND2X1  NAND2X1_71
timestamp 1743498307
transform 1 0 4216 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_79
timestamp 1743498307
transform 1 0 4264 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_182
timestamp 1743498307
transform 1 0 4312 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_181
timestamp 1743498307
transform -1 0 4440 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_53
timestamp 1743498307
transform 1 0 4440 0 1 4610
box -4 -6 100 206
use FILL  FILL_23_2_0
timestamp 1743498307
transform -1 0 4552 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_1
timestamp 1743498307
transform -1 0 4568 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_2
timestamp 1743498307
transform -1 0 4584 0 1 4610
box -4 -6 20 206
use MUX2X1  MUX2X1_73
timestamp 1743498307
transform -1 0 4680 0 1 4610
box -4 -6 100 206
use NAND2X1  NAND2X1_68
timestamp 1743498307
transform 1 0 4680 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_180
timestamp 1743498307
transform 1 0 4728 0 1 4610
box -4 -6 68 206
use BUFX4  BUFX4_65
timestamp 1743498307
transform -1 0 4856 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_63
timestamp 1743498307
transform 1 0 4856 0 1 4610
box -4 -6 100 206
use INVX1  INVX1_65
timestamp 1743498307
transform 1 0 4952 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_189
timestamp 1743498307
transform 1 0 4984 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_66
timestamp 1743498307
transform 1 0 5048 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_27
timestamp 1743498307
transform -1 0 5144 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_28
timestamp 1743498307
transform 1 0 5144 0 1 4610
box -4 -6 52 206
use MUX2X1  MUX2X1_56
timestamp 1743498307
transform 1 0 5192 0 1 4610
box -4 -6 100 206
use NOR2X1  NOR2X1_23
timestamp 1743498307
transform -1 0 5336 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_52
timestamp 1743498307
transform -1 0 5368 0 1 4610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_8
timestamp 1743498307
transform -1 0 5480 0 1 4610
box -4 -6 116 206
use NOR2X1  NOR2X1_30
timestamp 1743498307
transform -1 0 5528 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_53
timestamp 1743498307
transform -1 0 5560 0 1 4610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_13
timestamp 1743498307
transform 1 0 5560 0 1 4610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_7
timestamp 1743498307
transform 1 0 5672 0 1 4610
box -4 -6 116 206
use DFFSR  DFFSR_53
timestamp 1743498307
transform -1 0 6136 0 1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_326
timestamp 1743498307
transform -1 0 72 0 -1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_104
timestamp 1743498307
transform -1 0 168 0 -1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_325
timestamp 1743498307
transform -1 0 232 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_94
timestamp 1743498307
transform 1 0 232 0 -1 5010
box -4 -6 196 206
use OAI21X1  OAI21X1_280
timestamp 1743498307
transform 1 0 424 0 -1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_82
timestamp 1743498307
transform -1 0 584 0 -1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_279
timestamp 1743498307
transform -1 0 648 0 -1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_96
timestamp 1743498307
transform 1 0 648 0 -1 5010
box -4 -6 100 206
use NAND2X1  NAND2X1_107
timestamp 1743498307
transform 1 0 744 0 -1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_101
timestamp 1743498307
transform 1 0 792 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_92
timestamp 1743498307
transform 1 0 840 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_273
timestamp 1743498307
transform 1 0 872 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_274
timestamp 1743498307
transform -1 0 1000 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_349
timestamp 1743498307
transform -1 0 1064 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_26
timestamp 1743498307
transform 1 0 1064 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_337
timestamp 1743498307
transform -1 0 1192 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_94
timestamp 1743498307
transform 1 0 1192 0 -1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_37
timestamp 1743498307
transform -1 0 1288 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_73
timestamp 1743498307
transform -1 0 1640 0 -1 5010
box -4 -6 356 206
use FILL  FILL_24_0_0
timestamp 1743498307
transform -1 0 1656 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_1
timestamp 1743498307
transform -1 0 1672 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_2
timestamp 1743498307
transform -1 0 1688 0 -1 5010
box -4 -6 20 206
use NOR2X1  NOR2X1_33
timestamp 1743498307
transform -1 0 1736 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_71
timestamp 1743498307
transform -1 0 2088 0 -1 5010
box -4 -6 356 206
use DFFSR  DFFSR_70
timestamp 1743498307
transform -1 0 2440 0 -1 5010
box -4 -6 356 206
use BUFX4  BUFX4_86
timestamp 1743498307
transform 1 0 2440 0 -1 5010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_40
timestamp 1743498307
transform -1 0 2648 0 -1 5010
box -4 -6 148 206
use CLKBUF1  CLKBUF1_5
timestamp 1743498307
transform -1 0 2792 0 -1 5010
box -4 -6 148 206
use OAI21X1  OAI21X1_355
timestamp 1743498307
transform -1 0 2856 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_111
timestamp 1743498307
transform 1 0 2856 0 -1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_192
timestamp 1743498307
transform 1 0 2904 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_186
timestamp 1743498307
transform 1 0 2968 0 -1 5010
box -4 -6 68 206
use FILL  FILL_24_1_0
timestamp 1743498307
transform -1 0 3048 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_1
timestamp 1743498307
transform -1 0 3064 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_2
timestamp 1743498307
transform -1 0 3080 0 -1 5010
box -4 -6 20 206
use MUX2X1  MUX2X1_65
timestamp 1743498307
transform -1 0 3176 0 -1 5010
box -4 -6 100 206
use BUFX4  BUFX4_93
timestamp 1743498307
transform -1 0 3240 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_211
timestamp 1743498307
transform 1 0 3240 0 -1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_24
timestamp 1743498307
transform 1 0 3304 0 -1 5010
box -4 -6 52 206
use BUFX4  BUFX4_18
timestamp 1743498307
transform 1 0 3352 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_210
timestamp 1743498307
transform -1 0 3480 0 -1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_54
timestamp 1743498307
transform -1 0 3576 0 -1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_185
timestamp 1743498307
transform 1 0 3576 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_184
timestamp 1743498307
transform -1 0 3704 0 -1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_78
timestamp 1743498307
transform -1 0 3800 0 -1 5010
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_54
timestamp 1743498307
transform -1 0 3992 0 -1 5010
box -4 -6 196 206
use OAI21X1  OAI21X1_237
timestamp 1743498307
transform 1 0 3992 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_236
timestamp 1743498307
transform -1 0 4120 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_49
timestamp 1743498307
transform 1 0 4120 0 -1 5010
box -4 -6 196 206
use MUX2X1  MUX2X1_57
timestamp 1743498307
transform -1 0 4408 0 -1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_226
timestamp 1743498307
transform 1 0 4408 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_227
timestamp 1743498307
transform -1 0 4536 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_248
timestamp 1743498307
transform 1 0 4536 0 -1 5010
box -4 -6 68 206
use FILL  FILL_24_2_0
timestamp 1743498307
transform 1 0 4600 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_1
timestamp 1743498307
transform 1 0 4616 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_2
timestamp 1743498307
transform 1 0 4632 0 -1 5010
box -4 -6 20 206
use OAI21X1  OAI21X1_206
timestamp 1743498307
transform 1 0 4648 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_207
timestamp 1743498307
transform -1 0 4776 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_63
timestamp 1743498307
transform -1 0 4968 0 -1 5010
box -4 -6 196 206
use MUX2X1  MUX2X1_64
timestamp 1743498307
transform 1 0 4968 0 -1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_209
timestamp 1743498307
transform 1 0 5064 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_208
timestamp 1743498307
transform -1 0 5192 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_64
timestamp 1743498307
transform -1 0 5384 0 -1 5010
box -4 -6 196 206
use OAI21X1  OAI21X1_191
timestamp 1743498307
transform 1 0 5384 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_190
timestamp 1743498307
transform 1 0 5448 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_70
timestamp 1743498307
transform -1 0 5704 0 -1 5010
box -4 -6 196 206
use OAI21X1  OAI21X1_391
timestamp 1743498307
transform -1 0 5768 0 -1 5010
box -4 -6 68 206
use DFFSR  DFFSR_117
timestamp 1743498307
transform -1 0 6120 0 -1 5010
box -4 -6 356 206
use FILL  FILL_25_1
timestamp 1743498307
transform -1 0 6136 0 -1 5010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_78
timestamp 1743498307
transform 1 0 8 0 1 5010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_75
timestamp 1743498307
transform 1 0 200 0 1 5010
box -4 -6 196 206
use OAI21X1  OAI21X1_320
timestamp 1743498307
transform 1 0 392 0 1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_101
timestamp 1743498307
transform 1 0 456 0 1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_319
timestamp 1743498307
transform -1 0 616 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_309
timestamp 1743498307
transform 1 0 616 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_310
timestamp 1743498307
transform -1 0 744 0 1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_82
timestamp 1743498307
transform 1 0 744 0 1 5010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_92
timestamp 1743498307
transform 1 0 936 0 1 5010
box -4 -6 196 206
use INVX1  INVX1_96
timestamp 1743498307
transform -1 0 1160 0 1 5010
box -4 -6 36 206
use INVX1  INVX1_90
timestamp 1743498307
transform 1 0 1160 0 1 5010
box -4 -6 36 206
use MUX2X1  MUX2X1_95
timestamp 1743498307
transform -1 0 1288 0 1 5010
box -4 -6 100 206
use MUX2X1  MUX2X1_98
timestamp 1743498307
transform 1 0 1288 0 1 5010
box -4 -6 100 206
use NOR2X1  NOR2X1_38
timestamp 1743498307
transform 1 0 1384 0 1 5010
box -4 -6 52 206
use INVX1  INVX1_77
timestamp 1743498307
transform 1 0 1432 0 1 5010
box -4 -6 36 206
use FILL  FILL_25_0_0
timestamp 1743498307
transform -1 0 1480 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_0_1
timestamp 1743498307
transform -1 0 1496 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_0_2
timestamp 1743498307
transform -1 0 1512 0 1 5010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_30
timestamp 1743498307
transform -1 0 1656 0 1 5010
box -4 -6 148 206
use INVX1  INVX1_76
timestamp 1743498307
transform 1 0 1656 0 1 5010
box -4 -6 36 206
use NOR2X1  NOR2X1_40
timestamp 1743498307
transform 1 0 1688 0 1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_11
timestamp 1743498307
transform -1 0 1848 0 1 5010
box -4 -6 116 206
use CLKBUF1  CLKBUF1_29
timestamp 1743498307
transform 1 0 1848 0 1 5010
box -4 -6 148 206
use DFFSR  DFFSR_60
timestamp 1743498307
transform 1 0 1992 0 1 5010
box -4 -6 356 206
use OAI21X1  OAI21X1_356
timestamp 1743498307
transform -1 0 2408 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_112
timestamp 1743498307
transform 1 0 2408 0 1 5010
box -4 -6 52 206
use INVX1  INVX1_144
timestamp 1743498307
transform 1 0 2456 0 1 5010
box -4 -6 36 206
use DFFSR  DFFSR_130
timestamp 1743498307
transform 1 0 2488 0 1 5010
box -4 -6 356 206
use DFFSR  DFFSR_62
timestamp 1743498307
transform 1 0 2840 0 1 5010
box -4 -6 356 206
use FILL  FILL_25_1_0
timestamp 1743498307
transform -1 0 3208 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_1_1
timestamp 1743498307
transform -1 0 3224 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_1_2
timestamp 1743498307
transform -1 0 3240 0 1 5010
box -4 -6 20 206
use NAND2X1  NAND2X1_59
timestamp 1743498307
transform -1 0 3288 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_62
timestamp 1743498307
transform -1 0 3336 0 1 5010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_65
timestamp 1743498307
transform 1 0 3336 0 1 5010
box -4 -6 196 206
use NAND2X1  NAND2X1_61
timestamp 1743498307
transform 1 0 3528 0 1 5010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_59
timestamp 1743498307
transform 1 0 3576 0 1 5010
box -4 -6 196 206
use MUX2X1  MUX2X1_71
timestamp 1743498307
transform 1 0 3768 0 1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_223
timestamp 1743498307
transform 1 0 3864 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_58
timestamp 1743498307
transform -1 0 3976 0 1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_222
timestamp 1743498307
transform -1 0 4040 0 1 5010
box -4 -6 68 206
use BUFX4  BUFX4_64
timestamp 1743498307
transform -1 0 4104 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_70
timestamp 1743498307
transform 1 0 4104 0 1 5010
box -4 -6 36 206
use MUX2X1  MUX2X1_74
timestamp 1743498307
transform -1 0 4232 0 1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_256
timestamp 1743498307
transform 1 0 4232 0 1 5010
box -4 -6 68 206
use BUFX4  BUFX4_17
timestamp 1743498307
transform -1 0 4360 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_77
timestamp 1743498307
transform -1 0 4408 0 1 5010
box -4 -6 52 206
use BUFX4  BUFX4_16
timestamp 1743498307
transform 1 0 4408 0 1 5010
box -4 -6 68 206
use MUX2X1  MUX2X1_77
timestamp 1743498307
transform -1 0 4568 0 1 5010
box -4 -6 100 206
use FILL  FILL_25_2_0
timestamp 1743498307
transform -1 0 4584 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_2_1
timestamp 1743498307
transform -1 0 4600 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_2_2
timestamp 1743498307
transform -1 0 4616 0 1 5010
box -4 -6 20 206
use INVX1  INVX1_66
timestamp 1743498307
transform -1 0 4648 0 1 5010
box -4 -6 36 206
use NAND2X1  NAND2X1_73
timestamp 1743498307
transform -1 0 4696 0 1 5010
box -4 -6 52 206
use MUX2X1  MUX2X1_69
timestamp 1743498307
transform 1 0 4696 0 1 5010
box -4 -6 100 206
use NAND2X1  NAND2X1_57
timestamp 1743498307
transform 1 0 4792 0 1 5010
box -4 -6 52 206
use MUX2X1  MUX2X1_75
timestamp 1743498307
transform -1 0 4936 0 1 5010
box -4 -6 100 206
use BUFX4  BUFX4_96
timestamp 1743498307
transform -1 0 5000 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_60
timestamp 1743498307
transform 1 0 5000 0 1 5010
box -4 -6 52 206
use BUFX4  BUFX4_63
timestamp 1743498307
transform 1 0 5048 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_252
timestamp 1743498307
transform 1 0 5112 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_68
timestamp 1743498307
transform -1 0 5208 0 1 5010
box -4 -6 36 206
use MUX2X1  MUX2X1_70
timestamp 1743498307
transform 1 0 5208 0 1 5010
box -4 -6 100 206
use OAI21X1  OAI21X1_221
timestamp 1743498307
transform 1 0 5304 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_396
timestamp 1743498307
transform 1 0 5368 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_220
timestamp 1743498307
transform 1 0 5432 0 1 5010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_58
timestamp 1743498307
transform -1 0 5688 0 1 5010
box -4 -6 196 206
use NAND2X1  NAND2X1_123
timestamp 1743498307
transform -1 0 5736 0 1 5010
box -4 -6 52 206
use DFFSR  DFFSR_112
timestamp 1743498307
transform -1 0 6088 0 1 5010
box -4 -6 356 206
use FILL  FILL_26_1
timestamp 1743498307
transform 1 0 6088 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_2
timestamp 1743498307
transform 1 0 6104 0 1 5010
box -4 -6 20 206
use FILL  FILL_26_3
timestamp 1743498307
transform 1 0 6120 0 1 5010
box -4 -6 20 206
use DFFSR  DFFSR_131
timestamp 1743498307
transform 1 0 8 0 -1 5410
box -4 -6 356 206
use OAI21X1  OAI21X1_408
timestamp 1743498307
transform -1 0 424 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_128
timestamp 1743498307
transform -1 0 472 0 -1 5410
box -4 -6 52 206
use INVX1  INVX1_138
timestamp 1743498307
transform 1 0 472 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_414
timestamp 1743498307
transform 1 0 504 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_413
timestamp 1743498307
transform 1 0 568 0 -1 5410
box -4 -6 68 206
use DFFSR  DFFSR_123
timestamp 1743498307
transform -1 0 984 0 -1 5410
box -4 -6 356 206
use OAI21X1  OAI21X1_314
timestamp 1743498307
transform 1 0 984 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_313
timestamp 1743498307
transform 1 0 1048 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_307
timestamp 1743498307
transform 1 0 1112 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_308
timestamp 1743498307
transform -1 0 1240 0 -1 5410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_10
timestamp 1743498307
transform 1 0 1240 0 -1 5410
box -4 -6 116 206
use FILL  FILL_26_0_0
timestamp 1743498307
transform -1 0 1368 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_0_1
timestamp 1743498307
transform -1 0 1384 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_0_2
timestamp 1743498307
transform -1 0 1400 0 -1 5410
box -4 -6 20 206
use DFFSR  DFFSR_72
timestamp 1743498307
transform -1 0 1752 0 -1 5410
box -4 -6 356 206
use DFFSR  DFFSR_119
timestamp 1743498307
transform 1 0 1752 0 -1 5410
box -4 -6 356 206
use INVX1  INVX1_134
timestamp 1743498307
transform 1 0 2104 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_409
timestamp 1743498307
transform 1 0 2136 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_129
timestamp 1743498307
transform -1 0 2248 0 -1 5410
box -4 -6 52 206
use DFFSR  DFFSR_63
timestamp 1743498307
transform -1 0 2600 0 -1 5410
box -4 -6 356 206
use DFFSR  DFFSR_132
timestamp 1743498307
transform 1 0 2600 0 -1 5410
box -4 -6 356 206
use INVX1  INVX1_136
timestamp 1743498307
transform 1 0 2952 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_411
timestamp 1743498307
transform 1 0 2984 0 -1 5410
box -4 -6 68 206
use FILL  FILL_26_1_0
timestamp 1743498307
transform 1 0 3048 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_1_1
timestamp 1743498307
transform 1 0 3064 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_1_2
timestamp 1743498307
transform 1 0 3080 0 -1 5410
box -4 -6 20 206
use NAND2X1  NAND2X1_131
timestamp 1743498307
transform 1 0 3096 0 -1 5410
box -4 -6 52 206
use DFFSR  DFFSR_111
timestamp 1743498307
transform -1 0 3496 0 -1 5410
box -4 -6 356 206
use OAI21X1  OAI21X1_401
timestamp 1743498307
transform -1 0 3560 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_128
timestamp 1743498307
transform -1 0 3592 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_400
timestamp 1743498307
transform -1 0 3656 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_404
timestamp 1743498307
transform 1 0 3656 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_130
timestamp 1743498307
transform 1 0 3720 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_405
timestamp 1743498307
transform 1 0 3752 0 -1 5410
box -4 -6 68 206
use DFFSR  DFFSR_113
timestamp 1743498307
transform -1 0 4168 0 -1 5410
box -4 -6 356 206
use CLKBUF1  CLKBUF1_6
timestamp 1743498307
transform -1 0 4312 0 -1 5410
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_71
timestamp 1743498307
transform -1 0 4504 0 -1 5410
box -4 -6 196 206
use OAI21X1  OAI21X1_194
timestamp 1743498307
transform 1 0 4504 0 -1 5410
box -4 -6 68 206
use FILL  FILL_26_2_0
timestamp 1743498307
transform -1 0 4584 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_2_1
timestamp 1743498307
transform -1 0 4600 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_2_2
timestamp 1743498307
transform -1 0 4616 0 -1 5410
box -4 -6 20 206
use OAI21X1  OAI21X1_193
timestamp 1743498307
transform -1 0 4680 0 -1 5410
box -4 -6 68 206
use BUFX4  BUFX4_15
timestamp 1743498307
transform 1 0 4680 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_235
timestamp 1743498307
transform 1 0 4744 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_234
timestamp 1743498307
transform -1 0 4872 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_231
timestamp 1743498307
transform 1 0 4872 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_230
timestamp 1743498307
transform -1 0 5000 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_51
timestamp 1743498307
transform 1 0 5000 0 -1 5410
box -4 -6 196 206
use NAND2X1  NAND2X1_75
timestamp 1743498307
transform -1 0 5240 0 -1 5410
box -4 -6 52 206
use BUFX4  BUFX4_61
timestamp 1743498307
transform 1 0 5240 0 -1 5410
box -4 -6 68 206
use BUFX4  BUFX4_94
timestamp 1743498307
transform 1 0 5304 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_397
timestamp 1743498307
transform 1 0 5368 0 -1 5410
box -4 -6 68 206
use DFFSR  DFFSR_109
timestamp 1743498307
transform -1 0 5784 0 -1 5410
box -4 -6 356 206
use OAI21X1  OAI21X1_266
timestamp 1743498307
transform 1 0 5784 0 -1 5410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_23
timestamp 1743498307
transform -1 0 5992 0 -1 5410
box -4 -6 148 206
use OAI21X1  OAI21X1_403
timestamp 1743498307
transform -1 0 6056 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_129
timestamp 1743498307
transform -1 0 6088 0 -1 5410
box -4 -6 36 206
use FILL  FILL_27_1
timestamp 1743498307
transform -1 0 6104 0 -1 5410
box -4 -6 20 206
use FILL  FILL_27_2
timestamp 1743498307
transform -1 0 6120 0 -1 5410
box -4 -6 20 206
use FILL  FILL_27_3
timestamp 1743498307
transform -1 0 6136 0 -1 5410
box -4 -6 20 206
use INVX1  INVX1_133
timestamp 1743498307
transform -1 0 40 0 1 5410
box -4 -6 36 206
use DFFSR  DFFSR_129
timestamp 1743498307
transform 1 0 40 0 1 5410
box -4 -6 356 206
use BUFX2  BUFX2_25
timestamp 1743498307
transform -1 0 440 0 1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_88
timestamp 1743498307
transform 1 0 440 0 1 5410
box -4 -6 52 206
use INVX1  INVX1_141
timestamp 1743498307
transform -1 0 520 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_420
timestamp 1743498307
transform 1 0 520 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_419
timestamp 1743498307
transform 1 0 584 0 1 5410
box -4 -6 68 206
use DFFSR  DFFSR_126
timestamp 1743498307
transform -1 0 1000 0 1 5410
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_84
timestamp 1743498307
transform 1 0 1000 0 1 5410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_81
timestamp 1743498307
transform 1 0 1192 0 1 5410
box -4 -6 196 206
use FILL  FILL_27_0_0
timestamp 1743498307
transform 1 0 1384 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_0_1
timestamp 1743498307
transform 1 0 1400 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_0_2
timestamp 1743498307
transform 1 0 1416 0 1 5410
box -4 -6 20 206
use DFFSR  DFFSR_122
timestamp 1743498307
transform 1 0 1432 0 1 5410
box -4 -6 356 206
use BUFX2  BUFX2_21
timestamp 1743498307
transform -1 0 1832 0 1 5410
box -4 -6 52 206
use INVX1  INVX1_137
timestamp 1743498307
transform 1 0 1832 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_412
timestamp 1743498307
transform -1 0 1928 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_132
timestamp 1743498307
transform 1 0 1928 0 1 5410
box -4 -6 52 206
use BUFX2  BUFX2_18
timestamp 1743498307
transform -1 0 2024 0 1 5410
box -4 -6 52 206
use DFFSR  DFFSR_120
timestamp 1743498307
transform 1 0 2024 0 1 5410
box -4 -6 356 206
use INVX1  INVX1_135
timestamp 1743498307
transform 1 0 2376 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_410
timestamp 1743498307
transform 1 0 2408 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_130
timestamp 1743498307
transform 1 0 2472 0 1 5410
box -4 -6 52 206
use BUFX2  BUFX2_19
timestamp 1743498307
transform -1 0 2568 0 1 5410
box -4 -6 52 206
use DFFSR  DFFSR_121
timestamp 1743498307
transform 1 0 2568 0 1 5410
box -4 -6 356 206
use BUFX2  BUFX2_20
timestamp 1743498307
transform 1 0 2920 0 1 5410
box -4 -6 52 206
use FILL  FILL_27_1_0
timestamp 1743498307
transform -1 0 2984 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_1_1
timestamp 1743498307
transform -1 0 3000 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_1_2
timestamp 1743498307
transform -1 0 3016 0 1 5410
box -4 -6 20 206
use DFFSR  DFFSR_114
timestamp 1743498307
transform -1 0 3368 0 1 5410
box -4 -6 356 206
use INVX1  INVX1_131
timestamp 1743498307
transform 1 0 3368 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_407
timestamp 1743498307
transform 1 0 3400 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_406
timestamp 1743498307
transform -1 0 3528 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_127
timestamp 1743498307
transform 1 0 3528 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_399
timestamp 1743498307
transform 1 0 3560 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_398
timestamp 1743498307
transform 1 0 3624 0 1 5410
box -4 -6 68 206
use DFFSR  DFFSR_110
timestamp 1743498307
transform -1 0 4040 0 1 5410
box -4 -6 356 206
use CLKBUF1  CLKBUF1_27
timestamp 1743498307
transform -1 0 4184 0 1 5410
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_50
timestamp 1743498307
transform -1 0 4376 0 1 5410
box -4 -6 196 206
use OAI21X1  OAI21X1_229
timestamp 1743498307
transform 1 0 4376 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_228
timestamp 1743498307
transform -1 0 4504 0 1 5410
box -4 -6 68 206
use OR2X2  OR2X2_11
timestamp 1743498307
transform -1 0 4568 0 1 5410
box -4 -6 68 206
use FILL  FILL_27_2_0
timestamp 1743498307
transform -1 0 4584 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_2_1
timestamp 1743498307
transform -1 0 4600 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_2_2
timestamp 1743498307
transform -1 0 4616 0 1 5410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_53
timestamp 1743498307
transform -1 0 4808 0 1 5410
box -4 -6 196 206
use OAI21X1  OAI21X1_219
timestamp 1743498307
transform 1 0 4808 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_218
timestamp 1743498307
transform -1 0 4936 0 1 5410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_57
timestamp 1743498307
transform -1 0 5128 0 1 5410
box -4 -6 196 206
use OAI21X1  OAI21X1_232
timestamp 1743498307
transform 1 0 5128 0 1 5410
box -4 -6 68 206
use MUX2X1  MUX2X1_76
timestamp 1743498307
transform 1 0 5192 0 1 5410
box -4 -6 100 206
use OAI21X1  OAI21X1_233
timestamp 1743498307
transform -1 0 5352 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_126
timestamp 1743498307
transform 1 0 5352 0 1 5410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_52
timestamp 1743498307
transform -1 0 5576 0 1 5410
box -4 -6 196 206
use DFFSR  DFFSR_115
timestamp 1743498307
transform -1 0 5928 0 1 5410
box -4 -6 356 206
use INVX1  INVX1_121
timestamp 1743498307
transform -1 0 5960 0 1 5410
box -4 -6 36 206
use CLKBUF1  CLKBUF1_10
timestamp 1743498307
transform 1 0 5960 0 1 5410
box -4 -6 148 206
use FILL  FILL_28_1
timestamp 1743498307
transform 1 0 6104 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_2
timestamp 1743498307
transform 1 0 6120 0 1 5410
box -4 -6 20 206
<< labels >>
flabel metal4 s 1496 -40 1544 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 3032 -40 3080 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -19 3317 -13 3323 7 FreeSans 24 0 0 0 clk
port 2 nsew
flabel metal3 s 6157 3337 6163 3343 3 FreeSans 24 0 0 0 rst
port 3 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 dest[0]
port 4 nsew
flabel metal3 s -19 2337 -13 2343 7 FreeSans 24 0 0 0 dest[1]
port 5 nsew
flabel metal3 s 6157 1477 6163 1483 3 FreeSans 24 0 0 0 dest[2]
port 6 nsew
flabel metal3 s 6157 97 6163 103 3 FreeSans 24 0 0 0 dest[3]
port 7 nsew
flabel metal2 s 3725 5637 3731 5643 3 FreeSans 24 90 0 0 dest[4]
port 8 nsew
flabel metal2 s 3373 5637 3379 5643 3 FreeSans 24 90 0 0 dest[5]
port 9 nsew
flabel metal3 s -19 3497 -13 3503 7 FreeSans 24 0 0 0 dest[6]
port 10 nsew
flabel metal3 s -19 4297 -13 4303 7 FreeSans 24 0 0 0 dest[7]
port 11 nsew
flabel metal2 s 509 -23 515 -17 7 FreeSans 24 270 0 0 ext_data_in[0]
port 12 nsew
flabel metal3 s -19 2297 -13 2303 7 FreeSans 24 0 0 0 ext_data_in[1]
port 13 nsew
flabel metal2 s 477 -23 483 -17 7 FreeSans 24 270 0 0 ext_data_in[2]
port 14 nsew
flabel metal3 s -19 2097 -13 2103 7 FreeSans 24 0 0 0 ext_data_in[3]
port 15 nsew
flabel metal3 s 6157 1697 6163 1703 3 FreeSans 24 0 0 0 ext_data_in[4]
port 16 nsew
flabel metal2 s 5661 -23 5667 -17 7 FreeSans 24 270 0 0 ext_data_in[5]
port 17 nsew
flabel metal2 s 5629 -23 5635 -17 7 FreeSans 24 270 0 0 ext_data_in[6]
port 18 nsew
flabel metal3 s 6157 277 6163 283 3 FreeSans 24 0 0 0 ext_data_in[7]
port 19 nsew
flabel metal2 s 5357 5637 5363 5643 3 FreeSans 24 90 0 0 ext_data_in[8]
port 20 nsew
flabel metal2 s 3533 5637 3539 5643 3 FreeSans 24 90 0 0 ext_data_in[9]
port 21 nsew
flabel metal2 s 3565 5637 3571 5643 3 FreeSans 24 90 0 0 ext_data_in[10]
port 22 nsew
flabel metal2 s 6061 5637 6067 5643 3 FreeSans 24 90 0 0 ext_data_in[11]
port 23 nsew
flabel metal2 s 477 5637 483 5643 3 FreeSans 24 90 0 0 ext_data_in[12]
port 24 nsew
flabel metal3 s -19 3697 -13 3703 7 FreeSans 24 0 0 0 ext_data_in[13]
port 25 nsew
flabel metal3 s -19 3737 -13 3743 7 FreeSans 24 0 0 0 ext_data_in[14]
port 26 nsew
flabel metal2 s 509 5637 515 5643 3 FreeSans 24 90 0 0 ext_data_in[15]
port 27 nsew
flabel metal2 s 2173 -23 2179 -17 7 FreeSans 24 270 0 0 ext_data_out[0]
port 28 nsew
flabel metal2 s 1373 -23 1379 -17 7 FreeSans 24 270 0 0 ext_data_out[1]
port 29 nsew
flabel metal2 s 2621 -23 2627 -17 7 FreeSans 24 270 0 0 ext_data_out[2]
port 30 nsew
flabel metal2 s 2573 -23 2579 -17 7 FreeSans 24 270 0 0 ext_data_out[3]
port 31 nsew
flabel metal2 s 4013 -23 4019 -17 7 FreeSans 24 270 0 0 ext_data_out[4]
port 32 nsew
flabel metal2 s 2669 -23 2675 -17 7 FreeSans 24 270 0 0 ext_data_out[5]
port 33 nsew
flabel metal3 s 6157 1897 6163 1903 3 FreeSans 24 0 0 0 ext_data_out[6]
port 34 nsew
flabel metal2 s 3117 -23 3123 -17 7 FreeSans 24 270 0 0 ext_data_out[7]
port 35 nsew
flabel metal3 s 6157 1517 6163 1523 3 FreeSans 24 0 0 0 ext_data_out[8]
port 36 nsew
flabel metal3 s 6157 3497 6163 3503 3 FreeSans 24 0 0 0 ext_data_out[9]
port 37 nsew
flabel metal3 s 6157 3697 6163 3703 3 FreeSans 24 0 0 0 ext_data_out[10]
port 38 nsew
flabel metal3 s 6157 3097 6163 3103 3 FreeSans 24 0 0 0 ext_data_out[11]
port 39 nsew
flabel metal2 s 1997 5637 2003 5643 3 FreeSans 24 90 0 0 ext_data_out[12]
port 40 nsew
flabel metal2 s 2541 5637 2547 5643 3 FreeSans 24 90 0 0 ext_data_out[13]
port 41 nsew
flabel metal2 s 2941 5637 2947 5643 3 FreeSans 24 90 0 0 ext_data_out[14]
port 42 nsew
flabel metal2 s 1805 5637 1811 5643 3 FreeSans 24 90 0 0 ext_data_out[15]
port 43 nsew
flabel metal3 s -19 297 -13 303 7 FreeSans 24 0 0 0 pe_busy[0]
port 44 nsew
flabel metal3 s 6157 317 6163 323 3 FreeSans 24 0 0 0 pe_busy[1]
port 45 nsew
flabel metal2 s 6093 5637 6099 5643 3 FreeSans 24 90 0 0 pe_busy[2]
port 46 nsew
flabel metal2 s 413 5637 419 5643 3 FreeSans 24 90 0 0 pe_busy[3]
port 47 nsew
<< end >>

magic
tech scmos
magscale 1 2
timestamp 1743127117
<< metal1 >>
rect 2632 5006 2638 5014
rect 2646 5006 2652 5014
rect 2660 5006 2666 5014
rect 2674 5006 2680 5014
rect 5720 5006 5726 5014
rect 5734 5006 5740 5014
rect 5748 5006 5754 5014
rect 5762 5006 5768 5014
rect 6312 4976 6316 4984
rect 4893 4957 4908 4963
rect 5485 4957 5523 4963
rect 356 4937 371 4943
rect 413 4937 435 4943
rect 829 4937 851 4943
rect 1581 4937 1603 4943
rect 2029 4937 2044 4943
rect 3437 4937 3474 4943
rect 397 4917 412 4923
rect 893 4917 931 4923
rect 893 4897 899 4917
rect 1229 4917 1244 4923
rect 1533 4917 1564 4923
rect 1629 4917 1660 4923
rect 2910 4917 2940 4923
rect 3405 4917 3452 4923
rect 3837 4917 3874 4923
rect 4228 4917 4259 4923
rect 4317 4917 4355 4923
rect 5277 4917 5315 4923
rect 5341 4917 5379 4923
rect 4381 4897 4419 4903
rect 4436 4897 4467 4903
rect 5341 4897 5347 4917
rect 5437 4917 5475 4923
rect 5396 4897 5411 4903
rect 1112 4806 1118 4814
rect 1126 4806 1132 4814
rect 1140 4806 1146 4814
rect 1154 4806 1160 4814
rect 4152 4806 4158 4814
rect 4166 4806 4172 4814
rect 4180 4806 4186 4814
rect 4194 4806 4200 4814
rect 394 4776 396 4784
rect 2740 4776 2742 4784
rect 3034 4776 3036 4784
rect 614 4736 620 4744
rect 714 4736 716 4744
rect 892 4732 900 4736
rect 1628 4737 1644 4743
rect 1628 4732 1636 4737
rect 2989 4737 3012 4743
rect 5117 4737 5156 4743
rect 5308 4737 5347 4743
rect 5308 4732 5316 4737
rect 813 4703 819 4723
rect 813 4697 851 4703
rect 1245 4703 1251 4723
rect 1677 4704 1683 4723
rect 1812 4717 1827 4723
rect 3204 4717 3219 4723
rect 3421 4717 3459 4723
rect 1213 4697 1251 4703
rect 1636 4697 1667 4703
rect 1684 4697 1692 4703
rect 2269 4697 2316 4703
rect 2772 4697 2787 4703
rect 3037 4697 3091 4703
rect 3124 4697 3139 4703
rect 3149 4697 3164 4703
rect 3405 4697 3436 4703
rect 3645 4703 3651 4723
rect 3732 4717 3747 4723
rect 4308 4717 4323 4723
rect 3645 4697 3683 4703
rect 4141 4697 4204 4703
rect 4356 4697 4403 4703
rect 5188 4697 5235 4703
rect 5764 4697 5811 4703
rect 5821 4697 5852 4703
rect 5885 4703 5891 4723
rect 5885 4697 5923 4703
rect 5949 4697 5971 4703
rect 1821 4677 1852 4683
rect 2308 4677 2338 4683
rect 3364 4677 3379 4683
rect 3476 4677 3491 4683
rect 3565 4677 3587 4683
rect 3604 4677 3619 4683
rect 3716 4677 3731 4683
rect 4164 4677 4211 4683
rect 4253 4677 4268 4683
rect 4365 4677 4380 4683
rect 5197 4677 5212 4683
rect 5780 4677 5795 4683
rect 5949 4677 5955 4697
rect 6157 4703 6163 4723
rect 6157 4697 6195 4703
rect 6397 4677 6412 4683
rect 6813 4677 6876 4683
rect 1844 4657 1875 4663
rect 3108 4657 3123 4663
rect 3156 4657 3180 4663
rect 4093 4657 4131 4663
rect 5725 4657 5772 4663
rect 6045 4657 6067 4663
rect 906 4636 908 4644
rect 1348 4636 1350 4644
rect 3546 4636 3548 4644
rect 6148 4636 6150 4644
rect 2632 4606 2638 4614
rect 2646 4606 2652 4614
rect 2660 4606 2666 4614
rect 2674 4606 2680 4614
rect 5720 4606 5726 4614
rect 5734 4606 5740 4614
rect 5748 4606 5754 4614
rect 5762 4606 5768 4614
rect 2056 4576 2060 4584
rect 5444 4576 5446 4584
rect 2221 4557 2243 4563
rect 2989 4557 3004 4563
rect 5316 4557 5331 4563
rect 324 4537 339 4543
rect 436 4537 451 4543
rect 573 4537 595 4543
rect 253 4517 291 4523
rect 228 4496 236 4504
rect 253 4497 259 4517
rect 381 4517 419 4523
rect 381 4497 387 4517
rect 573 4523 579 4537
rect 1613 4537 1644 4543
rect 452 4517 467 4523
rect 477 4517 515 4523
rect 541 4517 579 4523
rect 509 4497 515 4517
rect 740 4517 755 4523
rect 1021 4517 1059 4523
rect 692 4496 700 4504
rect 1053 4497 1059 4517
rect 1453 4517 1468 4523
rect 1636 4517 1667 4523
rect 1725 4517 1740 4523
rect 2173 4523 2179 4543
rect 3012 4537 3027 4543
rect 3069 4537 3084 4543
rect 3133 4537 3148 4543
rect 2156 4517 2179 4523
rect 2156 4512 2164 4517
rect 3053 4517 3091 4523
rect 3133 4517 3139 4537
rect 3204 4536 3208 4544
rect 3373 4537 3388 4543
rect 3508 4537 3523 4543
rect 3581 4537 3603 4543
rect 3836 4543 3844 4544
rect 3828 4537 3844 4543
rect 4324 4537 4339 4543
rect 5373 4537 5395 4543
rect 6237 4543 6243 4563
rect 6237 4537 6275 4543
rect 3524 4517 3539 4523
rect 4804 4517 4828 4523
rect 5357 4517 5372 4523
rect 5549 4517 5596 4523
rect 6189 4517 6204 4523
rect 3012 4497 3027 4503
rect 3236 4497 3251 4503
rect 5316 4497 5331 4503
rect 5453 4497 5468 4503
rect 6340 4497 6371 4503
rect 1894 4476 1900 4484
rect 2125 4477 2140 4483
rect 2276 4477 2291 4483
rect 4877 4477 4892 4483
rect 5293 4477 5308 4483
rect 5620 4477 5635 4483
rect 1112 4406 1118 4414
rect 1126 4406 1132 4414
rect 1140 4406 1146 4414
rect 1154 4406 1160 4414
rect 4152 4406 4158 4414
rect 4166 4406 4172 4414
rect 4180 4406 4186 4414
rect 4194 4406 4200 4414
rect 1850 4376 1852 4384
rect 3012 4376 3014 4384
rect 3082 4376 3084 4384
rect 5300 4376 5302 4384
rect 5498 4376 5500 4384
rect 1690 4336 1692 4344
rect 2796 4332 2804 4336
rect 253 4303 259 4323
rect 253 4297 291 4303
rect 436 4297 451 4303
rect 621 4297 636 4303
rect 813 4303 819 4323
rect 836 4316 844 4324
rect 4973 4317 5011 4323
rect 781 4297 819 4303
rect 941 4297 956 4303
rect 1076 4297 1139 4303
rect 1604 4297 1619 4303
rect 3140 4297 3171 4303
rect 3380 4297 3395 4303
rect 4996 4297 5027 4303
rect 621 4277 652 4283
rect 1092 4277 1139 4283
rect 1245 4277 1260 4283
rect 2212 4277 2227 4283
rect 2180 4257 2195 4263
rect 2221 4257 2227 4277
rect 3101 4277 3123 4283
rect 3229 4277 3244 4283
rect 2333 4257 2348 4263
rect 3229 4257 3235 4277
rect 3261 4277 3292 4283
rect 3332 4277 3347 4283
rect 3357 4277 3372 4283
rect 4429 4277 4467 4283
rect 4429 4264 4435 4277
rect 4973 4257 4988 4263
rect 2632 4206 2638 4214
rect 2646 4206 2652 4214
rect 2660 4206 2666 4214
rect 2674 4206 2680 4214
rect 5720 4206 5726 4214
rect 5734 4206 5740 4214
rect 5748 4206 5754 4214
rect 5762 4206 5768 4214
rect 2292 4176 2294 4184
rect 3108 4176 3110 4184
rect 6184 4176 6188 4184
rect 6440 4176 6444 4184
rect 1380 4156 1382 4164
rect 276 4137 291 4143
rect 397 4137 419 4143
rect 276 4117 291 4123
rect 413 4123 419 4137
rect 541 4137 556 4143
rect 1172 4137 1219 4143
rect 1597 4137 1619 4143
rect 413 4117 444 4123
rect 461 4117 499 4123
rect 493 4097 499 4117
rect 1613 4123 1619 4137
rect 1556 4117 1571 4123
rect 1613 4117 1644 4123
rect 1757 4117 1788 4123
rect 1821 4117 1859 4123
rect 1853 4097 1859 4117
rect 2301 4117 2339 4123
rect 2301 4097 2307 4117
rect 2429 4123 2435 4143
rect 2525 4137 2547 4143
rect 3037 4137 3059 4143
rect 2413 4117 2435 4123
rect 2461 4117 2499 4123
rect 2493 4097 2499 4117
rect 3117 4117 3139 4123
rect 3149 4117 3187 4123
rect 3117 4104 3123 4117
rect 3389 4123 3395 4143
rect 3453 4137 3468 4143
rect 4045 4137 4083 4143
rect 3389 4117 3404 4123
rect 3540 4117 3555 4123
rect 4045 4117 4051 4137
rect 4973 4137 4995 4143
rect 6301 4137 6316 4143
rect 6228 4117 6259 4123
rect 2532 4097 2547 4103
rect 3021 4097 3036 4103
rect 3396 4097 3411 4103
rect 1284 4077 1315 4083
rect 1533 4077 1548 4083
rect 3677 4083 3683 4103
rect 3677 4077 3708 4083
rect 4132 4077 4179 4083
rect 5764 4077 5795 4083
rect 1149 4037 1196 4043
rect 6340 4036 6342 4044
rect 1112 4006 1118 4014
rect 1126 4006 1132 4014
rect 1140 4006 1146 4014
rect 1154 4006 1160 4014
rect 4152 4006 4158 4014
rect 4166 4006 4172 4014
rect 4180 4006 4186 4014
rect 4194 4006 4200 4014
rect 282 3976 284 3984
rect 1220 3976 1222 3984
rect 2746 3976 2748 3984
rect 3338 3976 3340 3984
rect 5210 3976 5212 3984
rect 5834 3976 5836 3984
rect 474 3936 476 3944
rect 2260 3936 2268 3944
rect 4460 3937 4499 3943
rect 4876 3932 4884 3936
rect 5004 3932 5012 3936
rect 5308 3932 5316 3936
rect 5756 3932 5764 3936
rect 125 3897 140 3903
rect 285 3897 323 3903
rect 317 3883 323 3897
rect 445 3903 451 3923
rect 1364 3917 1379 3923
rect 1412 3916 1420 3924
rect 1469 3917 1507 3923
rect 413 3897 451 3903
rect 500 3897 531 3903
rect 612 3897 627 3903
rect 941 3897 972 3903
rect 1021 3897 1036 3903
rect 1092 3897 1171 3903
rect 1421 3897 1436 3903
rect 1492 3897 1523 3903
rect 1709 3903 1715 3923
rect 3140 3917 3155 3923
rect 3277 3917 3315 3923
rect 5044 3917 5059 3923
rect 1645 3897 1683 3903
rect 1709 3897 1747 3903
rect 317 3877 332 3883
rect 493 3877 508 3883
rect 1645 3883 1651 3897
rect 1892 3897 1907 3903
rect 1917 3897 1948 3903
rect 2077 3897 2092 3903
rect 2116 3897 2131 3903
rect 3118 3897 3148 3903
rect 3549 3897 3580 3903
rect 3677 3897 3692 3903
rect 4174 3897 4259 3903
rect 5108 3897 5139 3903
rect 5421 3903 5427 3923
rect 5444 3916 5452 3924
rect 5389 3897 5427 3903
rect 5453 3897 5468 3903
rect 6173 3903 6179 3923
rect 6173 3897 6211 3903
rect 1629 3877 1651 3883
rect 1853 3877 1868 3883
rect 2381 3877 2396 3883
rect 3421 3877 3436 3883
rect 3572 3877 3587 3883
rect 3661 3877 3715 3883
rect 3581 3857 3587 3877
rect 4461 3877 4476 3883
rect 5972 3876 5974 3884
rect 6173 3877 6188 3883
rect 5644 3872 5652 3876
rect 4292 3856 4294 3864
rect 1085 3837 1116 3843
rect 4852 3836 4854 3844
rect 5716 3837 5763 3843
rect 2632 3806 2638 3814
rect 2646 3806 2652 3814
rect 2660 3806 2666 3814
rect 2674 3806 2680 3814
rect 5720 3806 5726 3814
rect 5734 3806 5740 3814
rect 5748 3806 5754 3814
rect 5762 3806 5768 3814
rect 5162 3776 5164 3784
rect 5725 3777 5772 3783
rect 3172 3756 3180 3764
rect 3416 3756 3420 3764
rect 6116 3757 6124 3763
rect 349 3737 364 3743
rect 468 3737 483 3743
rect 1005 3737 1027 3743
rect 1725 3737 1756 3743
rect 2148 3737 2163 3743
rect 2724 3737 2787 3743
rect 3252 3737 3315 3743
rect 3645 3737 3731 3743
rect 5101 3737 5116 3743
rect 5924 3737 5939 3743
rect 6333 3737 6348 3743
rect 269 3717 307 3723
rect 301 3697 307 3717
rect 356 3717 380 3723
rect 740 3717 755 3723
rect 765 3717 796 3723
rect 1748 3717 1763 3723
rect 685 3697 700 3703
rect 1069 3697 1084 3703
rect 1757 3697 1763 3717
rect 2189 3717 2204 3723
rect 3069 3717 3084 3723
rect 3213 3717 3260 3723
rect 4013 3717 4028 3723
rect 5021 3717 5059 3723
rect 2125 3697 2163 3703
rect 2701 3697 2787 3703
rect 618 3676 620 3684
rect 804 3677 819 3683
rect 1460 3677 1475 3683
rect 3460 3677 3475 3683
rect 3517 3677 3564 3683
rect 3837 3683 3843 3703
rect 5053 3697 5059 3717
rect 5108 3717 5139 3723
rect 5245 3717 5283 3723
rect 5076 3696 5084 3704
rect 5277 3697 5283 3717
rect 5412 3717 5427 3723
rect 5780 3717 5811 3723
rect 5837 3717 5875 3723
rect 5837 3697 5843 3717
rect 5965 3717 5980 3723
rect 6212 3717 6227 3723
rect 6141 3697 6163 3703
rect 3837 3677 3875 3683
rect 1226 3656 1228 3664
rect 3869 3657 3875 3677
rect 6228 3676 6230 3684
rect 916 3636 918 3644
rect 1044 3636 1046 3644
rect 1112 3606 1118 3614
rect 1126 3606 1132 3614
rect 1140 3606 1146 3614
rect 1154 3606 1160 3614
rect 4152 3606 4158 3614
rect 4166 3606 4172 3614
rect 4180 3606 4186 3614
rect 4194 3606 4200 3614
rect 922 3576 924 3584
rect 3066 3576 3068 3584
rect 5770 3576 5772 3584
rect 1156 3536 1158 3544
rect 2348 3537 2364 3543
rect 4228 3537 4260 3543
rect 5158 3536 5164 3544
rect 4748 3532 4756 3536
rect 188 3517 211 3523
rect 188 3512 196 3517
rect 228 3516 236 3524
rect 397 3503 403 3523
rect 365 3497 403 3503
rect 468 3497 483 3503
rect 813 3503 819 3523
rect 1309 3517 1331 3523
rect 1540 3516 1548 3524
rect 2957 3517 2972 3523
rect 5492 3516 5500 3524
rect 6060 3506 6068 3516
rect 813 3497 851 3503
rect 1261 3497 1276 3503
rect 1332 3497 1347 3503
rect 1549 3497 1564 3503
rect 3620 3497 3635 3503
rect 5085 3497 5100 3503
rect 5373 3497 5388 3503
rect 5524 3497 5555 3503
rect 5981 3497 5996 3503
rect 6157 3503 6163 3523
rect 6157 3497 6195 3503
rect 6301 3497 6332 3503
rect 6397 3503 6403 3523
rect 6365 3497 6403 3503
rect 6740 3497 6755 3503
rect 941 3477 956 3483
rect 2030 3477 2060 3483
rect 2157 3477 2179 3483
rect 2221 3477 2252 3483
rect 2349 3477 2371 3483
rect 3476 3477 3491 3483
rect 5453 3477 5475 3483
rect 5581 3477 5603 3483
rect 5636 3477 5651 3483
rect 6445 3477 6460 3483
rect 6781 3477 6819 3483
rect 6781 3464 6787 3477
rect 3860 3457 3875 3463
rect 5348 3456 5350 3464
rect 1069 3437 1116 3443
rect 1236 3436 1238 3444
rect 2100 3436 2104 3444
rect 4740 3436 4742 3444
rect 6276 3436 6278 3444
rect 2632 3406 2638 3414
rect 2646 3406 2652 3414
rect 2660 3406 2666 3414
rect 2674 3406 2680 3414
rect 5720 3406 5726 3414
rect 5734 3406 5740 3414
rect 5748 3406 5754 3414
rect 5762 3406 5768 3414
rect 1316 3376 1318 3384
rect 1364 3376 1366 3384
rect 1578 3376 1580 3384
rect 3194 3376 3196 3384
rect 3332 3376 3334 3384
rect 3492 3376 3494 3384
rect 3652 3376 3654 3384
rect 4148 3376 4150 3384
rect 4724 3376 4726 3384
rect 4772 3376 4774 3384
rect 2285 3357 2300 3363
rect 3588 3356 3596 3364
rect 340 3337 355 3343
rect 724 3337 740 3343
rect 973 3337 995 3343
rect 1276 3343 1284 3348
rect 1276 3337 1299 3343
rect 260 3317 291 3323
rect 324 3317 348 3323
rect 797 3317 812 3323
rect 996 3317 1011 3323
rect 1021 3317 1084 3323
rect 1517 3323 1523 3343
rect 1549 3337 1564 3343
rect 2292 3337 2322 3343
rect 3044 3337 3059 3343
rect 3101 3337 3123 3343
rect 3357 3337 3404 3343
rect 3620 3337 3635 3343
rect 3684 3337 3699 3343
rect 3924 3337 3955 3343
rect 4333 3337 4348 3343
rect 4900 3337 4915 3343
rect 5828 3337 5843 3343
rect 6061 3337 6076 3343
rect 6189 3337 6204 3343
rect 1517 3317 1555 3323
rect 1668 3317 1698 3323
rect 2189 3317 2227 3323
rect 3837 3323 3843 3336
rect 3837 3317 3859 3323
rect 4813 3317 4851 3323
rect 5021 3317 5036 3323
rect 5101 3317 5139 3323
rect 1373 3297 1395 3303
rect 1549 3297 1571 3303
rect 1661 3297 1676 3303
rect 3044 3297 3059 3303
rect 4733 3297 4748 3303
rect 5101 3297 5107 3317
rect 5892 3317 5907 3323
rect 5469 3297 5484 3303
rect 5901 3297 5907 3317
rect 6125 3317 6140 3323
rect 6605 3317 6620 3323
rect 5965 3297 5980 3303
rect 6269 3297 6291 3303
rect 189 3277 212 3283
rect 234 3276 236 3284
rect 5972 3277 5987 3283
rect 5981 3257 5987 3277
rect 6500 3276 6502 3284
rect 6580 3276 6582 3284
rect 6666 3276 6668 3284
rect 1460 3236 1464 3244
rect 1636 3236 1638 3244
rect 4852 3236 4854 3244
rect 1112 3206 1118 3214
rect 1126 3206 1132 3214
rect 1140 3206 1146 3214
rect 1154 3206 1160 3214
rect 4152 3206 4158 3214
rect 4166 3206 4172 3214
rect 4180 3206 4186 3214
rect 4194 3206 4200 3214
rect 4868 3176 4870 3184
rect 5396 3176 5398 3184
rect 5530 3176 5532 3184
rect 6330 3176 6332 3184
rect 1437 3137 1476 3143
rect 2116 3137 2132 3143
rect 2476 3137 2524 3143
rect 4637 3137 4652 3143
rect 429 3103 435 3123
rect 516 3117 531 3123
rect 2068 3117 2083 3123
rect 3012 3116 3020 3124
rect 3636 3116 3644 3124
rect 3661 3117 3699 3123
rect 356 3097 387 3103
rect 397 3097 435 3103
rect 2228 3097 2243 3103
rect 2397 3097 2428 3103
rect 3044 3097 3059 3103
rect 3101 3097 3116 3103
rect 477 3077 499 3083
rect 2068 3077 2099 3083
rect 2109 3077 2131 3083
rect 3325 3083 3331 3103
rect 3453 3097 3484 3103
rect 3501 3097 3555 3103
rect 4756 3097 4771 3103
rect 4893 3103 4899 3123
rect 4893 3097 4931 3103
rect 5101 3097 5132 3103
rect 5661 3097 5676 3103
rect 6029 3103 6035 3123
rect 5997 3097 6035 3103
rect 6301 3103 6307 3123
rect 6269 3097 6307 3103
rect 6468 3097 6483 3103
rect 6621 3103 6627 3123
rect 6589 3097 6627 3103
rect 3309 3077 3331 3083
rect 3380 3077 3395 3083
rect 3476 3077 3491 3083
rect 4733 3077 4748 3083
rect 5124 3077 5139 3083
rect 5213 3077 5228 3083
rect 4420 3057 4435 3063
rect 4794 3056 4796 3064
rect 5133 3057 5139 3077
rect 5357 3077 5379 3083
rect 5677 3077 5699 3083
rect 6132 3056 6134 3064
rect 6506 3056 6508 3064
rect 538 3036 540 3044
rect 596 3036 598 3044
rect 2052 3036 2054 3044
rect 3332 3037 3347 3043
rect 2632 3006 2638 3014
rect 2646 3006 2652 3014
rect 2660 3006 2666 3014
rect 2674 3006 2680 3014
rect 5720 3006 5726 3014
rect 5734 3006 5740 3014
rect 5748 3006 5754 3014
rect 5762 3006 5768 3014
rect 1098 2976 1100 2984
rect 5757 2977 5804 2983
rect 3594 2956 3596 2964
rect 3661 2957 3699 2963
rect 4762 2956 4764 2964
rect 29 2937 51 2943
rect 397 2937 419 2943
rect 964 2937 995 2943
rect 1005 2937 1027 2943
rect 1540 2937 1555 2943
rect 1565 2937 1587 2943
rect 2382 2937 2412 2943
rect 2461 2937 2499 2943
rect 93 2917 131 2923
rect 93 2897 99 2917
rect 253 2917 268 2923
rect 317 2917 355 2923
rect 189 2897 227 2903
rect 349 2897 355 2917
rect 461 2917 499 2923
rect 493 2897 499 2917
rect 589 2917 604 2923
rect 2941 2912 2947 2943
rect 3101 2912 3107 2943
rect 3165 2912 3171 2943
rect 3325 2937 3347 2943
rect 3357 2937 3379 2943
rect 3485 2937 3507 2943
rect 3325 2917 3331 2937
rect 3373 2917 3379 2937
rect 3501 2917 3507 2937
rect 4548 2937 4563 2943
rect 4605 2937 4627 2943
rect 4701 2937 4716 2943
rect 5245 2937 5260 2943
rect 5469 2937 5491 2943
rect 5981 2937 6003 2943
rect 4093 2917 4131 2923
rect 4644 2917 4675 2923
rect 4980 2917 4995 2923
rect 5236 2917 5283 2923
rect 5997 2923 6003 2937
rect 5997 2917 6035 2923
rect 6061 2917 6099 2923
rect 1012 2897 1027 2903
rect 3341 2897 3372 2903
rect 3476 2897 3491 2903
rect 6061 2897 6067 2917
rect 6260 2917 6291 2923
rect 6508 2903 6516 2908
rect 6493 2897 6516 2903
rect 172 2884 180 2888
rect 1572 2877 1588 2883
rect 3197 2877 3228 2883
rect 3309 2877 3324 2883
rect 3453 2877 3484 2883
rect 3453 2857 3459 2877
rect 6036 2856 6038 2864
rect 68 2836 70 2844
rect 378 2836 380 2844
rect 5146 2836 5148 2844
rect 5284 2836 5286 2844
rect 5364 2836 5366 2844
rect 1112 2806 1118 2814
rect 1126 2806 1132 2814
rect 1140 2806 1146 2814
rect 1154 2806 1160 2814
rect 4152 2806 4158 2814
rect 4166 2806 4172 2814
rect 4180 2806 4186 2814
rect 4194 2806 4200 2814
rect 2900 2776 2902 2784
rect 3588 2776 3590 2784
rect 5834 2756 5836 2764
rect 4013 2737 4035 2743
rect 3804 2724 3812 2728
rect 1748 2717 1763 2723
rect 2836 2716 2844 2724
rect 4029 2717 4035 2737
rect 6468 2736 6470 2744
rect 6634 2736 6636 2744
rect 5908 2716 5916 2724
rect 589 2697 627 2703
rect 1869 2697 1884 2703
rect 1716 2677 1731 2683
rect 1741 2677 1763 2683
rect 2797 2677 2803 2708
rect 2868 2697 2899 2703
rect 3620 2697 3651 2703
rect 3661 2697 3676 2703
rect 3908 2697 3923 2703
rect 3364 2677 3379 2683
rect 3389 2677 3427 2683
rect 3517 2677 3539 2683
rect 3556 2677 3571 2683
rect 3677 2677 3699 2683
rect 3716 2677 3731 2683
rect 4045 2683 4051 2703
rect 4157 2697 4243 2703
rect 5373 2697 5388 2703
rect 5636 2697 5667 2703
rect 5917 2697 5948 2703
rect 6004 2697 6019 2703
rect 6141 2703 6147 2723
rect 6109 2697 6147 2703
rect 6772 2697 6787 2703
rect 4029 2677 4051 2683
rect 5261 2677 5292 2683
rect 6372 2677 6387 2683
rect 1092 2656 1100 2664
rect 2269 2657 2284 2663
rect 4589 2657 4620 2663
rect 4973 2657 5011 2663
rect 3748 2636 3750 2644
rect 4052 2637 4067 2643
rect 6324 2636 6326 2644
rect 2632 2606 2638 2614
rect 2646 2606 2652 2614
rect 2660 2606 2666 2614
rect 2674 2606 2680 2614
rect 5720 2606 5726 2614
rect 5734 2606 5740 2614
rect 5748 2606 5754 2614
rect 5762 2606 5768 2614
rect 4900 2576 4902 2584
rect 148 2557 163 2563
rect 861 2557 899 2563
rect 1405 2537 1420 2543
rect 1604 2537 1619 2543
rect 2605 2537 2675 2543
rect 93 2517 108 2523
rect 1581 2517 1619 2523
rect 1709 2517 1747 2523
rect 3085 2512 3091 2543
rect 3149 2512 3155 2543
rect 3812 2537 3827 2543
rect 4093 2537 4147 2543
rect 3604 2517 3635 2523
rect 3732 2517 3763 2523
rect 4141 2517 4147 2537
rect 5053 2537 5068 2543
rect 5709 2537 5756 2543
rect 4580 2517 4595 2523
rect 4653 2517 4691 2523
rect 4925 2517 4963 2523
rect 5053 2517 5091 2523
rect 5709 2517 5795 2523
rect 3236 2496 3244 2504
rect 3572 2496 3580 2504
rect 3940 2497 3955 2503
rect 5709 2497 5715 2517
rect 6132 2517 6147 2523
rect 6468 2517 6499 2523
rect 6509 2517 6524 2523
rect 6669 2517 6684 2523
rect 6442 2476 6444 2484
rect 3636 2436 3638 2444
rect 3764 2436 3766 2444
rect 1112 2406 1118 2414
rect 1126 2406 1132 2414
rect 1140 2406 1146 2414
rect 1154 2406 1160 2414
rect 4152 2406 4158 2414
rect 4166 2406 4172 2414
rect 4180 2406 4186 2414
rect 4194 2406 4200 2414
rect 2266 2376 2268 2384
rect 2893 2337 2908 2343
rect 157 2297 188 2303
rect 1757 2297 1795 2303
rect 2228 2297 2243 2303
rect 2989 2297 3004 2303
rect 3149 2297 3164 2303
rect 3597 2303 3603 2323
rect 3597 2297 3635 2303
rect 4244 2297 4275 2303
rect 4333 2297 4387 2303
rect 4957 2297 4995 2303
rect 5645 2303 5651 2323
rect 5645 2297 5683 2303
rect 5732 2297 5778 2303
rect 6173 2297 6188 2303
rect 580 2277 595 2283
rect 1293 2277 1331 2283
rect 173 2257 188 2263
rect 685 2257 723 2263
rect 1325 2257 1331 2277
rect 3037 2277 3059 2283
rect 3709 2277 3724 2283
rect 3501 2257 3516 2263
rect 4189 2257 4252 2263
rect 4932 2256 4934 2264
rect 6644 2257 6659 2263
rect 2740 2237 2787 2243
rect 3444 2237 3459 2243
rect 5636 2236 5638 2244
rect 2632 2206 2638 2214
rect 2646 2206 2652 2214
rect 2660 2206 2666 2214
rect 2674 2206 2680 2214
rect 5720 2206 5726 2214
rect 5734 2206 5740 2214
rect 5748 2206 5754 2214
rect 5762 2206 5768 2214
rect 2372 2176 2374 2184
rect 3028 2176 3030 2184
rect 5864 2176 5868 2184
rect 6500 2176 6504 2184
rect 1165 2157 1203 2163
rect 2205 2157 2243 2163
rect 2253 2157 2291 2163
rect 3348 2156 3356 2164
rect 29 2137 51 2143
rect 2276 2137 2307 2143
rect 2388 2137 2419 2143
rect 2452 2137 2467 2143
rect 2996 2137 3011 2143
rect 2974 2117 2988 2123
rect 3044 2117 3075 2123
rect 3117 2123 3123 2143
rect 3540 2137 3570 2143
rect 5325 2137 5347 2143
rect 5444 2137 5475 2143
rect 5492 2137 5507 2143
rect 5597 2137 5640 2143
rect 5981 2137 5996 2143
rect 6077 2137 6108 2143
rect 3108 2117 3123 2123
rect 3380 2117 3411 2123
rect 3949 2117 3964 2123
rect 3997 2117 4060 2123
rect 5380 2117 5427 2123
rect 5437 2117 5452 2123
rect 5556 2117 5571 2123
rect 5700 2117 5747 2123
rect 5908 2117 5923 2123
rect 6573 2123 6579 2143
rect 6564 2117 6579 2123
rect 3076 2096 3084 2104
rect 3101 2097 3107 2116
rect 1149 2077 1180 2083
rect 5524 2076 5526 2084
rect 3306 2036 3308 2044
rect 3460 2036 3462 2044
rect 1112 2006 1118 2014
rect 1126 2006 1132 2014
rect 1140 2006 1146 2014
rect 1154 2006 1160 2014
rect 4152 2006 4158 2014
rect 4166 2006 4172 2014
rect 4180 2006 4186 2014
rect 4194 2006 4200 2014
rect 138 1976 140 1984
rect 684 1932 692 1936
rect 5796 1936 5798 1944
rect 1052 1932 1060 1936
rect 493 1917 531 1923
rect 1069 1917 1155 1923
rect 3412 1917 3427 1923
rect 3940 1917 3955 1923
rect 516 1897 547 1903
rect 669 1897 700 1903
rect 1277 1897 1308 1903
rect 1501 1897 1532 1903
rect 3412 1897 3443 1903
rect 3869 1897 3923 1903
rect 4893 1897 4931 1903
rect 5629 1903 5635 1923
rect 5629 1897 5667 1903
rect 5901 1903 5907 1923
rect 5901 1897 5939 1903
rect 6269 1897 6300 1903
rect 6685 1897 6716 1903
rect 6749 1897 6764 1903
rect 29 1877 51 1883
rect 573 1877 595 1883
rect 589 1864 595 1877
rect 2189 1877 2227 1883
rect 2221 1857 2227 1877
rect 3453 1877 3491 1883
rect 3508 1877 3523 1883
rect 3741 1877 3779 1883
rect 5245 1877 5283 1883
rect 6308 1877 6323 1883
rect 3564 1864 3572 1868
rect 4700 1864 4708 1868
rect 6628 1857 6643 1863
rect 6653 1857 6668 1863
rect 5316 1836 5320 1844
rect 6820 1836 6824 1844
rect 2632 1806 2638 1814
rect 2646 1806 2652 1814
rect 2660 1806 2666 1814
rect 2674 1806 2680 1814
rect 5720 1806 5726 1814
rect 5734 1806 5740 1814
rect 5748 1806 5754 1814
rect 5762 1806 5768 1814
rect 570 1776 572 1784
rect 4532 1776 4534 1784
rect 5770 1776 5772 1784
rect 1412 1756 1414 1764
rect 2077 1757 2115 1763
rect 717 1737 739 1743
rect 1565 1724 1571 1743
rect 1741 1737 1763 1743
rect 637 1717 675 1723
rect 669 1697 675 1717
rect 1572 1717 1603 1723
rect 1757 1723 1763 1737
rect 2605 1743 2611 1763
rect 5901 1757 5924 1763
rect 5916 1754 5924 1757
rect 6308 1756 6310 1764
rect 6493 1757 6515 1763
rect 6525 1757 6563 1763
rect 2573 1737 2611 1743
rect 3101 1737 3132 1743
rect 4909 1737 4931 1743
rect 5556 1737 5571 1743
rect 5869 1737 5891 1743
rect 6413 1743 6419 1756
rect 6397 1737 6419 1743
rect 1757 1717 1795 1723
rect 1885 1717 1923 1723
rect 1933 1717 1948 1723
rect 1188 1697 1203 1703
rect 1629 1697 1651 1703
rect 1796 1696 1804 1704
rect 1885 1697 1891 1717
rect 2029 1717 2060 1723
rect 3060 1717 3075 1723
rect 4701 1717 4716 1723
rect 4797 1717 4835 1723
rect 5668 1717 5708 1723
rect 5828 1717 5843 1723
rect 6173 1717 6211 1723
rect 1988 1697 2003 1703
rect 4852 1697 4867 1703
rect 6205 1697 6211 1717
rect 6404 1717 6435 1723
rect 6445 1717 6460 1723
rect 556 1684 564 1688
rect 1546 1676 1548 1684
rect 2026 1676 2028 1684
rect 2212 1677 2227 1683
rect 6234 1676 6236 1684
rect 6381 1677 6396 1683
rect 1124 1657 1171 1663
rect 3988 1636 3990 1644
rect 4676 1636 4678 1644
rect 4772 1636 4774 1644
rect 4890 1636 4892 1644
rect 1112 1606 1118 1614
rect 1126 1606 1132 1614
rect 1140 1606 1146 1614
rect 1154 1606 1160 1614
rect 4152 1606 4158 1614
rect 4166 1606 4172 1614
rect 4180 1606 4186 1614
rect 4194 1606 4200 1614
rect 68 1576 70 1584
rect 394 1576 396 1584
rect 906 1576 908 1584
rect 1892 1576 1894 1584
rect 4228 1577 4243 1583
rect 5178 1576 5180 1584
rect 1805 1537 1820 1543
rect 3037 1537 3052 1543
rect 3492 1537 3507 1543
rect 93 1503 99 1523
rect 93 1497 131 1503
rect 365 1503 371 1523
rect 333 1497 371 1503
rect 420 1497 451 1503
rect 532 1497 547 1503
rect 669 1503 675 1523
rect 669 1497 707 1503
rect 877 1503 883 1523
rect 845 1497 883 1503
rect 1284 1497 1299 1503
rect 1469 1497 1484 1503
rect 1549 1503 1555 1523
rect 1549 1497 1587 1503
rect 2109 1503 2115 1523
rect 2077 1497 2115 1503
rect 2532 1497 2563 1503
rect 13 1477 51 1483
rect 157 1477 188 1483
rect 436 1477 451 1483
rect 756 1477 771 1483
rect 1373 1477 1388 1483
rect 2013 1477 2028 1483
rect 2557 1477 2563 1497
rect 3076 1497 3091 1503
rect 5133 1497 5148 1503
rect 5261 1503 5267 1523
rect 5261 1497 5299 1503
rect 5373 1497 5388 1503
rect 5517 1503 5523 1523
rect 5428 1497 5443 1503
rect 5485 1497 5523 1503
rect 5636 1497 5651 1503
rect 5661 1497 5763 1503
rect 5869 1503 5875 1523
rect 5837 1497 5875 1503
rect 6020 1497 6035 1503
rect 6621 1497 6659 1503
rect 6669 1497 6684 1503
rect 3060 1477 3075 1483
rect 4317 1477 4339 1483
rect 5549 1477 5564 1483
rect 6509 1477 6524 1483
rect 6621 1483 6627 1497
rect 6765 1497 6780 1503
rect 6804 1497 6819 1503
rect 6605 1477 6627 1483
rect 972 1463 980 1472
rect 972 1457 1004 1463
rect 1220 1456 1222 1464
rect 2500 1456 2502 1464
rect 3476 1457 3507 1463
rect 5108 1457 5123 1463
rect 4356 1436 4358 1444
rect 5972 1436 5974 1444
rect 2632 1406 2638 1414
rect 2646 1406 2652 1414
rect 2660 1406 2666 1414
rect 2674 1406 2680 1414
rect 5720 1406 5726 1414
rect 5734 1406 5740 1414
rect 5748 1406 5754 1414
rect 5762 1406 5768 1414
rect 3034 1376 3036 1384
rect 5789 1377 5836 1383
rect 2477 1357 2492 1363
rect 653 1337 675 1343
rect 237 1317 268 1323
rect 653 1323 659 1337
rect 893 1337 908 1343
rect 1277 1337 1299 1343
rect 1405 1337 1427 1343
rect 1720 1336 1724 1344
rect 1821 1337 1836 1343
rect 2605 1337 2652 1343
rect 2829 1337 2851 1343
rect 6093 1337 6115 1343
rect 557 1317 595 1323
rect 621 1317 659 1323
rect 188 1303 196 1308
rect 188 1297 211 1303
rect 228 1296 236 1304
rect 589 1297 595 1317
rect 756 1317 771 1323
rect 797 1317 835 1323
rect 797 1297 803 1317
rect 1197 1317 1235 1323
rect 1053 1297 1075 1303
rect 1229 1297 1235 1317
rect 1453 1317 1484 1323
rect 1636 1317 1651 1323
rect 1940 1317 1971 1323
rect 2781 1317 2796 1323
rect 2964 1317 2979 1323
rect 5485 1317 5523 1323
rect 1853 1297 1891 1303
rect 1908 1296 1916 1304
rect 2980 1296 2988 1304
rect 5108 1297 5123 1303
rect 5485 1297 5491 1317
rect 6020 1317 6035 1323
rect 6109 1323 6115 1337
rect 6605 1337 6636 1343
rect 6109 1317 6147 1323
rect 6340 1317 6371 1323
rect 6669 1317 6684 1323
rect 6804 1317 6819 1323
rect 6212 1296 6220 1304
rect 6252 1303 6260 1308
rect 6237 1297 6260 1303
rect 470 1276 476 1284
rect 2925 1277 2940 1283
rect 5917 1277 5948 1283
rect 1972 1256 1974 1264
rect 772 1236 774 1244
rect 954 1236 956 1244
rect 1258 1236 1260 1244
rect 2506 1236 2508 1244
rect 4308 1237 4339 1243
rect 5588 1236 5590 1244
rect 1112 1206 1118 1214
rect 1126 1206 1132 1214
rect 1140 1206 1146 1214
rect 1154 1206 1160 1214
rect 4152 1206 4158 1214
rect 4166 1206 4172 1214
rect 4180 1206 4186 1214
rect 4194 1206 4200 1214
rect 308 1176 310 1184
rect 1994 1176 1996 1184
rect 2234 1176 2236 1184
rect 5866 1176 5868 1184
rect 6404 1176 6406 1184
rect 1828 1156 1830 1164
rect 1252 1137 1267 1143
rect 2556 1137 2572 1143
rect 3212 1137 3228 1143
rect 4700 1137 4716 1143
rect 5258 1136 5260 1144
rect 6084 1136 6090 1144
rect 6260 1136 6262 1144
rect 1028 1116 1036 1124
rect 333 1097 348 1103
rect 749 1097 780 1103
rect 1053 1103 1059 1123
rect 1924 1116 1932 1124
rect 2157 1117 2172 1123
rect 5789 1117 5811 1123
rect 5924 1116 5932 1124
rect 1053 1097 1091 1103
rect 1101 1097 1148 1103
rect 1485 1097 1500 1103
rect 1773 1097 1827 1103
rect 2061 1097 2083 1103
rect 2180 1097 2195 1103
rect 2317 1097 2355 1103
rect 2365 1097 2396 1103
rect 5428 1097 5459 1103
rect 5949 1103 5955 1123
rect 5908 1097 5923 1103
rect 5949 1097 5987 1103
rect 6285 1103 6291 1123
rect 6285 1097 6323 1103
rect 6333 1097 6348 1103
rect 6509 1097 6524 1103
rect 397 1077 412 1083
rect 1213 1077 1228 1083
rect 1284 1077 1299 1083
rect 1725 1077 1747 1083
rect 2445 1077 2467 1083
rect 2557 1077 2579 1083
rect 2589 1077 2668 1083
rect 3053 1077 3068 1083
rect 3213 1077 3235 1083
rect 3245 1077 3276 1083
rect 4596 1077 4611 1083
rect 4781 1077 4812 1083
rect 5172 1077 5187 1083
rect 5540 1077 5571 1083
rect 5748 1077 5763 1083
rect 1692 1063 1700 1066
rect 1692 1057 1715 1063
rect 6044 1063 6052 1066
rect 6029 1057 6052 1063
rect 5780 1036 5782 1044
rect 6836 1036 6838 1044
rect 2632 1006 2638 1014
rect 2646 1006 2652 1014
rect 2660 1006 2666 1014
rect 2674 1006 2680 1014
rect 5720 1006 5726 1014
rect 5734 1006 5740 1014
rect 5748 1006 5754 1014
rect 5762 1006 5768 1014
rect 596 976 598 984
rect 4452 976 4454 984
rect 5108 976 5110 984
rect 2205 957 2227 963
rect 3892 956 3900 964
rect 5764 957 5811 963
rect 5821 957 5844 963
rect 5836 954 5844 957
rect 77 937 99 943
rect 77 923 83 937
rect 285 937 300 943
rect 644 937 675 943
rect 1692 943 1700 948
rect 1692 937 1715 943
rect 2148 937 2163 943
rect 2413 937 2435 943
rect 2484 937 2508 943
rect 3005 937 3027 943
rect 3037 937 3052 943
rect 3853 937 3875 943
rect 3965 937 3987 943
rect 5165 937 5180 943
rect 5325 937 5347 943
rect 5485 937 5507 943
rect 6093 937 6108 943
rect 6372 937 6387 943
rect 6684 937 6708 943
rect 45 917 83 923
rect 180 917 195 923
rect 420 917 451 923
rect 461 917 499 923
rect 493 897 499 917
rect 548 917 563 923
rect 621 917 652 923
rect 1348 917 1363 923
rect 1373 917 1411 923
rect 1053 897 1075 903
rect 1405 897 1411 917
rect 1453 917 1468 923
rect 2141 917 2172 923
rect 1428 896 1436 904
rect 2141 897 2147 917
rect 2461 917 2524 923
rect 4612 917 4627 923
rect 5197 917 5235 923
rect 5364 917 5395 923
rect 5405 917 5459 923
rect 5565 917 5619 923
rect 6237 917 6275 923
rect 6285 917 6300 923
rect 3005 897 3020 903
rect 3853 897 3868 903
rect 4653 897 4691 903
rect 6212 896 6220 904
rect 6237 897 6243 917
rect 6372 917 6403 923
rect 6765 917 6796 923
rect 6508 903 6516 908
rect 6493 897 6516 903
rect 5116 884 5124 888
rect 522 876 524 884
rect 1482 876 1484 884
rect 3964 877 3980 883
rect 5132 884 5140 888
rect 266 856 268 864
rect 5236 856 5238 864
rect 388 836 390 844
rect 1098 836 1100 844
rect 1290 836 1292 844
rect 2376 836 2380 844
rect 4570 836 4572 844
rect 5562 836 5564 844
rect 5706 836 5708 844
rect 6468 836 6470 844
rect 1112 806 1118 814
rect 1126 806 1132 814
rect 1140 806 1146 814
rect 1154 806 1160 814
rect 4152 806 4158 814
rect 4166 806 4172 814
rect 4180 806 4186 814
rect 4194 806 4200 814
rect 1636 776 1638 784
rect 6180 776 6182 784
rect 6666 776 6668 784
rect 5802 756 5804 764
rect 1700 736 1702 744
rect 4044 737 4131 743
rect 4044 732 4052 737
rect 77 697 92 703
rect 269 703 275 723
rect 452 716 460 724
rect 1885 717 1907 723
rect 212 697 227 703
rect 237 697 275 703
rect 397 697 428 703
rect 461 697 499 703
rect 493 683 499 697
rect 573 697 588 703
rect 1156 697 1219 703
rect 1389 697 1404 703
rect 1684 697 1699 703
rect 1796 697 1827 703
rect 3949 703 3955 723
rect 5092 716 5100 724
rect 3885 697 3923 703
rect 3949 697 3987 703
rect 5117 703 5123 723
rect 5117 697 5155 703
rect 5661 703 5667 723
rect 5684 716 5692 724
rect 6205 717 6227 723
rect 5629 697 5667 703
rect 5693 697 5708 703
rect 6164 697 6179 703
rect 6349 697 6364 703
rect 6413 697 6428 703
rect 6532 697 6563 703
rect 493 677 515 683
rect 1309 677 1324 683
rect 1341 677 1363 683
rect 3997 677 4012 683
rect 4557 677 4572 683
rect 5053 677 5075 683
rect 4996 657 5011 663
rect 1828 636 1830 644
rect 1972 636 1976 644
rect 4045 637 4076 643
rect 2632 606 2638 614
rect 2646 606 2652 614
rect 2660 606 2666 614
rect 2674 606 2680 614
rect 5720 606 5726 614
rect 5734 606 5740 614
rect 5748 606 5754 614
rect 5762 606 5768 614
rect 346 576 348 584
rect 404 576 406 584
rect 868 576 870 584
rect 4564 576 4566 584
rect 5268 576 5270 584
rect 5800 576 5804 584
rect 1412 556 1414 564
rect 1764 557 1779 563
rect 372 537 380 543
rect 420 537 451 543
rect 1613 537 1635 543
rect 2980 537 3011 543
rect 3021 537 3043 543
rect 4932 537 4947 543
rect 5165 537 5203 543
rect 5700 537 5747 543
rect 6253 537 6268 543
rect 6756 537 6771 543
rect 77 517 92 523
rect 237 517 275 523
rect 269 497 275 517
rect 557 517 595 523
rect 589 497 595 517
rect 1124 517 1180 523
rect 3548 517 3580 523
rect 3548 516 3556 517
rect 4356 517 4403 523
rect 4973 517 4988 523
rect 5325 517 5363 523
rect 2493 497 2531 503
rect 3028 497 3043 503
rect 3133 497 3171 503
rect 3965 497 4003 503
rect 5357 497 5363 517
rect 5412 517 5420 523
rect 5428 517 5443 523
rect 6484 517 6508 523
rect 6733 517 6764 523
rect 6797 517 6835 523
rect 6829 497 6835 517
rect 332 484 340 488
rect 412 484 420 488
rect 3132 484 3140 488
rect 1332 476 1334 484
rect 4380 483 4388 488
rect 4340 477 4388 483
rect 4524 483 4532 488
rect 4572 484 4580 488
rect 4524 477 4540 483
rect 5068 484 5076 488
rect 5276 484 5284 488
rect 6474 476 6476 484
rect 5146 436 5148 444
rect 5658 436 5660 444
rect 6618 436 6620 444
rect 1112 406 1118 414
rect 1126 406 1132 414
rect 1140 406 1146 414
rect 1154 406 1160 414
rect 4152 406 4158 414
rect 4166 406 4172 414
rect 4180 406 4186 414
rect 4194 406 4200 414
rect 1764 376 1766 384
rect 1844 376 1846 384
rect 6714 376 6716 384
rect 6808 376 6812 384
rect 1034 356 1036 364
rect 4138 336 4140 344
rect 5732 337 5763 343
rect 6266 336 6268 344
rect 445 303 451 323
rect 1092 316 1100 324
rect 445 297 483 303
rect 493 297 508 303
rect 516 297 547 303
rect 557 297 588 303
rect 1380 297 1395 303
rect 1405 297 1436 303
rect 1517 297 1532 303
rect 1773 297 1795 303
rect 1928 297 1980 303
rect 2724 297 2755 303
rect 2781 303 2787 323
rect 2781 297 2819 303
rect 3092 297 3107 303
rect 3645 297 3683 303
rect 4093 297 4108 303
rect 4253 297 4291 303
rect 4717 303 4723 323
rect 4820 316 4828 324
rect 4676 297 4691 303
rect 4717 297 4755 303
rect 5316 297 5331 303
rect 5421 303 5427 323
rect 5348 297 5395 303
rect 5421 297 5459 303
rect 5549 303 5555 323
rect 5549 297 5587 303
rect 5604 297 5635 303
rect 5844 297 5875 303
rect 6237 303 6243 323
rect 6205 297 6243 303
rect 6269 297 6307 303
rect 381 277 403 283
rect 509 277 524 283
rect 781 277 796 283
rect 1972 277 2002 283
rect 2829 277 2844 283
rect 4660 277 4675 283
rect 4909 277 4931 283
rect 5485 277 5500 283
rect 6301 283 6307 297
rect 6388 297 6403 303
rect 6461 297 6476 303
rect 6557 303 6563 323
rect 6525 297 6563 303
rect 6685 303 6691 323
rect 6612 297 6643 303
rect 6653 297 6691 303
rect 6301 277 6323 283
rect 6461 277 6476 283
rect 3117 257 3155 263
rect 4045 257 4083 263
rect 5980 263 5988 266
rect 5965 257 5988 263
rect 2868 236 2870 244
rect 4180 237 4227 243
rect 2632 206 2638 214
rect 2646 206 2652 214
rect 2660 206 2666 214
rect 2674 206 2680 214
rect 5720 206 5726 214
rect 5734 206 5740 214
rect 5748 206 5754 214
rect 5762 206 5768 214
rect 2621 177 2668 183
rect 365 157 380 163
rect 1613 143 1619 163
rect 2333 157 2364 163
rect 2813 157 2828 163
rect 4573 157 4588 163
rect 5373 157 5388 163
rect 1437 137 1475 143
rect 1565 137 1619 143
rect 2493 137 2508 143
rect 2836 137 2850 143
rect 4596 137 4611 143
rect 6196 137 6211 143
rect 6861 137 6876 143
rect 429 117 444 123
rect 1528 117 1564 123
rect 2589 117 2604 123
rect 2717 117 2732 123
rect 2749 117 2787 123
rect 3341 117 3378 123
rect 5758 117 5843 123
rect 6125 117 6163 123
rect 6173 117 6204 123
rect 2516 97 2531 103
rect 6100 96 6108 104
rect 6125 97 6131 117
rect 6212 117 6227 123
rect 6237 117 6275 123
rect 6269 97 6275 117
rect 6685 117 6700 123
rect 6292 96 6300 104
rect 1112 6 1118 14
rect 1126 6 1132 14
rect 1140 6 1146 14
rect 1154 6 1160 14
rect 4152 6 4158 14
rect 4166 6 4172 14
rect 4180 6 4186 14
rect 4194 6 4200 14
<< m2contact >>
rect 2638 5006 2646 5014
rect 2652 5006 2660 5014
rect 2666 5006 2674 5014
rect 5726 5006 5734 5014
rect 5740 5006 5748 5014
rect 5754 5006 5762 5014
rect 2972 4976 2980 4984
rect 3804 4976 3812 4984
rect 4284 4976 4292 4984
rect 6316 4976 6324 4984
rect 172 4956 180 4964
rect 444 4956 452 4964
rect 620 4956 628 4964
rect 812 4956 820 4964
rect 1564 4956 1572 4964
rect 1836 4956 1844 4964
rect 2012 4956 2020 4964
rect 2220 4956 2228 4964
rect 2748 4956 2756 4964
rect 3148 4956 3156 4964
rect 3628 4956 3636 4964
rect 3868 4956 3876 4964
rect 4028 4956 4036 4964
rect 4300 4956 4308 4964
rect 4620 4956 4628 4964
rect 4796 4956 4804 4964
rect 4844 4956 4852 4964
rect 4908 4956 4916 4964
rect 5084 4956 5092 4964
rect 5260 4956 5268 4964
rect 5676 4956 5684 4964
rect 6060 4956 6068 4964
rect 6684 4956 6692 4964
rect 140 4936 148 4944
rect 348 4936 356 4944
rect 588 4936 596 4944
rect 876 4936 884 4944
rect 956 4936 964 4944
rect 1100 4936 1108 4944
rect 1484 4936 1492 4944
rect 1500 4936 1508 4944
rect 1868 4936 1876 4944
rect 2044 4936 2052 4944
rect 2252 4936 2260 4944
rect 2396 4936 2404 4944
rect 2524 4936 2532 4944
rect 2716 4936 2724 4944
rect 3116 4936 3124 4944
rect 3340 4936 3348 4944
rect 3660 4936 3668 4944
rect 4060 4936 4068 4944
rect 4332 4936 4340 4944
rect 4396 4936 4404 4944
rect 4652 4936 4660 4944
rect 5116 4936 5124 4944
rect 5292 4936 5300 4944
rect 5324 4936 5332 4944
rect 5388 4936 5396 4944
rect 5452 4936 5460 4944
rect 5708 4936 5716 4944
rect 6028 4936 6036 4944
rect 6252 4936 6260 4944
rect 6348 4936 6356 4944
rect 6364 4936 6372 4944
rect 6716 4936 6724 4944
rect 140 4916 148 4924
rect 252 4916 260 4924
rect 412 4916 420 4924
rect 492 4916 500 4924
rect 700 4916 708 4924
rect 860 4916 868 4924
rect 44 4896 52 4904
rect 364 4896 372 4904
rect 524 4900 532 4908
rect 940 4916 948 4924
rect 1244 4916 1252 4924
rect 1276 4916 1284 4924
rect 1356 4916 1364 4924
rect 1516 4916 1524 4924
rect 1564 4916 1572 4924
rect 1612 4916 1620 4924
rect 1660 4916 1668 4924
rect 1756 4916 1764 4924
rect 1980 4916 1988 4924
rect 2140 4916 2148 4924
rect 2364 4916 2372 4924
rect 2620 4916 2628 4924
rect 2940 4916 2948 4924
rect 3020 4916 3028 4924
rect 3228 4916 3236 4924
rect 3452 4916 3460 4924
rect 3548 4916 3556 4924
rect 4060 4916 4068 4924
rect 4220 4916 4228 4924
rect 4364 4916 4372 4924
rect 4716 4916 4724 4924
rect 4860 4916 4868 4924
rect 4922 4916 4930 4924
rect 5004 4916 5012 4924
rect 5228 4916 5236 4924
rect 908 4896 916 4904
rect 1548 4896 1556 4904
rect 1644 4896 1652 4904
rect 1964 4896 1972 4904
rect 2348 4896 2356 4904
rect 2620 4896 2628 4904
rect 3020 4896 3028 4904
rect 3724 4900 3732 4908
rect 4124 4900 4132 4908
rect 4428 4896 4436 4904
rect 4748 4896 4756 4904
rect 5180 4900 5188 4908
rect 5420 4916 5428 4924
rect 5596 4916 5604 4924
rect 5948 4916 5956 4924
rect 6604 4916 6612 4924
rect 5356 4896 5364 4904
rect 5388 4896 5396 4904
rect 5772 4900 5780 4908
rect 5932 4896 5940 4904
rect 6812 4896 6820 4904
rect 3724 4854 3732 4862
rect 4124 4854 4132 4862
rect 5180 4854 5188 4862
rect 5772 4854 5780 4862
rect 44 4836 52 4844
rect 332 4836 340 4844
rect 524 4836 532 4844
rect 780 4836 788 4844
rect 988 4836 996 4844
rect 1340 4836 1348 4844
rect 1676 4836 1684 4844
rect 1964 4836 1972 4844
rect 2060 4836 2068 4844
rect 2348 4836 2356 4844
rect 2620 4836 2628 4844
rect 3020 4836 3028 4844
rect 3308 4836 3316 4844
rect 3468 4836 3476 4844
rect 4748 4836 4756 4844
rect 4812 4836 4820 4844
rect 4828 4836 4836 4844
rect 5516 4836 5524 4844
rect 5932 4836 5940 4844
rect 6220 4836 6228 4844
rect 6476 4836 6484 4844
rect 6524 4836 6532 4844
rect 6812 4836 6820 4844
rect 1118 4806 1126 4814
rect 1132 4806 1140 4814
rect 1146 4806 1154 4814
rect 4158 4806 4166 4814
rect 4172 4806 4180 4814
rect 4186 4806 4194 4814
rect 316 4776 324 4784
rect 396 4776 404 4784
rect 2156 4776 2164 4784
rect 2732 4776 2740 4784
rect 2924 4776 2932 4784
rect 3036 4776 3044 4784
rect 3804 4776 3812 4784
rect 4092 4776 4100 4784
rect 4748 4776 4756 4784
rect 5116 4776 5124 4784
rect 5292 4776 5300 4784
rect 5628 4776 5636 4784
rect 5868 4776 5876 4784
rect 2588 4758 2596 4766
rect 4860 4758 4868 4766
rect 620 4736 628 4744
rect 716 4736 724 4744
rect 892 4736 900 4744
rect 1644 4736 1652 4744
rect 4428 4736 4436 4744
rect 316 4716 324 4724
rect 364 4716 372 4724
rect 428 4716 436 4724
rect 108 4696 116 4704
rect 396 4696 404 4704
rect 524 4694 532 4702
rect 684 4696 692 4704
rect 732 4696 740 4704
rect 748 4696 756 4704
rect 780 4696 788 4704
rect 828 4716 836 4724
rect 1228 4716 1236 4724
rect 860 4696 868 4704
rect 988 4694 996 4702
rect 1052 4696 1060 4704
rect 1196 4696 1204 4704
rect 1804 4716 1812 4724
rect 2156 4716 2164 4724
rect 2588 4712 2596 4720
rect 2764 4716 2772 4724
rect 3164 4716 3172 4724
rect 3196 4716 3204 4724
rect 3308 4716 3316 4724
rect 3356 4716 3364 4724
rect 3468 4716 3476 4724
rect 3532 4716 3540 4724
rect 1276 4696 1284 4704
rect 1308 4696 1316 4704
rect 1324 4696 1332 4704
rect 1372 4696 1380 4704
rect 1532 4694 1540 4702
rect 1628 4696 1636 4704
rect 1676 4696 1684 4704
rect 1692 4696 1700 4704
rect 1772 4696 1780 4704
rect 1788 4696 1796 4704
rect 2156 4696 2164 4704
rect 2316 4696 2324 4704
rect 2412 4696 2420 4704
rect 2604 4696 2612 4704
rect 2732 4696 2740 4704
rect 2764 4696 2772 4704
rect 2988 4696 2996 4704
rect 3100 4696 3108 4704
rect 3116 4696 3124 4704
rect 3164 4696 3172 4704
rect 3260 4696 3268 4704
rect 3388 4696 3396 4704
rect 3436 4696 3444 4704
rect 3660 4716 3668 4724
rect 3724 4716 3732 4724
rect 3756 4716 3764 4724
rect 3804 4716 3812 4724
rect 4204 4716 4212 4724
rect 4268 4716 4276 4724
rect 4284 4716 4292 4724
rect 4300 4716 4308 4724
rect 4748 4716 4756 4724
rect 4860 4712 4868 4720
rect 5260 4716 5268 4724
rect 5308 4716 5316 4724
rect 5628 4716 5636 4724
rect 5836 4716 5844 4724
rect 3692 4696 3700 4704
rect 4012 4696 4020 4704
rect 4204 4696 4212 4704
rect 4236 4696 4244 4704
rect 4348 4696 4356 4704
rect 4458 4696 4466 4704
rect 4540 4696 4548 4704
rect 4716 4696 4724 4704
rect 4748 4696 4756 4704
rect 4844 4696 4852 4704
rect 5180 4696 5188 4704
rect 5628 4696 5636 4704
rect 5756 4696 5764 4704
rect 5852 4696 5860 4704
rect 5900 4716 5908 4724
rect 6060 4716 6068 4724
rect 5932 4696 5940 4704
rect 220 4676 228 4684
rect 412 4676 420 4684
rect 460 4676 468 4684
rect 556 4676 564 4684
rect 764 4676 772 4684
rect 876 4676 884 4684
rect 924 4676 932 4684
rect 956 4676 964 4684
rect 1180 4676 1188 4684
rect 1244 4676 1252 4684
rect 1292 4676 1300 4684
rect 1564 4676 1572 4684
rect 1596 4676 1604 4684
rect 1644 4676 1652 4684
rect 1852 4676 1860 4684
rect 2060 4676 2068 4684
rect 2204 4676 2212 4684
rect 2300 4676 2308 4684
rect 2524 4676 2532 4684
rect 2716 4676 2724 4684
rect 2812 4676 2820 4684
rect 3052 4676 3060 4684
rect 3196 4676 3204 4684
rect 3244 4676 3252 4684
rect 3276 4676 3284 4684
rect 3324 4676 3332 4684
rect 3356 4676 3364 4684
rect 3436 4676 3444 4684
rect 3468 4676 3476 4684
rect 3596 4676 3604 4684
rect 3708 4676 3716 4684
rect 3900 4676 3908 4684
rect 4156 4676 4164 4684
rect 4268 4676 4276 4684
rect 4300 4676 4308 4684
rect 4380 4676 4388 4684
rect 4652 4676 4660 4684
rect 4924 4676 4932 4684
rect 5212 4676 5220 4684
rect 5276 4676 5284 4684
rect 5532 4676 5540 4684
rect 5692 4676 5700 4684
rect 5772 4676 5780 4684
rect 5852 4676 5860 4684
rect 5996 4696 6004 4704
rect 6092 4696 6100 4704
rect 6172 4716 6180 4724
rect 6524 4716 6532 4724
rect 6268 4696 6276 4704
rect 6332 4696 6340 4704
rect 6348 4696 6356 4704
rect 6396 4696 6404 4704
rect 6428 4696 6436 4704
rect 6444 4696 6452 4704
rect 6492 4696 6500 4704
rect 6556 4696 6564 4704
rect 6700 4696 6708 4704
rect 6780 4696 6788 4704
rect 6012 4676 6020 4684
rect 6108 4676 6116 4684
rect 6124 4676 6132 4684
rect 6204 4676 6212 4684
rect 6220 4676 6228 4684
rect 6316 4676 6324 4684
rect 6412 4676 6420 4684
rect 6572 4676 6580 4684
rect 6748 4676 6756 4684
rect 6876 4676 6884 4684
rect 188 4656 196 4664
rect 1724 4656 1732 4664
rect 1740 4656 1748 4664
rect 1804 4656 1812 4664
rect 1836 4656 1844 4664
rect 2028 4656 2036 4664
rect 2492 4656 2500 4664
rect 2796 4656 2804 4664
rect 2956 4656 2964 4664
rect 3068 4656 3076 4664
rect 3100 4656 3108 4664
rect 3148 4656 3156 4664
rect 3212 4656 3220 4664
rect 3932 4656 3940 4664
rect 4620 4656 4628 4664
rect 4956 4656 4964 4664
rect 5500 4656 5508 4664
rect 5676 4656 5684 4664
rect 5772 4656 5780 4664
rect 28 4636 36 4644
rect 428 4636 436 4644
rect 652 4636 660 4644
rect 812 4636 820 4644
rect 908 4636 916 4644
rect 1116 4636 1124 4644
rect 1340 4636 1348 4644
rect 1404 4636 1412 4644
rect 1628 4636 1636 4644
rect 1708 4636 1716 4644
rect 1756 4636 1764 4644
rect 2924 4636 2932 4644
rect 3308 4636 3316 4644
rect 3356 4636 3364 4644
rect 3500 4636 3508 4644
rect 3548 4636 3556 4644
rect 3580 4636 3588 4644
rect 3644 4636 3652 4644
rect 4316 4636 4324 4644
rect 4428 4636 4436 4644
rect 5148 4636 5156 4644
rect 5260 4636 5268 4644
rect 6028 4636 6036 4644
rect 6140 4636 6148 4644
rect 6476 4636 6484 4644
rect 6524 4636 6532 4644
rect 6588 4636 6596 4644
rect 2638 4606 2646 4614
rect 2652 4606 2660 4614
rect 2666 4606 2674 4614
rect 5726 4606 5734 4614
rect 5740 4606 5748 4614
rect 5754 4606 5762 4614
rect 380 4576 388 4584
rect 1532 4576 1540 4584
rect 2060 4576 2068 4584
rect 3164 4576 3172 4584
rect 3404 4576 3412 4584
rect 3772 4576 3780 4584
rect 4364 4576 4372 4584
rect 4764 4576 4772 4584
rect 4924 4576 4932 4584
rect 5436 4576 5444 4584
rect 5500 4576 5508 4584
rect 5964 4576 5972 4584
rect 6108 4576 6116 4584
rect 6364 4576 6372 4584
rect 6812 4576 6820 4584
rect 844 4556 852 4564
rect 1372 4556 1380 4564
rect 1644 4556 1652 4564
rect 1948 4556 1956 4564
rect 2444 4556 2452 4564
rect 2828 4556 2836 4564
rect 3004 4556 3012 4564
rect 3084 4556 3092 4564
rect 3180 4556 3188 4564
rect 3388 4556 3396 4564
rect 3564 4556 3572 4564
rect 3612 4556 3620 4564
rect 3756 4556 3764 4564
rect 4108 4556 4116 4564
rect 4540 4556 4548 4564
rect 4780 4556 4788 4564
rect 4796 4556 4804 4564
rect 4892 4556 4900 4564
rect 5132 4556 5140 4564
rect 5308 4556 5316 4564
rect 5404 4556 5412 4564
rect 5516 4556 5524 4564
rect 5788 4556 5796 4564
rect 6092 4556 6100 4564
rect 6156 4556 6164 4564
rect 172 4536 180 4544
rect 204 4536 212 4544
rect 316 4536 324 4544
rect 428 4536 436 4544
rect 524 4536 532 4544
rect 556 4536 564 4544
rect 140 4518 148 4526
rect 220 4516 228 4524
rect 220 4496 228 4504
rect 300 4516 308 4524
rect 348 4516 356 4524
rect 268 4496 276 4504
rect 444 4516 452 4524
rect 716 4536 724 4544
rect 780 4536 788 4544
rect 988 4536 996 4544
rect 1100 4536 1108 4544
rect 1260 4536 1268 4544
rect 1452 4536 1460 4544
rect 1484 4536 1492 4544
rect 1644 4536 1652 4544
rect 1692 4536 1700 4544
rect 1820 4536 1828 4544
rect 1996 4536 2004 4544
rect 2092 4536 2100 4544
rect 396 4496 404 4504
rect 492 4496 500 4504
rect 588 4516 596 4524
rect 636 4516 644 4524
rect 652 4516 660 4524
rect 700 4516 708 4524
rect 732 4516 740 4524
rect 764 4516 772 4524
rect 844 4518 852 4526
rect 1004 4516 1012 4524
rect 668 4496 676 4504
rect 700 4496 708 4504
rect 732 4496 740 4504
rect 1036 4496 1044 4504
rect 1068 4516 1076 4524
rect 1084 4516 1092 4524
rect 1276 4516 1284 4524
rect 1388 4516 1396 4524
rect 1404 4516 1412 4524
rect 1468 4516 1476 4524
rect 1500 4516 1508 4524
rect 1548 4516 1556 4524
rect 1564 4516 1572 4524
rect 1612 4516 1620 4524
rect 1628 4516 1636 4524
rect 1676 4516 1684 4524
rect 1708 4516 1716 4524
rect 1740 4516 1748 4524
rect 1804 4518 1812 4526
rect 1964 4516 1972 4524
rect 1980 4516 1988 4524
rect 2140 4516 2148 4524
rect 2476 4536 2484 4544
rect 2796 4536 2804 4544
rect 3004 4536 3012 4544
rect 3084 4536 3092 4544
rect 3116 4536 3124 4544
rect 2188 4516 2196 4524
rect 2572 4516 2580 4524
rect 2908 4516 2916 4524
rect 3148 4536 3156 4544
rect 3196 4536 3204 4544
rect 3308 4536 3316 4544
rect 3324 4536 3332 4544
rect 3388 4536 3396 4544
rect 3436 4536 3444 4544
rect 3468 4536 3476 4544
rect 3500 4536 3508 4544
rect 3820 4536 3828 4544
rect 4140 4536 4148 4544
rect 4316 4536 4324 4544
rect 4508 4536 4516 4544
rect 4732 4536 4740 4544
rect 4812 4536 4820 4544
rect 5100 4536 5108 4544
rect 5420 4536 5428 4544
rect 5468 4536 5476 4544
rect 5820 4536 5828 4544
rect 6012 4536 6020 4544
rect 6060 4536 6068 4544
rect 6124 4536 6132 4544
rect 6252 4556 6260 4564
rect 6524 4556 6532 4564
rect 6556 4536 6564 4544
rect 6700 4536 6708 4544
rect 3148 4516 3156 4524
rect 3228 4516 3236 4524
rect 3276 4516 3284 4524
rect 3292 4516 3300 4524
rect 3356 4516 3364 4524
rect 3420 4516 3428 4524
rect 3452 4516 3460 4524
rect 3484 4516 3492 4524
rect 3516 4516 3524 4524
rect 3564 4516 3572 4524
rect 3660 4516 3668 4524
rect 3724 4516 3732 4524
rect 3788 4516 3796 4524
rect 3820 4516 3828 4524
rect 3884 4516 3892 4524
rect 4236 4516 4244 4524
rect 4508 4516 4516 4524
rect 4796 4516 4804 4524
rect 4828 4516 4836 4524
rect 4844 4516 4852 4524
rect 4956 4516 4964 4524
rect 5020 4516 5028 4524
rect 5036 4516 5044 4524
rect 5372 4516 5380 4524
rect 5596 4516 5604 4524
rect 5708 4516 5716 4524
rect 5916 4516 5924 4524
rect 5996 4516 6004 4524
rect 6028 4516 6036 4524
rect 6140 4516 6148 4524
rect 6204 4516 6212 4524
rect 6220 4516 6228 4524
rect 6316 4516 6324 4524
rect 6444 4516 6452 4524
rect 6620 4516 6628 4524
rect 1532 4496 1540 4504
rect 1740 4496 1748 4504
rect 2156 4496 2164 4504
rect 2220 4496 2228 4504
rect 2540 4500 2548 4508
rect 2732 4500 2740 4508
rect 3004 4496 3012 4504
rect 3228 4496 3236 4504
rect 3260 4496 3268 4504
rect 3324 4496 3332 4504
rect 3676 4496 3684 4504
rect 3740 4496 3748 4504
rect 3804 4496 3812 4504
rect 3868 4496 3876 4504
rect 4204 4500 4212 4508
rect 4364 4496 4372 4504
rect 4444 4500 4452 4508
rect 4764 4496 4772 4504
rect 4860 4496 4868 4504
rect 5004 4496 5012 4504
rect 5308 4496 5316 4504
rect 5468 4496 5476 4504
rect 5500 4496 5508 4504
rect 5884 4500 5892 4508
rect 5964 4496 5972 4504
rect 6172 4496 6180 4504
rect 6332 4496 6340 4504
rect 6652 4496 6660 4504
rect 1900 4476 1908 4484
rect 1932 4476 1940 4484
rect 2140 4476 2148 4484
rect 2268 4476 2276 4484
rect 3212 4476 3220 4484
rect 3644 4476 3652 4484
rect 3708 4476 3716 4484
rect 3836 4476 3844 4484
rect 3900 4476 3908 4484
rect 4892 4476 4900 4484
rect 5308 4476 5316 4484
rect 5612 4476 5620 4484
rect 6268 4476 6276 4484
rect 6300 4476 6308 4484
rect 2540 4454 2548 4462
rect 3628 4456 3636 4464
rect 3724 4456 3732 4464
rect 3884 4456 3892 4464
rect 4204 4454 4212 4462
rect 4444 4454 4452 4462
rect 5884 4454 5892 4462
rect 6284 4456 6292 4464
rect 12 4436 20 4444
rect 972 4436 980 4444
rect 1164 4436 1172 4444
rect 1356 4436 1364 4444
rect 2108 4436 2116 4444
rect 2252 4436 2260 4444
rect 2732 4436 2740 4444
rect 2988 4436 2996 4444
rect 3596 4436 3604 4444
rect 3660 4436 3668 4444
rect 3788 4436 3796 4444
rect 3948 4436 3956 4444
rect 4700 4436 4708 4444
rect 5004 4436 5012 4444
rect 5548 4436 5556 4444
rect 6652 4436 6660 4444
rect 6812 4436 6820 4444
rect 1118 4406 1126 4414
rect 1132 4406 1140 4414
rect 1146 4406 1154 4414
rect 4158 4406 4166 4414
rect 4172 4406 4180 4414
rect 4186 4406 4194 4414
rect 364 4376 372 4384
rect 684 4376 692 4384
rect 1244 4376 1252 4384
rect 1292 4376 1300 4384
rect 1372 4376 1380 4384
rect 1852 4376 1860 4384
rect 2812 4376 2820 4384
rect 3004 4376 3012 4384
rect 3084 4376 3092 4384
rect 3308 4376 3316 4384
rect 3516 4376 3524 4384
rect 3628 4376 3636 4384
rect 3692 4376 3700 4384
rect 3724 4376 3732 4384
rect 3980 4376 3988 4384
rect 4380 4376 4388 4384
rect 4460 4376 4468 4384
rect 4524 4376 4532 4384
rect 4684 4376 4692 4384
rect 5180 4376 5188 4384
rect 5292 4376 5300 4384
rect 5388 4376 5396 4384
rect 5436 4376 5444 4384
rect 5500 4376 5508 4384
rect 6300 4376 6308 4384
rect 6364 4376 6372 4384
rect 2668 4358 2676 4366
rect 4124 4358 4132 4366
rect 5628 4358 5636 4366
rect 6764 4358 6772 4366
rect 12 4336 20 4344
rect 1692 4336 1700 4344
rect 2796 4336 2804 4344
rect 3420 4336 3428 4344
rect 3644 4336 3652 4344
rect 3740 4336 3748 4344
rect 3900 4336 3908 4344
rect 140 4294 148 4302
rect 220 4296 228 4304
rect 236 4296 244 4304
rect 268 4316 276 4324
rect 428 4316 436 4324
rect 796 4316 804 4324
rect 300 4296 308 4304
rect 348 4296 356 4304
rect 396 4296 404 4304
rect 412 4296 420 4304
rect 428 4296 436 4304
rect 460 4296 468 4304
rect 540 4296 548 4304
rect 556 4296 564 4304
rect 572 4296 580 4304
rect 636 4296 644 4304
rect 668 4296 676 4304
rect 716 4296 724 4304
rect 732 4296 740 4304
rect 764 4296 772 4304
rect 844 4316 852 4324
rect 1596 4316 1604 4324
rect 1660 4316 1668 4324
rect 1772 4316 1780 4324
rect 1820 4316 1828 4324
rect 2284 4316 2292 4324
rect 2668 4312 2676 4320
rect 3036 4316 3044 4324
rect 3052 4316 3060 4324
rect 3276 4316 3284 4324
rect 3324 4316 3332 4324
rect 3676 4316 3684 4324
rect 3772 4316 3780 4324
rect 3996 4316 4004 4324
rect 4124 4312 4132 4320
rect 4684 4316 4692 4324
rect 5324 4316 5332 4324
rect 5468 4316 5476 4324
rect 5836 4316 5844 4324
rect 5964 4316 5972 4324
rect 6300 4316 6308 4324
rect 6764 4312 6772 4320
rect 844 4296 852 4304
rect 956 4296 964 4304
rect 988 4296 996 4304
rect 1068 4296 1076 4304
rect 1180 4296 1188 4304
rect 1196 4296 1204 4304
rect 1212 4296 1220 4304
rect 1324 4296 1332 4304
rect 1340 4296 1348 4304
rect 1516 4296 1524 4304
rect 1596 4296 1604 4304
rect 1628 4296 1636 4304
rect 1692 4296 1700 4304
rect 1724 4296 1732 4304
rect 1740 4296 1748 4304
rect 1788 4296 1796 4304
rect 1852 4296 1860 4304
rect 1884 4296 1892 4304
rect 2012 4296 2020 4304
rect 2060 4296 2068 4304
rect 2172 4296 2180 4304
rect 2268 4296 2276 4304
rect 2348 4296 2356 4304
rect 2604 4296 2612 4304
rect 2700 4296 2708 4304
rect 3004 4296 3012 4304
rect 3084 4296 3092 4304
rect 3132 4296 3140 4304
rect 3180 4296 3188 4304
rect 3196 4296 3204 4304
rect 3372 4296 3380 4304
rect 3404 4296 3412 4304
rect 3452 4296 3460 4304
rect 3484 4296 3492 4304
rect 3564 4296 3572 4304
rect 3596 4296 3604 4304
rect 3660 4296 3668 4304
rect 3756 4296 3764 4304
rect 3820 4296 3828 4304
rect 3884 4296 3892 4304
rect 3932 4296 3940 4304
rect 4076 4296 4084 4304
rect 4300 4296 4308 4304
rect 4492 4296 4500 4304
rect 4684 4296 4692 4304
rect 4988 4296 4996 4304
rect 5036 4296 5044 4304
rect 5260 4296 5268 4304
rect 5292 4296 5300 4304
rect 5404 4296 5412 4304
rect 5500 4296 5508 4304
rect 5628 4296 5636 4304
rect 5932 4296 5940 4304
rect 6092 4296 6100 4304
rect 6316 4296 6324 4304
rect 6588 4296 6596 4304
rect 172 4276 180 4284
rect 204 4276 212 4284
rect 316 4276 324 4284
rect 476 4276 484 4284
rect 652 4276 660 4284
rect 748 4276 756 4284
rect 860 4276 868 4284
rect 988 4276 996 4284
rect 1084 4276 1092 4284
rect 1260 4276 1268 4284
rect 1532 4276 1540 4284
rect 1644 4276 1652 4284
rect 1708 4276 1716 4284
rect 1868 4276 1876 4284
rect 1916 4276 1924 4284
rect 2204 4276 2212 4284
rect 2140 4256 2148 4264
rect 2172 4256 2180 4264
rect 2204 4256 2212 4264
rect 2252 4276 2260 4284
rect 2316 4276 2324 4284
rect 2604 4276 2612 4284
rect 2828 4276 2836 4284
rect 2972 4276 2980 4284
rect 2988 4276 2996 4284
rect 2348 4256 2356 4264
rect 2380 4256 2388 4264
rect 2412 4256 2420 4264
rect 2572 4256 2580 4264
rect 3132 4256 3140 4264
rect 3148 4256 3156 4264
rect 3212 4256 3220 4264
rect 3244 4276 3252 4284
rect 3292 4276 3300 4284
rect 3324 4276 3332 4284
rect 3372 4276 3380 4284
rect 3436 4276 3444 4284
rect 3468 4276 3476 4284
rect 3500 4276 3508 4284
rect 3548 4276 3556 4284
rect 3580 4276 3588 4284
rect 3612 4276 3620 4284
rect 3836 4276 3844 4284
rect 3916 4276 3924 4284
rect 3948 4276 3956 4284
rect 3964 4276 3972 4284
rect 4188 4276 4196 4284
rect 4636 4276 4644 4284
rect 4780 4276 4788 4284
rect 5052 4276 5060 4284
rect 5068 4276 5076 4284
rect 5196 4276 5204 4284
rect 5228 4276 5236 4284
rect 5276 4276 5284 4284
rect 5356 4276 5364 4284
rect 5516 4276 5524 4284
rect 5740 4276 5748 4284
rect 6204 4276 6212 4284
rect 6476 4276 6484 4284
rect 6700 4276 6708 4284
rect 3532 4256 3540 4264
rect 3708 4256 3716 4264
rect 4220 4256 4228 4264
rect 4428 4256 4436 4264
rect 4812 4256 4820 4264
rect 4988 4256 4996 4264
rect 5340 4256 5348 4264
rect 5708 4256 5716 4264
rect 6172 4256 6180 4264
rect 6668 4256 6676 4264
rect 508 4236 516 4244
rect 876 4236 884 4244
rect 1404 4236 1412 4244
rect 1948 4236 1956 4244
rect 2156 4236 2164 4244
rect 2236 4236 2244 4244
rect 2364 4236 2372 4244
rect 2860 4236 2868 4244
rect 3788 4236 3796 4244
rect 3852 4236 3860 4244
rect 4412 4236 4420 4244
rect 4524 4236 4532 4244
rect 5388 4236 5396 4244
rect 5548 4236 5556 4244
rect 6012 4236 6020 4244
rect 6508 4236 6516 4244
rect 2638 4206 2646 4214
rect 2652 4206 2660 4214
rect 2666 4206 2674 4214
rect 5726 4206 5734 4214
rect 5740 4206 5748 4214
rect 5754 4206 5762 4214
rect 1852 4176 1860 4184
rect 1932 4176 1940 4184
rect 2284 4176 2292 4184
rect 2492 4176 2500 4184
rect 3100 4176 3108 4184
rect 3196 4176 3204 4184
rect 3228 4176 3236 4184
rect 3308 4176 3316 4184
rect 3404 4176 3412 4184
rect 3484 4176 3492 4184
rect 4172 4176 4180 4184
rect 4924 4176 4932 4184
rect 5548 4176 5556 4184
rect 6188 4176 6196 4184
rect 6444 4176 6452 4184
rect 652 4156 660 4164
rect 876 4156 884 4164
rect 1372 4156 1380 4164
rect 1452 4156 1460 4164
rect 1548 4156 1556 4164
rect 2092 4156 2100 4164
rect 2812 4156 2820 4164
rect 3068 4156 3076 4164
rect 3164 4156 3172 4164
rect 3212 4156 3220 4164
rect 3292 4156 3300 4164
rect 3468 4156 3476 4164
rect 3532 4156 3540 4164
rect 3996 4156 4004 4164
rect 4012 4156 4020 4164
rect 4092 4156 4100 4164
rect 4332 4156 4340 4164
rect 4668 4156 4676 4164
rect 5004 4156 5012 4164
rect 5260 4156 5268 4164
rect 5580 4156 5588 4164
rect 5948 4156 5956 4164
rect 6668 4156 6676 4164
rect 204 4136 212 4144
rect 268 4136 276 4144
rect 76 4116 84 4124
rect 124 4116 132 4124
rect 220 4116 228 4124
rect 236 4116 244 4124
rect 268 4116 276 4124
rect 332 4116 340 4124
rect 348 4116 356 4124
rect 364 4116 372 4124
rect 428 4136 436 4144
rect 508 4136 516 4144
rect 556 4136 564 4144
rect 844 4136 852 4144
rect 988 4136 996 4144
rect 1164 4136 1172 4144
rect 1260 4136 1268 4144
rect 444 4116 452 4124
rect 252 4096 260 4104
rect 476 4096 484 4104
rect 524 4116 532 4124
rect 572 4116 580 4124
rect 588 4116 596 4124
rect 620 4116 628 4124
rect 636 4116 644 4124
rect 796 4116 804 4124
rect 924 4116 932 4124
rect 1036 4116 1044 4124
rect 1244 4116 1252 4124
rect 1292 4116 1300 4124
rect 1340 4116 1348 4124
rect 1356 4116 1364 4124
rect 1404 4116 1412 4124
rect 1500 4116 1508 4124
rect 1548 4116 1556 4124
rect 1628 4136 1636 4144
rect 1660 4136 1668 4144
rect 1788 4136 1796 4144
rect 1900 4136 1908 4144
rect 2124 4136 2132 4144
rect 2268 4136 2276 4144
rect 2348 4136 2356 4144
rect 2364 4136 2372 4144
rect 1644 4116 1652 4124
rect 1692 4116 1700 4124
rect 1708 4116 1716 4124
rect 1788 4116 1796 4124
rect 1804 4116 1812 4124
rect 908 4096 916 4104
rect 1212 4096 1220 4104
rect 1276 4096 1284 4104
rect 1516 4096 1524 4104
rect 1676 4096 1684 4104
rect 1740 4096 1748 4104
rect 1836 4096 1844 4104
rect 1884 4116 1892 4124
rect 2012 4116 2020 4124
rect 2188 4100 2196 4108
rect 2380 4116 2388 4124
rect 2588 4136 2596 4144
rect 2780 4136 2788 4144
rect 3084 4136 3092 4144
rect 3276 4136 3284 4144
rect 3324 4136 3332 4144
rect 2444 4116 2452 4124
rect 2316 4096 2324 4104
rect 2476 4096 2484 4104
rect 2572 4116 2580 4124
rect 2780 4116 2788 4124
rect 3260 4116 3268 4124
rect 3340 4116 3348 4124
rect 3468 4136 3476 4144
rect 3500 4136 3508 4144
rect 3580 4136 3588 4144
rect 3836 4136 3844 4144
rect 3868 4136 3876 4144
rect 3900 4136 3908 4144
rect 4028 4136 4036 4144
rect 3404 4116 3412 4124
rect 3436 4116 3444 4124
rect 3516 4116 3524 4124
rect 3532 4116 3540 4124
rect 3564 4116 3572 4124
rect 3660 4116 3668 4124
rect 3708 4116 3716 4124
rect 3788 4116 3796 4124
rect 3820 4116 3828 4124
rect 3852 4116 3860 4124
rect 3916 4116 3924 4124
rect 3948 4116 3956 4124
rect 4364 4136 4372 4144
rect 4636 4136 4644 4144
rect 4860 4136 4868 4144
rect 5020 4136 5028 4144
rect 5068 4136 5076 4144
rect 5292 4136 5300 4144
rect 5500 4136 5508 4144
rect 5596 4136 5604 4144
rect 5644 4136 5652 4144
rect 5660 4136 5668 4144
rect 5692 4136 5700 4144
rect 5980 4136 5988 4144
rect 6124 4136 6132 4144
rect 6220 4136 6228 4144
rect 6268 4136 6276 4144
rect 6284 4136 6292 4144
rect 6316 4136 6324 4144
rect 6380 4136 6388 4144
rect 6476 4136 6484 4144
rect 6700 4136 6708 4144
rect 4060 4116 4068 4124
rect 4252 4116 4260 4124
rect 4476 4116 4484 4124
rect 4540 4116 4548 4124
rect 4556 4116 4564 4124
rect 4876 4116 4884 4124
rect 4892 4116 4900 4124
rect 4956 4116 4964 4124
rect 5036 4116 5044 4124
rect 5180 4116 5188 4124
rect 5404 4116 5412 4124
rect 5484 4116 5492 4124
rect 5516 4116 5524 4124
rect 5628 4116 5636 4124
rect 5676 4116 5684 4124
rect 5868 4116 5876 4124
rect 6092 4116 6100 4124
rect 6220 4116 6228 4124
rect 6332 4116 6340 4124
rect 6588 4116 6596 4124
rect 6796 4116 6804 4124
rect 2524 4096 2532 4104
rect 2684 4096 2692 4104
rect 3004 4096 3012 4104
rect 3036 4096 3044 4104
rect 3116 4096 3124 4104
rect 3228 4096 3236 4104
rect 3356 4096 3364 4104
rect 3388 4096 3396 4104
rect 3612 4096 3620 4104
rect 188 4076 196 4084
rect 684 4076 692 4084
rect 940 4076 948 4084
rect 1276 4076 1284 4084
rect 1484 4076 1492 4084
rect 1548 4076 1556 4084
rect 3372 4076 3380 4084
rect 3596 4076 3604 4084
rect 3644 4076 3652 4084
rect 3692 4096 3700 4104
rect 3804 4096 3812 4104
rect 3932 4096 3940 4104
rect 4428 4100 4436 4108
rect 4540 4096 4548 4104
rect 4908 4096 4916 4104
rect 4924 4096 4932 4104
rect 5068 4096 5076 4104
rect 5388 4096 5396 4104
rect 5548 4096 5556 4104
rect 5564 4096 5572 4104
rect 5596 4096 5604 4104
rect 5708 4096 5716 4104
rect 6044 4100 6052 4108
rect 6236 4096 6244 4104
rect 6364 4096 6372 4104
rect 6508 4096 6516 4104
rect 6764 4100 6772 4108
rect 3708 4076 3716 4084
rect 3724 4076 3732 4084
rect 3772 4076 3780 4084
rect 3964 4076 3972 4084
rect 4124 4076 4132 4084
rect 5100 4076 5108 4084
rect 5756 4076 5764 4084
rect 2188 4054 2196 4062
rect 2780 4056 2788 4064
rect 3708 4056 3716 4064
rect 3788 4056 3796 4064
rect 3868 4056 3876 4064
rect 6044 4054 6052 4062
rect 6764 4054 6772 4062
rect 668 4036 676 4044
rect 892 4036 900 4044
rect 924 4036 932 4044
rect 1196 4036 1204 4044
rect 1292 4036 1300 4044
rect 1436 4036 1444 4044
rect 1500 4036 1508 4044
rect 1932 4036 1940 4044
rect 2972 4036 2980 4044
rect 3628 4036 3636 4044
rect 3948 4036 3956 4044
rect 4060 4036 4068 4044
rect 4428 4036 4436 4044
rect 4540 4036 4548 4044
rect 4828 4036 4836 4044
rect 5388 4036 5396 4044
rect 5452 4036 5460 4044
rect 6332 4036 6340 4044
rect 1118 4006 1126 4014
rect 1132 4006 1140 4014
rect 1146 4006 1154 4014
rect 4158 4006 4166 4014
rect 4172 4006 4180 4014
rect 4186 4006 4194 4014
rect 236 3976 244 3984
rect 284 3976 292 3984
rect 636 3976 644 3984
rect 988 3976 996 3984
rect 1212 3976 1220 3984
rect 2460 3976 2468 3984
rect 2540 3976 2548 3984
rect 2748 3976 2756 3984
rect 3340 3976 3348 3984
rect 3756 3976 3764 3984
rect 3820 3976 3828 3984
rect 3884 3976 3892 3984
rect 4780 3976 4788 3984
rect 4940 3976 4948 3984
rect 5212 3976 5220 3984
rect 5676 3976 5684 3984
rect 5836 3976 5844 3984
rect 6060 3976 6068 3984
rect 6524 3976 6532 3984
rect 6812 3976 6820 3984
rect 1324 3956 1332 3964
rect 2860 3958 2868 3966
rect 476 3936 484 3944
rect 812 3936 820 3944
rect 1340 3936 1348 3944
rect 2012 3936 2020 3944
rect 2268 3936 2276 3944
rect 2588 3936 2596 3944
rect 3436 3936 3444 3944
rect 3772 3936 3780 3944
rect 4172 3936 4180 3944
rect 4876 3936 4884 3944
rect 5004 3936 5012 3944
rect 5308 3936 5316 3944
rect 5756 3936 5764 3944
rect 6044 3936 6052 3944
rect 6076 3936 6084 3944
rect 252 3916 260 3924
rect 428 3916 436 3924
rect 44 3896 52 3904
rect 140 3896 148 3904
rect 12 3876 20 3884
rect 124 3876 132 3884
rect 300 3876 308 3884
rect 364 3896 372 3904
rect 396 3896 404 3904
rect 828 3916 836 3924
rect 908 3916 916 3924
rect 1084 3916 1092 3924
rect 1244 3916 1252 3924
rect 1260 3916 1268 3924
rect 1356 3916 1364 3924
rect 1388 3916 1396 3924
rect 1420 3916 1428 3924
rect 1452 3916 1460 3924
rect 476 3896 484 3904
rect 492 3896 500 3904
rect 572 3896 580 3904
rect 588 3896 596 3904
rect 604 3896 612 3904
rect 668 3896 676 3904
rect 684 3896 692 3904
rect 780 3896 788 3904
rect 844 3896 852 3904
rect 972 3896 980 3904
rect 1036 3896 1044 3904
rect 1052 3896 1060 3904
rect 1084 3896 1092 3904
rect 1180 3896 1188 3904
rect 1212 3896 1220 3904
rect 1292 3896 1300 3904
rect 1356 3896 1364 3904
rect 1436 3896 1444 3904
rect 1484 3896 1492 3904
rect 1532 3896 1540 3904
rect 1564 3896 1572 3904
rect 1580 3896 1588 3904
rect 1628 3896 1636 3904
rect 1724 3916 1732 3924
rect 1932 3916 1940 3924
rect 1996 3916 2004 3924
rect 2860 3912 2868 3920
rect 3132 3916 3140 3924
rect 3244 3916 3252 3924
rect 3260 3916 3268 3924
rect 3372 3916 3380 3924
rect 3628 3916 3636 3924
rect 3692 3916 3700 3924
rect 3740 3916 3748 3924
rect 3836 3916 3844 3924
rect 3884 3916 3892 3924
rect 4780 3916 4788 3924
rect 4860 3916 4868 3924
rect 5036 3916 5044 3924
rect 5116 3916 5124 3924
rect 5180 3916 5188 3924
rect 5404 3916 5412 3924
rect 332 3876 340 3884
rect 380 3876 388 3884
rect 508 3876 516 3884
rect 524 3876 532 3884
rect 796 3876 804 3884
rect 956 3876 964 3884
rect 1036 3876 1044 3884
rect 1196 3876 1204 3884
rect 1308 3876 1316 3884
rect 1436 3876 1444 3884
rect 1484 3876 1492 3884
rect 1548 3876 1556 3884
rect 1756 3896 1764 3904
rect 1788 3896 1796 3904
rect 1804 3896 1812 3904
rect 1852 3896 1860 3904
rect 1884 3896 1892 3904
rect 1948 3896 1956 3904
rect 1964 3896 1972 3904
rect 2092 3896 2100 3904
rect 2108 3896 2116 3904
rect 2316 3896 2324 3904
rect 2332 3896 2340 3904
rect 2380 3896 2388 3904
rect 2412 3896 2420 3904
rect 2428 3896 2436 3904
rect 2476 3896 2484 3904
rect 2508 3896 2516 3904
rect 2716 3896 2724 3904
rect 2764 3896 2772 3904
rect 2780 3896 2788 3904
rect 2844 3896 2852 3904
rect 3036 3896 3044 3904
rect 3148 3896 3156 3904
rect 3212 3896 3220 3904
rect 3340 3896 3348 3904
rect 3404 3896 3412 3904
rect 3484 3896 3492 3904
rect 3516 3896 3524 3904
rect 3580 3896 3588 3904
rect 3612 3896 3620 3904
rect 3692 3896 3700 3904
rect 3756 3896 3764 3904
rect 3884 3896 3892 3904
rect 4268 3896 4276 3904
rect 4316 3896 4324 3904
rect 4396 3896 4404 3904
rect 4428 3896 4436 3904
rect 4572 3896 4580 3904
rect 4780 3896 4788 3904
rect 5068 3896 5076 3904
rect 5084 3896 5092 3904
rect 5100 3896 5108 3904
rect 5148 3896 5156 3904
rect 5212 3896 5220 3904
rect 5292 3896 5300 3904
rect 5372 3896 5380 3904
rect 5452 3916 5460 3924
rect 5804 3916 5812 3924
rect 6108 3916 6116 3924
rect 5468 3896 5476 3904
rect 5548 3896 5556 3904
rect 5836 3896 5844 3904
rect 5916 3894 5924 3902
rect 6092 3896 6100 3904
rect 6140 3896 6148 3904
rect 6188 3916 6196 3924
rect 6428 3916 6436 3924
rect 6524 3916 6532 3924
rect 6364 3894 6372 3902
rect 6460 3896 6468 3904
rect 6540 3896 6548 3904
rect 1660 3876 1668 3884
rect 1772 3876 1780 3884
rect 1868 3876 1876 3884
rect 1884 3876 1892 3884
rect 1948 3876 1956 3884
rect 1996 3876 2004 3884
rect 2204 3876 2212 3884
rect 2300 3876 2308 3884
rect 2396 3876 2404 3884
rect 2572 3876 2580 3884
rect 2924 3876 2932 3884
rect 3180 3876 3188 3884
rect 3196 3876 3204 3884
rect 3292 3876 3300 3884
rect 3356 3876 3364 3884
rect 3436 3876 3444 3884
rect 3468 3876 3476 3884
rect 3500 3876 3508 3884
rect 3564 3876 3572 3884
rect 700 3856 708 3864
rect 1148 3856 1156 3864
rect 2956 3856 2964 3864
rect 3244 3856 3252 3864
rect 3436 3856 3444 3864
rect 3724 3876 3732 3884
rect 3804 3876 3812 3884
rect 3980 3876 3988 3884
rect 4364 3876 4372 3884
rect 4412 3876 4420 3884
rect 4476 3876 4484 3884
rect 4684 3876 4692 3884
rect 4828 3876 4836 3884
rect 4908 3876 4916 3884
rect 4924 3876 4932 3884
rect 5036 3876 5044 3884
rect 5100 3876 5108 3884
rect 5164 3876 5172 3884
rect 5228 3876 5236 3884
rect 5340 3876 5348 3884
rect 5356 3876 5364 3884
rect 5468 3876 5476 3884
rect 5564 3876 5572 3884
rect 5644 3876 5652 3884
rect 5788 3876 5796 3884
rect 5852 3876 5860 3884
rect 5884 3876 5892 3884
rect 5964 3876 5972 3884
rect 6124 3876 6132 3884
rect 6188 3876 6196 3884
rect 6220 3876 6228 3884
rect 6396 3876 6404 3884
rect 6476 3876 6484 3884
rect 6620 3876 6628 3884
rect 3596 3856 3604 3864
rect 3628 3856 3636 3864
rect 4012 3856 4020 3864
rect 4284 3856 4292 3864
rect 4652 3856 4660 3864
rect 5692 3856 5700 3864
rect 6652 3856 6660 3864
rect 716 3836 724 3844
rect 748 3836 756 3844
rect 876 3836 884 3844
rect 908 3836 916 3844
rect 1116 3836 1124 3844
rect 1164 3836 1172 3844
rect 1260 3836 1268 3844
rect 1708 3836 1716 3844
rect 3116 3836 3124 3844
rect 3148 3836 3156 3844
rect 3372 3836 3380 3844
rect 3516 3836 3524 3844
rect 4492 3836 4500 3844
rect 4844 3836 4852 3844
rect 4876 3836 4884 3844
rect 5004 3836 5012 3844
rect 5260 3836 5268 3844
rect 5308 3836 5316 3844
rect 5708 3836 5716 3844
rect 6236 3836 6244 3844
rect 6428 3836 6436 3844
rect 2638 3806 2646 3814
rect 2652 3806 2660 3814
rect 2666 3806 2674 3814
rect 5726 3806 5734 3814
rect 5740 3806 5748 3814
rect 5754 3806 5762 3814
rect 188 3776 196 3784
rect 220 3776 228 3784
rect 1292 3776 1300 3784
rect 1500 3776 1508 3784
rect 2252 3776 2260 3784
rect 3132 3776 3140 3784
rect 3324 3776 3332 3784
rect 3628 3776 3636 3784
rect 3996 3776 4004 3784
rect 4076 3776 4084 3784
rect 5164 3776 5172 3784
rect 5276 3776 5284 3784
rect 5436 3776 5444 3784
rect 5772 3776 5780 3784
rect 6044 3776 6052 3784
rect 6156 3776 6164 3784
rect 6364 3776 6372 3784
rect 204 3756 212 3764
rect 556 3756 564 3764
rect 572 3756 580 3764
rect 700 3756 708 3764
rect 796 3756 804 3764
rect 1340 3756 1348 3764
rect 1356 3756 1364 3764
rect 1452 3756 1460 3764
rect 1484 3756 1492 3764
rect 1772 3756 1780 3764
rect 1964 3756 1972 3764
rect 2348 3756 2356 3764
rect 2540 3756 2548 3764
rect 2876 3756 2884 3764
rect 3052 3756 3060 3764
rect 3164 3756 3172 3764
rect 3244 3756 3252 3764
rect 3260 3756 3268 3764
rect 3420 3756 3428 3764
rect 3564 3756 3572 3764
rect 3676 3756 3684 3764
rect 3980 3756 3988 3764
rect 4332 3756 4340 3764
rect 4668 3756 4676 3764
rect 5996 3756 6004 3764
rect 6060 3756 6068 3764
rect 6108 3756 6116 3764
rect 6124 3756 6132 3764
rect 6476 3756 6484 3764
rect 6700 3756 6708 3764
rect 236 3736 244 3744
rect 300 3736 308 3744
rect 364 3736 372 3744
rect 460 3736 468 3744
rect 636 3736 644 3744
rect 652 3736 660 3744
rect 732 3736 740 3744
rect 892 3736 900 3744
rect 956 3736 964 3744
rect 1244 3736 1252 3744
rect 1388 3736 1396 3744
rect 1420 3736 1428 3744
rect 1628 3736 1636 3744
rect 1756 3736 1764 3744
rect 1788 3736 1796 3744
rect 1932 3736 1940 3744
rect 2140 3736 2148 3744
rect 2204 3736 2212 3744
rect 2300 3736 2308 3744
rect 2364 3736 2372 3744
rect 2508 3736 2516 3744
rect 2716 3736 2724 3744
rect 2828 3736 2836 3744
rect 2908 3736 2916 3744
rect 3084 3736 3092 3744
rect 3164 3736 3172 3744
rect 3196 3736 3204 3744
rect 3244 3736 3252 3744
rect 3340 3736 3348 3744
rect 3612 3736 3620 3744
rect 3756 3736 3764 3744
rect 4028 3736 4036 3744
rect 4364 3736 4372 3744
rect 4636 3736 4644 3744
rect 4860 3736 4868 3744
rect 5004 3736 5012 3744
rect 5116 3736 5124 3744
rect 5212 3736 5220 3744
rect 5324 3736 5332 3744
rect 5692 3736 5700 3744
rect 5788 3736 5796 3744
rect 5820 3736 5828 3744
rect 5900 3736 5908 3744
rect 5916 3736 5924 3744
rect 6188 3736 6196 3744
rect 6204 3736 6212 3744
rect 6348 3736 6356 3744
rect 6412 3736 6420 3744
rect 6428 3736 6436 3744
rect 6732 3736 6740 3744
rect 76 3716 84 3724
rect 124 3716 132 3724
rect 252 3716 260 3724
rect 284 3696 292 3704
rect 332 3716 340 3724
rect 348 3716 356 3724
rect 380 3716 388 3724
rect 428 3716 436 3724
rect 444 3716 452 3724
rect 476 3716 484 3724
rect 524 3716 532 3724
rect 540 3716 548 3724
rect 620 3716 628 3724
rect 732 3716 740 3724
rect 796 3716 804 3724
rect 828 3716 836 3724
rect 908 3716 916 3724
rect 972 3716 980 3724
rect 1036 3716 1044 3724
rect 1148 3716 1156 3724
rect 1228 3716 1236 3724
rect 1260 3716 1268 3724
rect 1324 3716 1332 3724
rect 1404 3716 1412 3724
rect 1612 3716 1620 3724
rect 1692 3716 1700 3724
rect 1740 3716 1748 3724
rect 588 3696 596 3704
rect 700 3696 708 3704
rect 780 3696 788 3704
rect 940 3696 948 3704
rect 1004 3696 1012 3704
rect 1084 3696 1092 3704
rect 1132 3696 1140 3704
rect 1196 3696 1204 3704
rect 1372 3696 1380 3704
rect 1836 3716 1844 3724
rect 2044 3716 2052 3724
rect 2204 3716 2212 3724
rect 2220 3716 2228 3724
rect 2268 3716 2276 3724
rect 2412 3716 2420 3724
rect 2812 3716 2820 3724
rect 2844 3716 2852 3724
rect 3084 3716 3092 3724
rect 3100 3716 3108 3724
rect 3148 3716 3156 3724
rect 3260 3716 3268 3724
rect 3292 3716 3300 3724
rect 3356 3716 3364 3724
rect 3388 3716 3396 3724
rect 3468 3716 3476 3724
rect 3532 3716 3540 3724
rect 3596 3716 3604 3724
rect 3660 3716 3668 3724
rect 3708 3716 3716 3724
rect 3772 3716 3780 3724
rect 3820 3716 3828 3724
rect 3868 3716 3876 3724
rect 3932 3716 3940 3724
rect 4028 3716 4036 3724
rect 4252 3716 4260 3724
rect 4460 3716 4468 3724
rect 4556 3716 4564 3724
rect 1836 3696 1844 3704
rect 2332 3696 2340 3704
rect 2444 3700 2452 3708
rect 3132 3696 3140 3704
rect 3372 3696 3380 3704
rect 3436 3696 3444 3704
rect 3500 3696 3508 3704
rect 3548 3696 3556 3704
rect 3580 3696 3588 3704
rect 3788 3696 3796 3704
rect 620 3676 628 3684
rect 796 3676 804 3684
rect 1164 3676 1172 3684
rect 1452 3676 1460 3684
rect 2780 3676 2788 3684
rect 3404 3676 3412 3684
rect 3452 3676 3460 3684
rect 3564 3676 3572 3684
rect 3804 3676 3812 3684
rect 3852 3696 3860 3704
rect 3916 3696 3924 3704
rect 4460 3696 4468 3704
rect 4540 3696 4548 3704
rect 4828 3696 4836 3704
rect 5036 3696 5044 3704
rect 5084 3716 5092 3724
rect 5100 3716 5108 3724
rect 5180 3716 5188 3724
rect 5196 3716 5204 3724
rect 5228 3716 5236 3724
rect 5084 3696 5092 3704
rect 5260 3696 5268 3704
rect 5308 3716 5316 3724
rect 5356 3716 5364 3724
rect 5404 3716 5412 3724
rect 5468 3716 5476 3724
rect 5484 3716 5492 3724
rect 5564 3716 5572 3724
rect 5628 3718 5636 3726
rect 5772 3716 5780 3724
rect 5340 3696 5348 3704
rect 5724 3696 5732 3704
rect 5884 3716 5892 3724
rect 5980 3716 5988 3724
rect 6028 3716 6036 3724
rect 6076 3716 6084 3724
rect 6204 3716 6212 3724
rect 6268 3716 6276 3724
rect 6284 3716 6292 3724
rect 6332 3716 6340 3724
rect 6396 3716 6404 3724
rect 6508 3716 6516 3724
rect 6812 3716 6820 3724
rect 5852 3696 5860 3704
rect 6092 3696 6100 3704
rect 6252 3696 6260 3704
rect 6364 3696 6372 3704
rect 6460 3696 6468 3704
rect 6796 3700 6804 3708
rect 668 3656 676 3664
rect 1148 3656 1156 3664
rect 1228 3656 1236 3664
rect 2444 3654 2452 3662
rect 3484 3656 3492 3664
rect 3756 3656 3764 3664
rect 3884 3676 3892 3684
rect 3948 3676 3956 3684
rect 5372 3676 5380 3684
rect 6220 3676 6228 3684
rect 3932 3656 3940 3664
rect 4172 3656 4180 3664
rect 396 3636 404 3644
rect 716 3636 724 3644
rect 860 3636 868 3644
rect 908 3636 916 3644
rect 1036 3636 1044 3644
rect 1436 3636 1444 3644
rect 1836 3636 1844 3644
rect 2124 3636 2132 3644
rect 2300 3636 2308 3644
rect 3020 3636 3028 3644
rect 4012 3636 4020 3644
rect 4460 3636 4468 3644
rect 4540 3636 4548 3644
rect 4972 3636 4980 3644
rect 5388 3636 5396 3644
rect 5500 3636 5508 3644
rect 6444 3636 6452 3644
rect 6508 3636 6516 3644
rect 6540 3636 6548 3644
rect 6796 3636 6804 3644
rect 1118 3606 1126 3614
rect 1132 3606 1140 3614
rect 1146 3606 1154 3614
rect 4158 3606 4166 3614
rect 4172 3606 4180 3614
rect 4186 3606 4194 3614
rect 188 3576 196 3584
rect 572 3576 580 3584
rect 924 3576 932 3584
rect 1740 3576 1748 3584
rect 2284 3576 2292 3584
rect 2924 3576 2932 3584
rect 3068 3576 3076 3584
rect 3132 3576 3140 3584
rect 3292 3576 3300 3584
rect 3420 3576 3428 3584
rect 3580 3576 3588 3584
rect 3804 3576 3812 3584
rect 4332 3576 4340 3584
rect 4668 3576 4676 3584
rect 5772 3576 5780 3584
rect 2476 3558 2484 3566
rect 3484 3556 3492 3564
rect 4124 3558 4132 3566
rect 5196 3556 5204 3564
rect 1148 3536 1156 3544
rect 2364 3536 2372 3544
rect 2732 3536 2740 3544
rect 3116 3536 3124 3544
rect 3372 3536 3380 3544
rect 3436 3536 3444 3544
rect 3564 3536 3572 3544
rect 3756 3536 3764 3544
rect 3820 3536 3828 3544
rect 4220 3536 4228 3544
rect 4748 3536 4756 3544
rect 5164 3536 5172 3544
rect 236 3516 244 3524
rect 268 3516 276 3524
rect 380 3516 388 3524
rect 76 3496 84 3504
rect 124 3496 132 3504
rect 236 3496 244 3504
rect 300 3496 308 3504
rect 348 3496 356 3504
rect 588 3516 596 3524
rect 700 3516 708 3524
rect 428 3496 436 3504
rect 460 3496 468 3504
rect 524 3496 532 3504
rect 540 3496 548 3504
rect 620 3496 628 3504
rect 636 3496 644 3504
rect 668 3496 676 3504
rect 684 3496 692 3504
rect 732 3496 740 3504
rect 780 3496 788 3504
rect 828 3516 836 3524
rect 892 3516 900 3524
rect 1068 3516 1076 3524
rect 1180 3516 1188 3524
rect 1388 3516 1396 3524
rect 1500 3516 1508 3524
rect 1516 3516 1524 3524
rect 1548 3516 1556 3524
rect 1580 3516 1588 3524
rect 1644 3516 1652 3524
rect 1740 3516 1748 3524
rect 2172 3516 2180 3524
rect 2396 3516 2404 3524
rect 2476 3512 2484 3520
rect 2972 3516 2980 3524
rect 3020 3516 3028 3524
rect 3036 3516 3044 3524
rect 3148 3516 3156 3524
rect 3212 3516 3220 3524
rect 3404 3516 3412 3524
rect 3596 3516 3604 3524
rect 3612 3516 3620 3524
rect 3660 3516 3668 3524
rect 3788 3516 3796 3524
rect 4124 3512 4132 3520
rect 4348 3516 4356 3524
rect 4668 3516 4676 3524
rect 4812 3516 4820 3524
rect 5244 3516 5252 3524
rect 5452 3516 5460 3524
rect 5484 3516 5492 3524
rect 5516 3516 5524 3524
rect 5532 3516 5540 3524
rect 5628 3516 5636 3524
rect 6060 3516 6068 3524
rect 860 3496 868 3504
rect 924 3496 932 3504
rect 1004 3496 1012 3504
rect 1036 3496 1044 3504
rect 1148 3496 1156 3504
rect 1196 3496 1204 3504
rect 1212 3496 1220 3504
rect 1276 3496 1284 3504
rect 1324 3496 1332 3504
rect 1356 3496 1364 3504
rect 1420 3496 1428 3504
rect 1468 3496 1476 3504
rect 1564 3496 1572 3504
rect 1612 3496 1620 3504
rect 1660 3496 1668 3504
rect 1676 3496 1684 3504
rect 1756 3496 1764 3504
rect 2204 3496 2212 3504
rect 2316 3496 2324 3504
rect 2444 3496 2452 3504
rect 3068 3496 3076 3504
rect 3132 3496 3140 3504
rect 3164 3496 3172 3504
rect 3228 3496 3236 3504
rect 3244 3496 3252 3504
rect 3308 3496 3316 3504
rect 3324 3496 3332 3504
rect 3388 3496 3396 3504
rect 3420 3496 3428 3504
rect 3468 3496 3476 3504
rect 3532 3496 3540 3504
rect 3580 3496 3588 3504
rect 3612 3496 3620 3504
rect 3708 3496 3716 3504
rect 3772 3496 3780 3504
rect 3804 3496 3812 3504
rect 4156 3496 4164 3504
rect 4284 3496 4292 3504
rect 4572 3496 4580 3504
rect 4636 3496 4644 3504
rect 4780 3496 4788 3504
rect 4940 3496 4948 3504
rect 5100 3496 5108 3504
rect 5260 3496 5268 3504
rect 5276 3496 5284 3504
rect 5308 3496 5316 3504
rect 5324 3496 5332 3504
rect 5388 3496 5396 3504
rect 5420 3496 5428 3504
rect 5484 3496 5492 3504
rect 5516 3496 5524 3504
rect 5564 3496 5572 3504
rect 5740 3496 5748 3504
rect 5788 3496 5796 3504
rect 5804 3496 5812 3504
rect 5836 3496 5844 3504
rect 5884 3496 5892 3504
rect 5900 3496 5908 3504
rect 5996 3496 6004 3504
rect 6124 3496 6132 3504
rect 6140 3496 6148 3504
rect 6172 3516 6180 3524
rect 6380 3516 6388 3524
rect 6204 3496 6212 3504
rect 6236 3496 6244 3504
rect 6252 3496 6260 3504
rect 6332 3496 6340 3504
rect 6348 3496 6356 3504
rect 6428 3496 6436 3504
rect 6460 3496 6468 3504
rect 6476 3496 6484 3504
rect 6620 3496 6628 3504
rect 6700 3496 6708 3504
rect 6732 3496 6740 3504
rect 252 3476 260 3484
rect 268 3476 276 3484
rect 316 3476 324 3484
rect 332 3476 340 3484
rect 444 3476 452 3484
rect 476 3476 484 3484
rect 556 3476 564 3484
rect 748 3476 756 3484
rect 764 3476 772 3484
rect 876 3476 884 3484
rect 956 3476 964 3484
rect 1020 3476 1028 3484
rect 1132 3476 1140 3484
rect 1372 3476 1380 3484
rect 1404 3476 1412 3484
rect 1436 3476 1444 3484
rect 1452 3476 1460 3484
rect 1564 3476 1572 3484
rect 1596 3476 1604 3484
rect 1628 3476 1636 3484
rect 1692 3476 1700 3484
rect 1836 3476 1844 3484
rect 2060 3476 2068 3484
rect 2252 3476 2260 3484
rect 2300 3476 2308 3484
rect 2380 3476 2388 3484
rect 2540 3476 2548 3484
rect 2812 3476 2820 3484
rect 2988 3476 2996 3484
rect 3084 3476 3092 3484
rect 3180 3476 3188 3484
rect 3212 3476 3220 3484
rect 3260 3476 3268 3484
rect 3292 3476 3300 3484
rect 3340 3476 3348 3484
rect 3372 3476 3380 3484
rect 3468 3476 3476 3484
rect 3516 3476 3524 3484
rect 3644 3476 3652 3484
rect 3692 3476 3700 3484
rect 3724 3476 3732 3484
rect 3756 3476 3764 3484
rect 4060 3476 4068 3484
rect 4268 3476 4276 3484
rect 4300 3476 4308 3484
rect 4316 3476 4324 3484
rect 4572 3476 4580 3484
rect 4716 3476 4724 3484
rect 4764 3476 4772 3484
rect 4956 3476 4964 3484
rect 5036 3476 5044 3484
rect 5292 3476 5300 3484
rect 5404 3476 5412 3484
rect 5628 3476 5636 3484
rect 5660 3476 5668 3484
rect 5964 3476 5972 3484
rect 6108 3476 6116 3484
rect 6220 3476 6228 3484
rect 6332 3476 6340 3484
rect 6412 3476 6420 3484
rect 6460 3476 6468 3484
rect 6668 3476 6676 3484
rect 1292 3456 1300 3464
rect 1868 3456 1876 3464
rect 2236 3456 2244 3464
rect 2572 3456 2580 3464
rect 2972 3456 2980 3464
rect 3852 3456 3860 3464
rect 4028 3456 4036 3464
rect 4540 3456 4548 3464
rect 5212 3456 5220 3464
rect 5340 3456 5348 3464
rect 5612 3456 5620 3464
rect 6492 3456 6500 3464
rect 6732 3456 6740 3464
rect 6780 3456 6788 3464
rect 6796 3456 6804 3464
rect 396 3436 404 3444
rect 700 3436 708 3444
rect 812 3436 820 3444
rect 972 3436 980 3444
rect 1116 3436 1124 3444
rect 1228 3436 1236 3444
rect 1500 3436 1508 3444
rect 2092 3436 2100 3444
rect 3020 3436 3028 3444
rect 3660 3436 3668 3444
rect 4380 3436 4388 3444
rect 4732 3436 4740 3444
rect 4812 3436 4820 3444
rect 4828 3436 4836 3444
rect 5228 3436 5236 3444
rect 5852 3436 5860 3444
rect 6092 3436 6100 3444
rect 6268 3436 6276 3444
rect 6508 3436 6516 3444
rect 6716 3436 6724 3444
rect 6764 3436 6772 3444
rect 2638 3406 2646 3414
rect 2652 3406 2660 3414
rect 2666 3406 2674 3414
rect 5726 3406 5734 3414
rect 5740 3406 5748 3414
rect 5754 3406 5762 3414
rect 604 3376 612 3384
rect 652 3376 660 3384
rect 908 3376 916 3384
rect 1276 3376 1284 3384
rect 1308 3376 1316 3384
rect 1356 3376 1364 3384
rect 1580 3376 1588 3384
rect 2044 3376 2052 3384
rect 2268 3376 2276 3384
rect 3196 3376 3204 3384
rect 3324 3376 3332 3384
rect 3484 3376 3492 3384
rect 3644 3376 3652 3384
rect 3788 3376 3796 3384
rect 3804 3376 3812 3384
rect 4140 3376 4148 3384
rect 4716 3376 4724 3384
rect 4764 3376 4772 3384
rect 4908 3376 4916 3384
rect 5100 3376 5108 3384
rect 5596 3376 5604 3384
rect 6092 3376 6100 3384
rect 6428 3376 6436 3384
rect 6876 3376 6884 3384
rect 716 3356 724 3364
rect 1404 3356 1412 3364
rect 1852 3356 1860 3364
rect 2236 3356 2244 3364
rect 2300 3356 2308 3364
rect 2476 3356 2484 3364
rect 2860 3356 2868 3364
rect 3596 3356 3604 3364
rect 4268 3356 4276 3364
rect 4524 3356 4532 3364
rect 4796 3356 4804 3364
rect 5180 3356 5188 3364
rect 5196 3356 5204 3364
rect 6348 3356 6356 3364
rect 6364 3356 6372 3364
rect 252 3336 260 3344
rect 316 3336 324 3344
rect 332 3336 340 3344
rect 620 3336 628 3344
rect 700 3336 708 3344
rect 716 3336 724 3344
rect 924 3336 932 3344
rect 1180 3336 1188 3344
rect 1340 3336 1348 3344
rect 1420 3336 1428 3344
rect 76 3316 84 3324
rect 124 3316 132 3324
rect 236 3316 244 3324
rect 252 3316 260 3324
rect 300 3316 308 3324
rect 316 3316 324 3324
rect 348 3316 356 3324
rect 396 3316 404 3324
rect 412 3316 420 3324
rect 476 3318 484 3326
rect 540 3316 548 3324
rect 812 3316 820 3324
rect 844 3316 852 3324
rect 940 3316 948 3324
rect 988 3316 996 3324
rect 1084 3316 1092 3324
rect 1148 3318 1156 3326
rect 1532 3336 1540 3344
rect 1564 3336 1572 3344
rect 1596 3336 1604 3344
rect 1612 3336 1620 3344
rect 1884 3336 1892 3344
rect 2172 3336 2180 3344
rect 2204 3336 2212 3344
rect 2284 3336 2292 3344
rect 2508 3336 2516 3344
rect 2828 3336 2836 3344
rect 3036 3336 3044 3344
rect 3164 3336 3172 3344
rect 3212 3336 3220 3344
rect 3244 3336 3252 3344
rect 3276 3336 3284 3344
rect 3324 3336 3332 3344
rect 3404 3336 3412 3344
rect 3436 3336 3444 3344
rect 3484 3336 3492 3344
rect 3516 3336 3524 3344
rect 3564 3336 3572 3344
rect 3596 3336 3604 3344
rect 3612 3336 3620 3344
rect 3676 3336 3684 3344
rect 3724 3336 3732 3344
rect 3756 3336 3764 3344
rect 3836 3336 3844 3344
rect 3868 3336 3876 3344
rect 3900 3336 3908 3344
rect 3916 3336 3924 3344
rect 3964 3336 3972 3344
rect 3996 3336 4004 3344
rect 4012 3336 4020 3344
rect 4028 3336 4036 3344
rect 4076 3336 4084 3344
rect 4108 3336 4116 3344
rect 4124 3336 4132 3344
rect 4220 3336 4228 3344
rect 4284 3336 4292 3344
rect 4348 3336 4356 3344
rect 4556 3336 4564 3344
rect 4700 3336 4708 3344
rect 4748 3336 4756 3344
rect 4828 3336 4836 3344
rect 4892 3336 4900 3344
rect 5020 3336 5028 3344
rect 5052 3336 5060 3344
rect 5164 3336 5172 3344
rect 5212 3336 5220 3344
rect 5244 3336 5252 3344
rect 5308 3336 5316 3344
rect 5404 3336 5412 3344
rect 5452 3336 5460 3344
rect 5532 3336 5540 3344
rect 5564 3336 5572 3344
rect 5692 3336 5700 3344
rect 5820 3336 5828 3344
rect 5900 3336 5908 3344
rect 5948 3336 5956 3344
rect 6076 3336 6084 3344
rect 6140 3336 6148 3344
rect 6204 3336 6212 3344
rect 6220 3336 6228 3344
rect 6252 3336 6260 3344
rect 6476 3336 6484 3344
rect 6684 3336 6692 3344
rect 6716 3336 6724 3344
rect 1628 3316 1636 3324
rect 1660 3316 1668 3324
rect 1980 3316 1988 3324
rect 2076 3316 2084 3324
rect 2092 3316 2100 3324
rect 2252 3316 2260 3324
rect 2396 3316 2404 3324
rect 2940 3316 2948 3324
rect 3084 3316 3092 3324
rect 3148 3316 3156 3324
rect 3228 3316 3236 3324
rect 3292 3316 3300 3324
rect 3308 3316 3316 3324
rect 3372 3316 3380 3324
rect 3388 3316 3396 3324
rect 3452 3316 3460 3324
rect 3468 3316 3476 3324
rect 3532 3316 3540 3324
rect 3548 3316 3556 3324
rect 3612 3316 3620 3324
rect 3676 3316 3684 3324
rect 3740 3316 3748 3324
rect 3884 3316 3892 3324
rect 3916 3316 3924 3324
rect 3980 3316 3988 3324
rect 4044 3316 4052 3324
rect 4092 3316 4100 3324
rect 4236 3316 4244 3324
rect 4300 3316 4308 3324
rect 4636 3316 4644 3324
rect 4940 3316 4948 3324
rect 4956 3316 4964 3324
rect 4972 3316 4980 3324
rect 5036 3316 5044 3324
rect 5068 3316 5076 3324
rect 204 3296 212 3304
rect 268 3296 276 3304
rect 652 3296 660 3304
rect 972 3296 980 3304
rect 1036 3296 1044 3304
rect 1324 3296 1332 3304
rect 1676 3296 1684 3304
rect 1948 3300 1956 3308
rect 2124 3296 2132 3304
rect 2156 3296 2164 3304
rect 2604 3296 2612 3304
rect 2764 3300 2772 3308
rect 3036 3296 3044 3304
rect 3116 3296 3124 3304
rect 3180 3296 3188 3304
rect 3660 3296 3668 3304
rect 3788 3296 3796 3304
rect 3804 3296 3812 3304
rect 3932 3296 3940 3304
rect 4060 3296 4068 3304
rect 4156 3296 4164 3304
rect 4268 3296 4276 3304
rect 4332 3296 4340 3304
rect 4364 3296 4372 3304
rect 4620 3300 4628 3308
rect 4748 3296 4756 3304
rect 4780 3296 4788 3304
rect 4876 3296 4884 3304
rect 5148 3316 5156 3324
rect 5228 3316 5236 3324
rect 5276 3316 5284 3324
rect 5356 3316 5364 3324
rect 5420 3316 5428 3324
rect 5484 3316 5492 3324
rect 5548 3316 5556 3324
rect 5724 3318 5732 3326
rect 5852 3316 5860 3324
rect 5868 3316 5876 3324
rect 5884 3316 5892 3324
rect 5116 3296 5124 3304
rect 5260 3296 5268 3304
rect 5340 3296 5348 3304
rect 5452 3296 5460 3304
rect 5484 3296 5492 3304
rect 5516 3296 5524 3304
rect 5580 3296 5588 3304
rect 5884 3296 5892 3304
rect 5932 3316 5940 3324
rect 5980 3316 5988 3324
rect 6028 3316 6036 3324
rect 6140 3316 6148 3324
rect 6156 3316 6164 3324
rect 6236 3316 6244 3324
rect 6316 3316 6324 3324
rect 6380 3316 6388 3324
rect 6396 3316 6404 3324
rect 6444 3316 6452 3324
rect 6492 3316 6500 3324
rect 6540 3316 6548 3324
rect 6556 3316 6564 3324
rect 6620 3316 6628 3324
rect 6668 3316 6676 3324
rect 6748 3318 6756 3326
rect 6812 3316 6820 3324
rect 5980 3296 5988 3304
rect 6092 3296 6100 3304
rect 6332 3296 6340 3304
rect 6524 3296 6532 3304
rect 6636 3296 6644 3304
rect 236 3276 244 3284
rect 3244 3276 3252 3284
rect 5372 3276 5380 3284
rect 5500 3276 5508 3284
rect 5964 3276 5972 3284
rect 1948 3254 1956 3262
rect 2764 3254 2772 3262
rect 3692 3256 3700 3264
rect 4620 3254 4628 3262
rect 5996 3276 6004 3284
rect 6300 3276 6308 3284
rect 6492 3276 6500 3284
rect 6572 3276 6580 3284
rect 6668 3276 6676 3284
rect 668 3236 676 3244
rect 908 3236 916 3244
rect 1452 3236 1460 3244
rect 1628 3236 1636 3244
rect 2604 3236 2612 3244
rect 3020 3236 3028 3244
rect 3404 3236 3412 3244
rect 4844 3236 4852 3244
rect 5356 3236 5364 3244
rect 1118 3206 1126 3214
rect 1132 3206 1140 3214
rect 1146 3206 1154 3214
rect 4158 3206 4166 3214
rect 4172 3206 4180 3214
rect 4186 3206 4194 3214
rect 44 3176 52 3184
rect 652 3176 660 3184
rect 940 3176 948 3184
rect 972 3176 980 3184
rect 1020 3176 1028 3184
rect 1148 3176 1156 3184
rect 1548 3176 1556 3184
rect 1596 3176 1604 3184
rect 2348 3176 2356 3184
rect 2908 3176 2916 3184
rect 2956 3176 2964 3184
rect 3132 3176 3140 3184
rect 3692 3176 3700 3184
rect 3980 3176 3988 3184
rect 4396 3176 4404 3184
rect 4668 3176 4676 3184
rect 4860 3176 4868 3184
rect 5052 3176 5060 3184
rect 5388 3176 5396 3184
rect 5468 3176 5476 3184
rect 5532 3176 5540 3184
rect 6332 3176 6340 3184
rect 6364 3176 6372 3184
rect 1692 3156 1700 3164
rect 1948 3158 1956 3166
rect 2604 3158 2612 3166
rect 3212 3156 3220 3164
rect 4140 3158 4148 3166
rect 332 3136 340 3144
rect 1036 3136 1044 3144
rect 2108 3136 2116 3144
rect 2524 3136 2532 3144
rect 2860 3136 2868 3144
rect 3148 3136 3156 3144
rect 3340 3136 3348 3144
rect 4652 3136 4660 3144
rect 5164 3136 5172 3144
rect 5948 3136 5956 3144
rect 6860 3136 6868 3144
rect 44 3116 52 3124
rect 412 3116 420 3124
rect 76 3096 84 3104
rect 252 3096 260 3104
rect 348 3096 356 3104
rect 508 3116 516 3124
rect 604 3116 612 3124
rect 652 3116 660 3124
rect 1004 3116 1012 3124
rect 1148 3116 1156 3124
rect 1468 3116 1476 3124
rect 1532 3116 1540 3124
rect 1948 3112 1956 3120
rect 2060 3116 2068 3124
rect 2380 3116 2388 3124
rect 2604 3112 2612 3120
rect 2940 3116 2948 3124
rect 3004 3116 3012 3124
rect 3036 3116 3044 3124
rect 3116 3116 3124 3124
rect 3180 3116 3188 3124
rect 3196 3116 3204 3124
rect 3276 3116 3284 3124
rect 3308 3116 3316 3124
rect 3516 3116 3524 3124
rect 3628 3116 3636 3124
rect 3980 3116 3988 3124
rect 4140 3112 4148 3120
rect 4732 3116 4740 3124
rect 460 3096 468 3104
rect 860 3096 868 3104
rect 1020 3096 1028 3104
rect 1132 3096 1140 3104
rect 1356 3096 1364 3104
rect 1500 3096 1508 3104
rect 1660 3096 1668 3104
rect 1772 3096 1780 3104
rect 1980 3096 1988 3104
rect 2156 3096 2164 3104
rect 2220 3096 2228 3104
rect 2428 3096 2436 3104
rect 2444 3096 2452 3104
rect 2572 3096 2580 3104
rect 3004 3096 3012 3104
rect 3036 3096 3044 3104
rect 3116 3096 3124 3104
rect 3164 3096 3172 3104
rect 3244 3096 3252 3104
rect 140 3076 148 3084
rect 364 3076 372 3084
rect 428 3076 436 3084
rect 556 3076 564 3084
rect 572 3076 580 3084
rect 748 3076 756 3084
rect 1244 3076 1252 3084
rect 1516 3076 1524 3084
rect 1564 3076 1572 3084
rect 1884 3076 1892 3084
rect 2028 3076 2036 3084
rect 2060 3076 2068 3084
rect 2172 3076 2180 3084
rect 2268 3076 2276 3084
rect 2364 3076 2372 3084
rect 2412 3076 2420 3084
rect 2428 3076 2436 3084
rect 2460 3076 2468 3084
rect 2668 3076 2676 3084
rect 2892 3076 2900 3084
rect 2972 3076 2980 3084
rect 2988 3076 2996 3084
rect 3084 3076 3092 3084
rect 3228 3076 3236 3084
rect 3420 3096 3428 3104
rect 3484 3096 3492 3104
rect 3580 3096 3588 3104
rect 3628 3096 3636 3104
rect 3948 3096 3956 3104
rect 4108 3096 4116 3104
rect 4316 3096 4324 3104
rect 4524 3096 4532 3104
rect 4700 3096 4708 3104
rect 4748 3096 4756 3104
rect 4812 3096 4820 3104
rect 4828 3096 4836 3104
rect 4860 3096 4868 3104
rect 4908 3116 4916 3124
rect 4972 3116 4980 3124
rect 5068 3116 5076 3124
rect 5356 3116 5364 3124
rect 5420 3116 5428 3124
rect 5500 3116 5508 3124
rect 5612 3116 5620 3124
rect 5628 3116 5636 3124
rect 6012 3116 6020 3124
rect 4940 3096 4948 3104
rect 5004 3096 5012 3104
rect 5084 3096 5092 3104
rect 5132 3096 5140 3104
rect 5164 3096 5172 3104
rect 5180 3096 5188 3104
rect 5292 3096 5300 3104
rect 5324 3096 5332 3104
rect 5388 3096 5396 3104
rect 5436 3096 5444 3104
rect 5532 3096 5540 3104
rect 5580 3096 5588 3104
rect 5676 3096 5684 3104
rect 5836 3096 5844 3104
rect 5980 3096 5988 3104
rect 6284 3116 6292 3124
rect 6060 3096 6068 3104
rect 6092 3096 6100 3104
rect 6108 3096 6116 3104
rect 6156 3096 6164 3104
rect 6188 3096 6196 3104
rect 6604 3116 6612 3124
rect 6332 3096 6340 3104
rect 6428 3096 6436 3104
rect 6460 3096 6468 3104
rect 6524 3096 6532 3104
rect 6540 3096 6548 3104
rect 6572 3096 6580 3104
rect 6636 3096 6644 3104
rect 6652 3096 6660 3104
rect 6732 3094 6740 3102
rect 3372 3076 3380 3084
rect 3436 3076 3444 3084
rect 3468 3076 3476 3084
rect 3532 3076 3540 3084
rect 3596 3076 3604 3084
rect 3612 3076 3620 3084
rect 3884 3076 3892 3084
rect 4204 3076 4212 3084
rect 4444 3076 4452 3084
rect 4476 3076 4484 3084
rect 4684 3076 4692 3084
rect 4748 3076 4756 3084
rect 4844 3076 4852 3084
rect 4956 3076 4964 3084
rect 4988 3076 4996 3084
rect 5020 3076 5028 3084
rect 5116 3076 5124 3084
rect 172 3056 180 3064
rect 508 3056 516 3064
rect 780 3056 788 3064
rect 988 3056 996 3064
rect 1276 3056 1284 3064
rect 1580 3056 1588 3064
rect 1852 3056 1860 3064
rect 2700 3056 2708 3064
rect 3068 3056 3076 3064
rect 3580 3056 3588 3064
rect 3852 3056 3860 3064
rect 4236 3056 4244 3064
rect 4412 3056 4420 3064
rect 4652 3056 4660 3064
rect 4796 3056 4804 3064
rect 5036 3056 5044 3064
rect 5228 3076 5236 3084
rect 5308 3076 5316 3084
rect 5548 3076 5556 3084
rect 5564 3076 5572 3084
rect 5596 3076 5604 3084
rect 5628 3076 5636 3084
rect 5788 3076 5796 3084
rect 5964 3076 5972 3084
rect 6076 3076 6084 3084
rect 6252 3076 6260 3084
rect 6348 3076 6356 3084
rect 6396 3076 6404 3084
rect 6556 3076 6564 3084
rect 6668 3076 6676 3084
rect 6764 3076 6772 3084
rect 5708 3056 5716 3064
rect 6124 3056 6132 3064
rect 6412 3056 6420 3064
rect 6444 3056 6452 3064
rect 6508 3056 6516 3064
rect 540 3036 548 3044
rect 588 3036 596 3044
rect 1468 3036 1476 3044
rect 1628 3036 1636 3044
rect 2044 3036 2052 3044
rect 2188 3036 2196 3044
rect 2316 3036 2324 3044
rect 3324 3036 3332 3044
rect 3452 3036 3460 3044
rect 3548 3036 3556 3044
rect 4396 3036 4404 3044
rect 5260 3036 5268 3044
rect 6028 3036 6036 3044
rect 6220 3036 6228 3044
rect 2638 3006 2646 3014
rect 2652 3006 2660 3014
rect 2666 3006 2674 3014
rect 5726 3006 5734 3014
rect 5740 3006 5748 3014
rect 5754 3006 5762 3014
rect 492 2976 500 2984
rect 556 2976 564 2984
rect 1100 2976 1108 2984
rect 2908 2976 2916 2984
rect 3308 2976 3316 2984
rect 3692 2976 3700 2984
rect 4076 2976 4084 2984
rect 4524 2976 4532 2984
rect 4876 2976 4884 2984
rect 5084 2976 5092 2984
rect 5420 2976 5428 2984
rect 5804 2976 5812 2984
rect 6140 2976 6148 2984
rect 6396 2976 6404 2984
rect 6492 2976 6500 2984
rect 6508 2976 6516 2984
rect 6812 2976 6820 2984
rect 12 2956 20 2964
rect 428 2956 436 2964
rect 780 2956 788 2964
rect 1340 2956 1348 2964
rect 1804 2956 1812 2964
rect 2220 2956 2228 2964
rect 2508 2956 2516 2964
rect 2748 2956 2756 2964
rect 3596 2956 3604 2964
rect 3644 2956 3652 2964
rect 3852 2956 3860 2964
rect 4140 2956 4148 2964
rect 4364 2956 4372 2964
rect 4636 2956 4644 2964
rect 4764 2956 4772 2964
rect 5068 2956 5076 2964
rect 5500 2956 5508 2964
rect 6204 2956 6212 2964
rect 6316 2956 6324 2964
rect 6332 2956 6340 2964
rect 156 2936 164 2944
rect 204 2936 212 2944
rect 236 2936 244 2944
rect 268 2936 276 2944
rect 284 2936 292 2944
rect 444 2936 452 2944
rect 540 2936 548 2944
rect 604 2936 612 2944
rect 748 2936 756 2944
rect 956 2936 964 2944
rect 1068 2936 1076 2944
rect 1116 2936 1124 2944
rect 1308 2936 1316 2944
rect 1532 2936 1540 2944
rect 1628 2936 1636 2944
rect 1772 2936 1780 2944
rect 1996 2936 2004 2944
rect 2028 2936 2036 2944
rect 2188 2936 2196 2944
rect 2412 2936 2420 2944
rect 2444 2936 2452 2944
rect 2716 2936 2724 2944
rect 60 2916 68 2924
rect 140 2916 148 2924
rect 268 2916 276 2924
rect 300 2916 308 2924
rect 108 2896 116 2904
rect 332 2896 340 2904
rect 380 2916 388 2924
rect 476 2896 484 2904
rect 524 2916 532 2924
rect 604 2916 612 2924
rect 860 2916 868 2924
rect 1052 2916 1060 2924
rect 1420 2916 1428 2924
rect 1612 2916 1620 2924
rect 1708 2916 1716 2924
rect 2012 2916 2020 2924
rect 2188 2916 2196 2924
rect 2828 2916 2836 2924
rect 2956 2916 2964 2924
rect 3004 2916 3012 2924
rect 3084 2916 3092 2924
rect 3148 2916 3156 2924
rect 3276 2936 3284 2944
rect 3212 2916 3220 2924
rect 3452 2916 3460 2924
rect 3884 2936 3892 2944
rect 4332 2936 4340 2944
rect 4540 2936 4548 2944
rect 4652 2936 4660 2944
rect 4716 2936 4724 2944
rect 4812 2936 4820 2944
rect 4860 2936 4868 2944
rect 5004 2936 5012 2944
rect 5260 2936 5268 2944
rect 3564 2916 3572 2924
rect 3612 2916 3620 2924
rect 3628 2916 3636 2924
rect 3948 2916 3956 2924
rect 4028 2916 4036 2924
rect 4044 2916 4052 2924
rect 4268 2916 4276 2924
rect 4332 2916 4340 2924
rect 4588 2916 4596 2924
rect 4636 2916 4644 2924
rect 4732 2916 4740 2924
rect 4780 2916 4788 2924
rect 4796 2916 4804 2924
rect 4828 2916 4836 2924
rect 4972 2916 4980 2924
rect 5116 2916 5124 2924
rect 5164 2916 5172 2924
rect 5180 2916 5188 2924
rect 5212 2916 5220 2924
rect 5228 2916 5236 2924
rect 5324 2916 5332 2924
rect 5340 2916 5348 2924
rect 5388 2916 5396 2924
rect 5452 2916 5460 2924
rect 5516 2916 5524 2924
rect 5644 2916 5652 2924
rect 5692 2916 5700 2924
rect 5820 2916 5828 2924
rect 5836 2916 5844 2924
rect 5884 2916 5892 2924
rect 5916 2916 5924 2924
rect 5932 2916 5940 2924
rect 5980 2916 5988 2924
rect 6012 2936 6020 2944
rect 6124 2936 6132 2944
rect 6188 2936 6196 2944
rect 6252 2936 6260 2944
rect 6300 2936 6308 2944
rect 6444 2936 6452 2944
rect 6668 2936 6676 2944
rect 6700 2936 6708 2944
rect 556 2896 564 2904
rect 684 2900 692 2908
rect 940 2896 948 2904
rect 972 2896 980 2904
rect 1004 2896 1012 2904
rect 1084 2896 1092 2904
rect 1212 2896 1220 2904
rect 1532 2896 1540 2904
rect 1676 2896 1684 2904
rect 1964 2896 1972 2904
rect 2044 2896 2052 2904
rect 2124 2900 2132 2908
rect 2476 2896 2484 2904
rect 2524 2896 2532 2904
rect 2652 2900 2660 2908
rect 3228 2896 3236 2904
rect 3244 2896 3252 2904
rect 3372 2896 3380 2904
rect 3468 2896 3476 2904
rect 3980 2896 3988 2904
rect 4236 2896 4244 2904
rect 4556 2896 4564 2904
rect 4700 2896 4708 2904
rect 4860 2896 4868 2904
rect 5196 2896 5204 2904
rect 5308 2896 5316 2904
rect 5420 2896 5428 2904
rect 6108 2916 6116 2924
rect 6172 2916 6180 2924
rect 6236 2916 6244 2924
rect 6252 2916 6260 2924
rect 6348 2916 6356 2924
rect 6364 2916 6372 2924
rect 6412 2916 6420 2924
rect 6460 2916 6468 2924
rect 6620 2916 6628 2924
rect 6076 2896 6084 2904
rect 6140 2896 6148 2904
rect 6204 2896 6212 2904
rect 6268 2896 6276 2904
rect 172 2876 180 2884
rect 1500 2876 1508 2884
rect 1564 2876 1572 2884
rect 2972 2876 2980 2884
rect 3068 2876 3076 2884
rect 3132 2876 3140 2884
rect 3228 2876 3236 2884
rect 3324 2876 3332 2884
rect 3388 2876 3396 2884
rect 3436 2876 3444 2884
rect 2124 2854 2132 2862
rect 3212 2856 3220 2864
rect 3484 2876 3492 2884
rect 3516 2876 3524 2884
rect 5868 2876 5876 2884
rect 6028 2856 6036 2864
rect 60 2836 68 2844
rect 380 2836 388 2844
rect 684 2836 692 2844
rect 1212 2836 1220 2844
rect 1676 2836 1684 2844
rect 2428 2836 2436 2844
rect 2652 2836 2660 2844
rect 2956 2836 2964 2844
rect 3084 2836 3092 2844
rect 3148 2836 3156 2844
rect 3260 2836 3268 2844
rect 3372 2836 3380 2844
rect 3500 2836 3508 2844
rect 3980 2836 3988 2844
rect 4236 2836 4244 2844
rect 5148 2836 5156 2844
rect 5276 2836 5284 2844
rect 5356 2836 5364 2844
rect 5548 2836 5556 2844
rect 1118 2806 1126 2814
rect 1132 2806 1140 2814
rect 1146 2806 1154 2814
rect 4158 2806 4166 2814
rect 4172 2806 4180 2814
rect 4186 2806 4194 2814
rect 44 2776 52 2784
rect 332 2776 340 2784
rect 684 2776 692 2784
rect 972 2776 980 2784
rect 1020 2776 1028 2784
rect 1052 2776 1060 2784
rect 1196 2776 1204 2784
rect 1324 2776 1332 2784
rect 1900 2776 1908 2784
rect 2188 2776 2196 2784
rect 2236 2776 2244 2784
rect 2300 2776 2308 2784
rect 2588 2776 2596 2784
rect 2892 2776 2900 2784
rect 3580 2776 3588 2784
rect 3788 2776 3796 2784
rect 3948 2776 3956 2784
rect 4300 2776 4308 2784
rect 4636 2776 4644 2784
rect 4684 2776 4692 2784
rect 5020 2776 5028 2784
rect 5036 2776 5044 2784
rect 5292 2776 5300 2784
rect 5580 2776 5588 2784
rect 5612 2776 5620 2784
rect 6204 2776 6212 2784
rect 6252 2776 6260 2784
rect 1628 2758 1636 2766
rect 3004 2758 3012 2766
rect 3340 2756 3348 2764
rect 5836 2756 5844 2764
rect 6668 2756 6676 2764
rect 1372 2736 1380 2744
rect 2764 2736 2772 2744
rect 44 2716 52 2724
rect 508 2716 516 2724
rect 652 2716 660 2724
rect 972 2716 980 2724
rect 1084 2716 1092 2724
rect 1628 2712 1636 2720
rect 1708 2716 1716 2724
rect 1740 2716 1748 2724
rect 2188 2716 2196 2724
rect 2588 2716 2596 2724
rect 2748 2716 2756 2724
rect 2812 2716 2820 2724
rect 2844 2716 2852 2724
rect 2924 2716 2932 2724
rect 3004 2712 3012 2720
rect 3324 2716 3332 2724
rect 3404 2716 3412 2724
rect 3452 2716 3460 2724
rect 3468 2716 3476 2724
rect 3612 2716 3620 2724
rect 3628 2716 3636 2724
rect 3756 2716 3764 2724
rect 3772 2716 3780 2724
rect 3804 2716 3812 2724
rect 4060 2736 4068 2744
rect 6460 2736 6468 2744
rect 6636 2736 6644 2744
rect 4300 2716 4308 2724
rect 4684 2716 4692 2724
rect 5212 2716 5220 2724
rect 5388 2716 5396 2724
rect 5596 2716 5604 2724
rect 5884 2716 5892 2724
rect 5916 2716 5924 2724
rect 5948 2716 5956 2724
rect 6124 2716 6132 2724
rect 252 2696 260 2704
rect 540 2696 548 2704
rect 764 2696 772 2704
rect 972 2696 980 2704
rect 1644 2696 1652 2704
rect 1788 2696 1796 2704
rect 1884 2696 1892 2704
rect 2188 2696 2196 2704
rect 2236 2696 2244 2704
rect 2380 2696 2388 2704
rect 2588 2696 2596 2704
rect 2684 2696 2692 2704
rect 2780 2696 2788 2704
rect 140 2676 148 2684
rect 364 2676 372 2684
rect 492 2676 500 2684
rect 556 2676 564 2684
rect 604 2676 612 2684
rect 876 2676 884 2684
rect 1116 2676 1124 2684
rect 1308 2676 1316 2684
rect 1564 2676 1572 2684
rect 1708 2676 1716 2684
rect 1804 2676 1812 2684
rect 2092 2676 2100 2684
rect 2492 2676 2500 2684
rect 2716 2676 2724 2684
rect 2844 2696 2852 2704
rect 2860 2696 2868 2704
rect 2972 2696 2980 2704
rect 3500 2696 3508 2704
rect 3580 2696 3588 2704
rect 3612 2696 3620 2704
rect 3676 2696 3684 2704
rect 3788 2696 3796 2704
rect 3884 2696 3892 2704
rect 3900 2696 3908 2704
rect 3980 2696 3988 2704
rect 2860 2676 2868 2684
rect 2876 2676 2884 2684
rect 3068 2676 3076 2684
rect 3262 2676 3270 2684
rect 3292 2676 3300 2684
rect 3356 2676 3364 2684
rect 3548 2676 3556 2684
rect 3708 2676 3716 2684
rect 3836 2676 3844 2684
rect 4092 2696 4100 2704
rect 4108 2696 4116 2704
rect 4332 2696 4340 2704
rect 4508 2696 4516 2704
rect 4684 2696 4692 2704
rect 5244 2696 5252 2704
rect 5324 2696 5332 2704
rect 5356 2696 5364 2704
rect 5388 2696 5396 2704
rect 5452 2694 5460 2702
rect 5628 2696 5636 2704
rect 5708 2696 5716 2704
rect 5724 2696 5732 2704
rect 5804 2696 5812 2704
rect 5852 2696 5860 2704
rect 5868 2696 5876 2704
rect 5948 2696 5956 2704
rect 5980 2696 5988 2704
rect 5996 2696 6004 2704
rect 6092 2696 6100 2704
rect 6236 2716 6244 2724
rect 6428 2716 6436 2724
rect 6492 2716 6500 2724
rect 6540 2716 6548 2724
rect 6604 2716 6612 2724
rect 6172 2696 6180 2704
rect 6284 2696 6292 2704
rect 6300 2696 6308 2704
rect 6348 2696 6356 2704
rect 6396 2696 6404 2704
rect 6460 2696 6468 2704
rect 6524 2696 6532 2704
rect 6572 2696 6580 2704
rect 6588 2696 6596 2704
rect 6636 2696 6644 2704
rect 6732 2696 6740 2704
rect 6764 2696 6772 2704
rect 4396 2676 4404 2684
rect 4780 2676 4788 2684
rect 5068 2676 5076 2684
rect 5196 2676 5204 2684
rect 5292 2676 5300 2684
rect 5340 2676 5348 2684
rect 5420 2676 5428 2684
rect 5628 2676 5636 2684
rect 5932 2676 5940 2684
rect 5996 2676 6004 2684
rect 6044 2676 6052 2684
rect 6076 2676 6084 2684
rect 6188 2676 6196 2684
rect 6268 2676 6276 2684
rect 6364 2676 6372 2684
rect 6412 2676 6420 2684
rect 6444 2676 6452 2684
rect 6652 2676 6660 2684
rect 172 2656 180 2664
rect 572 2656 580 2664
rect 844 2656 852 2664
rect 1036 2656 1044 2664
rect 1068 2656 1076 2664
rect 1084 2656 1092 2664
rect 1340 2656 1348 2664
rect 1532 2656 1540 2664
rect 2060 2656 2068 2664
rect 2284 2656 2292 2664
rect 2460 2656 2468 2664
rect 3100 2656 3108 2664
rect 3436 2656 3444 2664
rect 3548 2656 3556 2664
rect 3708 2656 3716 2664
rect 4252 2656 4260 2664
rect 4428 2656 4436 2664
rect 4620 2656 4628 2664
rect 4812 2656 4820 2664
rect 5052 2656 5060 2664
rect 6220 2656 6228 2664
rect 508 2636 516 2644
rect 652 2636 660 2644
rect 1836 2636 1844 2644
rect 2300 2636 2308 2644
rect 3292 2636 3300 2644
rect 3324 2636 3332 2644
rect 3468 2636 3476 2644
rect 3740 2636 3748 2644
rect 3852 2636 3860 2644
rect 4012 2636 4020 2644
rect 4044 2636 4052 2644
rect 4140 2636 4148 2644
rect 4972 2636 4980 2644
rect 5212 2636 5220 2644
rect 5676 2636 5684 2644
rect 5948 2636 5956 2644
rect 6140 2636 6148 2644
rect 6316 2636 6324 2644
rect 2638 2606 2646 2614
rect 2652 2606 2660 2614
rect 2666 2606 2674 2614
rect 5726 2606 5734 2614
rect 5740 2606 5748 2614
rect 5754 2606 5762 2614
rect 3804 2596 3812 2604
rect 3932 2596 3940 2604
rect 124 2576 132 2584
rect 892 2576 900 2584
rect 1292 2576 1300 2584
rect 2172 2576 2180 2584
rect 2252 2576 2260 2584
rect 2748 2576 2756 2584
rect 3580 2576 3588 2584
rect 3948 2576 3956 2584
rect 4028 2576 4036 2584
rect 4060 2576 4068 2584
rect 4556 2576 4564 2584
rect 4636 2576 4644 2584
rect 4892 2576 4900 2584
rect 5468 2576 5476 2584
rect 6012 2576 6020 2584
rect 6028 2576 6036 2584
rect 6220 2576 6228 2584
rect 6876 2576 6884 2584
rect 108 2556 116 2564
rect 140 2556 148 2564
rect 316 2556 324 2564
rect 668 2556 676 2564
rect 1052 2556 1060 2564
rect 1564 2556 1572 2564
rect 1692 2556 1700 2564
rect 1820 2556 1828 2564
rect 2012 2556 2020 2564
rect 2204 2556 2212 2564
rect 2412 2556 2420 2564
rect 2588 2556 2596 2564
rect 2908 2556 2916 2564
rect 3292 2556 3300 2564
rect 3804 2556 3812 2564
rect 3932 2556 3940 2564
rect 4108 2556 4116 2564
rect 4396 2556 4404 2564
rect 4700 2556 4708 2564
rect 4972 2556 4980 2564
rect 5100 2556 5108 2564
rect 5276 2556 5284 2564
rect 5436 2556 5444 2564
rect 5596 2556 5604 2564
rect 5884 2556 5892 2564
rect 60 2536 68 2544
rect 348 2536 356 2544
rect 700 2536 708 2544
rect 1084 2536 1092 2544
rect 1420 2536 1428 2544
rect 1596 2536 1604 2544
rect 1836 2536 1844 2544
rect 1980 2536 1988 2544
rect 2444 2536 2452 2544
rect 2700 2536 2708 2544
rect 2940 2536 2948 2544
rect 44 2516 52 2524
rect 108 2516 116 2524
rect 236 2516 244 2524
rect 444 2516 452 2524
rect 588 2516 596 2524
rect 764 2516 772 2524
rect 1180 2516 1188 2524
rect 1660 2516 1668 2524
rect 1676 2516 1684 2524
rect 1788 2516 1796 2524
rect 1804 2516 1812 2524
rect 1868 2516 1876 2524
rect 2092 2516 2100 2524
rect 2444 2516 2452 2524
rect 2684 2516 2692 2524
rect 3020 2516 3028 2524
rect 3100 2516 3108 2524
rect 3260 2536 3268 2544
rect 3276 2536 3284 2544
rect 3340 2536 3348 2544
rect 3356 2536 3364 2544
rect 3404 2536 3412 2544
rect 3532 2536 3540 2544
rect 3596 2536 3604 2544
rect 3612 2536 3620 2544
rect 3676 2536 3684 2544
rect 3692 2536 3700 2544
rect 3740 2536 3748 2544
rect 3804 2536 3812 2544
rect 3980 2536 3988 2544
rect 3164 2516 3172 2524
rect 3244 2516 3252 2524
rect 3292 2516 3300 2524
rect 3324 2516 3332 2524
rect 3580 2516 3588 2524
rect 3596 2516 3604 2524
rect 3660 2516 3668 2524
rect 3724 2516 3732 2524
rect 3836 2516 3844 2524
rect 3868 2516 3876 2524
rect 3996 2516 4004 2524
rect 4364 2536 4372 2544
rect 4716 2536 4724 2544
rect 4844 2536 4852 2544
rect 5068 2536 5076 2544
rect 5244 2536 5252 2544
rect 5660 2536 5668 2544
rect 5756 2536 5764 2544
rect 5820 2536 5828 2544
rect 6188 2536 6196 2544
rect 6460 2536 6468 2544
rect 6524 2536 6532 2544
rect 6636 2536 6644 2544
rect 6716 2536 6724 2544
rect 4268 2516 4276 2524
rect 4572 2516 4580 2524
rect 4604 2516 4612 2524
rect 4860 2516 4868 2524
rect 4876 2516 4884 2524
rect 4988 2516 4996 2524
rect 5004 2516 5012 2524
rect 5148 2516 5156 2524
rect 5580 2516 5588 2524
rect 5676 2516 5684 2524
rect 444 2496 452 2504
rect 508 2496 516 2504
rect 796 2496 804 2504
rect 1148 2500 1156 2508
rect 1916 2500 1924 2508
rect 2508 2500 2516 2508
rect 2716 2496 2724 2504
rect 3004 2500 3012 2508
rect 3212 2496 3220 2504
rect 3244 2496 3252 2504
rect 3388 2496 3396 2504
rect 3548 2496 3556 2504
rect 3580 2496 3588 2504
rect 3724 2496 3732 2504
rect 3788 2496 3796 2504
rect 3852 2496 3860 2504
rect 3916 2496 3924 2504
rect 3932 2496 3940 2504
rect 4124 2496 4132 2504
rect 4300 2500 4308 2508
rect 5180 2500 5188 2508
rect 5804 2516 5812 2524
rect 5884 2518 5892 2526
rect 6124 2516 6132 2524
rect 6284 2516 6292 2524
rect 6332 2516 6340 2524
rect 6444 2516 6452 2524
rect 6460 2516 6468 2524
rect 6524 2516 6532 2524
rect 6556 2516 6564 2524
rect 6572 2516 6580 2524
rect 6604 2516 6612 2524
rect 6620 2516 6628 2524
rect 6652 2516 6660 2524
rect 6684 2516 6692 2524
rect 6748 2518 6756 2526
rect 5772 2496 5780 2504
rect 6412 2496 6420 2504
rect 6476 2496 6484 2504
rect 6684 2496 6692 2504
rect 12 2476 20 2484
rect 3116 2476 3124 2484
rect 3180 2476 3188 2484
rect 3884 2476 3892 2484
rect 4156 2476 4164 2484
rect 6444 2476 6452 2484
rect 1148 2454 1156 2462
rect 1916 2454 1924 2462
rect 2508 2454 2516 2462
rect 3004 2454 3012 2462
rect 3900 2456 3908 2464
rect 4140 2456 4148 2464
rect 4300 2454 4308 2462
rect 5180 2454 5188 2462
rect 444 2436 452 2444
rect 796 2436 804 2444
rect 844 2436 852 2444
rect 1532 2436 1540 2444
rect 1756 2436 1764 2444
rect 2220 2436 2228 2444
rect 3100 2436 3108 2444
rect 3164 2436 3172 2444
rect 3372 2436 3380 2444
rect 3628 2436 3636 2444
rect 3708 2436 3716 2444
rect 3756 2436 3764 2444
rect 3868 2436 3876 2444
rect 4028 2436 4036 2444
rect 1118 2406 1126 2414
rect 1132 2406 1140 2414
rect 1146 2406 1154 2414
rect 4158 2406 4166 2414
rect 4172 2406 4180 2414
rect 4186 2406 4194 2414
rect 204 2376 212 2384
rect 524 2376 532 2384
rect 828 2376 836 2384
rect 908 2376 916 2384
rect 1196 2376 1204 2384
rect 1404 2376 1412 2384
rect 2268 2376 2276 2384
rect 2844 2376 2852 2384
rect 3548 2376 3556 2384
rect 3740 2376 3748 2384
rect 3836 2376 3844 2384
rect 3900 2376 3908 2384
rect 4508 2376 4516 2384
rect 5500 2376 5508 2384
rect 6060 2376 6068 2384
rect 6108 2376 6116 2384
rect 6332 2376 6340 2384
rect 6668 2376 6676 2384
rect 1660 2358 1668 2366
rect 2140 2358 2148 2366
rect 2444 2358 2452 2366
rect 3244 2358 3252 2366
rect 4604 2358 4612 2366
rect 5084 2358 5092 2366
rect 2908 2336 2916 2344
rect 3756 2336 3764 2344
rect 3820 2336 3828 2344
rect 524 2316 532 2324
rect 908 2316 916 2324
rect 1660 2312 1668 2320
rect 2140 2312 2148 2320
rect 2316 2316 2324 2324
rect 2444 2312 2452 2320
rect 2940 2316 2948 2324
rect 2956 2316 2964 2324
rect 3100 2316 3108 2324
rect 3164 2316 3172 2324
rect 3244 2312 3252 2320
rect 188 2296 196 2304
rect 524 2296 532 2304
rect 588 2296 596 2304
rect 636 2296 644 2304
rect 652 2296 660 2304
rect 700 2296 708 2304
rect 764 2296 772 2304
rect 780 2296 788 2304
rect 796 2296 804 2304
rect 844 2296 852 2304
rect 908 2296 916 2304
rect 1116 2296 1124 2304
rect 1276 2296 1284 2304
rect 1372 2296 1380 2304
rect 1484 2296 1492 2304
rect 1676 2296 1684 2304
rect 1836 2296 1844 2304
rect 1852 2296 1860 2304
rect 2172 2296 2180 2304
rect 2220 2296 2228 2304
rect 2284 2296 2292 2304
rect 2300 2296 2308 2304
rect 2332 2296 2340 2304
rect 2348 2296 2356 2304
rect 2396 2296 2404 2304
rect 2620 2296 2628 2304
rect 2702 2296 2710 2304
rect 3004 2296 3012 2304
rect 3068 2296 3076 2304
rect 3132 2296 3140 2304
rect 3164 2296 3172 2304
rect 3228 2296 3236 2304
rect 3612 2316 3620 2324
rect 3788 2316 3796 2324
rect 3852 2316 3860 2324
rect 3900 2316 3908 2324
rect 4604 2312 4612 2320
rect 5084 2312 5092 2320
rect 5548 2316 5556 2324
rect 3644 2296 3652 2304
rect 3676 2296 3684 2304
rect 3772 2296 3780 2304
rect 3836 2296 3844 2304
rect 3900 2296 3908 2304
rect 4108 2296 4116 2304
rect 4236 2296 4244 2304
rect 4284 2296 4292 2304
rect 4316 2296 4324 2304
rect 4572 2296 4580 2304
rect 4780 2296 4788 2304
rect 4892 2296 4900 2304
rect 4908 2296 4916 2304
rect 5068 2296 5076 2304
rect 5420 2296 5428 2304
rect 5532 2296 5540 2304
rect 5564 2296 5572 2304
rect 5580 2296 5588 2304
rect 5660 2316 5668 2324
rect 6060 2316 6068 2324
rect 6332 2316 6340 2324
rect 5724 2296 5732 2304
rect 5852 2296 5860 2304
rect 6076 2296 6084 2304
rect 6188 2296 6196 2304
rect 6236 2294 6244 2302
rect 6332 2296 6340 2304
rect 6748 2296 6756 2304
rect 140 2276 148 2284
rect 428 2276 436 2284
rect 572 2276 580 2284
rect 748 2276 756 2284
rect 1004 2276 1012 2284
rect 188 2256 196 2264
rect 236 2256 244 2264
rect 396 2256 404 2264
rect 668 2256 676 2264
rect 1036 2256 1044 2264
rect 1308 2256 1316 2264
rect 1356 2276 1364 2284
rect 1596 2276 1604 2284
rect 2076 2276 2084 2284
rect 2364 2276 2372 2284
rect 2508 2276 2516 2284
rect 2812 2276 2820 2284
rect 2876 2276 2884 2284
rect 2908 2276 2916 2284
rect 3004 2276 3012 2284
rect 3116 2276 3124 2284
rect 3308 2276 3316 2284
rect 3532 2276 3540 2284
rect 3564 2276 3572 2284
rect 3660 2276 3668 2284
rect 3724 2276 3732 2284
rect 3996 2276 4004 2284
rect 4396 2276 4404 2284
rect 4668 2276 4676 2284
rect 5148 2276 5156 2284
rect 5404 2276 5412 2284
rect 5596 2276 5604 2284
rect 5612 2276 5620 2284
rect 5692 2276 5700 2284
rect 5964 2276 5972 2284
rect 6268 2276 6276 2284
rect 6428 2276 6436 2284
rect 6748 2276 6756 2284
rect 1564 2256 1572 2264
rect 1740 2256 1748 2264
rect 2044 2256 2052 2264
rect 2540 2256 2548 2264
rect 2828 2256 2836 2264
rect 2860 2256 2868 2264
rect 3020 2256 3028 2264
rect 3340 2256 3348 2264
rect 3516 2256 3524 2264
rect 4028 2256 4036 2264
rect 4252 2256 4260 2264
rect 4364 2256 4372 2264
rect 4700 2256 4708 2264
rect 4924 2256 4932 2264
rect 5004 2256 5012 2264
rect 5180 2256 5188 2264
rect 5340 2256 5348 2264
rect 5388 2256 5396 2264
rect 5468 2256 5476 2264
rect 5932 2256 5940 2264
rect 6460 2256 6468 2264
rect 6636 2256 6644 2264
rect 28 2236 36 2244
rect 732 2236 740 2244
rect 1340 2236 1348 2244
rect 1804 2236 1812 2244
rect 1884 2236 1892 2244
rect 2732 2236 2740 2244
rect 2940 2236 2948 2244
rect 2956 2236 2964 2244
rect 3100 2236 3108 2244
rect 3436 2236 3444 2244
rect 3596 2236 3604 2244
rect 4508 2236 4516 2244
rect 4860 2236 4868 2244
rect 5372 2236 5380 2244
rect 5452 2236 5460 2244
rect 5484 2236 5492 2244
rect 5628 2236 5636 2244
rect 6620 2236 6628 2244
rect 6860 2236 6868 2244
rect 2638 2206 2646 2214
rect 2652 2206 2660 2214
rect 2666 2206 2674 2214
rect 5726 2206 5734 2214
rect 5740 2206 5748 2214
rect 5754 2206 5762 2214
rect 2812 2196 2820 2204
rect 620 2176 628 2184
rect 1196 2176 1204 2184
rect 1548 2176 1556 2184
rect 2364 2176 2372 2184
rect 3020 2176 3028 2184
rect 3132 2176 3140 2184
rect 3180 2176 3188 2184
rect 3196 2176 3204 2184
rect 3244 2176 3252 2184
rect 3500 2176 3508 2184
rect 5276 2176 5284 2184
rect 5292 2176 5300 2184
rect 5868 2176 5876 2184
rect 6492 2176 6500 2184
rect 6684 2176 6692 2184
rect 12 2156 20 2164
rect 268 2156 276 2164
rect 780 2156 788 2164
rect 1356 2156 1364 2164
rect 1708 2156 1716 2164
rect 2044 2156 2052 2164
rect 2396 2156 2404 2164
rect 2588 2156 2596 2164
rect 2812 2156 2820 2164
rect 3340 2156 3348 2164
rect 3724 2156 3732 2164
rect 4236 2156 4244 2164
rect 4668 2156 4676 2164
rect 4844 2156 4852 2164
rect 5036 2156 5044 2164
rect 5404 2156 5412 2164
rect 5484 2156 5492 2164
rect 5564 2156 5572 2164
rect 5788 2156 5796 2164
rect 6284 2156 6292 2164
rect 92 2136 100 2144
rect 236 2136 244 2144
rect 588 2136 596 2144
rect 812 2136 820 2144
rect 956 2136 964 2144
rect 1084 2136 1092 2144
rect 1388 2136 1396 2144
rect 1740 2136 1748 2144
rect 2012 2136 2020 2144
rect 2268 2136 2276 2144
rect 2316 2136 2324 2144
rect 2348 2136 2356 2144
rect 2380 2136 2388 2144
rect 2444 2136 2452 2144
rect 2780 2136 2788 2144
rect 2988 2136 2996 2144
rect 3052 2136 3060 2144
rect 60 2116 68 2124
rect 236 2116 244 2124
rect 700 2116 708 2124
rect 908 2116 916 2124
rect 1484 2116 1492 2124
rect 1836 2116 1844 2124
rect 1900 2116 1908 2124
rect 2124 2116 2132 2124
rect 2268 2116 2276 2124
rect 2332 2116 2340 2124
rect 2428 2116 2436 2124
rect 2492 2116 2500 2124
rect 2556 2116 2564 2124
rect 2700 2116 2708 2124
rect 2988 2116 2996 2124
rect 3036 2116 3044 2124
rect 3100 2116 3108 2124
rect 3196 2136 3204 2144
rect 3324 2136 3332 2144
rect 3372 2136 3380 2144
rect 3420 2136 3428 2144
rect 3436 2136 3444 2144
rect 3532 2136 3540 2144
rect 3756 2136 3764 2144
rect 3916 2136 3924 2144
rect 3964 2136 3972 2144
rect 4204 2136 4212 2144
rect 4700 2136 4708 2144
rect 5004 2136 5012 2144
rect 5228 2136 5236 2144
rect 5388 2136 5396 2144
rect 5436 2136 5444 2144
rect 5484 2136 5492 2144
rect 5772 2136 5780 2144
rect 5804 2136 5812 2144
rect 5900 2136 5908 2144
rect 5996 2136 6004 2144
rect 6108 2136 6116 2144
rect 6316 2136 6324 2144
rect 6460 2136 6468 2144
rect 6556 2136 6564 2144
rect 3212 2116 3220 2124
rect 3308 2116 3316 2124
rect 3372 2116 3380 2124
rect 3452 2116 3460 2124
rect 3852 2116 3860 2124
rect 3964 2116 3972 2124
rect 3980 2116 3988 2124
rect 4060 2116 4068 2124
rect 4108 2116 4116 2124
rect 4428 2116 4436 2124
rect 4506 2116 4514 2124
rect 4700 2116 4708 2124
rect 4892 2116 4900 2124
rect 5004 2116 5012 2124
rect 5116 2116 5124 2124
rect 5244 2116 5252 2124
rect 5372 2116 5380 2124
rect 5452 2116 5460 2124
rect 5516 2116 5524 2124
rect 5548 2116 5556 2124
rect 5612 2116 5620 2124
rect 5660 2116 5668 2124
rect 5692 2116 5700 2124
rect 5900 2116 5908 2124
rect 5932 2116 5940 2124
rect 5980 2116 5988 2124
rect 6012 2116 6020 2124
rect 6028 2116 6036 2124
rect 6076 2116 6084 2124
rect 6122 2116 6130 2124
rect 6204 2116 6212 2124
rect 6428 2116 6436 2124
rect 6556 2116 6564 2124
rect 6716 2136 6724 2144
rect 92 2096 100 2104
rect 140 2096 148 2104
rect 908 2096 916 2104
rect 1452 2100 1460 2108
rect 1836 2096 1844 2104
rect 1916 2096 1924 2104
rect 2380 2096 2388 2104
rect 2572 2096 2580 2104
rect 2684 2096 2692 2104
rect 3036 2096 3044 2104
rect 3068 2096 3076 2104
rect 3276 2096 3284 2104
rect 3340 2096 3348 2104
rect 3388 2096 3396 2104
rect 3484 2096 3492 2104
rect 3500 2096 3508 2104
rect 3820 2100 3828 2108
rect 4012 2096 4020 2104
rect 4140 2100 4148 2108
rect 4796 2096 4804 2104
rect 4940 2100 4948 2108
rect 5276 2096 5284 2104
rect 5292 2096 5300 2104
rect 5340 2096 5348 2104
rect 5548 2096 5556 2104
rect 5676 2096 5684 2104
rect 6412 2096 6420 2104
rect 1180 2076 1188 2084
rect 5516 2076 5524 2084
rect 5644 2076 5652 2084
rect 1452 2054 1460 2062
rect 3820 2054 3828 2062
rect 4140 2054 4148 2062
rect 4700 2056 4708 2064
rect 4940 2054 4948 2062
rect 140 2036 148 2044
rect 428 2036 436 2044
rect 476 2036 484 2044
rect 620 2036 628 2044
rect 908 2036 916 2044
rect 1068 2036 1076 2044
rect 1836 2036 1844 2044
rect 1916 2036 1924 2044
rect 2204 2036 2212 2044
rect 2524 2036 2532 2044
rect 2684 2036 2692 2044
rect 3244 2036 3252 2044
rect 3308 2036 3316 2044
rect 3452 2036 3460 2044
rect 4396 2036 4404 2044
rect 4460 2036 4468 2044
rect 4860 2036 4868 2044
rect 5196 2036 5204 2044
rect 6412 2036 6420 2044
rect 6828 2036 6836 2044
rect 1118 2006 1126 2014
rect 1132 2006 1140 2014
rect 1146 2006 1154 2014
rect 4158 2006 4166 2014
rect 4172 2006 4180 2014
rect 4186 2006 4194 2014
rect 140 1976 148 1984
rect 204 1976 212 1984
rect 2124 1976 2132 1984
rect 2588 1976 2596 1984
rect 2988 1976 2996 1984
rect 3036 1976 3044 1984
rect 3100 1976 3108 1984
rect 3964 1976 3972 1984
rect 4028 1976 4036 1984
rect 4284 1976 4292 1984
rect 5068 1976 5076 1984
rect 5260 1976 5268 1984
rect 492 1956 500 1964
rect 3708 1956 3716 1964
rect 4540 1958 4548 1966
rect 684 1936 692 1944
rect 1052 1936 1060 1944
rect 3980 1936 3988 1944
rect 4044 1936 4052 1944
rect 5788 1936 5796 1944
rect 6396 1936 6404 1944
rect 92 1916 100 1924
rect 108 1916 116 1924
rect 204 1916 212 1924
rect 716 1916 724 1924
rect 732 1916 740 1924
rect 796 1916 804 1924
rect 1404 1916 1412 1924
rect 2124 1916 2132 1924
rect 2588 1916 2596 1924
rect 2988 1916 2996 1924
rect 3100 1916 3108 1924
rect 3404 1916 3412 1924
rect 3468 1916 3476 1924
rect 3756 1916 3764 1924
rect 3804 1916 3812 1924
rect 3900 1916 3908 1924
rect 3932 1916 3940 1924
rect 4012 1916 4020 1924
rect 4540 1912 4548 1920
rect 4620 1916 4628 1924
rect 60 1896 68 1904
rect 140 1896 148 1904
rect 236 1896 244 1904
rect 508 1896 516 1904
rect 556 1896 564 1904
rect 700 1896 708 1904
rect 764 1896 772 1904
rect 828 1896 836 1904
rect 908 1894 916 1902
rect 1180 1896 1188 1904
rect 1308 1896 1316 1904
rect 1532 1896 1540 1904
rect 1692 1896 1700 1904
rect 2108 1896 2116 1904
rect 2172 1896 2180 1904
rect 2268 1896 2276 1904
rect 2380 1896 2388 1904
rect 2556 1896 2564 1904
rect 2780 1896 2788 1904
rect 3004 1896 3012 1904
rect 3100 1896 3108 1904
rect 3404 1896 3412 1904
rect 3836 1896 3844 1904
rect 3964 1896 3972 1904
rect 4028 1896 4036 1904
rect 4572 1896 4580 1904
rect 4652 1896 4660 1904
rect 4828 1896 4836 1904
rect 4844 1896 4852 1904
rect 4876 1896 4884 1904
rect 5100 1896 5108 1904
rect 5260 1896 5268 1904
rect 5452 1896 5460 1904
rect 5596 1896 5604 1904
rect 5612 1896 5620 1904
rect 5644 1916 5652 1924
rect 5676 1896 5684 1904
rect 5756 1896 5764 1904
rect 5772 1896 5780 1904
rect 5820 1896 5828 1904
rect 5868 1896 5876 1904
rect 5884 1896 5892 1904
rect 5916 1916 5924 1924
rect 6220 1916 6228 1924
rect 6284 1916 6292 1924
rect 6716 1916 6724 1924
rect 5948 1896 5956 1904
rect 6092 1896 6100 1904
rect 6188 1896 6196 1904
rect 6204 1896 6212 1904
rect 6252 1896 6260 1904
rect 6300 1896 6308 1904
rect 6316 1896 6324 1904
rect 6364 1896 6372 1904
rect 6380 1896 6388 1904
rect 6508 1896 6516 1904
rect 6620 1896 6628 1904
rect 6668 1896 6676 1904
rect 6716 1896 6724 1904
rect 6764 1896 6772 1904
rect 156 1876 164 1884
rect 300 1876 308 1884
rect 604 1876 612 1884
rect 652 1876 660 1884
rect 780 1876 788 1884
rect 844 1876 852 1884
rect 876 1876 884 1884
rect 924 1876 932 1884
rect 1084 1876 1092 1884
rect 1196 1876 1204 1884
rect 1228 1876 1236 1884
rect 1500 1876 1508 1884
rect 1644 1876 1652 1884
rect 2028 1876 2036 1884
rect 12 1856 20 1864
rect 92 1856 100 1864
rect 332 1856 340 1864
rect 588 1856 596 1864
rect 700 1856 708 1864
rect 1420 1856 1428 1864
rect 1996 1856 2004 1864
rect 2204 1856 2212 1864
rect 2252 1876 2260 1884
rect 2298 1876 2306 1884
rect 2492 1876 2500 1884
rect 2892 1876 2900 1884
rect 3196 1876 3204 1884
rect 3390 1876 3398 1884
rect 3500 1876 3508 1884
rect 3676 1876 3684 1884
rect 3692 1876 3700 1884
rect 3724 1876 3732 1884
rect 3820 1876 3828 1884
rect 3884 1876 3892 1884
rect 3932 1876 3940 1884
rect 4204 1876 4212 1884
rect 4476 1876 4484 1884
rect 4668 1876 4676 1884
rect 4812 1876 4820 1884
rect 4956 1876 4964 1884
rect 5180 1876 5188 1884
rect 5372 1876 5380 1884
rect 5404 1876 5412 1884
rect 5580 1876 5588 1884
rect 5692 1876 5700 1884
rect 5852 1876 5860 1884
rect 5964 1876 5972 1884
rect 6076 1876 6084 1884
rect 6172 1876 6180 1884
rect 6236 1876 6244 1884
rect 6300 1876 6308 1884
rect 6524 1876 6532 1884
rect 6764 1876 6772 1884
rect 6780 1876 6788 1884
rect 6876 1876 6884 1884
rect 2236 1856 2244 1864
rect 2460 1856 2468 1864
rect 2860 1856 2868 1864
rect 3052 1856 3060 1864
rect 3228 1856 3236 1864
rect 3564 1856 3572 1864
rect 4444 1856 4452 1864
rect 4700 1856 4708 1864
rect 4940 1856 4948 1864
rect 5164 1856 5172 1864
rect 5228 1856 5236 1864
rect 6588 1856 6596 1864
rect 6604 1856 6612 1864
rect 6620 1856 6628 1864
rect 6668 1856 6676 1864
rect 6700 1856 6708 1864
rect 636 1836 644 1844
rect 732 1836 740 1844
rect 796 1836 804 1844
rect 1036 1836 1044 1844
rect 1148 1836 1156 1844
rect 1388 1836 1396 1844
rect 1612 1836 1620 1844
rect 1804 1836 1812 1844
rect 1836 1836 1844 1844
rect 2700 1836 2708 1844
rect 3532 1836 3540 1844
rect 3804 1836 3812 1844
rect 3836 1836 3844 1844
rect 4092 1836 4100 1844
rect 4620 1836 4628 1844
rect 5068 1836 5076 1844
rect 5132 1836 5140 1844
rect 5212 1836 5220 1844
rect 5308 1836 5316 1844
rect 5564 1836 5572 1844
rect 5980 1836 5988 1844
rect 6716 1836 6724 1844
rect 6812 1836 6820 1844
rect 2638 1806 2646 1814
rect 2652 1806 2660 1814
rect 2666 1806 2674 1814
rect 5726 1806 5734 1814
rect 5740 1806 5748 1814
rect 5754 1806 5762 1814
rect 572 1776 580 1784
rect 1308 1776 1316 1784
rect 1884 1776 1892 1784
rect 2124 1776 2132 1784
rect 2172 1776 2180 1784
rect 2620 1776 2628 1784
rect 3612 1776 3620 1784
rect 4076 1776 4084 1784
rect 4172 1776 4180 1784
rect 4524 1776 4532 1784
rect 4588 1776 4596 1784
rect 5500 1776 5508 1784
rect 5772 1776 5780 1784
rect 5916 1776 5924 1784
rect 6364 1776 6372 1784
rect 6508 1776 6516 1784
rect 6556 1776 6564 1784
rect 172 1756 180 1764
rect 412 1756 420 1764
rect 748 1756 756 1764
rect 924 1756 932 1764
rect 1180 1756 1188 1764
rect 1404 1756 1412 1764
rect 1500 1756 1508 1764
rect 1660 1756 1668 1764
rect 1980 1756 1988 1764
rect 2060 1756 2068 1764
rect 2188 1756 2196 1764
rect 2380 1756 2388 1764
rect 2588 1756 2596 1764
rect 140 1736 148 1744
rect 588 1736 596 1744
rect 604 1736 612 1744
rect 684 1736 692 1744
rect 892 1736 900 1744
rect 1228 1736 1236 1744
rect 1356 1736 1364 1744
rect 140 1716 148 1724
rect 252 1716 260 1724
rect 412 1718 420 1726
rect 1580 1736 1588 1744
rect 1628 1736 1636 1744
rect 620 1716 628 1724
rect 44 1696 52 1704
rect 652 1696 660 1704
rect 700 1716 708 1724
rect 796 1716 804 1724
rect 1244 1716 1252 1724
rect 1340 1716 1348 1724
rect 1372 1716 1380 1724
rect 1388 1716 1396 1724
rect 1436 1716 1444 1724
rect 1468 1716 1476 1724
rect 1548 1716 1556 1724
rect 1564 1716 1572 1724
rect 1676 1716 1684 1724
rect 1692 1716 1700 1724
rect 1740 1716 1748 1724
rect 1772 1736 1780 1744
rect 1836 1736 1844 1744
rect 1948 1736 1956 1744
rect 2044 1736 2052 1744
rect 2140 1736 2148 1744
rect 2412 1736 2420 1744
rect 2876 1756 2884 1764
rect 3148 1756 3156 1764
rect 3404 1756 3412 1764
rect 3772 1756 3780 1764
rect 4332 1756 4340 1764
rect 4556 1756 4564 1764
rect 4844 1756 4852 1764
rect 4940 1756 4948 1764
rect 4956 1756 4964 1764
rect 5212 1756 5220 1764
rect 5420 1756 5428 1764
rect 5548 1756 5556 1764
rect 6124 1756 6132 1764
rect 6300 1756 6308 1764
rect 6412 1756 6420 1764
rect 6716 1756 6724 1764
rect 2636 1736 2644 1744
rect 2844 1736 2852 1744
rect 3132 1736 3140 1744
rect 3164 1736 3172 1744
rect 3180 1736 3188 1744
rect 3372 1736 3380 1744
rect 3804 1736 3812 1744
rect 4364 1736 4372 1744
rect 4508 1736 4516 1744
rect 4620 1736 4628 1744
rect 5004 1736 5012 1744
rect 5180 1736 5188 1744
rect 5548 1736 5556 1744
rect 5612 1736 5620 1744
rect 5628 1736 5636 1744
rect 6076 1736 6084 1744
rect 6140 1736 6148 1744
rect 6252 1736 6260 1744
rect 6748 1736 6756 1744
rect 1852 1716 1860 1724
rect 796 1696 804 1704
rect 1084 1696 1092 1704
rect 1180 1696 1188 1704
rect 1308 1696 1316 1704
rect 1484 1696 1492 1704
rect 1516 1696 1524 1704
rect 1788 1696 1796 1704
rect 1820 1696 1828 1704
rect 1948 1716 1956 1724
rect 2060 1716 2068 1724
rect 2092 1716 2100 1724
rect 2156 1716 2164 1724
rect 2300 1716 2308 1724
rect 2508 1716 2516 1724
rect 2556 1716 2564 1724
rect 2652 1716 2660 1724
rect 2748 1716 2756 1724
rect 2956 1716 2964 1724
rect 3052 1716 3060 1724
rect 3196 1716 3204 1724
rect 3212 1716 3220 1724
rect 3292 1716 3300 1724
rect 3804 1716 3812 1724
rect 3948 1716 3956 1724
rect 3964 1716 3972 1724
rect 4012 1716 4020 1724
rect 4044 1716 4052 1724
rect 4252 1716 4260 1724
rect 4476 1716 4484 1724
rect 4636 1716 4644 1724
rect 4652 1716 4660 1724
rect 4716 1716 4724 1724
rect 4732 1716 4740 1724
rect 4748 1716 4756 1724
rect 4892 1716 4900 1724
rect 5036 1716 5044 1724
rect 5084 1716 5092 1724
rect 5452 1716 5460 1724
rect 5468 1716 5476 1724
rect 5596 1716 5604 1724
rect 5660 1716 5668 1724
rect 5708 1716 5716 1724
rect 5740 1716 5748 1724
rect 5788 1716 5796 1724
rect 5804 1716 5812 1724
rect 5820 1716 5828 1724
rect 5852 1716 5860 1724
rect 6044 1718 6052 1726
rect 6156 1716 6164 1724
rect 1900 1696 1908 1704
rect 1980 1696 1988 1704
rect 2508 1696 2516 1704
rect 2780 1700 2788 1708
rect 3132 1696 3140 1704
rect 3228 1696 3236 1704
rect 3276 1696 3284 1704
rect 3564 1696 3572 1704
rect 3868 1700 3876 1708
rect 4428 1700 4436 1708
rect 4540 1696 4548 1704
rect 4588 1696 4596 1704
rect 4844 1696 4852 1704
rect 5084 1696 5092 1704
rect 5564 1696 5572 1704
rect 5660 1696 5668 1704
rect 5820 1696 5828 1704
rect 6188 1696 6196 1704
rect 6236 1716 6244 1724
rect 6268 1716 6276 1724
rect 6284 1716 6292 1724
rect 6332 1716 6340 1724
rect 6396 1716 6404 1724
rect 6460 1716 6468 1724
rect 6748 1716 6756 1724
rect 6364 1696 6372 1704
rect 6812 1700 6820 1708
rect 332 1676 340 1684
rect 556 1676 564 1684
rect 1212 1676 1220 1684
rect 1548 1676 1556 1684
rect 2028 1676 2036 1684
rect 2204 1676 2212 1684
rect 6236 1676 6244 1684
rect 6396 1676 6404 1684
rect 1116 1656 1124 1664
rect 2780 1654 2788 1662
rect 6812 1654 6820 1662
rect 44 1636 52 1644
rect 540 1636 548 1644
rect 796 1636 804 1644
rect 1276 1636 1284 1644
rect 1964 1636 1972 1644
rect 2508 1636 2516 1644
rect 3036 1636 3044 1644
rect 3276 1636 3284 1644
rect 3868 1636 3876 1644
rect 3980 1636 3988 1644
rect 4428 1636 4436 1644
rect 4572 1636 4580 1644
rect 4668 1636 4676 1644
rect 4764 1636 4772 1644
rect 4892 1636 4900 1644
rect 4972 1636 4980 1644
rect 5084 1636 5092 1644
rect 5372 1636 5380 1644
rect 5420 1636 5428 1644
rect 5532 1636 5540 1644
rect 5644 1636 5652 1644
rect 6108 1636 6116 1644
rect 6444 1636 6452 1644
rect 6460 1636 6468 1644
rect 1118 1606 1126 1614
rect 1132 1606 1140 1614
rect 1146 1606 1154 1614
rect 4158 1606 4166 1614
rect 4172 1606 4180 1614
rect 4186 1606 4194 1614
rect 60 1576 68 1584
rect 396 1576 404 1584
rect 908 1576 916 1584
rect 1372 1576 1380 1584
rect 1884 1576 1892 1584
rect 2412 1576 2420 1584
rect 3164 1576 3172 1584
rect 3788 1576 3796 1584
rect 4220 1576 4228 1584
rect 4732 1576 4740 1584
rect 4796 1576 4804 1584
rect 5084 1576 5092 1584
rect 5180 1576 5188 1584
rect 5404 1576 5412 1584
rect 5580 1576 5588 1584
rect 6172 1576 6180 1584
rect 6316 1576 6324 1584
rect 6380 1576 6388 1584
rect 2956 1558 2964 1566
rect 3900 1558 3908 1566
rect 4444 1558 4452 1566
rect 6412 1556 6420 1564
rect 940 1536 948 1544
rect 1820 1536 1828 1544
rect 2172 1536 2180 1544
rect 3052 1536 3060 1544
rect 3116 1536 3124 1544
rect 3452 1536 3460 1544
rect 3484 1536 3492 1544
rect 6220 1536 6228 1544
rect 6236 1536 6244 1544
rect 6700 1536 6708 1544
rect 60 1496 68 1504
rect 108 1516 116 1524
rect 348 1516 356 1524
rect 140 1496 148 1504
rect 220 1496 228 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 396 1496 404 1504
rect 412 1496 420 1504
rect 492 1496 500 1504
rect 508 1496 516 1504
rect 524 1496 532 1504
rect 556 1496 564 1504
rect 588 1496 596 1504
rect 604 1496 612 1504
rect 636 1496 644 1504
rect 684 1516 692 1524
rect 860 1516 868 1524
rect 716 1496 724 1504
rect 796 1496 804 1504
rect 828 1496 836 1504
rect 1324 1516 1332 1524
rect 908 1496 916 1504
rect 1052 1496 1060 1504
rect 1180 1496 1188 1504
rect 1196 1496 1204 1504
rect 1244 1496 1252 1504
rect 1276 1496 1284 1504
rect 1308 1496 1316 1504
rect 1340 1496 1348 1504
rect 1404 1496 1412 1504
rect 1420 1496 1428 1504
rect 1484 1496 1492 1504
rect 1516 1496 1524 1504
rect 1564 1516 1572 1524
rect 2092 1516 2100 1524
rect 1596 1496 1604 1504
rect 1676 1494 1684 1502
rect 1852 1496 1860 1504
rect 1868 1496 1876 1504
rect 1916 1496 1924 1504
rect 1948 1496 1956 1504
rect 1964 1496 1972 1504
rect 2012 1496 2020 1504
rect 2060 1496 2068 1504
rect 2748 1516 2756 1524
rect 3164 1516 3172 1524
rect 3788 1516 3796 1524
rect 3900 1512 3908 1520
rect 4316 1516 4324 1524
rect 4364 1516 4372 1524
rect 4444 1512 4452 1520
rect 4796 1516 4804 1524
rect 5148 1516 5156 1524
rect 2124 1496 2132 1504
rect 2140 1496 2148 1504
rect 2284 1496 2292 1504
rect 2364 1496 2372 1504
rect 2380 1496 2388 1504
rect 2428 1496 2436 1504
rect 2460 1496 2468 1504
rect 2476 1496 2484 1504
rect 2524 1496 2532 1504
rect 188 1476 196 1484
rect 300 1476 308 1484
rect 412 1476 420 1484
rect 428 1476 436 1484
rect 620 1476 628 1484
rect 668 1476 676 1484
rect 732 1476 740 1484
rect 748 1476 756 1484
rect 812 1476 820 1484
rect 924 1476 932 1484
rect 1068 1476 1076 1484
rect 1276 1476 1284 1484
rect 1388 1476 1396 1484
rect 1468 1476 1476 1484
rect 1500 1476 1508 1484
rect 1548 1476 1556 1484
rect 1612 1476 1620 1484
rect 1644 1476 1652 1484
rect 2028 1476 2036 1484
rect 2044 1476 2052 1484
rect 2156 1476 2164 1484
rect 2332 1476 2340 1484
rect 2604 1496 2612 1504
rect 2956 1496 2964 1504
rect 3068 1496 3076 1504
rect 3372 1496 3380 1504
rect 3580 1496 3588 1504
rect 3804 1496 3812 1504
rect 3868 1496 3876 1504
rect 4076 1496 4084 1504
rect 4284 1496 4292 1504
rect 4412 1496 4420 1504
rect 4620 1496 4628 1504
rect 4796 1496 4804 1504
rect 5148 1496 5156 1504
rect 5180 1496 5188 1504
rect 5228 1496 5236 1504
rect 5276 1516 5284 1524
rect 5468 1516 5476 1524
rect 5308 1496 5316 1504
rect 5388 1496 5396 1504
rect 5420 1496 5428 1504
rect 5628 1516 5636 1524
rect 5740 1516 5748 1524
rect 5852 1516 5860 1524
rect 5612 1496 5620 1504
rect 5628 1496 5636 1504
rect 5772 1496 5780 1504
rect 5820 1496 5828 1504
rect 6140 1516 6148 1524
rect 6268 1516 6276 1524
rect 6684 1516 6692 1524
rect 5900 1496 5908 1504
rect 5932 1496 5940 1504
rect 5948 1496 5956 1504
rect 5996 1496 6004 1504
rect 6012 1496 6020 1504
rect 6108 1496 6116 1504
rect 6204 1496 6212 1504
rect 6252 1496 6260 1504
rect 6284 1496 6292 1504
rect 6348 1496 6356 1504
rect 6444 1496 6452 1504
rect 6460 1496 6468 1504
rect 6508 1496 6516 1504
rect 6540 1496 6548 1504
rect 6556 1496 6564 1504
rect 6604 1496 6612 1504
rect 2652 1476 2660 1484
rect 2844 1476 2852 1484
rect 3038 1476 3046 1484
rect 3052 1476 3060 1484
rect 3260 1476 3268 1484
rect 3692 1476 3700 1484
rect 3964 1476 3972 1484
rect 4268 1476 4276 1484
rect 4508 1476 4516 1484
rect 4892 1476 4900 1484
rect 5196 1476 5204 1484
rect 5212 1476 5220 1484
rect 5324 1476 5332 1484
rect 5420 1476 5428 1484
rect 5500 1476 5508 1484
rect 5564 1476 5572 1484
rect 5676 1476 5684 1484
rect 5788 1476 5796 1484
rect 5804 1476 5812 1484
rect 5916 1476 5924 1484
rect 6092 1476 6100 1484
rect 6524 1476 6532 1484
rect 6684 1496 6692 1504
rect 6780 1496 6788 1504
rect 6796 1496 6804 1504
rect 6636 1476 6644 1484
rect 28 1456 36 1464
rect 1004 1456 1012 1464
rect 1212 1456 1220 1464
rect 1820 1456 1828 1464
rect 2492 1456 2500 1464
rect 2876 1456 2884 1464
rect 3292 1456 3300 1464
rect 3468 1456 3476 1464
rect 3660 1456 3668 1464
rect 3996 1456 4004 1464
rect 4156 1456 4164 1464
rect 4252 1456 4260 1464
rect 4540 1456 4548 1464
rect 4700 1456 4708 1464
rect 4748 1456 4756 1464
rect 4924 1456 4932 1464
rect 5100 1456 5108 1464
rect 5340 1456 5348 1464
rect 5388 1456 5396 1464
rect 5484 1456 5492 1464
rect 6428 1456 6436 1464
rect 6828 1456 6836 1464
rect 252 1436 260 1444
rect 1836 1436 1844 1444
rect 3116 1436 3124 1444
rect 4348 1436 4356 1444
rect 5260 1436 5268 1444
rect 5356 1436 5364 1444
rect 5468 1436 5476 1444
rect 5516 1436 5524 1444
rect 5868 1436 5876 1444
rect 5964 1436 5972 1444
rect 6060 1436 6068 1444
rect 6140 1436 6148 1444
rect 6172 1436 6180 1444
rect 6316 1436 6324 1444
rect 6380 1436 6388 1444
rect 2638 1406 2646 1414
rect 2652 1406 2660 1414
rect 2666 1406 2674 1414
rect 5726 1406 5734 1414
rect 5740 1406 5748 1414
rect 5754 1406 5762 1414
rect 268 1376 276 1384
rect 508 1376 516 1384
rect 1596 1376 1604 1384
rect 1676 1376 1684 1384
rect 2428 1376 2436 1384
rect 2684 1376 2692 1384
rect 2796 1376 2804 1384
rect 3036 1376 3044 1384
rect 3948 1376 3956 1384
rect 4732 1376 4740 1384
rect 5084 1376 5092 1384
rect 5116 1376 5124 1384
rect 5836 1376 5844 1384
rect 5852 1376 5860 1384
rect 5964 1376 5972 1384
rect 6252 1376 6260 1384
rect 6700 1376 6708 1384
rect 380 1356 388 1364
rect 876 1356 884 1364
rect 1308 1356 1316 1364
rect 1388 1356 1396 1364
rect 1628 1356 1636 1364
rect 2188 1356 2196 1364
rect 2492 1356 2500 1364
rect 2524 1356 2532 1364
rect 2748 1356 2756 1364
rect 3244 1356 3252 1364
rect 3452 1356 3460 1364
rect 3468 1356 3476 1364
rect 3676 1356 3684 1364
rect 4108 1356 4116 1364
rect 4380 1356 4388 1364
rect 4572 1356 4580 1364
rect 4924 1356 4932 1364
rect 5404 1356 5412 1364
rect 5564 1356 5572 1364
rect 6460 1356 6468 1364
rect 6828 1356 6836 1364
rect 252 1336 260 1344
rect 316 1336 324 1344
rect 524 1336 532 1344
rect 588 1336 596 1344
rect 636 1336 644 1344
rect 76 1316 84 1324
rect 124 1316 132 1324
rect 268 1316 276 1324
rect 300 1316 308 1324
rect 396 1316 404 1324
rect 540 1316 548 1324
rect 748 1336 756 1344
rect 860 1336 868 1344
rect 908 1336 916 1344
rect 1084 1336 1092 1344
rect 1116 1336 1124 1344
rect 1180 1336 1188 1344
rect 1532 1336 1540 1344
rect 1548 1336 1556 1344
rect 1612 1336 1620 1344
rect 1724 1336 1732 1344
rect 1788 1336 1796 1344
rect 1836 1336 1844 1344
rect 1868 1336 1876 1344
rect 1932 1336 1940 1344
rect 1948 1336 1956 1344
rect 2220 1336 2228 1344
rect 2460 1336 2468 1344
rect 2652 1336 2660 1344
rect 2892 1336 2900 1344
rect 2940 1336 2948 1344
rect 2956 1336 2964 1344
rect 3052 1336 3060 1344
rect 3276 1336 3284 1344
rect 3644 1336 3652 1344
rect 4140 1336 4148 1344
rect 4540 1336 4548 1344
rect 4892 1336 4900 1344
rect 5164 1336 5172 1344
rect 5340 1336 5348 1344
rect 5436 1336 5444 1344
rect 5548 1336 5556 1344
rect 5884 1336 5892 1344
rect 6012 1336 6020 1344
rect 236 1296 244 1304
rect 268 1296 276 1304
rect 572 1296 580 1304
rect 668 1316 676 1324
rect 716 1316 724 1324
rect 732 1316 740 1324
rect 748 1316 756 1324
rect 844 1316 852 1324
rect 924 1316 932 1324
rect 972 1316 980 1324
rect 988 1316 996 1324
rect 1020 1316 1028 1324
rect 1100 1316 1108 1324
rect 812 1296 820 1304
rect 1004 1296 1012 1304
rect 1212 1296 1220 1304
rect 1260 1316 1268 1324
rect 1340 1316 1348 1324
rect 1436 1316 1444 1324
rect 1484 1316 1492 1324
rect 1500 1316 1508 1324
rect 1516 1316 1524 1324
rect 1564 1316 1572 1324
rect 1628 1316 1636 1324
rect 1740 1316 1748 1324
rect 1804 1316 1812 1324
rect 1916 1316 1924 1324
rect 1932 1316 1940 1324
rect 2300 1316 2308 1324
rect 2396 1316 2404 1324
rect 2492 1316 2500 1324
rect 2556 1316 2564 1324
rect 2716 1316 2724 1324
rect 2796 1316 2804 1324
rect 2876 1316 2884 1324
rect 2956 1316 2964 1324
rect 3372 1316 3380 1324
rect 3420 1316 3428 1324
rect 3500 1316 3508 1324
rect 3756 1316 3764 1324
rect 3916 1316 3924 1324
rect 4028 1316 4036 1324
rect 4236 1316 4244 1324
rect 4364 1316 4372 1324
rect 4444 1316 4452 1324
rect 5004 1316 5012 1324
rect 5148 1316 5156 1324
rect 5308 1318 5316 1326
rect 5372 1316 5380 1324
rect 5452 1316 5460 1324
rect 5468 1316 5476 1324
rect 1324 1296 1332 1304
rect 1468 1296 1476 1304
rect 1484 1296 1492 1304
rect 1596 1296 1604 1304
rect 1756 1296 1764 1304
rect 1772 1296 1780 1304
rect 1836 1296 1844 1304
rect 1916 1296 1924 1304
rect 1996 1296 2004 1304
rect 2284 1300 2292 1308
rect 2412 1296 2420 1304
rect 2796 1296 2804 1304
rect 2844 1296 2852 1304
rect 2908 1296 2916 1304
rect 2972 1296 2980 1304
rect 3004 1296 3012 1304
rect 3020 1296 3028 1304
rect 3084 1296 3092 1304
rect 3340 1300 3348 1308
rect 3580 1300 3588 1308
rect 4204 1300 4212 1308
rect 4476 1300 4484 1308
rect 4796 1296 4804 1304
rect 5100 1296 5108 1304
rect 5532 1316 5540 1324
rect 5596 1316 5604 1324
rect 5676 1316 5684 1324
rect 5724 1316 5732 1324
rect 5932 1316 5940 1324
rect 5996 1316 6004 1324
rect 6012 1316 6020 1324
rect 6044 1316 6052 1324
rect 6092 1316 6100 1324
rect 6124 1336 6132 1344
rect 6172 1336 6180 1344
rect 6188 1336 6196 1344
rect 6412 1336 6420 1344
rect 6636 1336 6644 1344
rect 6204 1316 6212 1324
rect 6332 1316 6340 1324
rect 6476 1316 6484 1324
rect 6492 1316 6500 1324
rect 6540 1316 6548 1324
rect 6572 1316 6580 1324
rect 6652 1316 6660 1324
rect 6684 1316 6692 1324
rect 6796 1316 6804 1324
rect 5500 1296 5508 1304
rect 5852 1296 5860 1304
rect 5900 1296 5908 1304
rect 5948 1296 5956 1304
rect 5964 1296 5972 1304
rect 6172 1296 6180 1304
rect 6204 1296 6212 1304
rect 6684 1296 6692 1304
rect 476 1276 484 1284
rect 1036 1276 1044 1284
rect 1356 1276 1364 1284
rect 1724 1276 1732 1284
rect 2380 1276 2388 1284
rect 2940 1276 2948 1284
rect 5180 1276 5188 1284
rect 5948 1276 5956 1284
rect 6444 1276 6452 1284
rect 1964 1256 1972 1264
rect 3340 1254 3348 1262
rect 3580 1254 3588 1262
rect 4204 1254 4212 1262
rect 188 1236 196 1244
rect 764 1236 772 1244
rect 956 1236 964 1244
rect 1260 1236 1268 1244
rect 1340 1236 1348 1244
rect 2028 1236 2036 1244
rect 2284 1236 2292 1244
rect 2364 1236 2372 1244
rect 2428 1236 2436 1244
rect 2508 1236 2516 1244
rect 3420 1236 3428 1244
rect 3500 1236 3508 1244
rect 3836 1236 3844 1244
rect 3884 1236 3892 1244
rect 4300 1236 4308 1244
rect 4396 1236 4404 1244
rect 4476 1236 4484 1244
rect 4732 1236 4740 1244
rect 4796 1236 4804 1244
rect 5580 1236 5588 1244
rect 6524 1236 6532 1244
rect 1118 1206 1126 1214
rect 1132 1206 1140 1214
rect 1146 1206 1154 1214
rect 4158 1206 4166 1214
rect 4172 1206 4180 1214
rect 4186 1206 4194 1214
rect 300 1176 308 1184
rect 460 1176 468 1184
rect 732 1176 740 1184
rect 988 1176 996 1184
rect 1692 1176 1700 1184
rect 1996 1176 2004 1184
rect 2188 1176 2196 1184
rect 2236 1176 2244 1184
rect 3132 1176 3140 1184
rect 3580 1176 3588 1184
rect 3644 1176 3652 1184
rect 4092 1176 4100 1184
rect 4540 1176 4548 1184
rect 5772 1176 5780 1184
rect 5868 1176 5876 1184
rect 6396 1176 6404 1184
rect 6604 1176 6612 1184
rect 1820 1156 1828 1164
rect 2940 1158 2948 1166
rect 3900 1158 3908 1166
rect 4252 1156 4260 1164
rect 4828 1156 4836 1164
rect 5084 1158 5092 1166
rect 6044 1156 6052 1164
rect 668 1136 676 1144
rect 1244 1136 1252 1144
rect 2572 1136 2580 1144
rect 2684 1136 2692 1144
rect 3228 1136 3236 1144
rect 3292 1136 3300 1144
rect 4012 1136 4020 1144
rect 4124 1136 4132 1144
rect 4716 1136 4724 1144
rect 5260 1136 5268 1144
rect 6076 1136 6084 1144
rect 6252 1136 6260 1144
rect 1020 1116 1028 1124
rect 60 1094 68 1102
rect 124 1096 132 1104
rect 252 1096 260 1104
rect 268 1096 276 1104
rect 284 1096 292 1104
rect 348 1096 356 1104
rect 364 1096 372 1104
rect 428 1096 436 1104
rect 556 1096 564 1104
rect 684 1096 692 1104
rect 700 1096 708 1104
rect 780 1096 788 1104
rect 876 1096 884 1104
rect 1020 1096 1028 1104
rect 1068 1116 1076 1124
rect 1212 1116 1220 1124
rect 1276 1116 1284 1124
rect 1340 1116 1348 1124
rect 1500 1116 1508 1124
rect 1788 1116 1796 1124
rect 1852 1116 1860 1124
rect 1900 1116 1908 1124
rect 1932 1116 1940 1124
rect 1964 1116 1972 1124
rect 2076 1116 2084 1124
rect 2140 1116 2148 1124
rect 2172 1116 2180 1124
rect 2380 1116 2388 1124
rect 2444 1116 2452 1124
rect 2492 1116 2500 1124
rect 2604 1116 2612 1124
rect 2940 1112 2948 1120
rect 3260 1116 3268 1124
rect 3580 1116 3588 1124
rect 3900 1112 3908 1120
rect 4108 1116 4116 1124
rect 4540 1116 4548 1124
rect 4748 1116 4756 1124
rect 4796 1116 4804 1124
rect 5084 1112 5092 1120
rect 5228 1116 5236 1124
rect 5436 1116 5444 1124
rect 5516 1116 5524 1124
rect 5532 1116 5540 1124
rect 5836 1116 5844 1124
rect 5916 1116 5924 1124
rect 1148 1096 1156 1104
rect 1180 1096 1188 1104
rect 1308 1096 1316 1104
rect 1372 1096 1380 1104
rect 1388 1096 1396 1104
rect 1420 1096 1428 1104
rect 1436 1096 1444 1104
rect 1468 1096 1476 1104
rect 1500 1096 1508 1104
rect 1564 1094 1572 1102
rect 1756 1096 1764 1104
rect 1932 1096 1940 1104
rect 1996 1096 2004 1104
rect 2172 1096 2180 1104
rect 2220 1096 2228 1104
rect 2268 1096 2276 1104
rect 2396 1096 2404 1104
rect 2412 1096 2420 1104
rect 2524 1096 2532 1104
rect 2956 1096 2964 1104
rect 3020 1096 3028 1104
rect 3084 1096 3092 1104
rect 3180 1096 3188 1104
rect 3372 1096 3380 1104
rect 3724 1096 3732 1104
rect 4044 1096 4052 1104
rect 4156 1096 4164 1104
rect 4332 1096 4340 1104
rect 4540 1096 4548 1104
rect 4636 1096 4644 1104
rect 4668 1096 4676 1104
rect 4908 1096 4916 1104
rect 5116 1096 5124 1104
rect 5212 1096 5220 1104
rect 5260 1096 5268 1104
rect 5420 1096 5428 1104
rect 5468 1096 5476 1104
rect 5564 1096 5572 1104
rect 5612 1096 5620 1104
rect 5628 1096 5636 1104
rect 5644 1096 5652 1104
rect 5868 1096 5876 1104
rect 5900 1096 5908 1104
rect 5964 1116 5972 1124
rect 6172 1094 6180 1102
rect 6252 1096 6260 1104
rect 6300 1116 6308 1124
rect 6780 1116 6788 1124
rect 6348 1096 6356 1104
rect 6364 1096 6372 1104
rect 6380 1096 6388 1104
rect 6428 1096 6436 1104
rect 6524 1096 6532 1104
rect 6572 1096 6580 1104
rect 6748 1096 6756 1104
rect 6796 1096 6804 1104
rect 6812 1096 6820 1104
rect 6860 1096 6868 1104
rect 412 1076 420 1084
rect 508 1076 516 1084
rect 876 1076 884 1084
rect 1004 1076 1012 1084
rect 1116 1076 1124 1084
rect 1228 1076 1236 1084
rect 1244 1076 1252 1084
rect 1276 1076 1284 1084
rect 1452 1076 1460 1084
rect 1532 1076 1540 1084
rect 1804 1076 1812 1084
rect 1884 1076 1892 1084
rect 1948 1076 1956 1084
rect 2012 1076 2020 1084
rect 2108 1076 2116 1084
rect 2172 1076 2180 1084
rect 2284 1076 2292 1084
rect 2332 1076 2340 1084
rect 2396 1076 2404 1084
rect 2508 1076 2516 1084
rect 2668 1076 2676 1084
rect 2876 1076 2884 1084
rect 3068 1076 3076 1084
rect 3116 1076 3124 1084
rect 3164 1076 3172 1084
rect 3276 1076 3284 1084
rect 3484 1076 3492 1084
rect 3836 1076 3844 1084
rect 3980 1076 3988 1084
rect 4028 1076 4036 1084
rect 4060 1076 4068 1084
rect 4076 1076 4084 1084
rect 4172 1076 4180 1084
rect 4444 1076 4452 1084
rect 4588 1076 4596 1084
rect 4652 1076 4660 1084
rect 4700 1076 4708 1084
rect 4716 1076 4724 1084
rect 4764 1076 4772 1084
rect 4812 1076 4820 1084
rect 5020 1076 5028 1084
rect 5164 1076 5172 1084
rect 5276 1076 5284 1084
rect 5292 1076 5300 1084
rect 5420 1076 5428 1084
rect 5484 1076 5492 1084
rect 5500 1076 5508 1084
rect 5532 1076 5540 1084
rect 5740 1076 5748 1084
rect 5884 1076 5892 1084
rect 5900 1076 5908 1084
rect 5996 1076 6004 1084
rect 6204 1076 6212 1084
rect 6236 1076 6244 1084
rect 6348 1076 6356 1084
rect 6716 1076 6724 1084
rect 6732 1076 6740 1084
rect 780 1056 788 1064
rect 1340 1056 1348 1064
rect 1868 1056 1876 1064
rect 2028 1056 2036 1064
rect 2124 1056 2132 1064
rect 2204 1056 2212 1064
rect 2252 1056 2260 1064
rect 2316 1056 2324 1064
rect 2844 1056 2852 1064
rect 3148 1056 3156 1064
rect 3452 1056 3460 1064
rect 3804 1056 3812 1064
rect 3996 1056 4004 1064
rect 4412 1056 4420 1064
rect 4988 1056 4996 1064
rect 5820 1056 5828 1064
rect 6476 1056 6484 1064
rect 188 1036 196 1044
rect 220 1036 228 1044
rect 460 1036 468 1044
rect 796 1036 804 1044
rect 2044 1036 2052 1044
rect 2492 1036 2500 1044
rect 3644 1036 3652 1044
rect 4124 1036 4132 1044
rect 4748 1036 4756 1044
rect 5676 1036 5684 1044
rect 5772 1036 5780 1044
rect 6012 1036 6020 1044
rect 6540 1036 6548 1044
rect 6780 1036 6788 1044
rect 6828 1036 6836 1044
rect 2638 1006 2646 1014
rect 2652 1006 2660 1014
rect 2666 1006 2674 1014
rect 5726 1006 5734 1014
rect 5740 1006 5748 1014
rect 5754 1006 5762 1014
rect 12 976 20 984
rect 348 976 356 984
rect 588 976 596 984
rect 716 976 724 984
rect 1212 976 1220 984
rect 1484 976 1492 984
rect 1740 976 1748 984
rect 1772 976 1780 984
rect 2140 976 2148 984
rect 2236 976 2244 984
rect 2300 976 2308 984
rect 2556 976 2564 984
rect 2924 976 2932 984
rect 4444 976 4452 984
rect 4652 976 4660 984
rect 5068 976 5076 984
rect 5100 976 5108 984
rect 5132 976 5140 984
rect 5276 976 5284 984
rect 5836 976 5844 984
rect 6124 976 6132 984
rect 6508 976 6516 984
rect 6876 976 6884 984
rect 908 956 916 964
rect 1500 956 1508 964
rect 1932 956 1940 964
rect 2716 956 2724 964
rect 3244 956 3252 964
rect 3420 956 3428 964
rect 3612 956 3620 964
rect 3900 956 3908 964
rect 4252 956 4260 964
rect 4844 956 4852 964
rect 5180 956 5188 964
rect 5356 956 5364 964
rect 5516 956 5524 964
rect 5756 956 5764 964
rect 60 936 68 944
rect 220 936 228 944
rect 236 936 244 944
rect 300 936 308 944
rect 364 936 372 944
rect 428 936 436 944
rect 540 936 548 944
rect 636 936 644 944
rect 876 936 884 944
rect 1116 936 1124 944
rect 1340 936 1348 944
rect 1452 936 1460 944
rect 1964 936 1972 944
rect 2108 936 2116 944
rect 2140 936 2148 944
rect 2252 936 2260 944
rect 2316 936 2324 944
rect 2476 936 2484 944
rect 2508 936 2516 944
rect 2748 936 2756 944
rect 2956 936 2964 944
rect 3052 936 3060 944
rect 3276 936 3284 944
rect 3580 936 3588 944
rect 3804 936 3812 944
rect 3916 936 3924 944
rect 4284 936 4292 944
rect 4428 936 4436 944
rect 4524 936 4532 944
rect 4588 936 4596 944
rect 4604 936 4612 944
rect 4876 936 4884 944
rect 5020 936 5028 944
rect 5084 936 5092 944
rect 5180 936 5188 944
rect 5212 936 5220 944
rect 5420 936 5428 944
rect 5580 936 5588 944
rect 5644 936 5652 944
rect 5996 936 6004 944
rect 6108 936 6116 944
rect 6172 936 6180 944
rect 6188 936 6196 944
rect 6300 936 6308 944
rect 6348 936 6356 944
rect 6364 936 6372 944
rect 6444 936 6452 944
rect 92 916 100 924
rect 140 916 148 924
rect 156 916 164 924
rect 172 916 180 924
rect 204 916 212 924
rect 268 916 276 924
rect 316 916 324 924
rect 380 916 388 924
rect 412 916 420 924
rect 12 896 20 904
rect 172 896 180 904
rect 236 896 244 904
rect 348 896 356 904
rect 412 896 420 904
rect 476 896 484 904
rect 524 916 532 924
rect 540 916 548 924
rect 572 916 580 924
rect 652 916 660 924
rect 700 916 708 924
rect 828 916 836 924
rect 924 916 932 924
rect 940 916 948 924
rect 1020 916 1028 924
rect 1100 916 1108 924
rect 1180 916 1188 924
rect 1260 916 1268 924
rect 1308 916 1316 924
rect 1324 916 1332 924
rect 1340 916 1348 924
rect 1004 896 1012 904
rect 1388 896 1396 904
rect 1436 916 1444 924
rect 1468 916 1476 924
rect 1564 918 1572 926
rect 1628 916 1636 924
rect 2060 916 2068 924
rect 1436 896 1444 904
rect 1740 896 1748 904
rect 2028 900 2036 908
rect 2172 916 2180 924
rect 2268 916 2276 924
rect 2524 916 2532 924
rect 2636 916 2644 924
rect 2892 916 2900 924
rect 2972 916 2980 924
rect 3164 916 3172 924
rect 3372 916 3380 924
rect 3692 916 3700 924
rect 3820 916 3828 924
rect 3932 916 3940 924
rect 4380 916 4388 924
rect 4492 916 4500 924
rect 4508 916 4516 924
rect 4572 916 4580 924
rect 4604 916 4612 924
rect 4764 916 4772 924
rect 4956 916 4964 924
rect 5036 916 5044 924
rect 5308 916 5316 924
rect 5356 916 5364 924
rect 5468 916 5476 924
rect 5628 916 5636 924
rect 5676 916 5684 924
rect 5724 916 5732 924
rect 5740 916 5748 924
rect 5964 918 5972 926
rect 6028 916 6036 924
rect 6044 916 6052 924
rect 6092 916 6100 924
rect 6156 916 6164 924
rect 6204 916 6212 924
rect 2204 896 2212 904
rect 2428 896 2436 904
rect 2844 896 2852 904
rect 3020 896 3028 904
rect 3052 896 3060 904
rect 3084 896 3092 904
rect 3340 900 3348 908
rect 3516 900 3524 908
rect 3868 896 3876 904
rect 3900 896 3908 904
rect 4012 896 4020 904
rect 4092 896 4100 904
rect 4348 900 4356 908
rect 4460 896 4468 904
rect 4540 896 4548 904
rect 4940 900 4948 908
rect 5068 896 5076 904
rect 5260 896 5268 904
rect 5276 896 5284 904
rect 5372 896 5380 904
rect 5436 896 5444 904
rect 5532 896 5540 904
rect 5596 896 5604 904
rect 6124 896 6132 904
rect 6204 896 6212 904
rect 6300 916 6308 924
rect 6316 916 6324 924
rect 6364 916 6372 924
rect 6412 916 6420 924
rect 6460 916 6468 924
rect 6572 916 6580 924
rect 6636 918 6644 926
rect 6796 916 6804 924
rect 6252 896 6260 904
rect 6428 896 6436 904
rect 524 876 532 884
rect 972 876 980 884
rect 1036 876 1044 884
rect 1484 876 1492 884
rect 3980 876 3988 884
rect 4476 876 4484 884
rect 4652 876 4660 884
rect 5116 876 5124 884
rect 5132 876 5140 884
rect 268 856 276 864
rect 2028 854 2036 862
rect 3340 854 3348 862
rect 4940 854 4948 862
rect 5228 856 5236 864
rect 380 836 388 844
rect 1100 836 1108 844
rect 1292 836 1300 844
rect 1692 836 1700 844
rect 2380 836 2388 844
rect 2844 836 2852 844
rect 3436 836 3444 844
rect 3516 836 3524 844
rect 3772 836 3780 844
rect 3996 836 4004 844
rect 4348 836 4356 844
rect 4572 836 4580 844
rect 5564 836 5572 844
rect 5708 836 5716 844
rect 6460 836 6468 844
rect 1118 806 1126 814
rect 1132 806 1140 814
rect 1146 806 1154 814
rect 4158 806 4166 814
rect 4172 806 4180 814
rect 4186 806 4194 814
rect 860 776 868 784
rect 1628 776 1636 784
rect 1868 776 1876 784
rect 2396 776 2404 784
rect 2684 776 2692 784
rect 2780 776 2788 784
rect 3404 776 3412 784
rect 3836 776 3844 784
rect 4620 776 4628 784
rect 4684 776 4692 784
rect 5532 776 5540 784
rect 5900 776 5908 784
rect 6124 776 6132 784
rect 6172 776 6180 784
rect 6668 776 6676 784
rect 6700 776 6708 784
rect 3084 758 3092 766
rect 4380 758 4388 766
rect 5804 756 5812 764
rect 6844 756 6852 764
rect 188 736 196 744
rect 1452 736 1460 744
rect 1692 736 1700 744
rect 3004 736 3012 744
rect 3340 736 3348 744
rect 5548 736 5556 744
rect 5836 736 5844 744
rect 5852 736 5860 744
rect 6108 736 6116 744
rect 6236 736 6244 744
rect 6444 736 6452 744
rect 252 716 260 724
rect 92 696 100 704
rect 204 696 212 704
rect 428 716 436 724
rect 460 716 468 724
rect 940 716 948 724
rect 1196 716 1204 724
rect 1308 716 1316 724
rect 1404 716 1412 724
rect 1420 716 1428 724
rect 1468 716 1476 724
rect 1532 716 1540 724
rect 1596 716 1604 724
rect 1660 716 1668 724
rect 1724 716 1732 724
rect 1836 716 1844 724
rect 2316 716 2324 724
rect 2396 716 2404 724
rect 2908 716 2916 724
rect 3084 712 3092 720
rect 3404 716 3412 724
rect 300 696 308 704
rect 332 696 340 704
rect 348 696 356 704
rect 380 696 388 704
rect 428 696 436 704
rect 204 676 212 684
rect 316 676 324 684
rect 476 676 484 684
rect 508 696 516 704
rect 556 696 564 704
rect 588 696 596 704
rect 604 696 612 704
rect 652 696 660 704
rect 668 696 676 704
rect 732 694 740 702
rect 1020 696 1028 704
rect 1148 696 1156 704
rect 1228 696 1236 704
rect 1276 696 1284 704
rect 1372 696 1380 704
rect 1404 696 1412 704
rect 1436 696 1444 704
rect 1500 696 1508 704
rect 1564 696 1572 704
rect 1628 696 1636 704
rect 1676 696 1684 704
rect 1740 696 1748 704
rect 1788 696 1796 704
rect 2236 696 2244 704
rect 2300 696 2308 704
rect 2396 696 2404 704
rect 2604 696 2612 704
rect 2972 696 2980 704
rect 2988 696 2996 704
rect 3052 696 3060 704
rect 3436 696 3444 704
rect 3964 716 3972 724
rect 4044 716 4052 724
rect 4380 712 4388 720
rect 4460 716 4468 724
rect 4508 716 4516 724
rect 4684 716 4692 724
rect 5084 716 5092 724
rect 4396 696 4404 704
rect 4540 696 4548 704
rect 4684 696 4692 704
rect 5084 696 5092 704
rect 5132 716 5140 724
rect 5580 716 5588 724
rect 5644 716 5652 724
rect 5164 696 5172 704
rect 5388 694 5396 702
rect 5564 696 5572 704
rect 5612 696 5620 704
rect 5692 716 5700 724
rect 5772 716 5780 724
rect 5884 716 5892 724
rect 6140 716 6148 724
rect 6268 716 6276 724
rect 6428 716 6436 724
rect 6636 716 6644 724
rect 5708 696 5716 704
rect 5804 696 5812 704
rect 5868 696 5876 704
rect 6012 696 6020 704
rect 6124 696 6132 704
rect 6156 696 6164 704
rect 6252 696 6260 704
rect 6284 696 6292 704
rect 6300 696 6308 704
rect 6364 696 6372 704
rect 6396 696 6404 704
rect 6428 696 6436 704
rect 6524 696 6532 704
rect 6668 696 6676 704
rect 700 676 708 684
rect 908 676 916 684
rect 972 676 980 684
rect 1244 676 1252 684
rect 1260 676 1268 684
rect 1324 676 1332 684
rect 1484 676 1492 684
rect 1548 676 1556 684
rect 1612 676 1620 684
rect 1676 676 1684 684
rect 1804 676 1812 684
rect 1852 676 1860 684
rect 1932 676 1940 684
rect 2028 676 2036 684
rect 2044 676 2052 684
rect 2348 676 2356 684
rect 2492 676 2500 684
rect 2892 676 2900 684
rect 2940 676 2948 684
rect 2956 676 2964 684
rect 3148 676 3156 684
rect 3500 676 3508 684
rect 3724 676 3732 684
rect 3900 676 3908 684
rect 4012 676 4020 684
rect 4316 676 4324 684
rect 4492 676 4500 684
rect 4572 676 4580 684
rect 4636 676 4644 684
rect 4780 676 4788 684
rect 5180 676 5188 684
rect 5324 676 5332 684
rect 5420 676 5428 684
rect 5596 676 5604 684
rect 5708 676 5716 684
rect 5820 676 5828 684
rect 6060 676 6068 684
rect 6156 676 6164 684
rect 6348 676 6356 684
rect 6380 676 6388 684
rect 6572 676 6580 684
rect 6684 676 6692 684
rect 6732 676 6740 684
rect 60 656 68 664
rect 268 656 276 664
rect 876 656 884 664
rect 1324 656 1332 664
rect 1532 656 1540 664
rect 1916 656 1924 664
rect 2268 656 2276 664
rect 2524 656 2532 664
rect 2924 656 2932 664
rect 3180 656 3188 664
rect 3532 656 3540 664
rect 3868 656 3876 664
rect 4284 656 4292 664
rect 4812 656 4820 664
rect 4972 656 4980 664
rect 4988 656 4996 664
rect 5020 656 5028 664
rect 5036 656 5044 664
rect 6716 656 6724 664
rect 620 636 628 644
rect 892 636 900 644
rect 940 636 948 644
rect 1132 636 1140 644
rect 1596 636 1604 644
rect 1772 636 1780 644
rect 1820 636 1828 644
rect 1964 636 1972 644
rect 2156 636 2164 644
rect 2204 636 2212 644
rect 2316 636 2324 644
rect 3692 636 3700 644
rect 3948 636 3956 644
rect 4076 636 4084 644
rect 4460 636 4468 644
rect 4508 636 4516 644
rect 5212 636 5220 644
rect 5516 636 5524 644
rect 2638 606 2646 614
rect 2652 606 2660 614
rect 2666 606 2674 614
rect 5726 606 5734 614
rect 5740 606 5748 614
rect 5754 606 5762 614
rect 188 576 196 584
rect 348 576 356 584
rect 396 576 404 584
rect 828 576 836 584
rect 860 576 868 584
rect 1068 576 1076 584
rect 1228 576 1236 584
rect 1484 576 1492 584
rect 1676 576 1684 584
rect 2124 576 2132 584
rect 2524 576 2532 584
rect 3596 576 3604 584
rect 3996 576 4004 584
rect 4524 576 4532 584
rect 4556 576 4564 584
rect 4908 576 4916 584
rect 5068 576 5076 584
rect 5260 576 5268 584
rect 5356 576 5364 584
rect 5612 576 5620 584
rect 5804 576 5812 584
rect 5852 576 5860 584
rect 5996 576 6004 584
rect 6828 576 6836 584
rect 60 556 68 564
rect 700 556 708 564
rect 1404 556 1412 564
rect 1468 556 1476 564
rect 1596 556 1604 564
rect 1756 556 1764 564
rect 1932 556 1940 564
rect 2332 556 2340 564
rect 2796 556 2804 564
rect 3324 556 3332 564
rect 3756 556 3764 564
rect 4156 556 4164 564
rect 4428 556 4436 564
rect 4748 556 4756 564
rect 5196 556 5204 564
rect 6124 556 6132 564
rect 204 536 212 544
rect 268 536 276 544
rect 316 536 324 544
rect 364 536 372 544
rect 380 536 388 544
rect 412 536 420 544
rect 524 536 532 544
rect 636 536 644 544
rect 668 536 676 544
rect 844 536 852 544
rect 924 536 932 544
rect 1180 536 1188 544
rect 1244 536 1252 544
rect 1308 536 1316 544
rect 1964 536 1972 544
rect 2300 536 2308 544
rect 2572 536 2580 544
rect 2764 536 2772 544
rect 2972 536 2980 544
rect 3084 536 3092 544
rect 3100 536 3108 544
rect 3356 536 3364 544
rect 3564 536 3572 544
rect 3788 536 3796 544
rect 3932 536 3940 544
rect 4188 536 4196 544
rect 4412 536 4420 544
rect 4444 536 4452 544
rect 4492 536 4500 544
rect 4540 536 4548 544
rect 4716 536 4724 544
rect 4924 536 4932 544
rect 4988 536 4996 544
rect 5004 536 5012 544
rect 5052 536 5060 544
rect 5100 536 5108 544
rect 5244 536 5252 544
rect 5292 536 5300 544
rect 5404 536 5412 544
rect 5436 536 5444 544
rect 5516 536 5524 544
rect 5580 536 5588 544
rect 5676 536 5684 544
rect 5692 536 5700 544
rect 5836 536 5844 544
rect 5884 536 5892 544
rect 6268 536 6276 544
rect 6492 536 6500 544
rect 6508 536 6516 544
rect 6556 536 6564 544
rect 6732 536 6740 544
rect 6748 536 6756 544
rect 6876 536 6884 544
rect 92 516 100 524
rect 124 516 132 524
rect 220 516 228 524
rect 252 496 260 504
rect 300 516 308 524
rect 444 516 452 524
rect 492 516 500 524
rect 508 516 516 524
rect 540 516 548 524
rect 572 496 580 504
rect 604 516 612 524
rect 620 516 628 524
rect 700 518 708 526
rect 940 516 948 524
rect 956 516 964 524
rect 1004 516 1012 524
rect 1052 516 1060 524
rect 1100 516 1108 524
rect 1116 516 1124 524
rect 1180 516 1188 524
rect 1196 516 1204 524
rect 1260 516 1268 524
rect 1276 516 1284 524
rect 1324 516 1332 524
rect 1372 516 1380 524
rect 1388 516 1396 524
rect 1436 516 1444 524
rect 1516 516 1524 524
rect 1564 516 1572 524
rect 1580 516 1588 524
rect 1644 516 1652 524
rect 1708 516 1716 524
rect 2060 516 2068 524
rect 2156 516 2164 524
rect 2188 516 2196 524
rect 2204 516 2212 524
rect 2556 516 2564 524
rect 2668 516 2676 524
rect 2876 516 2884 524
rect 3068 516 3076 524
rect 3436 516 3444 524
rect 3580 516 3588 524
rect 3676 516 3684 524
rect 3788 516 3796 524
rect 4284 516 4292 524
rect 4348 516 4356 524
rect 4620 516 4628 524
rect 4988 516 4996 524
rect 5036 516 5044 524
rect 5148 516 5156 524
rect 5228 516 5236 524
rect 5308 516 5316 524
rect 876 496 884 504
rect 892 496 900 504
rect 1228 496 1236 504
rect 1292 496 1300 504
rect 1356 496 1364 504
rect 1676 496 1684 504
rect 1692 496 1700 504
rect 2028 500 2036 508
rect 2236 500 2244 508
rect 2700 500 2708 508
rect 2956 496 2964 504
rect 2988 496 2996 504
rect 3020 496 3028 504
rect 3420 500 3428 508
rect 3884 496 3892 504
rect 4252 500 4260 508
rect 4652 500 4660 508
rect 4940 496 4948 504
rect 5004 496 5012 504
rect 5116 496 5124 504
rect 5340 496 5348 504
rect 5388 516 5396 524
rect 5404 516 5412 524
rect 5420 516 5428 524
rect 5484 516 5492 524
rect 5500 516 5508 524
rect 5532 516 5540 524
rect 5548 516 5556 524
rect 5660 516 5668 524
rect 5916 516 5924 524
rect 5964 516 5972 524
rect 5980 516 5988 524
rect 6124 518 6132 526
rect 6188 516 6196 524
rect 6204 516 6212 524
rect 6252 516 6260 524
rect 6332 516 6340 524
rect 6348 516 6356 524
rect 6364 516 6372 524
rect 6412 516 6420 524
rect 6476 516 6484 524
rect 6508 516 6516 524
rect 6540 516 6548 524
rect 6588 516 6596 524
rect 6636 516 6644 524
rect 6652 516 6660 524
rect 6668 516 6676 524
rect 6684 516 6692 524
rect 6764 516 6772 524
rect 6780 516 6788 524
rect 5564 496 5572 504
rect 5612 496 5620 504
rect 5628 496 5636 504
rect 5852 496 5860 504
rect 6444 496 6452 504
rect 6508 496 6516 504
rect 6812 496 6820 504
rect 6860 516 6868 524
rect 332 476 340 484
rect 412 476 420 484
rect 1324 476 1332 484
rect 1724 476 1732 484
rect 2524 476 2532 484
rect 3132 476 3140 484
rect 4332 476 4340 484
rect 4540 476 4548 484
rect 4572 476 4580 484
rect 5068 476 5076 484
rect 5276 476 5284 484
rect 6476 476 6484 484
rect 1708 456 1716 464
rect 2028 454 2036 462
rect 2124 456 2132 464
rect 2236 454 2244 462
rect 2700 454 2708 462
rect 3420 454 3428 462
rect 908 436 916 444
rect 988 436 996 444
rect 1532 436 1540 444
rect 3116 436 3124 444
rect 3596 436 3604 444
rect 3884 436 3892 444
rect 3948 436 3956 444
rect 4252 436 4260 444
rect 4476 436 4484 444
rect 4652 436 4660 444
rect 5148 436 5156 444
rect 5660 436 5668 444
rect 5932 436 5940 444
rect 6300 436 6308 444
rect 6396 436 6404 444
rect 6620 436 6628 444
rect 1118 406 1126 414
rect 1132 406 1140 414
rect 1146 406 1154 414
rect 4158 406 4166 414
rect 4172 406 4180 414
rect 4186 406 4194 414
rect 44 376 52 384
rect 332 376 340 384
rect 668 376 676 384
rect 908 376 916 384
rect 1356 376 1364 384
rect 1452 376 1460 384
rect 1724 376 1732 384
rect 1756 376 1764 384
rect 1836 376 1844 384
rect 2284 376 2292 384
rect 2908 376 2916 384
rect 3756 376 3764 384
rect 4636 376 4644 384
rect 4972 376 4980 384
rect 5260 376 5268 384
rect 5644 376 5652 384
rect 5948 376 5956 384
rect 6716 376 6724 384
rect 6812 376 6820 384
rect 1036 356 1044 364
rect 2396 358 2404 366
rect 3404 358 3412 366
rect 4380 358 4388 366
rect 4140 336 4148 344
rect 5724 336 5732 344
rect 5980 336 5988 344
rect 6268 336 6276 344
rect 44 316 52 324
rect 76 296 84 304
rect 412 296 420 304
rect 460 316 468 324
rect 572 316 580 324
rect 636 316 644 324
rect 940 316 948 324
rect 1004 316 1012 324
rect 1068 316 1076 324
rect 1100 316 1108 324
rect 1420 316 1428 324
rect 1436 316 1444 324
rect 1484 316 1492 324
rect 2284 316 2292 324
rect 2396 312 2404 320
rect 508 296 516 304
rect 588 296 596 304
rect 604 296 612 304
rect 972 296 980 304
rect 1036 296 1044 304
rect 1100 296 1108 304
rect 1228 294 1236 302
rect 1372 296 1380 304
rect 1436 296 1444 304
rect 1500 296 1508 304
rect 1532 296 1540 304
rect 1596 294 1604 302
rect 1660 296 1668 304
rect 1852 296 1860 304
rect 1980 296 1988 304
rect 2076 296 2084 304
rect 2188 296 2196 304
rect 2348 296 2356 304
rect 2572 296 2580 304
rect 2716 296 2724 304
rect 2764 296 2772 304
rect 2796 316 2804 324
rect 2876 316 2884 324
rect 3084 316 3092 324
rect 3404 312 3412 320
rect 3708 316 3716 324
rect 3756 316 3764 324
rect 4108 316 4116 324
rect 4220 316 4228 324
rect 4380 312 4388 320
rect 3052 296 3060 304
rect 3084 296 3092 304
rect 3228 296 3236 304
rect 3436 296 3444 304
rect 3788 296 3796 304
rect 4108 296 4116 304
rect 4140 296 4148 304
rect 4348 296 4356 304
rect 4556 296 4564 304
rect 4668 296 4676 304
rect 4732 316 4740 324
rect 4796 316 4804 324
rect 4828 316 4836 324
rect 4860 316 4868 324
rect 5260 316 5268 324
rect 5308 316 5316 324
rect 4764 296 4772 304
rect 4828 296 4836 304
rect 4892 296 4900 304
rect 5052 296 5060 304
rect 5308 296 5316 304
rect 5340 296 5348 304
rect 5436 316 5444 324
rect 5468 296 5476 304
rect 5516 296 5524 304
rect 5564 316 5572 324
rect 6220 316 6228 324
rect 5596 296 5604 304
rect 5676 296 5684 304
rect 5692 296 5700 304
rect 5836 296 5844 304
rect 6108 294 6116 302
rect 6188 296 6196 304
rect 6540 316 6548 324
rect 140 276 148 284
rect 428 276 436 284
rect 524 276 532 284
rect 588 276 596 284
rect 652 276 660 284
rect 796 276 804 284
rect 988 276 996 284
rect 1052 276 1060 284
rect 1116 276 1124 284
rect 1244 276 1252 284
rect 1372 276 1380 284
rect 1468 276 1476 284
rect 1532 276 1540 284
rect 1868 276 1876 284
rect 1964 276 1972 284
rect 2188 276 2196 284
rect 2460 276 2468 284
rect 2732 276 2740 284
rect 2844 276 2852 284
rect 3020 276 3028 284
rect 3036 276 3044 284
rect 3340 276 3348 284
rect 3484 276 3492 284
rect 3660 276 3668 284
rect 3692 276 3700 284
rect 3852 276 3860 284
rect 4156 276 4164 284
rect 4268 276 4276 284
rect 4444 276 4452 284
rect 4652 276 4660 284
rect 4700 276 4708 284
rect 4780 276 4788 284
rect 4844 276 4852 284
rect 4876 276 4884 284
rect 5164 276 5172 284
rect 5356 276 5364 284
rect 5372 276 5380 284
rect 5404 276 5412 284
rect 5500 276 5508 284
rect 5596 276 5604 284
rect 5820 276 5828 284
rect 5916 276 5924 284
rect 6044 276 6052 284
rect 6140 276 6148 284
rect 6172 276 6180 284
rect 6284 276 6292 284
rect 6316 296 6324 304
rect 6364 296 6372 304
rect 6380 296 6388 304
rect 6412 296 6420 304
rect 6476 296 6484 304
rect 6508 296 6516 304
rect 6668 316 6676 324
rect 6588 296 6596 304
rect 6604 296 6612 304
rect 6716 296 6724 304
rect 6476 276 6484 284
rect 6492 276 6500 284
rect 6604 276 6612 284
rect 6620 276 6628 284
rect 6732 276 6740 284
rect 6748 276 6756 284
rect 6844 276 6852 284
rect 172 256 180 264
rect 364 256 372 264
rect 1740 256 1748 264
rect 1804 256 1812 264
rect 1820 256 1828 264
rect 2156 256 2164 264
rect 2492 256 2500 264
rect 3084 256 3092 264
rect 3308 256 3316 264
rect 3628 256 3636 264
rect 3884 256 3892 264
rect 4300 256 4308 264
rect 4476 256 4484 264
rect 4940 256 4948 264
rect 5132 256 5140 264
rect 636 236 644 244
rect 908 236 916 244
rect 940 236 948 244
rect 1788 236 1796 244
rect 2652 236 2660 244
rect 2860 236 2868 244
rect 2908 236 2916 244
rect 3148 236 3156 244
rect 3596 236 3604 244
rect 4044 236 4052 244
rect 4172 236 4180 244
rect 5548 236 5556 244
rect 6556 236 6564 244
rect 2638 206 2646 214
rect 2652 206 2660 214
rect 2666 206 2674 214
rect 5726 206 5734 214
rect 5740 206 5748 214
rect 5754 206 5762 214
rect 460 176 468 184
rect 492 176 500 184
rect 1404 176 1412 184
rect 1628 176 1636 184
rect 2668 176 2676 184
rect 3244 176 3252 184
rect 3372 176 3380 184
rect 4652 176 4660 184
rect 4684 176 4692 184
rect 5036 176 5044 184
rect 5404 176 5412 184
rect 5756 176 5764 184
rect 5884 176 5892 184
rect 6332 176 6340 184
rect 6364 176 6372 184
rect 6428 176 6436 184
rect 6620 176 6628 184
rect 6812 176 6820 184
rect 12 156 20 164
rect 204 156 212 164
rect 380 156 388 164
rect 444 156 452 164
rect 652 156 660 164
rect 1004 156 1012 164
rect 1452 156 1460 164
rect 1596 156 1604 164
rect 28 136 36 144
rect 172 136 180 144
rect 684 136 692 144
rect 842 136 850 144
rect 1036 136 1044 144
rect 1244 136 1252 144
rect 1676 156 1684 164
rect 1836 156 1844 164
rect 2172 156 2180 164
rect 2364 156 2372 164
rect 2444 156 2452 164
rect 2604 156 2612 164
rect 2732 156 2740 164
rect 2828 156 2836 164
rect 3004 156 3012 164
rect 3532 156 3540 164
rect 3964 156 3972 164
rect 4412 156 4420 164
rect 4588 156 4596 164
rect 4620 156 4628 164
rect 4636 156 4644 164
rect 4844 156 4852 164
rect 5020 156 5028 164
rect 5212 156 5220 164
rect 5388 156 5396 164
rect 5420 156 5428 164
rect 5596 156 5604 164
rect 6348 156 6356 164
rect 1868 136 1876 144
rect 2140 136 2148 144
rect 2508 136 2516 144
rect 2764 136 2772 144
rect 2828 136 2836 144
rect 3036 136 3044 144
rect 3292 136 3300 144
rect 3564 136 3572 144
rect 3932 136 3940 144
rect 4126 136 4134 144
rect 4380 136 4388 144
rect 4588 136 4596 144
rect 4876 136 4884 144
rect 5180 136 5188 144
rect 5564 136 5572 144
rect 6044 136 6052 144
rect 6076 136 6084 144
rect 6188 136 6196 144
rect 6316 136 6324 144
rect 6412 136 6420 144
rect 6492 136 6500 144
rect 6588 136 6596 144
rect 6876 136 6884 144
rect 76 116 84 124
rect 284 116 292 124
rect 444 116 452 124
rect 572 116 580 124
rect 780 116 788 124
rect 924 116 932 124
rect 1116 116 1124 124
rect 1276 118 1284 126
rect 1420 116 1428 124
rect 1564 116 1572 124
rect 1644 116 1652 124
rect 1964 116 1972 124
rect 2028 116 2036 124
rect 2252 116 2260 124
rect 2380 116 2388 124
rect 2396 116 2404 124
rect 2476 116 2484 124
rect 2604 116 2612 124
rect 2732 116 2740 124
rect 2924 116 2932 124
rect 3132 116 3140 124
rect 3212 116 3220 124
rect 3660 116 3668 124
rect 3708 116 3716 124
rect 3756 116 3764 124
rect 3836 116 3844 124
rect 4044 116 4052 124
rect 4188 116 4196 124
rect 4284 116 4292 124
rect 4492 116 4500 124
rect 4764 116 4772 124
rect 4988 116 4996 124
rect 5084 116 5092 124
rect 5292 116 5300 124
rect 5468 116 5476 124
rect 6012 118 6020 126
rect 6092 116 6100 124
rect 108 100 116 108
rect 780 96 788 104
rect 1132 96 1140 104
rect 1964 96 1972 104
rect 2076 100 2084 108
rect 2444 96 2452 104
rect 2508 96 2516 104
rect 2540 96 2548 104
rect 2812 96 2820 104
rect 3100 100 3108 108
rect 3660 96 3668 104
rect 3836 96 3844 104
rect 4284 96 4292 104
rect 4940 100 4948 108
rect 5084 96 5092 104
rect 5500 100 5508 108
rect 6092 96 6100 104
rect 6204 116 6212 124
rect 6140 96 6148 104
rect 6252 96 6260 104
rect 6300 116 6308 124
rect 6396 116 6404 124
rect 6540 116 6548 124
rect 6700 116 6708 124
rect 6732 116 6740 124
rect 6844 116 6852 124
rect 6300 96 6308 104
rect 6364 96 6372 104
rect 6812 96 6820 104
rect 2076 54 2084 62
rect 3100 54 3108 62
rect 4940 54 4948 62
rect 5500 54 5508 62
rect 108 36 116 44
rect 396 36 404 44
rect 780 36 788 44
rect 1132 36 1140 44
rect 1964 36 1972 44
rect 2428 36 2436 44
rect 2556 36 2564 44
rect 2684 36 2692 44
rect 3180 36 3188 44
rect 3308 36 3316 44
rect 3660 36 3668 44
rect 3740 36 3748 44
rect 3788 36 3796 44
rect 3836 36 3844 44
rect 4156 36 4164 44
rect 4284 36 4292 44
rect 5084 36 5092 44
rect 5868 36 5876 44
rect 1118 6 1126 14
rect 1132 6 1140 14
rect 1146 6 1154 14
rect 4158 6 4166 14
rect 4172 6 4180 14
rect 4186 6 4194 14
<< metal2 >>
rect 429 5037 451 5043
rect 445 4964 451 5037
rect 813 4964 819 5043
rect 1565 4964 1571 5043
rect 2237 5004 2243 5043
rect 2957 5037 2979 5043
rect 2632 5006 2638 5014
rect 2646 5006 2652 5014
rect 2660 5006 2666 5014
rect 2674 5006 2680 5014
rect 2973 4984 2979 5037
rect 3805 5037 3827 5043
rect 4269 5037 4291 5043
rect 3805 4984 3811 5037
rect 4285 4984 4291 5037
rect 4797 4964 4803 5043
rect 4845 5004 4851 5043
rect 4877 4984 4883 5043
rect 4845 4964 4851 4976
rect 4909 4964 4915 5043
rect 5389 5037 5411 5043
rect 45 4844 51 4896
rect 141 4824 147 4916
rect 173 4843 179 4956
rect 413 4904 419 4916
rect 173 4837 195 4843
rect 109 4704 115 4816
rect 29 4484 35 4636
rect 13 4324 19 4336
rect 29 4043 35 4476
rect 29 4037 51 4043
rect 13 3884 19 3896
rect 13 2904 19 2956
rect 29 2924 35 4037
rect 45 3904 51 4037
rect 77 3484 83 3496
rect 109 3304 115 4696
rect 189 4664 195 4837
rect 317 4724 323 4776
rect 333 4724 339 4836
rect 397 4784 403 4896
rect 525 4844 531 4900
rect 397 4704 403 4756
rect 621 4744 627 4956
rect 861 4924 867 4956
rect 1613 4944 1619 4956
rect 701 4864 707 4916
rect 861 4904 867 4916
rect 941 4904 947 4916
rect 893 4897 908 4903
rect 685 4704 691 4716
rect 781 4704 787 4736
rect 829 4704 835 4716
rect 189 4604 195 4656
rect 173 4597 188 4603
rect 173 4544 179 4597
rect 381 4584 387 4676
rect 141 4504 147 4518
rect 173 4284 179 4536
rect 205 4464 211 4536
rect 228 4517 243 4523
rect 205 4284 211 4456
rect 237 4424 243 4517
rect 269 4444 275 4496
rect 301 4304 307 4516
rect 317 4504 323 4536
rect 349 4524 355 4536
rect 397 4504 403 4696
rect 413 4504 419 4676
rect 429 4564 435 4636
rect 461 4544 467 4676
rect 525 4544 531 4694
rect 557 4604 563 4676
rect 685 4644 691 4696
rect 637 4637 652 4643
rect 468 4537 483 4543
rect 429 4504 435 4536
rect 205 4144 211 4276
rect 221 4164 227 4296
rect 317 4284 323 4496
rect 397 4484 403 4496
rect 365 4384 371 4416
rect 397 4304 403 4436
rect 413 4304 419 4376
rect 429 4324 435 4356
rect 445 4344 451 4516
rect 317 4164 323 4276
rect 125 3884 131 4116
rect 189 4084 195 4096
rect 205 4024 211 4136
rect 221 4124 227 4136
rect 349 4124 355 4176
rect 269 4104 275 4116
rect 253 4084 259 4096
rect 141 3904 147 3936
rect 269 3923 275 4096
rect 285 3984 291 4076
rect 333 4023 339 4116
rect 333 4017 355 4023
rect 260 3917 275 3923
rect 125 3724 131 3876
rect 189 3744 195 3776
rect 205 3764 211 3916
rect 221 3784 227 3796
rect 237 3744 243 3816
rect 125 3504 131 3716
rect 189 3584 195 3596
rect 237 3543 243 3736
rect 253 3724 259 3896
rect 333 3884 339 3896
rect 301 3824 307 3876
rect 253 3564 259 3716
rect 285 3704 291 3736
rect 301 3724 307 3736
rect 333 3724 339 3756
rect 349 3724 355 4017
rect 365 3964 371 4116
rect 397 4084 403 4296
rect 429 4144 435 4156
rect 445 4124 451 4336
rect 461 4244 467 4296
rect 477 4284 483 4537
rect 557 4464 563 4536
rect 589 4524 595 4636
rect 637 4524 643 4637
rect 717 4544 723 4656
rect 685 4517 700 4523
rect 557 4304 563 4356
rect 509 4164 515 4236
rect 477 4064 483 4096
rect 541 4044 547 4296
rect 557 4184 563 4296
rect 589 4283 595 4516
rect 637 4504 643 4516
rect 653 4384 659 4516
rect 669 4504 675 4516
rect 685 4384 691 4517
rect 717 4464 723 4536
rect 733 4444 739 4496
rect 717 4437 732 4443
rect 669 4304 675 4316
rect 573 4277 595 4283
rect 557 4024 563 4136
rect 573 4124 579 4277
rect 637 4264 643 4296
rect 653 4284 659 4296
rect 653 4164 659 4196
rect 573 4104 579 4116
rect 621 4064 627 4116
rect 637 4104 643 4116
rect 365 3904 371 3956
rect 429 3924 435 3976
rect 493 3904 499 3916
rect 493 3844 499 3896
rect 509 3884 515 4016
rect 637 3984 643 3996
rect 525 3884 531 3896
rect 573 3884 579 3896
rect 605 3884 611 3896
rect 461 3744 467 3756
rect 237 3537 259 3543
rect 125 3324 131 3496
rect 237 3324 243 3496
rect 253 3484 259 3537
rect 301 3504 307 3536
rect 349 3504 355 3556
rect 253 3464 259 3476
rect 253 3344 259 3456
rect 317 3444 323 3476
rect 333 3464 339 3476
rect 317 3344 323 3436
rect 333 3324 339 3336
rect 349 3324 355 3476
rect 365 3444 371 3736
rect 477 3724 483 3776
rect 525 3724 531 3736
rect 541 3724 547 3776
rect 381 3584 387 3716
rect 429 3704 435 3716
rect 397 3544 403 3636
rect 429 3604 435 3696
rect 461 3504 467 3576
rect 541 3504 547 3716
rect 557 3704 563 3756
rect 573 3697 588 3703
rect 573 3584 579 3697
rect 589 3524 595 3556
rect 477 3484 483 3496
rect 445 3444 451 3476
rect 397 3344 403 3436
rect 541 3384 547 3496
rect 557 3484 563 3496
rect 557 3404 563 3476
rect 413 3324 419 3376
rect 477 3326 483 3336
rect 125 3304 131 3316
rect 45 3124 51 3176
rect 77 3104 83 3296
rect 269 3284 275 3296
rect 157 2944 163 2956
rect 237 2944 243 3016
rect 61 2904 67 2916
rect 109 2884 115 2896
rect 45 2724 51 2776
rect 61 2684 67 2836
rect 173 2784 179 2876
rect 253 2704 259 3096
rect 285 2964 291 3096
rect 317 3024 323 3316
rect 397 3304 403 3316
rect 333 3124 339 3136
rect 349 3104 355 3276
rect 285 2944 291 2956
rect 349 2924 355 3096
rect 365 3084 371 3096
rect 381 2924 387 3156
rect 461 3104 467 3156
rect 493 2984 499 3356
rect 541 3324 547 3336
rect 589 3304 595 3516
rect 605 3503 611 3876
rect 653 3784 659 4096
rect 685 4084 691 4116
rect 669 4004 675 4036
rect 701 3903 707 4376
rect 717 4304 723 4437
rect 749 4303 755 4696
rect 765 4664 771 4676
rect 829 4664 835 4696
rect 845 4604 851 4736
rect 861 4624 867 4696
rect 877 4684 883 4876
rect 893 4844 899 4897
rect 893 4744 899 4836
rect 941 4764 947 4896
rect 957 4884 963 4936
rect 1261 4917 1276 4923
rect 989 4744 995 4836
rect 1112 4806 1118 4814
rect 1126 4806 1132 4814
rect 1140 4806 1146 4814
rect 1154 4806 1160 4814
rect 1229 4724 1235 4836
rect 845 4564 851 4596
rect 877 4564 883 4676
rect 781 4544 787 4556
rect 765 4344 771 4516
rect 765 4304 771 4336
rect 740 4297 755 4303
rect 733 4224 739 4296
rect 781 4284 787 4536
rect 845 4504 851 4518
rect 861 4464 867 4536
rect 797 4264 803 4316
rect 861 4284 867 4456
rect 877 4244 883 4256
rect 877 4164 883 4236
rect 909 4204 915 4636
rect 957 4304 963 4676
rect 989 4644 995 4694
rect 1117 4644 1123 4656
rect 989 4544 995 4556
rect 1005 4524 1011 4616
rect 973 4184 979 4436
rect 989 4304 995 4316
rect 797 4124 803 4136
rect 909 4104 915 4176
rect 989 4144 995 4276
rect 1005 4204 1011 4516
rect 1037 4444 1043 4496
rect 1037 4124 1043 4136
rect 781 3924 787 4036
rect 781 3904 787 3916
rect 692 3897 707 3903
rect 669 3864 675 3896
rect 669 3764 675 3856
rect 637 3744 643 3756
rect 685 3724 691 3896
rect 797 3884 803 4056
rect 893 3964 899 4036
rect 925 3923 931 4036
rect 989 3984 995 4016
rect 916 3917 931 3923
rect 829 3904 835 3916
rect 845 3904 851 3916
rect 813 3897 828 3903
rect 701 3864 707 3876
rect 717 3743 723 3836
rect 749 3824 755 3836
rect 797 3764 803 3836
rect 813 3744 819 3897
rect 957 3884 963 3956
rect 877 3844 883 3876
rect 973 3864 979 3896
rect 1021 3883 1027 3996
rect 1037 3904 1043 3956
rect 1021 3877 1036 3883
rect 717 3737 732 3743
rect 621 3704 627 3716
rect 701 3704 707 3736
rect 829 3724 835 3756
rect 733 3704 739 3716
rect 701 3564 707 3696
rect 605 3497 620 3503
rect 621 3484 627 3496
rect 605 3384 611 3396
rect 653 3384 659 3516
rect 685 3504 691 3536
rect 717 3524 723 3636
rect 733 3504 739 3696
rect 781 3664 787 3696
rect 669 3424 675 3496
rect 733 3484 739 3496
rect 749 3484 755 3516
rect 701 3364 707 3436
rect 717 3364 723 3456
rect 765 3444 771 3476
rect 797 3344 803 3676
rect 621 3324 627 3336
rect 701 3284 707 3336
rect 813 3324 819 3436
rect 829 3424 835 3516
rect 861 3504 867 3636
rect 877 3484 883 3836
rect 909 3743 915 3836
rect 957 3744 963 3796
rect 900 3737 915 3743
rect 973 3724 979 3856
rect 941 3664 947 3696
rect 877 3464 883 3476
rect 829 3384 835 3416
rect 845 3304 851 3316
rect 605 3124 611 3136
rect 653 3124 659 3176
rect 669 3164 675 3236
rect 509 3064 515 3116
rect 749 3084 755 3176
rect 877 3104 883 3456
rect 909 3404 915 3636
rect 925 3384 931 3496
rect 941 3424 947 3636
rect 957 3564 963 3716
rect 973 3644 979 3716
rect 1037 3704 1043 3716
rect 1005 3684 1011 3696
rect 957 3484 963 3556
rect 1005 3504 1011 3516
rect 941 3324 947 3416
rect 909 3124 915 3236
rect 941 3184 947 3236
rect 541 2963 547 3036
rect 557 2984 563 3056
rect 541 2957 563 2963
rect 429 2924 435 2956
rect 253 2623 259 2696
rect 269 2624 275 2916
rect 381 2904 387 2916
rect 333 2884 339 2896
rect 429 2884 435 2916
rect 477 2904 483 2916
rect 381 2704 387 2836
rect 477 2784 483 2896
rect 525 2884 531 2916
rect 557 2904 563 2957
rect 365 2664 371 2676
rect 237 2617 259 2623
rect 125 2584 131 2596
rect 109 2524 115 2556
rect 45 2504 51 2516
rect 13 2484 19 2496
rect 205 2384 211 2616
rect 237 2524 243 2617
rect 317 2564 323 2636
rect 445 2444 451 2496
rect 29 2184 35 2236
rect 141 2164 147 2276
rect 397 2184 403 2256
rect 404 2177 419 2183
rect 269 2164 275 2176
rect 13 2104 19 2156
rect 61 1904 67 2116
rect 93 2024 99 2096
rect 141 2044 147 2096
rect 109 1924 115 2036
rect 141 1984 147 2016
rect 205 1924 211 1976
rect 237 1904 243 2116
rect 13 1864 19 1896
rect 45 1644 51 1696
rect 61 1584 67 1736
rect 29 1464 35 1516
rect 77 1503 83 1896
rect 141 1844 147 1896
rect 237 1823 243 1896
rect 301 1864 307 1876
rect 237 1817 259 1823
rect 253 1724 259 1817
rect 333 1764 339 1856
rect 413 1764 419 2177
rect 493 2164 499 2676
rect 509 2664 515 2716
rect 509 2544 515 2636
rect 541 2604 547 2696
rect 573 2684 579 3076
rect 589 2724 595 3036
rect 605 2944 611 3076
rect 861 3064 867 3096
rect 957 3084 963 3476
rect 1021 3444 1027 3476
rect 1037 3444 1043 3496
rect 1053 3484 1059 3896
rect 1069 3584 1075 4296
rect 1085 4284 1091 4516
rect 1117 4464 1123 4636
rect 1181 4564 1187 4676
rect 1197 4624 1203 4696
rect 1245 4684 1251 4916
rect 1261 4704 1267 4917
rect 1325 4704 1331 4716
rect 1373 4704 1379 4836
rect 1485 4824 1491 4936
rect 1245 4544 1251 4656
rect 1261 4544 1267 4696
rect 1277 4644 1283 4696
rect 1293 4664 1299 4676
rect 1293 4564 1299 4616
rect 1373 4564 1379 4696
rect 1172 4437 1187 4443
rect 1112 4406 1118 4414
rect 1126 4406 1132 4414
rect 1140 4406 1146 4414
rect 1154 4406 1160 4414
rect 1181 4304 1187 4437
rect 1245 4384 1251 4536
rect 1149 4064 1155 4096
rect 1112 4006 1118 4014
rect 1126 4006 1132 4014
rect 1140 4006 1146 4014
rect 1154 4006 1160 4014
rect 1181 3944 1187 4296
rect 1197 4224 1203 4296
rect 1197 3944 1203 4036
rect 1213 3984 1219 4096
rect 1229 3964 1235 4296
rect 1261 4144 1267 4276
rect 1245 4124 1251 4136
rect 1277 4104 1283 4456
rect 1293 4384 1299 4556
rect 1389 4524 1395 4696
rect 1453 4524 1459 4536
rect 1469 4524 1475 4636
rect 1501 4624 1507 4936
rect 1613 4924 1619 4936
rect 1517 4904 1523 4916
rect 1565 4904 1571 4916
rect 1549 4884 1555 4896
rect 1677 4844 1683 4876
rect 1757 4864 1763 4916
rect 1533 4584 1539 4694
rect 1597 4684 1603 4836
rect 1677 4744 1683 4836
rect 1565 4644 1571 4676
rect 1645 4664 1651 4676
rect 1629 4544 1635 4636
rect 1645 4564 1651 4656
rect 1412 4517 1427 4523
rect 1085 3924 1091 3936
rect 1085 3704 1091 3716
rect 1117 3704 1123 3836
rect 1133 3704 1139 3936
rect 1213 3904 1219 3916
rect 1149 3824 1155 3856
rect 1149 3724 1155 3816
rect 1085 3664 1091 3696
rect 1181 3684 1187 3896
rect 1197 3704 1203 3716
rect 1149 3664 1155 3676
rect 1069 3524 1075 3536
rect 1085 3364 1091 3656
rect 1112 3606 1118 3614
rect 1126 3606 1132 3614
rect 1140 3606 1146 3614
rect 1154 3606 1160 3614
rect 1213 3584 1219 3896
rect 1229 3744 1235 3956
rect 1245 3924 1251 3936
rect 1261 3924 1267 3956
rect 1277 3904 1283 4076
rect 1293 3964 1299 4036
rect 1293 3904 1299 3916
rect 1277 3844 1283 3876
rect 1293 3864 1299 3896
rect 1309 3884 1315 4156
rect 1325 4044 1331 4296
rect 1341 4124 1347 4216
rect 1357 4164 1363 4436
rect 1373 4384 1379 4396
rect 1389 4364 1395 4516
rect 1421 4504 1427 4517
rect 1373 4144 1379 4156
rect 1357 3944 1363 4116
rect 1341 3904 1347 3936
rect 1357 3924 1363 3936
rect 1261 3763 1267 3836
rect 1293 3784 1299 3836
rect 1357 3824 1363 3896
rect 1373 3764 1379 4096
rect 1389 4004 1395 4356
rect 1405 4204 1411 4236
rect 1421 4123 1427 4496
rect 1469 4324 1475 4516
rect 1485 4404 1491 4536
rect 1645 4524 1651 4536
rect 1677 4524 1683 4696
rect 1725 4664 1731 4716
rect 1773 4684 1779 4696
rect 1837 4683 1843 4956
rect 2013 4944 2019 4956
rect 2397 4944 2403 4956
rect 2749 4944 2755 4956
rect 1869 4924 1875 4936
rect 1965 4844 1971 4896
rect 2349 4844 2355 4896
rect 2157 4724 2163 4776
rect 1821 4677 1843 4683
rect 1805 4664 1811 4676
rect 1821 4644 1827 4677
rect 1709 4544 1715 4636
rect 1757 4584 1763 4636
rect 1469 4163 1475 4316
rect 1517 4304 1523 4336
rect 1533 4304 1539 4496
rect 1549 4384 1555 4516
rect 1565 4484 1571 4516
rect 1613 4504 1619 4516
rect 1556 4377 1571 4383
rect 1549 4164 1555 4176
rect 1460 4157 1475 4163
rect 1412 4117 1427 4123
rect 1405 3984 1411 4116
rect 1501 4083 1507 4116
rect 1517 4104 1523 4136
rect 1549 4104 1555 4116
rect 1501 4077 1523 4083
rect 1389 3924 1395 3956
rect 1437 3944 1443 4036
rect 1245 3757 1267 3763
rect 1245 3744 1251 3757
rect 1261 3724 1267 3736
rect 1229 3704 1235 3716
rect 1165 3503 1171 3576
rect 1181 3504 1187 3516
rect 1197 3504 1203 3536
rect 1261 3524 1267 3716
rect 1261 3504 1267 3516
rect 1277 3504 1283 3616
rect 1325 3564 1331 3716
rect 1357 3683 1363 3756
rect 1405 3724 1411 3896
rect 1421 3744 1427 3916
rect 1437 3904 1443 3916
rect 1453 3884 1459 3916
rect 1437 3864 1443 3876
rect 1501 3864 1507 4036
rect 1517 3824 1523 4077
rect 1453 3764 1459 3796
rect 1501 3784 1507 3796
rect 1485 3764 1491 3776
rect 1373 3704 1379 3716
rect 1357 3677 1379 3683
rect 1156 3497 1171 3503
rect 1133 3464 1139 3476
rect 989 3324 995 3356
rect 1037 3304 1043 3356
rect 1117 3324 1123 3436
rect 1213 3384 1219 3496
rect 1309 3384 1315 3516
rect 973 3284 979 3296
rect 973 3184 979 3216
rect 1021 3184 1027 3276
rect 1037 3144 1043 3236
rect 781 2964 787 3056
rect 685 2844 691 2900
rect 781 2864 787 2956
rect 861 2924 867 3056
rect 973 2904 979 2936
rect 973 2724 979 2776
rect 573 2504 579 2656
rect 653 2604 659 2636
rect 669 2564 675 2636
rect 701 2544 707 2596
rect 765 2524 771 2696
rect 877 2684 883 2696
rect 845 2644 851 2656
rect 893 2584 899 2596
rect 973 2584 979 2696
rect 989 2604 995 3056
rect 1085 2944 1091 3316
rect 1181 3304 1187 3336
rect 1325 3304 1331 3456
rect 1341 3344 1347 3676
rect 1357 3504 1363 3556
rect 1373 3484 1379 3677
rect 1421 3484 1427 3496
rect 1437 3484 1443 3636
rect 1453 3484 1459 3676
rect 1501 3524 1507 3576
rect 1517 3524 1523 3816
rect 1357 3384 1363 3436
rect 1112 3206 1118 3214
rect 1126 3206 1132 3214
rect 1140 3206 1146 3214
rect 1154 3206 1160 3214
rect 1149 3124 1155 3176
rect 1101 2984 1107 3076
rect 1133 3064 1139 3096
rect 1117 2944 1123 2976
rect 1005 2744 1011 2896
rect 1021 2784 1027 2916
rect 1069 2904 1075 2936
rect 1085 2904 1091 2936
rect 1053 2784 1059 2876
rect 1112 2806 1118 2814
rect 1126 2806 1132 2814
rect 1140 2806 1146 2814
rect 1154 2806 1160 2814
rect 1117 2684 1123 2696
rect 1037 2604 1043 2656
rect 1069 2624 1075 2656
rect 1181 2644 1187 3296
rect 1341 3244 1347 3336
rect 1373 3144 1379 3476
rect 1405 3464 1411 3476
rect 1421 3444 1427 3476
rect 1469 3424 1475 3496
rect 1501 3384 1507 3436
rect 1405 3324 1411 3356
rect 1421 3344 1427 3356
rect 1517 3324 1523 3516
rect 1533 3484 1539 3896
rect 1549 3884 1555 4076
rect 1565 3904 1571 4377
rect 1613 4364 1619 4496
rect 1693 4404 1699 4536
rect 1700 4397 1715 4403
rect 1629 4277 1644 4283
rect 1581 3904 1587 3916
rect 1581 3804 1587 3896
rect 1565 3504 1571 3536
rect 1597 3524 1603 4236
rect 1629 4144 1635 4277
rect 1661 4144 1667 4316
rect 1693 4304 1699 4316
rect 1709 4284 1715 4397
rect 1725 4304 1731 4576
rect 1821 4544 1827 4636
rect 1853 4544 1859 4676
rect 1949 4564 1955 4696
rect 2317 4684 2323 4696
rect 1981 4524 1987 4616
rect 2029 4584 2035 4656
rect 2061 4584 2067 4676
rect 2205 4624 2211 4676
rect 2493 4664 2499 4936
rect 2525 4824 2531 4936
rect 2621 4844 2627 4896
rect 2717 4843 2723 4936
rect 2717 4837 2739 4843
rect 2733 4784 2739 4837
rect 2589 4720 2595 4758
rect 2093 4524 2099 4536
rect 1789 4304 1795 4356
rect 1821 4324 1827 4476
rect 1853 4384 1859 4496
rect 1677 4104 1683 4196
rect 1693 4124 1699 4156
rect 1709 4124 1715 4136
rect 1629 3824 1635 3896
rect 1677 3884 1683 4096
rect 1725 4064 1731 4296
rect 1741 4204 1747 4296
rect 1789 4144 1795 4276
rect 1805 4264 1811 4296
rect 1773 4137 1788 4143
rect 1773 3964 1779 4137
rect 1805 4124 1811 4256
rect 1821 4184 1827 4316
rect 1901 4304 1907 4476
rect 1981 4404 1987 4516
rect 2109 4304 2115 4436
rect 1853 4264 1859 4296
rect 1885 4264 1891 4296
rect 1853 4184 1859 4236
rect 1933 4184 1939 4256
rect 2061 4244 2067 4296
rect 2141 4264 2147 4476
rect 2157 4284 2163 4496
rect 2189 4384 2195 4516
rect 2173 4304 2179 4316
rect 2205 4284 2211 4616
rect 2445 4564 2451 4576
rect 2221 4484 2227 4496
rect 2221 4263 2227 4476
rect 2253 4344 2259 4436
rect 2276 4297 2291 4303
rect 2253 4284 2259 4296
rect 2212 4257 2227 4263
rect 1949 4144 1955 4236
rect 2093 4164 2099 4216
rect 2157 4204 2163 4236
rect 1789 4103 1795 4116
rect 1837 4104 1843 4136
rect 1885 4104 1891 4116
rect 1789 4097 1811 4103
rect 1757 3904 1763 3916
rect 1773 3884 1779 3956
rect 1789 3904 1795 3996
rect 1805 3904 1811 4097
rect 1869 3903 1875 3916
rect 1885 3904 1891 3936
rect 1860 3897 1875 3903
rect 1661 3844 1667 3876
rect 1629 3704 1635 3736
rect 1661 3624 1667 3816
rect 1693 3724 1699 3796
rect 1709 3724 1715 3836
rect 1805 3824 1811 3896
rect 1853 3784 1859 3896
rect 1869 3864 1875 3876
rect 1901 3844 1907 4136
rect 2013 4024 2019 4116
rect 2013 3924 2019 3936
rect 1997 3904 2003 3916
rect 1949 3844 1955 3876
rect 1965 3864 1971 3896
rect 1741 3724 1747 3736
rect 1757 3724 1763 3736
rect 1613 3484 1619 3496
rect 1629 3484 1635 3536
rect 1661 3504 1667 3616
rect 1693 3484 1699 3556
rect 1741 3524 1747 3576
rect 1757 3504 1763 3716
rect 1869 3704 1875 3776
rect 1965 3764 1971 3776
rect 1933 3744 1939 3756
rect 2045 3724 2051 4016
rect 2093 3904 2099 4156
rect 2125 4144 2131 4196
rect 2205 4144 2211 4256
rect 2237 4124 2243 4236
rect 2285 4184 2291 4297
rect 2317 4284 2323 4376
rect 2349 4304 2355 4316
rect 2317 4104 2323 4276
rect 2445 4264 2451 4556
rect 2477 4443 2483 4536
rect 2605 4524 2611 4696
rect 2813 4684 2819 4816
rect 2632 4606 2638 4614
rect 2646 4606 2652 4614
rect 2660 4606 2666 4614
rect 2674 4606 2680 4614
rect 2717 4524 2723 4676
rect 2813 4604 2819 4676
rect 2909 4524 2915 4916
rect 2925 4784 2931 4936
rect 2941 4664 2947 4916
rect 3021 4844 3027 4896
rect 3037 4784 3043 4936
rect 3117 4704 3123 4936
rect 3453 4924 3459 4936
rect 3629 4924 3635 4956
rect 4029 4924 4035 4956
rect 3725 4862 3731 4900
rect 3261 4704 3267 4736
rect 2989 4664 2995 4696
rect 2925 4564 2931 4636
rect 2541 4462 2547 4500
rect 2477 4437 2499 4443
rect 2349 4144 2355 4256
rect 2365 4164 2371 4236
rect 2381 4144 2387 4256
rect 2445 4224 2451 4256
rect 2189 4062 2195 4100
rect 2317 3923 2323 4096
rect 2301 3917 2323 3923
rect 2109 3884 2115 3896
rect 2205 3884 2211 3916
rect 2301 3884 2307 3917
rect 2333 3904 2339 3936
rect 2349 3924 2355 4136
rect 2045 3704 2051 3716
rect 1837 3644 1843 3696
rect 1565 3344 1571 3476
rect 1597 3424 1603 3476
rect 1581 3384 1587 3416
rect 1597 3324 1603 3336
rect 1629 3324 1635 3456
rect 1837 3444 1843 3476
rect 1869 3464 1875 3696
rect 1869 3403 1875 3456
rect 1853 3397 1875 3403
rect 1677 3364 1683 3376
rect 1853 3364 1859 3397
rect 1405 3104 1411 3316
rect 1677 3304 1683 3356
rect 1885 3344 1891 3416
rect 2045 3384 2051 3556
rect 2061 3484 2067 3756
rect 2125 3604 2131 3636
rect 2173 3524 2179 3836
rect 2253 3784 2259 3816
rect 2205 3664 2211 3716
rect 2205 3504 2211 3656
rect 2221 3524 2227 3716
rect 2212 3497 2236 3503
rect 2237 3464 2243 3496
rect 2244 3457 2259 3463
rect 1981 3304 1987 3316
rect 1453 3184 1459 3236
rect 1549 3184 1555 3276
rect 1597 3184 1603 3296
rect 1949 3262 1955 3300
rect 1357 3064 1363 3096
rect 1565 3084 1571 3176
rect 1277 3024 1283 3056
rect 1341 2964 1347 3016
rect 1469 2984 1475 3036
rect 1197 2784 1203 2856
rect 1213 2844 1219 2896
rect 1341 2864 1347 2956
rect 1421 2924 1427 2956
rect 1517 2904 1523 3076
rect 1549 2903 1555 3076
rect 1540 2897 1555 2903
rect 1325 2784 1331 2836
rect 1373 2724 1379 2736
rect 525 2324 531 2376
rect 653 2304 659 2316
rect 765 2304 771 2456
rect 781 2324 787 2516
rect 797 2444 803 2496
rect 829 2384 835 2536
rect 1149 2462 1155 2500
rect 781 2304 787 2316
rect 845 2304 851 2436
rect 1112 2406 1118 2414
rect 1126 2406 1132 2414
rect 1140 2406 1146 2414
rect 1154 2406 1160 2414
rect 909 2324 915 2376
rect 525 2244 531 2296
rect 621 2184 627 2256
rect 589 2144 595 2156
rect 477 1864 483 2036
rect 509 1904 515 1916
rect 557 1884 563 1896
rect 141 1624 147 1716
rect 68 1497 83 1503
rect 61 1124 67 1496
rect 77 1324 83 1376
rect 13 984 19 1036
rect 13 904 19 916
rect 29 304 35 1116
rect 61 1044 67 1094
rect 93 1023 99 1616
rect 285 1504 291 1576
rect 333 1524 339 1676
rect 125 1104 131 1316
rect 221 1124 227 1496
rect 317 1484 323 1496
rect 237 1343 243 1476
rect 253 1363 259 1436
rect 253 1357 275 1363
rect 269 1344 275 1357
rect 317 1344 323 1456
rect 349 1344 355 1476
rect 381 1364 387 1756
rect 413 1643 419 1718
rect 397 1637 419 1643
rect 397 1584 403 1637
rect 413 1524 419 1616
rect 413 1504 419 1516
rect 397 1484 403 1496
rect 413 1464 419 1476
rect 237 1337 252 1343
rect 269 1324 275 1336
rect 381 1324 387 1356
rect 253 1104 259 1116
rect 285 1104 291 1236
rect 301 1184 307 1316
rect 365 1104 371 1116
rect 77 1017 99 1023
rect 61 684 67 936
rect 61 564 67 656
rect 45 324 51 376
rect 77 304 83 1017
rect 93 924 99 936
rect 157 924 163 1096
rect 253 1084 259 1096
rect 141 904 147 916
rect 189 903 195 1036
rect 221 964 227 1036
rect 221 944 227 956
rect 180 897 195 903
rect 189 724 195 736
rect 205 704 211 916
rect 93 664 99 696
rect 221 683 227 936
rect 269 924 275 976
rect 317 924 323 996
rect 237 884 243 896
rect 333 704 339 1096
rect 349 1064 355 1096
rect 349 984 355 1056
rect 381 984 387 1276
rect 429 1084 435 1096
rect 365 944 371 956
rect 413 924 419 1076
rect 429 1024 435 1076
rect 429 944 435 976
rect 356 897 371 903
rect 349 704 355 716
rect 212 677 227 683
rect 365 683 371 897
rect 381 724 387 836
rect 349 677 371 683
rect 205 644 211 676
rect 93 524 99 536
rect 125 444 131 516
rect 189 504 195 576
rect 205 544 211 636
rect 221 524 227 556
rect 301 524 307 556
rect 317 544 323 676
rect 349 584 355 677
rect 397 584 403 876
rect 413 844 419 896
rect 445 703 451 1556
rect 525 1524 531 1776
rect 557 1704 563 1876
rect 573 1784 579 1936
rect 621 1864 627 2036
rect 637 1984 643 2296
rect 701 2284 707 2296
rect 701 2124 707 2236
rect 733 2204 739 2236
rect 781 2164 787 2176
rect 813 2144 819 2196
rect 685 1944 691 2036
rect 797 1924 803 1936
rect 733 1904 739 1916
rect 765 1904 771 1916
rect 829 1904 835 1916
rect 589 1824 595 1856
rect 637 1844 643 1896
rect 877 1884 883 2176
rect 909 2124 915 2296
rect 1005 2284 1011 2316
rect 1181 2304 1187 2516
rect 1197 2384 1203 2556
rect 1037 2244 1043 2256
rect 1197 2184 1203 2256
rect 1085 2144 1091 2156
rect 1245 2144 1251 2596
rect 1293 2584 1299 2636
rect 1309 2604 1315 2676
rect 1533 2664 1539 2856
rect 1549 2804 1555 2897
rect 1565 2764 1571 2876
rect 1581 2784 1587 3056
rect 1613 2924 1619 3096
rect 1629 3084 1635 3236
rect 1949 3120 1955 3158
rect 1981 3104 1987 3296
rect 2061 3124 2067 3396
rect 2205 3344 2211 3456
rect 1773 3064 1779 3096
rect 1629 3044 1635 3056
rect 1629 3023 1635 3036
rect 1629 3017 1651 3023
rect 1629 2944 1635 2996
rect 1613 2844 1619 2916
rect 1629 2720 1635 2758
rect 1645 2704 1651 3017
rect 1709 2964 1715 3056
rect 1709 2924 1715 2956
rect 1773 2944 1779 3036
rect 1805 2964 1811 3016
rect 1805 2904 1811 2936
rect 1677 2844 1683 2896
rect 1709 2724 1715 2796
rect 1789 2704 1795 2836
rect 1805 2684 1811 2896
rect 1812 2677 1827 2683
rect 1277 2284 1283 2296
rect 1341 2264 1347 2656
rect 1421 2544 1427 2596
rect 1821 2564 1827 2677
rect 1837 2604 1843 2636
rect 1693 2544 1699 2556
rect 1373 2304 1379 2416
rect 1405 2384 1411 2536
rect 1533 2404 1539 2436
rect 1565 2404 1571 2496
rect 1341 2204 1347 2236
rect 1357 2224 1363 2276
rect 1389 2144 1395 2196
rect 1485 2124 1491 2296
rect 1565 2264 1571 2396
rect 1597 2324 1603 2536
rect 1661 2503 1667 2516
rect 1661 2497 1683 2503
rect 1677 2424 1683 2497
rect 1677 2384 1683 2416
rect 1661 2320 1667 2358
rect 1677 2304 1683 2336
rect 1757 2284 1763 2436
rect 1565 2244 1571 2256
rect 1565 2164 1571 2236
rect 909 2044 915 2096
rect 1053 1944 1059 1956
rect 596 1817 611 1823
rect 605 1744 611 1817
rect 637 1764 643 1836
rect 653 1744 659 1876
rect 925 1864 931 1876
rect 701 1724 707 1756
rect 621 1704 627 1716
rect 541 1624 547 1636
rect 733 1564 739 1836
rect 797 1784 803 1836
rect 925 1764 931 1856
rect 749 1704 755 1756
rect 797 1644 803 1696
rect 493 1504 499 1516
rect 525 1504 531 1516
rect 589 1504 595 1516
rect 797 1504 803 1556
rect 493 1384 499 1496
rect 509 1404 515 1496
rect 509 1304 515 1376
rect 525 1344 531 1416
rect 541 1344 547 1436
rect 605 1364 611 1496
rect 669 1484 675 1496
rect 621 1464 627 1476
rect 461 1184 467 1196
rect 477 1084 483 1276
rect 525 1204 531 1336
rect 541 1324 547 1336
rect 589 1324 595 1336
rect 557 1104 563 1116
rect 605 1104 611 1356
rect 621 1343 627 1456
rect 717 1444 723 1496
rect 733 1424 739 1476
rect 749 1464 755 1476
rect 621 1337 636 1343
rect 669 1324 675 1376
rect 685 1104 691 1396
rect 717 1324 723 1376
rect 749 1344 755 1456
rect 717 1304 723 1316
rect 733 1283 739 1316
rect 717 1277 739 1283
rect 717 1104 723 1277
rect 749 1263 755 1316
rect 765 1304 771 1356
rect 733 1257 755 1263
rect 733 1184 739 1257
rect 765 1124 771 1236
rect 781 1104 787 1136
rect 461 984 467 1036
rect 477 904 483 956
rect 525 924 531 976
rect 509 704 515 856
rect 436 697 451 703
rect 413 544 419 556
rect 445 544 451 697
rect 29 163 35 296
rect 20 157 35 163
rect 77 124 83 296
rect 173 264 179 436
rect 333 384 339 476
rect 333 324 339 376
rect 381 264 387 536
rect 445 524 451 536
rect 493 524 499 576
rect 509 524 515 596
rect 525 544 531 636
rect 541 564 547 916
rect 573 864 579 916
rect 557 704 563 836
rect 589 704 595 856
rect 493 504 499 516
rect 413 344 419 476
rect 173 164 179 256
rect 109 44 115 100
rect 365 -23 371 256
rect 381 164 387 256
rect 461 184 467 276
rect 493 184 499 336
rect 509 304 515 496
rect 429 157 444 163
rect 397 -17 403 36
rect 429 -17 435 157
rect 509 144 515 296
rect 525 284 531 536
rect 573 504 579 616
rect 589 604 595 696
rect 637 684 643 936
rect 653 924 659 956
rect 669 704 675 1096
rect 685 924 691 1096
rect 701 1084 707 1096
rect 781 1064 787 1096
rect 797 1064 803 1496
rect 813 1424 819 1476
rect 829 1444 835 1496
rect 836 1437 851 1443
rect 845 1324 851 1437
rect 861 1344 867 1416
rect 877 1364 883 1616
rect 909 1584 915 1636
rect 1037 1524 1043 1836
rect 909 1484 915 1496
rect 1069 1484 1075 2036
rect 1112 2006 1118 2014
rect 1126 2006 1132 2014
rect 1140 2006 1146 2014
rect 1154 2006 1160 2014
rect 1181 1904 1187 2076
rect 1453 2062 1459 2100
rect 1501 1904 1507 2156
rect 1149 1644 1155 1836
rect 1181 1764 1187 1776
rect 1197 1724 1203 1876
rect 1229 1864 1235 1876
rect 1309 1784 1315 1896
rect 1501 1884 1507 1896
rect 1421 1864 1427 1876
rect 1229 1724 1235 1736
rect 1341 1724 1347 1756
rect 1245 1704 1251 1716
rect 1229 1697 1244 1703
rect 1112 1606 1118 1614
rect 1126 1606 1132 1614
rect 1140 1606 1146 1614
rect 1154 1606 1160 1614
rect 1229 1584 1235 1697
rect 1357 1703 1363 1736
rect 1373 1724 1379 1736
rect 1389 1724 1395 1836
rect 1357 1697 1379 1703
rect 1197 1504 1203 1516
rect 925 1464 931 1476
rect 1181 1464 1187 1496
rect 813 1144 819 1296
rect 877 1104 883 1116
rect 957 1104 963 1236
rect 973 1183 979 1316
rect 1005 1304 1011 1456
rect 1021 1244 1027 1316
rect 973 1177 988 1183
rect 701 924 707 1056
rect 797 1004 803 1036
rect 717 964 723 976
rect 877 944 883 1076
rect 989 1024 995 1156
rect 1005 1024 1011 1076
rect 829 884 835 916
rect 861 784 867 836
rect 877 824 883 936
rect 941 924 947 1016
rect 973 884 979 936
rect 1021 924 1027 1056
rect 1037 924 1043 1276
rect 1053 1124 1059 1416
rect 1085 1344 1091 1356
rect 1197 1343 1203 1496
rect 1213 1464 1219 1476
rect 1188 1337 1203 1343
rect 1085 1317 1100 1323
rect 1069 1124 1075 1176
rect 1069 1104 1075 1116
rect 1085 983 1091 1317
rect 1112 1206 1118 1214
rect 1126 1206 1132 1214
rect 1140 1206 1146 1214
rect 1154 1206 1160 1214
rect 1117 1084 1123 1116
rect 1149 1104 1155 1116
rect 1181 1104 1187 1176
rect 1213 1144 1219 1296
rect 1229 1184 1235 1576
rect 1245 1504 1251 1636
rect 1277 1544 1283 1636
rect 1277 1504 1283 1536
rect 1309 1504 1315 1696
rect 1373 1584 1379 1697
rect 1389 1584 1395 1716
rect 1437 1644 1443 1716
rect 1533 1704 1539 1896
rect 1549 1724 1555 1796
rect 1581 1764 1587 2216
rect 1645 1884 1651 1896
rect 1613 1764 1619 1836
rect 1581 1744 1587 1756
rect 1517 1684 1523 1696
rect 1325 1524 1331 1576
rect 1277 1424 1283 1476
rect 1245 1144 1251 1276
rect 1261 1184 1267 1236
rect 1245 1084 1251 1096
rect 1213 984 1219 1016
rect 1085 977 1100 983
rect 1101 924 1107 976
rect 1037 884 1043 916
rect 1117 904 1123 936
rect 1181 924 1187 956
rect 1229 904 1235 1076
rect 1261 924 1267 1036
rect 1277 1004 1283 1076
rect 733 702 739 716
rect 621 524 627 636
rect 637 544 643 676
rect 653 624 659 696
rect 669 644 675 696
rect 701 564 707 676
rect 829 584 835 616
rect 861 584 867 756
rect 909 684 915 836
rect 877 624 883 656
rect 893 624 899 636
rect 845 544 851 576
rect 925 544 931 876
rect 1293 864 1299 1456
rect 1325 1363 1331 1516
rect 1341 1504 1347 1556
rect 1421 1504 1427 1596
rect 1389 1364 1395 1376
rect 1316 1357 1331 1363
rect 1325 1264 1331 1296
rect 1341 1264 1347 1316
rect 1341 1124 1347 1236
rect 1309 984 1315 1096
rect 1357 924 1363 1276
rect 1373 1044 1379 1096
rect 1405 1083 1411 1496
rect 1469 1484 1475 1496
rect 1485 1464 1491 1496
rect 1501 1484 1507 1636
rect 1549 1604 1555 1676
rect 1549 1484 1555 1496
rect 1565 1464 1571 1516
rect 1597 1504 1603 1536
rect 1517 1324 1523 1436
rect 1533 1344 1539 1416
rect 1549 1344 1555 1356
rect 1421 1104 1427 1236
rect 1437 1204 1443 1316
rect 1469 1284 1475 1296
rect 1485 1244 1491 1296
rect 1501 1124 1507 1316
rect 1581 1304 1587 1476
rect 1597 1444 1603 1496
rect 1613 1484 1619 1596
rect 1629 1564 1635 1736
rect 1645 1484 1651 1876
rect 1693 1824 1699 1896
rect 1709 1864 1715 2156
rect 1741 2144 1747 2236
rect 1789 2223 1795 2516
rect 1805 2404 1811 2516
rect 1853 2423 1859 2796
rect 1885 2704 1891 3056
rect 1901 2784 1907 2976
rect 1997 2944 2003 2996
rect 2029 2944 2035 3076
rect 2077 3064 2083 3316
rect 2093 3104 2099 3316
rect 2157 3284 2163 3296
rect 2109 3144 2115 3156
rect 2157 3104 2163 3256
rect 2205 3184 2211 3336
rect 2221 3104 2227 3396
rect 2253 3324 2259 3457
rect 2269 3404 2275 3716
rect 2285 3584 2291 3816
rect 2301 3764 2307 3876
rect 2317 3844 2323 3896
rect 2365 3844 2371 4136
rect 2381 4124 2387 4136
rect 2381 3904 2387 3916
rect 2413 3904 2419 4096
rect 2461 3984 2467 4276
rect 2477 4144 2483 4336
rect 2493 4184 2499 4437
rect 2605 4304 2611 4516
rect 2733 4444 2739 4500
rect 2669 4320 2675 4358
rect 2797 4344 2803 4516
rect 2813 4384 2819 4436
rect 2632 4206 2638 4214
rect 2646 4206 2652 4214
rect 2660 4206 2666 4214
rect 2674 4206 2680 4214
rect 2573 4124 2579 4156
rect 2429 3904 2435 3936
rect 2509 3904 2515 3936
rect 2413 3824 2419 3896
rect 2477 3884 2483 3896
rect 2509 3804 2515 3896
rect 2525 3864 2531 4096
rect 2685 4064 2691 4096
rect 2701 4063 2707 4296
rect 2797 4204 2803 4336
rect 2813 4204 2819 4256
rect 2861 4204 2867 4236
rect 2813 4164 2819 4196
rect 2781 4144 2787 4156
rect 2781 4064 2787 4116
rect 2692 4057 2707 4063
rect 2541 3984 2547 4056
rect 2909 4024 2915 4516
rect 2957 4304 2963 4656
rect 3005 4564 3011 4696
rect 3101 4684 3107 4696
rect 3053 4564 3059 4676
rect 2989 4324 2995 4436
rect 3005 4384 3011 4496
rect 3069 4464 3075 4656
rect 3085 4384 3091 4536
rect 3060 4317 3075 4323
rect 2989 4264 2995 4276
rect 2749 3984 2755 3996
rect 2717 3904 2723 3956
rect 2781 3904 2787 3976
rect 2845 3904 2851 4016
rect 2861 3920 2867 3958
rect 2541 3784 2547 3836
rect 2573 3824 2579 3876
rect 2632 3806 2638 3814
rect 2646 3806 2652 3814
rect 2660 3806 2666 3814
rect 2674 3806 2680 3814
rect 2541 3764 2547 3776
rect 2509 3744 2515 3756
rect 2413 3704 2419 3716
rect 2333 3684 2339 3696
rect 2285 3544 2291 3576
rect 2285 3364 2291 3516
rect 2301 3484 2307 3636
rect 2397 3524 2403 3636
rect 2301 3364 2307 3476
rect 2285 3344 2291 3356
rect 2397 3343 2403 3516
rect 2413 3504 2419 3696
rect 2445 3662 2451 3700
rect 2477 3520 2483 3558
rect 2541 3504 2547 3756
rect 2829 3744 2835 3756
rect 2845 3744 2851 3896
rect 2925 3884 2931 4256
rect 3037 4164 3043 4316
rect 3005 4004 3011 4096
rect 3053 3944 3059 4296
rect 3069 4264 3075 4317
rect 3085 4244 3091 4296
rect 3101 4184 3107 4656
rect 3149 4544 3155 4656
rect 3165 4584 3171 4696
rect 3277 4684 3283 4696
rect 3325 4684 3331 4816
rect 3197 4624 3203 4676
rect 3149 4484 3155 4516
rect 3181 4424 3187 4556
rect 3229 4364 3235 4496
rect 3197 4304 3203 4336
rect 3133 4264 3139 4276
rect 2957 3844 2963 3856
rect 2909 3744 2915 3816
rect 2781 3624 2787 3676
rect 2813 3664 2819 3716
rect 2909 3564 2915 3736
rect 2925 3584 2931 3836
rect 2573 3464 2579 3496
rect 2813 3484 2819 3556
rect 2632 3406 2638 3414
rect 2646 3406 2652 3414
rect 2660 3406 2666 3414
rect 2674 3406 2680 3414
rect 2381 3337 2403 3343
rect 2253 3264 2259 3316
rect 2253 3204 2259 3256
rect 2349 3184 2355 3316
rect 2157 3044 2163 3096
rect 2173 3004 2179 3076
rect 2269 3044 2275 3076
rect 2189 2964 2195 3036
rect 2221 2964 2227 3016
rect 2013 2844 2019 2916
rect 2189 2904 2195 2916
rect 2045 2824 2051 2896
rect 2125 2862 2131 2900
rect 2237 2784 2243 2836
rect 2301 2784 2307 3136
rect 2381 3124 2387 3337
rect 2477 3204 2483 3356
rect 2445 3104 2451 3196
rect 2413 3064 2419 3076
rect 2429 3044 2435 3076
rect 2461 3064 2467 3076
rect 1901 2704 1907 2776
rect 2189 2724 2195 2776
rect 2317 2704 2323 3036
rect 2477 3024 2483 3196
rect 2573 3104 2579 3296
rect 2605 3244 2611 3296
rect 2765 3262 2771 3300
rect 2605 3120 2611 3158
rect 2669 3084 2675 3096
rect 2701 3064 2707 3196
rect 2701 3024 2707 3056
rect 2632 3006 2638 3014
rect 2646 3006 2652 3014
rect 2660 3006 2666 3014
rect 2674 3006 2680 3014
rect 2477 2904 2483 2976
rect 2749 2964 2755 3016
rect 1869 2524 1875 2576
rect 1837 2417 1859 2423
rect 1837 2304 1843 2417
rect 1853 2304 1859 2396
rect 1789 2217 1811 2223
rect 1805 1964 1811 2217
rect 1837 2164 1843 2296
rect 1885 2264 1891 2696
rect 2093 2584 2099 2676
rect 2013 2504 2019 2556
rect 2189 2524 2195 2696
rect 2205 2564 2211 2616
rect 2237 2584 2243 2696
rect 2253 2584 2259 2616
rect 2285 2584 2291 2656
rect 2301 2624 2307 2636
rect 1917 2462 1923 2500
rect 2141 2320 2147 2358
rect 2173 2304 2179 2356
rect 2221 2304 2227 2436
rect 2269 2384 2275 2536
rect 2333 2524 2339 2736
rect 2381 2704 2387 2896
rect 2429 2844 2435 2856
rect 2429 2804 2435 2836
rect 2477 2784 2483 2896
rect 2653 2844 2659 2900
rect 2749 2784 2755 2956
rect 2829 2924 2835 3216
rect 2861 3204 2867 3356
rect 2941 3324 2947 3736
rect 2989 3484 2995 3756
rect 2973 3464 2979 3476
rect 2941 3224 2947 3316
rect 2989 3244 2995 3476
rect 2909 3184 2915 3216
rect 3005 3164 3011 3656
rect 3037 3524 3043 3836
rect 3053 3764 3059 3936
rect 3069 3764 3075 4156
rect 3085 3844 3091 4136
rect 3117 4084 3123 4096
rect 3133 4064 3139 4256
rect 3149 3964 3155 4256
rect 3181 4004 3187 4296
rect 3245 4284 3251 4676
rect 3309 4584 3315 4636
rect 3325 4524 3331 4536
rect 3261 4464 3267 4496
rect 3277 4484 3283 4516
rect 3293 4444 3299 4516
rect 3309 4497 3324 4503
rect 3309 4384 3315 4497
rect 3277 4324 3283 4336
rect 3197 4184 3203 4256
rect 3213 4164 3219 4216
rect 3229 4184 3235 4236
rect 3229 4084 3235 4096
rect 3133 3884 3139 3916
rect 3149 3904 3155 3916
rect 3181 3884 3187 3976
rect 3197 3884 3203 3956
rect 3213 3904 3219 3996
rect 3245 3924 3251 4276
rect 3261 4144 3267 4256
rect 3277 4163 3283 4316
rect 3293 4264 3299 4276
rect 3309 4184 3315 4356
rect 3277 4157 3292 4163
rect 3325 4163 3331 4276
rect 3341 4164 3347 4836
rect 3469 4824 3475 4836
rect 3437 4737 3491 4743
rect 3357 4704 3363 4716
rect 3437 4704 3443 4737
rect 3469 4704 3475 4716
rect 3485 4704 3491 4737
rect 3533 4704 3539 4716
rect 3357 4684 3363 4696
rect 3389 4644 3395 4696
rect 3469 4684 3475 4696
rect 3469 4664 3475 4676
rect 3357 4564 3363 4636
rect 3405 4584 3411 4656
rect 3389 4544 3395 4556
rect 3437 4544 3443 4636
rect 3501 4624 3507 4636
rect 3501 4604 3507 4616
rect 3357 4444 3363 4516
rect 3421 4444 3427 4516
rect 3405 4323 3411 4416
rect 3421 4344 3427 4376
rect 3405 4317 3427 4323
rect 3357 4297 3372 4303
rect 3357 4264 3363 4297
rect 3373 4264 3379 4276
rect 3405 4184 3411 4216
rect 3309 4157 3331 4163
rect 3261 4124 3267 4136
rect 3277 4124 3283 4136
rect 3261 3924 3267 3936
rect 3133 3784 3139 3836
rect 3069 3737 3084 3743
rect 3069 3584 3075 3737
rect 3101 3724 3107 3756
rect 3149 3743 3155 3836
rect 3197 3804 3203 3876
rect 3213 3764 3219 3896
rect 3245 3764 3251 3796
rect 3133 3737 3155 3743
rect 3037 3484 3043 3516
rect 3021 3303 3027 3436
rect 3021 3297 3036 3303
rect 2909 2984 2915 3056
rect 2941 2984 2947 3116
rect 2957 2924 2963 3136
rect 2973 3084 2979 3156
rect 2989 3084 2995 3136
rect 2589 2724 2595 2776
rect 2781 2704 2787 2816
rect 2493 2664 2499 2676
rect 2461 2604 2467 2656
rect 2413 2564 2419 2596
rect 2589 2564 2595 2616
rect 2301 2304 2307 2396
rect 2077 2284 2083 2296
rect 2285 2284 2291 2296
rect 1885 2224 1891 2236
rect 2045 2164 2051 2256
rect 2317 2184 2323 2316
rect 1837 2124 1843 2136
rect 1901 2124 1907 2136
rect 1837 2044 1843 2096
rect 1917 2044 1923 2096
rect 2125 2023 2131 2116
rect 2109 2017 2131 2023
rect 2029 1864 2035 1876
rect 1661 1744 1667 1756
rect 1661 1604 1667 1736
rect 1693 1724 1699 1756
rect 1741 1684 1747 1716
rect 1613 1424 1619 1476
rect 1629 1364 1635 1436
rect 1677 1384 1683 1416
rect 1405 1077 1427 1083
rect 1309 884 1315 916
rect 1325 864 1331 916
rect 1341 904 1347 916
rect 973 684 979 816
rect 1112 806 1118 814
rect 1126 806 1132 814
rect 1140 806 1146 814
rect 1154 806 1160 814
rect 1277 804 1283 836
rect 941 584 947 636
rect 669 384 675 536
rect 573 324 579 336
rect 589 304 595 316
rect 797 284 803 456
rect 637 204 643 236
rect 653 164 659 276
rect 685 144 691 196
rect 893 144 899 496
rect 909 384 915 416
rect 925 284 931 536
rect 941 524 947 556
rect 941 504 947 516
rect 941 324 947 436
rect 973 424 979 676
rect 1069 584 1075 676
rect 1133 644 1139 656
rect 1197 644 1203 716
rect 1229 684 1235 696
rect 1101 524 1107 596
rect 1117 524 1123 636
rect 1133 604 1139 636
rect 1133 564 1139 596
rect 1229 584 1235 636
rect 989 304 995 436
rect 1005 384 1011 516
rect 1181 424 1187 516
rect 1112 406 1118 414
rect 1126 406 1132 414
rect 1140 406 1146 414
rect 1154 406 1160 414
rect 1005 324 1011 376
rect 1037 304 1043 336
rect 1069 324 1075 356
rect 1197 344 1203 516
rect 1229 504 1235 556
rect 1245 544 1251 676
rect 1261 624 1267 676
rect 1309 584 1315 716
rect 1325 684 1331 716
rect 1245 503 1251 536
rect 1261 524 1267 556
rect 1341 523 1347 896
rect 1373 704 1379 956
rect 1389 884 1395 896
rect 1389 844 1395 876
rect 1421 784 1427 1077
rect 1437 1044 1443 1096
rect 1453 1024 1459 1076
rect 1453 944 1459 1016
rect 1485 984 1491 1116
rect 1437 924 1443 936
rect 1469 924 1475 936
rect 1460 917 1468 923
rect 1405 724 1411 756
rect 1421 724 1427 736
rect 1437 704 1443 816
rect 1453 744 1459 916
rect 1501 824 1507 956
rect 1565 904 1571 918
rect 1437 684 1443 696
rect 1485 584 1491 676
rect 1501 584 1507 696
rect 1549 684 1555 796
rect 1565 704 1571 736
rect 1332 517 1347 523
rect 1245 497 1267 503
rect 1229 302 1235 316
rect 973 264 979 296
rect 1117 264 1123 276
rect 909 164 915 236
rect 941 204 947 236
rect 1037 144 1043 196
rect 1245 164 1251 276
rect 1261 264 1267 497
rect 1245 144 1251 156
rect 445 124 451 136
rect 1277 126 1283 516
rect 1293 484 1299 496
rect 1341 304 1347 517
rect 1373 504 1379 516
rect 1357 484 1363 496
rect 1437 484 1443 516
rect 1405 184 1411 476
rect 1453 384 1459 496
rect 1469 384 1475 556
rect 1581 524 1587 1296
rect 1597 1284 1603 1296
rect 1597 724 1603 1276
rect 1629 1164 1635 1316
rect 1693 1184 1699 1236
rect 1629 784 1635 796
rect 1677 704 1683 1176
rect 1709 704 1715 1556
rect 1741 1504 1747 1676
rect 1773 1644 1779 1736
rect 1805 1704 1811 1836
rect 1885 1784 1891 1816
rect 2061 1764 2067 1816
rect 2093 1764 2099 1976
rect 2109 1924 2115 2017
rect 2125 1924 2131 1976
rect 2109 1904 2115 1916
rect 2125 1784 2131 1856
rect 1821 1684 1827 1696
rect 1837 1644 1843 1736
rect 1821 1464 1827 1536
rect 1869 1504 1875 1696
rect 1885 1584 1891 1716
rect 1853 1484 1859 1496
rect 1725 1304 1731 1336
rect 1725 1084 1731 1276
rect 1741 1264 1747 1316
rect 1757 1304 1763 1396
rect 1837 1344 1843 1436
rect 1869 1404 1875 1496
rect 1869 1344 1875 1356
rect 1933 1344 1939 1556
rect 1949 1544 1955 1716
rect 1981 1704 1987 1756
rect 2141 1744 2147 1896
rect 1965 1564 1971 1636
rect 2013 1504 2019 1516
rect 1949 1424 1955 1496
rect 1965 1364 1971 1496
rect 2045 1484 2051 1736
rect 2093 1724 2099 1736
rect 2157 1724 2163 2156
rect 2333 2124 2339 2276
rect 2349 2244 2355 2296
rect 2365 2284 2371 2316
rect 2397 2304 2403 2356
rect 2349 2144 2355 2216
rect 2365 2204 2371 2276
rect 2413 2264 2419 2556
rect 2445 2443 2451 2516
rect 2509 2462 2515 2500
rect 2429 2437 2451 2443
rect 2429 2344 2435 2437
rect 2605 2403 2611 2696
rect 2685 2684 2691 2696
rect 2717 2684 2723 2696
rect 2632 2606 2638 2614
rect 2646 2606 2652 2614
rect 2660 2606 2666 2614
rect 2674 2606 2680 2614
rect 2701 2544 2707 2656
rect 2685 2444 2691 2516
rect 2717 2404 2723 2496
rect 2605 2397 2627 2403
rect 2429 2283 2435 2336
rect 2445 2320 2451 2358
rect 2621 2304 2627 2397
rect 2429 2277 2451 2283
rect 2397 2164 2403 2196
rect 2429 2124 2435 2236
rect 2445 2144 2451 2277
rect 2509 2184 2515 2276
rect 2253 2117 2268 2123
rect 2189 2037 2204 2043
rect 2173 1784 2179 1796
rect 2189 1764 2195 2037
rect 2253 1904 2259 2117
rect 2541 2084 2547 2256
rect 2632 2206 2638 2214
rect 2646 2206 2652 2214
rect 2660 2206 2666 2214
rect 2674 2206 2680 2214
rect 2813 2204 2819 2276
rect 2829 2264 2835 2796
rect 2893 2784 2899 2896
rect 2973 2884 2979 2956
rect 3021 2923 3027 3236
rect 3053 3123 3059 3516
rect 3085 3503 3091 3716
rect 3133 3704 3139 3737
rect 3149 3683 3155 3716
rect 3165 3684 3171 3736
rect 3133 3677 3155 3683
rect 3076 3497 3091 3503
rect 3069 3324 3075 3496
rect 3085 3464 3091 3476
rect 3085 3324 3091 3396
rect 3044 3117 3059 3123
rect 3069 3064 3075 3096
rect 3085 3084 3091 3296
rect 3085 3024 3091 3076
rect 3012 2917 3027 2923
rect 2852 2717 2867 2723
rect 2861 2704 2867 2717
rect 2845 2624 2851 2696
rect 2877 2644 2883 2676
rect 2957 2604 2963 2836
rect 2973 2744 2979 2876
rect 3005 2804 3011 2916
rect 3069 2884 3075 2956
rect 3101 2923 3107 3596
rect 3133 3584 3139 3677
rect 3117 3544 3123 3556
rect 3149 3524 3155 3576
rect 3165 3504 3171 3536
rect 3197 3484 3203 3696
rect 3213 3504 3219 3516
rect 3229 3504 3235 3516
rect 3261 3484 3267 3616
rect 3117 3304 3123 3476
rect 3117 3144 3123 3296
rect 3133 3184 3139 3476
rect 3181 3424 3187 3476
rect 3197 3384 3203 3456
rect 3165 3344 3171 3356
rect 3181 3304 3187 3376
rect 3149 3144 3155 3156
rect 3181 3124 3187 3136
rect 3197 3124 3203 3336
rect 3213 3284 3219 3336
rect 3229 3324 3235 3436
rect 3245 3344 3251 3476
rect 3261 3404 3267 3476
rect 3277 3383 3283 3656
rect 3309 3584 3315 4157
rect 3325 4104 3331 4136
rect 3341 4064 3347 4116
rect 3341 3984 3347 3996
rect 3341 3904 3347 3936
rect 3389 3923 3395 4096
rect 3405 4064 3411 4116
rect 3380 3917 3395 3923
rect 3405 3904 3411 3996
rect 3357 3864 3363 3876
rect 3373 3824 3379 3836
rect 3421 3824 3427 4317
rect 3437 4284 3443 4536
rect 3453 4524 3459 4556
rect 3485 4524 3491 4576
rect 3453 4364 3459 4516
rect 3501 4503 3507 4536
rect 3517 4524 3523 4556
rect 3501 4497 3523 4503
rect 3453 4304 3459 4316
rect 3485 4304 3491 4356
rect 3485 4284 3491 4296
rect 3501 4284 3507 4416
rect 3517 4384 3523 4497
rect 3533 4283 3539 4656
rect 3581 4644 3587 4716
rect 3597 4684 3603 4816
rect 3549 4544 3555 4636
rect 3581 4524 3587 4636
rect 3597 4624 3603 4676
rect 3613 4564 3619 4676
rect 3549 4284 3555 4416
rect 3565 4324 3571 4516
rect 3597 4323 3603 4436
rect 3613 4343 3619 4556
rect 3645 4484 3651 4636
rect 3661 4524 3667 4536
rect 3629 4384 3635 4396
rect 3661 4384 3667 4436
rect 3693 4424 3699 4696
rect 3709 4664 3715 4676
rect 3709 4484 3715 4596
rect 3773 4584 3779 4736
rect 3805 4724 3811 4776
rect 4013 4704 4019 4836
rect 3933 4624 3939 4656
rect 3789 4524 3795 4536
rect 3741 4504 3747 4516
rect 3693 4384 3699 4416
rect 3613 4337 3635 4343
rect 3597 4317 3619 4323
rect 3565 4304 3571 4316
rect 3597 4284 3603 4296
rect 3613 4284 3619 4317
rect 3517 4277 3539 4283
rect 3437 4264 3443 4276
rect 3469 4264 3475 4276
rect 3437 4124 3443 4196
rect 3437 4084 3443 4116
rect 3453 3944 3459 4216
rect 3469 4164 3475 4216
rect 3485 4184 3491 4236
rect 3469 4024 3475 4136
rect 3437 3884 3443 3916
rect 3485 3904 3491 4156
rect 3501 4144 3507 4196
rect 3517 4163 3523 4277
rect 3533 4204 3539 4256
rect 3517 4157 3532 4163
rect 3517 4104 3523 4116
rect 3501 3964 3507 4016
rect 3469 3784 3475 3876
rect 3453 3777 3468 3783
rect 3341 3624 3347 3736
rect 3389 3724 3395 3776
rect 3357 3604 3363 3716
rect 3437 3664 3443 3696
rect 3453 3684 3459 3777
rect 3485 3684 3491 3896
rect 3501 3884 3507 3956
rect 3517 3904 3523 4076
rect 3549 4023 3555 4256
rect 3565 4124 3571 4236
rect 3581 4203 3587 4276
rect 3581 4197 3603 4203
rect 3581 4144 3587 4176
rect 3597 4103 3603 4197
rect 3613 4164 3619 4256
rect 3629 4184 3635 4337
rect 3661 4304 3667 4356
rect 3709 4344 3715 4476
rect 3732 4457 3747 4463
rect 3725 4384 3731 4436
rect 3741 4344 3747 4457
rect 3773 4324 3779 4496
rect 3821 4484 3827 4516
rect 3869 4504 3875 4616
rect 3661 4244 3667 4296
rect 3581 4097 3603 4103
rect 3581 4024 3587 4097
rect 3613 4024 3619 4096
rect 3629 4063 3635 4136
rect 3661 4084 3667 4116
rect 3629 4057 3651 4063
rect 3549 4017 3571 4023
rect 3517 3824 3523 3836
rect 3533 3724 3539 3756
rect 3549 3704 3555 3996
rect 3565 3884 3571 4017
rect 3581 3904 3587 3956
rect 3613 3943 3619 3956
rect 3629 3943 3635 4036
rect 3613 3937 3635 3943
rect 3613 3904 3619 3937
rect 3565 3764 3571 3876
rect 3581 3723 3587 3796
rect 3613 3764 3619 3896
rect 3629 3824 3635 3856
rect 3629 3784 3635 3796
rect 3613 3724 3619 3736
rect 3565 3717 3587 3723
rect 3565 3684 3571 3717
rect 3597 3683 3603 3716
rect 3581 3677 3603 3683
rect 3325 3544 3331 3596
rect 3421 3584 3427 3596
rect 3581 3584 3587 3677
rect 3437 3544 3443 3556
rect 3565 3544 3571 3556
rect 3380 3537 3411 3543
rect 3325 3504 3331 3536
rect 3405 3524 3411 3537
rect 3645 3523 3651 4057
rect 3661 3924 3667 4036
rect 3677 3804 3683 4296
rect 3709 4244 3715 4256
rect 3709 4124 3715 4196
rect 3725 4103 3731 4116
rect 3709 4097 3731 4103
rect 3709 4084 3715 4097
rect 3693 4063 3699 4076
rect 3693 4057 3708 4063
rect 3741 4044 3747 4316
rect 3757 4284 3763 4296
rect 3773 4223 3779 4316
rect 3789 4264 3795 4436
rect 3837 4404 3843 4476
rect 3757 4217 3779 4223
rect 3757 4124 3763 4217
rect 3789 4203 3795 4236
rect 3773 4197 3795 4203
rect 3773 4164 3779 4197
rect 3789 4124 3795 4176
rect 3805 4104 3811 4316
rect 3821 4304 3827 4356
rect 3869 4324 3875 4496
rect 3901 4484 3907 4596
rect 3885 4464 3891 4476
rect 3901 4344 3907 4436
rect 3837 4284 3843 4316
rect 3885 4304 3891 4316
rect 3901 4304 3907 4336
rect 3933 4304 3939 4596
rect 3981 4384 3987 4536
rect 3997 4324 4003 4456
rect 4013 4424 4019 4696
rect 4029 4564 4035 4916
rect 4061 4844 4067 4916
rect 4125 4862 4131 4900
rect 4152 4806 4158 4814
rect 4166 4806 4172 4814
rect 4180 4806 4186 4814
rect 4194 4806 4200 4814
rect 4221 4784 4227 4916
rect 4333 4784 4339 4936
rect 4269 4724 4275 4776
rect 4429 4744 4435 4896
rect 4269 4684 4275 4716
rect 4301 4704 4307 4716
rect 4717 4704 4723 4916
rect 4749 4844 4755 4896
rect 4749 4724 4755 4776
rect 4301 4684 4307 4696
rect 4237 4524 4243 4656
rect 4205 4462 4211 4500
rect 3837 4184 3843 4216
rect 3853 4204 3859 4236
rect 3837 4144 3843 4176
rect 3853 4124 3859 4196
rect 3901 4144 3907 4156
rect 3933 4144 3939 4296
rect 3949 4264 3955 4276
rect 3997 4164 4003 4176
rect 3949 4124 3955 4156
rect 4029 4124 4035 4136
rect 4061 4124 4067 4356
rect 4077 4304 4083 4416
rect 4152 4406 4158 4414
rect 4166 4406 4172 4414
rect 4180 4406 4186 4414
rect 4194 4406 4200 4414
rect 4269 4404 4275 4676
rect 4349 4644 4355 4696
rect 4317 4544 4323 4636
rect 4349 4604 4355 4636
rect 4365 4584 4371 4676
rect 4365 4464 4371 4496
rect 4381 4424 4387 4676
rect 4541 4664 4547 4696
rect 4749 4664 4755 4696
rect 4429 4544 4435 4636
rect 4621 4624 4627 4656
rect 4541 4564 4547 4616
rect 4765 4584 4771 4936
rect 4813 4564 4819 4836
rect 4509 4544 4515 4556
rect 4445 4462 4451 4500
rect 4381 4384 4387 4396
rect 4461 4384 4467 4416
rect 4125 4320 4131 4358
rect 4493 4304 4499 4316
rect 4509 4304 4515 4516
rect 4541 4443 4547 4556
rect 4797 4524 4803 4556
rect 4829 4543 4835 4836
rect 5005 4824 5011 4916
rect 4861 4720 4867 4758
rect 4845 4664 4851 4696
rect 4893 4564 4899 4616
rect 4925 4584 4931 4656
rect 4820 4537 4835 4543
rect 4525 4437 4547 4443
rect 4525 4384 4531 4437
rect 4685 4324 4691 4376
rect 4189 4223 4195 4276
rect 4173 4217 4195 4223
rect 4173 4184 4179 4217
rect 4221 4164 4227 4256
rect 4301 4224 4307 4296
rect 3789 4064 3795 4076
rect 3757 3984 3763 3996
rect 3741 3944 3747 3976
rect 3773 3944 3779 3996
rect 3821 3984 3827 4056
rect 3917 4044 3923 4116
rect 4093 4104 4099 4156
rect 4253 4124 4259 4216
rect 4413 4204 4419 4236
rect 4493 4204 4499 4296
rect 4365 4144 4371 4196
rect 3933 4084 3939 4096
rect 3965 4064 3971 4076
rect 3693 3924 3699 3936
rect 3741 3924 3747 3936
rect 3757 3904 3763 3916
rect 3661 3704 3667 3716
rect 3693 3664 3699 3896
rect 3773 3784 3779 3936
rect 3885 3924 3891 3976
rect 3837 3884 3843 3916
rect 3757 3724 3763 3736
rect 3709 3704 3715 3716
rect 3725 3624 3731 3696
rect 3773 3604 3779 3716
rect 3805 3704 3811 3876
rect 3869 3724 3875 3916
rect 3805 3664 3811 3676
rect 3821 3664 3827 3716
rect 3885 3684 3891 3696
rect 3805 3584 3811 3596
rect 3620 3517 3635 3523
rect 3645 3517 3660 3523
rect 3389 3504 3395 3516
rect 3453 3497 3468 3503
rect 3293 3464 3299 3476
rect 3309 3444 3315 3496
rect 3341 3484 3347 3496
rect 3341 3443 3347 3476
rect 3421 3464 3427 3496
rect 3341 3437 3363 3443
rect 3261 3377 3283 3383
rect 3133 3103 3139 3116
rect 3165 3104 3171 3116
rect 3124 3097 3139 3103
rect 3229 3084 3235 3296
rect 3261 3123 3267 3377
rect 3277 3324 3283 3336
rect 3293 3324 3299 3416
rect 3357 3324 3363 3437
rect 3373 3324 3379 3396
rect 3389 3324 3395 3416
rect 3405 3364 3411 3456
rect 3405 3344 3411 3356
rect 3437 3344 3443 3496
rect 3453 3404 3459 3497
rect 3597 3503 3603 3516
rect 3597 3497 3612 3503
rect 3469 3344 3475 3476
rect 3485 3384 3491 3456
rect 3517 3364 3523 3476
rect 3581 3444 3587 3496
rect 3517 3344 3523 3356
rect 3261 3117 3276 3123
rect 3092 2917 3107 2923
rect 3133 2884 3139 2956
rect 3149 2924 3155 2936
rect 3085 2824 3091 2836
rect 3149 2804 3155 2836
rect 3005 2720 3011 2758
rect 3101 2704 3107 2776
rect 2973 2604 2979 2696
rect 3069 2664 3075 2676
rect 3101 2664 3107 2696
rect 2909 2504 2915 2556
rect 2941 2544 2947 2556
rect 3021 2524 3027 2596
rect 3005 2462 3011 2500
rect 2845 2384 2851 2416
rect 2909 2344 2915 2456
rect 2957 2324 2963 2416
rect 3101 2324 3107 2436
rect 2877 2284 2883 2296
rect 2909 2284 2915 2296
rect 2941 2264 2947 2316
rect 3133 2304 3139 2616
rect 3181 2484 3187 2956
rect 3229 2944 3235 3076
rect 3245 3064 3251 3096
rect 3277 2984 3283 3116
rect 3245 2923 3251 2976
rect 3229 2917 3251 2923
rect 3229 2904 3235 2917
rect 3293 2904 3299 3316
rect 3309 3204 3315 3316
rect 3373 3304 3379 3316
rect 3437 3303 3443 3336
rect 3549 3324 3555 3376
rect 3604 3357 3619 3363
rect 3613 3344 3619 3357
rect 3565 3324 3571 3336
rect 3629 3324 3635 3517
rect 3661 3484 3667 3516
rect 3645 3464 3651 3476
rect 3645 3384 3651 3396
rect 3677 3344 3683 3476
rect 3693 3444 3699 3476
rect 3725 3364 3731 3476
rect 3741 3404 3747 3536
rect 3725 3344 3731 3356
rect 3741 3324 3747 3396
rect 3773 3384 3779 3496
rect 3789 3384 3795 3516
rect 3805 3384 3811 3496
rect 3437 3297 3459 3303
rect 3341 3144 3347 3156
rect 3213 2864 3219 2896
rect 3165 2324 3171 2436
rect 2941 2164 2947 2236
rect 2685 2044 2691 2096
rect 2525 2004 2531 2036
rect 2701 2004 2707 2116
rect 2781 2104 2787 2136
rect 2813 2004 2819 2156
rect 2957 2144 2963 2236
rect 2989 2144 2995 2156
rect 3005 2064 3011 2276
rect 3021 2244 3027 2256
rect 3053 2144 3059 2156
rect 3037 2124 3043 2136
rect 2269 1904 2275 1956
rect 2381 1904 2387 1916
rect 2557 1904 2563 1996
rect 2589 1924 2595 1976
rect 2781 1904 2787 1996
rect 3037 1984 3043 2056
rect 2989 1924 2995 1976
rect 2253 1884 2259 1896
rect 2205 1864 2211 1876
rect 2493 1864 2499 1876
rect 2461 1844 2467 1856
rect 2605 1783 2611 1876
rect 2632 1806 2638 1814
rect 2646 1806 2652 1814
rect 2660 1806 2666 1814
rect 2674 1806 2680 1814
rect 2701 1784 2707 1836
rect 2861 1823 2867 1856
rect 2861 1817 2883 1823
rect 2605 1777 2620 1783
rect 2589 1764 2595 1776
rect 2877 1764 2883 1817
rect 2061 1544 2067 1716
rect 2061 1504 2067 1536
rect 2093 1524 2099 1536
rect 2157 1524 2163 1636
rect 2093 1504 2099 1516
rect 2141 1484 2147 1496
rect 2157 1484 2163 1516
rect 1741 1244 1747 1256
rect 1725 944 1731 1076
rect 1741 984 1747 1116
rect 1757 1104 1763 1196
rect 1757 964 1763 1096
rect 1773 984 1779 1156
rect 1805 1103 1811 1316
rect 1933 1303 1939 1316
rect 1924 1297 1939 1303
rect 1789 1097 1811 1103
rect 1789 984 1795 1097
rect 1805 1064 1811 1076
rect 1725 764 1731 936
rect 1741 884 1747 896
rect 1757 824 1763 956
rect 1757 724 1763 756
rect 1725 684 1731 716
rect 1613 664 1619 676
rect 1677 584 1683 676
rect 1565 504 1571 516
rect 1444 317 1459 323
rect 1421 264 1427 276
rect 1421 124 1427 256
rect 1453 204 1459 317
rect 1485 304 1491 316
rect 1533 304 1539 436
rect 1565 324 1571 496
rect 1597 484 1603 556
rect 1645 524 1651 576
rect 1709 524 1715 656
rect 1757 564 1763 716
rect 1789 704 1795 976
rect 1837 884 1843 1296
rect 1997 1284 2003 1296
rect 1853 1124 1859 1276
rect 1901 1124 1907 1236
rect 1997 1184 2003 1196
rect 1933 1084 1939 1096
rect 1949 1064 1955 1076
rect 2029 1064 2035 1096
rect 1853 1057 1868 1063
rect 1821 683 1827 856
rect 1853 743 1859 1057
rect 1933 924 1939 956
rect 2045 944 2051 1036
rect 1869 784 1875 816
rect 1837 737 1859 743
rect 1837 724 1843 737
rect 1933 724 1939 916
rect 2029 862 2035 900
rect 1837 704 1843 716
rect 1853 684 1859 716
rect 1933 684 1939 696
rect 1821 677 1843 683
rect 1805 664 1811 676
rect 1453 164 1459 196
rect 1469 164 1475 276
rect 1629 184 1635 516
rect 1677 484 1683 496
rect 1693 384 1699 496
rect 1757 484 1763 556
rect 1709 464 1715 476
rect 1757 384 1763 416
rect 1773 304 1779 636
rect 1821 524 1827 636
rect 1837 384 1843 677
rect 2061 664 2067 916
rect 1965 544 1971 636
rect 2093 524 2099 1396
rect 2189 1364 2195 1456
rect 2205 1444 2211 1676
rect 2109 964 2115 1076
rect 2125 1064 2131 1216
rect 2221 1204 2227 1336
rect 2301 1324 2307 1716
rect 2381 1624 2387 1756
rect 2333 1484 2339 1616
rect 2413 1584 2419 1736
rect 2557 1724 2563 1736
rect 2653 1724 2659 1756
rect 2509 1644 2515 1696
rect 2461 1504 2467 1516
rect 2333 1464 2339 1476
rect 2365 1404 2371 1496
rect 2429 1484 2435 1496
rect 2493 1464 2499 1476
rect 2525 1444 2531 1496
rect 2397 1324 2403 1416
rect 2285 1244 2291 1300
rect 2237 1184 2243 1196
rect 2180 1117 2195 1123
rect 2125 943 2131 1056
rect 2141 984 2147 1116
rect 2189 1104 2195 1117
rect 2221 1104 2227 1116
rect 2301 1083 2307 1236
rect 2381 1223 2387 1276
rect 2365 1217 2387 1223
rect 2365 1184 2371 1217
rect 2381 1124 2387 1176
rect 2397 1144 2403 1316
rect 2413 1304 2419 1436
rect 2429 1384 2435 1396
rect 2557 1384 2563 1696
rect 2749 1524 2755 1716
rect 2781 1662 2787 1700
rect 2653 1444 2659 1476
rect 2632 1406 2638 1414
rect 2646 1406 2652 1414
rect 2660 1406 2666 1414
rect 2674 1406 2680 1414
rect 2461 1344 2467 1356
rect 2493 1324 2499 1356
rect 2413 1244 2419 1296
rect 2445 1244 2451 1276
rect 2381 1084 2387 1116
rect 2397 1104 2403 1116
rect 2413 1104 2419 1196
rect 2429 1184 2435 1236
rect 2445 1124 2451 1236
rect 2493 1204 2499 1316
rect 2525 1104 2531 1196
rect 2605 1164 2611 1296
rect 2292 1077 2307 1083
rect 2173 1064 2179 1076
rect 2260 1057 2275 1063
rect 2116 937 2140 943
rect 2173 924 2179 956
rect 2205 904 2211 1056
rect 2237 984 2243 996
rect 2253 944 2259 1016
rect 2269 924 2275 1057
rect 2317 1044 2323 1056
rect 2333 1024 2339 1076
rect 2301 984 2307 1016
rect 2397 1004 2403 1076
rect 2317 944 2323 956
rect 2429 904 2435 1036
rect 2493 944 2499 1036
rect 2509 944 2515 1076
rect 2525 924 2531 1096
rect 2557 984 2563 1056
rect 2317 724 2323 736
rect 2397 724 2403 776
rect 2125 584 2131 676
rect 2157 564 2163 636
rect 2061 504 2067 516
rect 2029 462 2035 500
rect 2141 383 2147 556
rect 2205 524 2211 636
rect 2317 603 2323 636
rect 2349 624 2355 676
rect 2397 664 2403 696
rect 2493 684 2499 836
rect 2589 804 2595 1136
rect 2605 1124 2611 1156
rect 2653 1044 2659 1336
rect 2733 1283 2739 1456
rect 2749 1384 2755 1516
rect 2845 1423 2851 1476
rect 2877 1464 2883 1756
rect 2957 1644 2963 1716
rect 3021 1637 3036 1643
rect 2957 1504 2963 1558
rect 2829 1417 2851 1423
rect 2797 1384 2803 1416
rect 2797 1324 2803 1336
rect 2797 1284 2803 1296
rect 2717 1277 2739 1283
rect 2632 1006 2638 1014
rect 2646 1006 2652 1014
rect 2660 1006 2666 1014
rect 2674 1006 2680 1014
rect 2717 964 2723 1277
rect 2829 1224 2835 1417
rect 2845 1304 2851 1396
rect 2893 1364 2899 1416
rect 3021 1404 3027 1637
rect 3053 1544 3059 1716
rect 3069 1504 3075 1516
rect 3037 1384 3043 1456
rect 3053 1424 3059 1476
rect 2893 1344 2899 1356
rect 2957 1344 2963 1356
rect 3053 1344 3059 1356
rect 2941 1304 2947 1336
rect 2957 1204 2963 1316
rect 3021 1264 3027 1296
rect 3069 1204 3075 1496
rect 3085 1304 3091 2236
rect 3101 2184 3107 2236
rect 3101 1924 3107 1976
rect 3117 1683 3123 2276
rect 3133 2184 3139 2256
rect 3181 2204 3187 2416
rect 3197 2284 3203 2756
rect 3213 2504 3219 2576
rect 3229 2523 3235 2876
rect 3309 2723 3315 2956
rect 3325 2944 3331 3036
rect 3357 2944 3363 3016
rect 3373 2904 3379 3076
rect 3325 2884 3331 2896
rect 3389 2884 3395 3216
rect 3405 3144 3411 3236
rect 3453 3204 3459 3297
rect 3469 3264 3475 3316
rect 3533 3284 3539 3316
rect 3549 3264 3555 3316
rect 3613 3304 3619 3316
rect 3677 3304 3683 3316
rect 3757 3304 3763 3336
rect 3789 3304 3795 3316
rect 3805 3304 3811 3336
rect 3821 3304 3827 3496
rect 3837 3344 3843 3396
rect 3869 3344 3875 3476
rect 3901 3344 3907 4016
rect 3949 4004 3955 4036
rect 4061 4024 4067 4036
rect 3917 3743 3923 3996
rect 3981 3844 3987 3876
rect 3997 3784 4003 3816
rect 3917 3737 3939 3743
rect 3933 3724 3939 3737
rect 3933 3704 3939 3716
rect 3917 3344 3923 3696
rect 3981 3624 3987 3756
rect 4013 3703 4019 3856
rect 4077 3784 4083 3816
rect 4029 3744 4035 3776
rect 4125 3724 4131 4076
rect 4152 4006 4158 4014
rect 4166 4006 4172 4014
rect 4180 4006 4186 4014
rect 4194 4006 4200 4014
rect 4253 3824 4259 4116
rect 4429 4044 4435 4100
rect 4317 3904 4323 3996
rect 4493 3904 4499 4196
rect 4509 4124 4515 4296
rect 4525 4164 4531 4236
rect 4701 4224 4707 4436
rect 4781 4284 4787 4396
rect 4829 4384 4835 4516
rect 4845 4404 4851 4516
rect 4861 4444 4867 4496
rect 4957 4484 4963 4516
rect 4941 4477 4956 4483
rect 4637 4144 4643 4176
rect 4541 4044 4547 4096
rect 4269 3804 4275 3896
rect 4285 3864 4291 3876
rect 4013 3697 4035 3703
rect 4029 3644 4035 3697
rect 4013 3584 4019 3636
rect 4029 3464 4035 3636
rect 4152 3606 4158 3614
rect 4166 3606 4172 3614
rect 4180 3606 4186 3614
rect 4194 3606 4200 3614
rect 4125 3520 4131 3558
rect 4221 3544 4227 3656
rect 3901 3324 3907 3336
rect 3981 3324 3987 3376
rect 3997 3344 4003 3356
rect 4029 3324 4035 3336
rect 3661 3264 3667 3296
rect 3757 3284 3763 3296
rect 3885 3283 3891 3316
rect 3917 3304 3923 3316
rect 3933 3283 3939 3296
rect 4045 3284 4051 3316
rect 4061 3304 4067 3456
rect 4141 3384 4147 3476
rect 4221 3384 4227 3536
rect 4077 3344 4083 3356
rect 4125 3344 4131 3356
rect 4237 3324 4243 3576
rect 4253 3504 4259 3716
rect 4333 3644 4339 3756
rect 4365 3624 4371 3736
rect 4333 3584 4339 3616
rect 4429 3584 4435 3896
rect 4461 3644 4467 3696
rect 4493 3684 4499 3836
rect 4525 3583 4531 3756
rect 4557 3724 4563 4116
rect 4573 3724 4579 3896
rect 4653 3823 4659 3856
rect 4685 3844 4691 3876
rect 4653 3817 4675 3823
rect 4637 3744 4643 3816
rect 4669 3764 4675 3817
rect 4541 3644 4547 3696
rect 4525 3577 4547 3583
rect 4285 3504 4291 3576
rect 4285 3477 4300 3483
rect 4269 3464 4275 3476
rect 4285 3344 4291 3477
rect 4317 3464 4323 3476
rect 4541 3464 4547 3577
rect 4573 3504 4579 3716
rect 4669 3524 4675 3576
rect 4749 3544 4755 4076
rect 4781 3924 4787 3976
rect 4781 3864 4787 3896
rect 4845 3884 4851 4216
rect 4893 4144 4899 4476
rect 4877 3964 4883 4036
rect 4877 3944 4883 3956
rect 4861 3924 4867 3936
rect 4861 3744 4867 3896
rect 4813 3524 4819 3576
rect 4573 3464 4579 3476
rect 4333 3304 4339 3436
rect 4541 3403 4547 3456
rect 4525 3397 4547 3403
rect 4525 3364 4531 3397
rect 4557 3344 4563 3376
rect 4637 3324 4643 3496
rect 3885 3277 3939 3283
rect 3421 3064 3427 3096
rect 3437 3084 3443 3116
rect 3453 3064 3459 3196
rect 3469 3164 3475 3256
rect 3309 2717 3324 2723
rect 3293 2644 3299 2676
rect 3277 2544 3283 2576
rect 3229 2517 3244 2523
rect 3229 2424 3235 2517
rect 3261 2503 3267 2516
rect 3252 2497 3267 2503
rect 3277 2484 3283 2536
rect 3325 2524 3331 2636
rect 3357 2464 3363 2536
rect 3373 2484 3379 2836
rect 3421 2824 3427 3056
rect 3437 2884 3443 3016
rect 3453 2964 3459 3036
rect 3453 2924 3459 2936
rect 3405 2744 3411 2816
rect 3421 2704 3427 2756
rect 3437 2723 3443 2776
rect 3453 2764 3459 2916
rect 3469 2904 3475 3076
rect 3517 3044 3523 3116
rect 3533 3084 3539 3176
rect 3581 3104 3587 3116
rect 3613 3084 3619 3096
rect 3629 3024 3635 3096
rect 3693 2984 3699 3016
rect 3565 2924 3571 2956
rect 3597 2944 3603 2956
rect 3485 2844 3491 2876
rect 3613 2864 3619 2916
rect 3469 2823 3475 2836
rect 3469 2817 3491 2823
rect 3469 2724 3475 2796
rect 3485 2783 3491 2817
rect 3501 2804 3507 2836
rect 3629 2784 3635 2916
rect 3485 2777 3507 2783
rect 3501 2763 3507 2777
rect 3501 2757 3523 2763
rect 3437 2717 3452 2723
rect 3405 2544 3411 2696
rect 3469 2564 3475 2636
rect 3389 2504 3395 2536
rect 3373 2404 3379 2436
rect 3245 2320 3251 2358
rect 3229 2283 3235 2296
rect 3309 2284 3315 2316
rect 3229 2277 3251 2283
rect 3181 2184 3187 2196
rect 3133 2104 3139 2176
rect 3197 2144 3203 2176
rect 3213 2124 3219 2216
rect 3245 2184 3251 2277
rect 3341 2203 3347 2256
rect 3341 2197 3363 2203
rect 3309 2124 3315 2176
rect 3325 2124 3331 2136
rect 3277 2104 3283 2116
rect 3341 2064 3347 2096
rect 3357 2084 3363 2197
rect 3421 2164 3427 2476
rect 3485 2244 3491 2656
rect 3501 2624 3507 2696
rect 3517 2683 3523 2757
rect 3629 2724 3635 2736
rect 3588 2697 3612 2703
rect 3517 2677 3548 2683
rect 3677 2624 3683 2696
rect 3709 2684 3715 2976
rect 3757 2924 3763 3276
rect 3981 3124 3987 3176
rect 3885 3064 3891 3076
rect 3853 2964 3859 3056
rect 3949 2924 3955 3096
rect 3757 2724 3763 2836
rect 3949 2784 3955 2916
rect 3981 2844 3987 2896
rect 3613 2617 3651 2623
rect 3373 2144 3379 2156
rect 3437 2144 3443 2236
rect 3501 2184 3507 2276
rect 3517 2264 3523 2476
rect 3533 2363 3539 2536
rect 3581 2524 3587 2576
rect 3613 2563 3619 2617
rect 3645 2604 3651 2617
rect 3597 2557 3619 2563
rect 3597 2544 3603 2557
rect 3677 2544 3683 2616
rect 3693 2544 3699 2576
rect 3597 2503 3603 2516
rect 3588 2497 3603 2503
rect 3549 2484 3555 2496
rect 3613 2424 3619 2536
rect 3725 2524 3731 2556
rect 3741 2544 3747 2636
rect 3661 2444 3667 2516
rect 3549 2384 3555 2396
rect 3533 2357 3555 2363
rect 3421 2124 3427 2136
rect 3453 2124 3459 2136
rect 3197 1884 3203 1896
rect 3229 1864 3235 1996
rect 3245 1984 3251 2036
rect 3309 1924 3315 2036
rect 3357 1804 3363 2076
rect 3389 2044 3395 2096
rect 3453 1904 3459 2036
rect 3469 1924 3475 2096
rect 3405 1764 3411 1796
rect 3373 1744 3379 1756
rect 3165 1724 3171 1736
rect 3117 1677 3139 1683
rect 3117 1364 3123 1436
rect 2941 1120 2947 1158
rect 2957 1024 2963 1096
rect 2925 984 2931 1016
rect 2637 764 2643 916
rect 2717 804 2723 956
rect 2957 944 2963 956
rect 2973 924 2979 1196
rect 3133 1184 3139 1677
rect 3165 1524 3171 1576
rect 3197 1524 3203 1716
rect 3277 1644 3283 1696
rect 3293 1644 3299 1716
rect 3261 1464 3267 1476
rect 3181 1104 3187 1196
rect 2845 844 2851 896
rect 2781 784 2787 796
rect 2605 704 2611 756
rect 2893 704 2899 916
rect 2909 724 2915 736
rect 2973 704 2979 916
rect 2301 597 2323 603
rect 2301 544 2307 597
rect 2189 504 2195 516
rect 2141 377 2163 383
rect 1565 124 1571 136
rect 1645 124 1651 196
rect 1661 184 1667 296
rect 1853 284 1859 296
rect 1869 284 1875 296
rect 1981 284 1987 296
rect 1805 264 1811 276
rect 1741 164 1747 256
rect 1789 204 1795 236
rect 1837 164 1843 176
rect 2077 164 2083 296
rect 2157 264 2163 377
rect 2189 304 2195 496
rect 2237 462 2243 500
rect 2333 384 2339 556
rect 2493 384 2499 656
rect 2525 584 2531 616
rect 2557 524 2563 576
rect 2573 544 2579 556
rect 2605 524 2611 696
rect 2941 684 2947 696
rect 2632 606 2638 614
rect 2646 606 2652 614
rect 2660 606 2666 614
rect 2674 606 2680 614
rect 2525 404 2531 476
rect 2701 462 2707 500
rect 2285 324 2291 376
rect 2397 320 2403 358
rect 2157 203 2163 256
rect 2157 197 2179 203
rect 2173 184 2179 197
rect 2173 164 2179 176
rect 1965 124 1971 156
rect 2141 144 2147 156
rect 2349 124 2355 296
rect 2461 284 2467 296
rect 2493 264 2499 376
rect 2781 343 2787 396
rect 2797 384 2803 556
rect 2877 524 2883 636
rect 2781 337 2803 343
rect 2797 324 2803 337
rect 2877 324 2883 496
rect 2893 304 2899 676
rect 2957 564 2963 676
rect 2973 584 2979 696
rect 2989 504 2995 616
rect 3021 564 3027 896
rect 3037 544 3043 1036
rect 3053 824 3059 896
rect 3053 644 3059 696
rect 3069 684 3075 1076
rect 3117 964 3123 1076
rect 3245 1064 3251 1356
rect 3277 1284 3283 1336
rect 3373 1324 3379 1496
rect 3405 1464 3411 1756
rect 3485 1544 3491 2096
rect 3517 1524 3523 2256
rect 3533 2144 3539 2276
rect 3533 1784 3539 1836
rect 3549 1824 3555 2357
rect 3613 2324 3619 2336
rect 3629 2324 3635 2436
rect 3677 2304 3683 2516
rect 3732 2497 3747 2503
rect 3597 2144 3603 2236
rect 3677 2224 3683 2296
rect 3709 2284 3715 2436
rect 3741 2384 3747 2497
rect 3773 2464 3779 2716
rect 3805 2604 3811 2716
rect 3981 2704 3987 2816
rect 4029 2784 4035 2916
rect 4061 2884 4067 3296
rect 4157 3244 4163 3296
rect 4621 3262 4627 3300
rect 4152 3206 4158 3214
rect 4166 3206 4172 3214
rect 4180 3206 4186 3214
rect 4194 3206 4200 3214
rect 4669 3184 4675 3496
rect 4861 3464 4867 3736
rect 4877 3584 4883 3836
rect 4893 3824 4899 4116
rect 4909 3984 4915 4096
rect 4925 3924 4931 4096
rect 4941 4044 4947 4477
rect 4957 4124 4963 4376
rect 4973 4144 4979 4556
rect 5037 4524 5043 4816
rect 5085 4664 5091 4956
rect 5117 4944 5123 4956
rect 5261 4924 5267 4956
rect 5325 4944 5331 4956
rect 5277 4937 5292 4943
rect 5181 4862 5187 4900
rect 5229 4884 5235 4916
rect 5117 4784 5123 4856
rect 5277 4784 5283 4937
rect 5293 4784 5299 4896
rect 5357 4864 5363 4896
rect 5181 4664 5187 4696
rect 5277 4684 5283 4776
rect 5133 4564 5139 4656
rect 5181 4644 5187 4656
rect 5149 4604 5155 4636
rect 5101 4544 5107 4556
rect 5005 4444 5011 4496
rect 4989 4304 4995 4436
rect 5021 4304 5027 4516
rect 5133 4384 5139 4556
rect 4989 4083 4995 4256
rect 5021 4244 5027 4296
rect 5069 4284 5075 4336
rect 5053 4224 5059 4276
rect 5005 4104 5011 4156
rect 4989 4077 5011 4083
rect 4941 3984 4947 4036
rect 5005 3944 5011 4077
rect 5037 3964 5043 4096
rect 5053 4004 5059 4216
rect 5069 4024 5075 4096
rect 4701 3344 4707 3356
rect 4141 3120 4147 3158
rect 4525 3104 4531 3156
rect 4653 3124 4659 3136
rect 4733 3124 4739 3436
rect 4765 3384 4771 3456
rect 4765 3303 4771 3356
rect 4781 3304 4787 3376
rect 4756 3297 4771 3303
rect 4749 3104 4755 3116
rect 4781 3104 4787 3276
rect 4797 3184 4803 3356
rect 4813 3324 4819 3436
rect 4893 3363 4899 3756
rect 4909 3724 4915 3876
rect 4925 3784 4931 3876
rect 4941 3784 4947 3856
rect 4909 3484 4915 3716
rect 4973 3583 4979 3636
rect 4957 3577 4979 3583
rect 4941 3464 4947 3496
rect 4957 3484 4963 3577
rect 4909 3384 4915 3456
rect 4877 3357 4899 3363
rect 4829 3284 4835 3336
rect 4877 3304 4883 3357
rect 4077 2984 4083 3076
rect 4141 2964 4147 3036
rect 4237 2964 4243 3056
rect 4317 3004 4323 3096
rect 4685 3084 4691 3096
rect 4701 3084 4707 3096
rect 4797 3083 4803 3116
rect 4829 3104 4835 3156
rect 4845 3124 4851 3236
rect 4813 3084 4819 3096
rect 4781 3077 4803 3083
rect 4413 3024 4419 3056
rect 4269 2924 4275 2996
rect 4477 2964 4483 3076
rect 4637 2964 4643 2976
rect 4653 2964 4659 3056
rect 4685 2944 4691 3076
rect 4717 2944 4723 3076
rect 4237 2844 4243 2896
rect 4152 2806 4158 2814
rect 4166 2806 4172 2814
rect 4180 2806 4186 2814
rect 4194 2806 4200 2814
rect 4093 2704 4099 2776
rect 4301 2724 4307 2776
rect 4333 2704 4339 2916
rect 4557 2784 4563 2896
rect 4564 2777 4579 2783
rect 3892 2697 3900 2703
rect 3853 2524 3859 2636
rect 3869 2564 3875 2696
rect 3933 2564 3939 2596
rect 3949 2584 3955 2636
rect 3981 2563 3987 2696
rect 4109 2664 4115 2696
rect 4013 2564 4019 2636
rect 4029 2584 4035 2596
rect 3981 2557 4003 2563
rect 3869 2524 3875 2556
rect 3997 2524 4003 2557
rect 3837 2504 3843 2516
rect 3789 2464 3795 2496
rect 3853 2464 3859 2496
rect 3885 2484 3891 2496
rect 3757 2364 3763 2436
rect 3837 2384 3843 2416
rect 3725 2284 3731 2296
rect 3757 2204 3763 2336
rect 3789 2324 3795 2376
rect 3773 2204 3779 2296
rect 3805 2244 3811 2356
rect 3853 2324 3859 2376
rect 3837 2284 3843 2296
rect 3453 1364 3459 1516
rect 3581 1504 3587 1976
rect 3725 1944 3731 2156
rect 3853 2124 3859 2296
rect 3821 2062 3827 2100
rect 3805 1924 3811 1976
rect 3821 1884 3827 1916
rect 3613 1784 3619 1876
rect 3677 1824 3683 1876
rect 3661 1464 3667 1796
rect 3693 1484 3699 1836
rect 3773 1764 3779 1796
rect 3805 1744 3811 1836
rect 3869 1744 3875 2436
rect 3885 1884 3891 2436
rect 3933 2424 3939 2496
rect 4013 2384 4019 2556
rect 4045 2544 4051 2636
rect 4061 2584 4067 2616
rect 4109 2584 4115 2656
rect 4116 2557 4131 2563
rect 4125 2504 4131 2557
rect 4141 2544 4147 2636
rect 4429 2604 4435 2656
rect 4141 2464 4147 2516
rect 4157 2484 4163 2496
rect 3901 2324 3907 2376
rect 4029 2324 4035 2436
rect 4152 2406 4158 2414
rect 4166 2406 4172 2414
rect 4180 2406 4186 2414
rect 4194 2406 4200 2414
rect 4237 2344 4243 2456
rect 3901 1944 3907 2176
rect 3901 1924 3907 1936
rect 3933 1924 3939 2316
rect 4109 2304 4115 2316
rect 4237 2304 4243 2336
rect 4269 2324 4275 2516
rect 4285 2384 4291 2496
rect 4301 2462 4307 2500
rect 4509 2384 4515 2596
rect 4573 2524 4579 2777
rect 4589 2444 4595 2916
rect 4637 2784 4643 2916
rect 4717 2884 4723 2936
rect 4733 2924 4739 2956
rect 4749 2904 4755 3076
rect 4781 3024 4787 3077
rect 4765 2924 4771 2956
rect 4781 2924 4787 3016
rect 4813 2944 4819 2996
rect 4829 2944 4835 3096
rect 4845 3004 4851 3076
rect 4861 3064 4867 3096
rect 4877 2984 4883 3056
rect 4877 2964 4883 2976
rect 4797 2924 4803 2936
rect 4813 2804 4819 2936
rect 4861 2904 4867 2916
rect 4685 2724 4691 2776
rect 4893 2684 4899 3336
rect 4973 3324 4979 3416
rect 4941 3184 4947 3316
rect 4957 3164 4963 3316
rect 4909 3124 4915 3136
rect 4973 3124 4979 3256
rect 4989 3184 4995 3936
rect 5037 3924 5043 3956
rect 5053 3884 5059 3996
rect 5069 3904 5075 3916
rect 5085 3904 5091 4296
rect 5101 3904 5107 3976
rect 5149 3944 5155 4436
rect 5213 4384 5219 4676
rect 5261 4544 5267 4636
rect 5405 4564 5411 5037
rect 5517 5004 5523 5043
rect 5720 5006 5726 5014
rect 5734 5006 5740 5014
rect 5748 5006 5754 5014
rect 5762 5006 5768 5014
rect 5709 4924 5715 4936
rect 5597 4884 5603 4916
rect 5773 4862 5779 4900
rect 5629 4724 5635 4776
rect 5789 4704 5795 4956
rect 6372 4937 6387 4943
rect 5853 4704 5859 4936
rect 6029 4924 6035 4936
rect 5869 4784 5875 4916
rect 5933 4844 5939 4896
rect 5421 4623 5427 4676
rect 5501 4664 5507 4696
rect 5533 4644 5539 4676
rect 5421 4617 5443 4623
rect 5421 4544 5427 4596
rect 5437 4584 5443 4617
rect 5501 4584 5507 4636
rect 5517 4564 5523 4596
rect 5380 4517 5395 4523
rect 5293 4497 5308 4503
rect 5293 4384 5299 4497
rect 5309 4323 5315 4476
rect 5389 4384 5395 4517
rect 5309 4317 5324 4323
rect 5197 4264 5203 4276
rect 5261 4264 5267 4296
rect 5197 4244 5203 4256
rect 5181 4124 5187 4236
rect 5261 4164 5267 4236
rect 5277 4224 5283 4276
rect 5293 4244 5299 4296
rect 5341 4264 5347 4276
rect 5357 4244 5363 4276
rect 5389 4124 5395 4236
rect 5405 4204 5411 4296
rect 5405 4124 5411 4156
rect 5181 3924 5187 4076
rect 5389 4044 5395 4096
rect 5213 3984 5219 4016
rect 5005 3764 5011 3836
rect 5117 3824 5123 3916
rect 5229 3884 5235 3956
rect 5293 3904 5299 4036
rect 5309 3944 5315 4036
rect 5005 3724 5011 3736
rect 5037 3704 5043 3816
rect 5165 3784 5171 3856
rect 5117 3724 5123 3736
rect 5181 3724 5187 3816
rect 5213 3744 5219 3856
rect 5229 3724 5235 3796
rect 5261 3784 5267 3836
rect 5277 3784 5283 3896
rect 5357 3884 5363 3956
rect 5069 3717 5084 3723
rect 5069 3683 5075 3717
rect 5101 3703 5107 3716
rect 5092 3697 5107 3703
rect 5101 3684 5107 3697
rect 5069 3677 5091 3683
rect 5021 3324 5027 3336
rect 5037 3304 5043 3316
rect 5053 3284 5059 3336
rect 5005 3124 5011 3216
rect 5053 3184 5059 3196
rect 5085 3144 5091 3677
rect 5165 3544 5171 3716
rect 5197 3624 5203 3716
rect 5229 3464 5235 3716
rect 5261 3704 5267 3756
rect 5309 3724 5315 3776
rect 5341 3744 5347 3876
rect 5373 3804 5379 3896
rect 5405 3824 5411 3916
rect 5325 3704 5331 3736
rect 5101 3384 5107 3456
rect 5117 3444 5123 3456
rect 5117 3304 5123 3436
rect 5204 3357 5235 3363
rect 5149 3224 5155 3316
rect 5181 3264 5187 3356
rect 5229 3344 5235 3357
rect 5245 3344 5251 3516
rect 5277 3484 5283 3496
rect 5293 3484 5299 3696
rect 5341 3683 5347 3696
rect 5325 3677 5347 3683
rect 5309 3544 5315 3636
rect 5325 3564 5331 3677
rect 5357 3664 5363 3716
rect 5373 3684 5379 3736
rect 5405 3724 5411 3756
rect 5309 3504 5315 3536
rect 5325 3504 5331 3556
rect 5309 3344 5315 3456
rect 5172 3137 5180 3143
rect 4941 3104 4947 3116
rect 4957 2964 4963 3076
rect 4973 3064 4979 3116
rect 5005 3104 5011 3116
rect 4973 2924 4979 2936
rect 4989 2924 4995 3076
rect 5037 3064 5043 3136
rect 5053 3043 5059 3136
rect 5069 3083 5075 3116
rect 5181 3104 5187 3136
rect 5092 3097 5107 3103
rect 5069 3077 5091 3083
rect 5037 3037 5059 3043
rect 4621 2584 4627 2656
rect 4637 2584 4643 2676
rect 4781 2664 4787 2676
rect 5005 2664 5011 2936
rect 5021 2784 5027 2836
rect 5037 2784 5043 3037
rect 5085 2984 5091 3077
rect 5101 2824 5107 3097
rect 5117 2984 5123 3076
rect 5197 2944 5203 3116
rect 5213 2964 5219 3336
rect 5309 3324 5315 3336
rect 5277 3224 5283 3316
rect 5325 3304 5331 3496
rect 5341 3464 5347 3476
rect 5357 3324 5363 3656
rect 5277 3144 5283 3216
rect 5229 2984 5235 3076
rect 5293 3064 5299 3096
rect 5309 3084 5315 3196
rect 5325 3104 5331 3136
rect 5341 3124 5347 3296
rect 5373 3284 5379 3676
rect 5389 3524 5395 3636
rect 5421 3604 5427 4496
rect 5469 4444 5475 4496
rect 5501 4384 5507 4456
rect 5517 4384 5523 4556
rect 5517 4224 5523 4276
rect 5485 4104 5491 4116
rect 5501 4104 5507 4136
rect 5453 3964 5459 4036
rect 5469 3904 5475 3936
rect 5453 3877 5468 3883
rect 5453 3704 5459 3877
rect 5469 3684 5475 3716
rect 5421 3504 5427 3536
rect 5389 3464 5395 3496
rect 5389 3424 5395 3456
rect 5405 3444 5411 3476
rect 5389 3244 5395 3396
rect 5421 3324 5427 3496
rect 5437 3444 5443 3616
rect 5469 3584 5475 3676
rect 5485 3604 5491 3716
rect 5501 3564 5507 3636
rect 5533 3624 5539 4616
rect 5597 4524 5603 4656
rect 5629 4524 5635 4696
rect 5693 4604 5699 4676
rect 5757 4664 5763 4696
rect 5720 4606 5726 4614
rect 5734 4606 5740 4614
rect 5748 4606 5754 4614
rect 5762 4606 5768 4614
rect 5789 4564 5795 4696
rect 5901 4664 5907 4716
rect 5933 4624 5939 4696
rect 5949 4544 5955 4916
rect 6349 4844 6355 4936
rect 6013 4684 6019 4716
rect 6061 4704 6067 4716
rect 6093 4704 6099 4716
rect 6125 4684 6131 4696
rect 5965 4584 5971 4676
rect 6029 4543 6035 4636
rect 6061 4544 6067 4576
rect 6093 4564 6099 4676
rect 6109 4664 6115 4676
rect 6109 4584 6115 4616
rect 6125 4564 6131 4676
rect 6093 4544 6099 4556
rect 6020 4537 6035 4543
rect 5821 4524 5827 4536
rect 5917 4524 5923 4536
rect 5997 4504 6003 4516
rect 5549 4444 5555 4496
rect 5549 4324 5555 4436
rect 5613 4264 5619 4476
rect 5885 4462 5891 4500
rect 5629 4304 5635 4358
rect 5933 4304 5939 4476
rect 5549 4204 5555 4236
rect 5549 4104 5555 4116
rect 5581 4103 5587 4156
rect 5597 4124 5603 4136
rect 5629 4124 5635 4236
rect 5693 4144 5699 4216
rect 5720 4206 5726 4214
rect 5734 4206 5740 4214
rect 5748 4206 5754 4214
rect 5762 4206 5768 4214
rect 5581 4097 5596 4103
rect 5629 3924 5635 4116
rect 5645 3964 5651 4136
rect 5661 4117 5676 4123
rect 5549 3904 5555 3916
rect 5565 3864 5571 3876
rect 5565 3724 5571 3856
rect 5645 3824 5651 3876
rect 5629 3684 5635 3718
rect 5533 3484 5539 3516
rect 5565 3424 5571 3496
rect 5565 3344 5571 3356
rect 5357 3124 5363 3236
rect 5389 3184 5395 3236
rect 5421 3144 5427 3316
rect 5437 3104 5443 3296
rect 5469 3184 5475 3256
rect 5389 3084 5395 3096
rect 5165 2924 5171 2936
rect 5117 2884 5123 2916
rect 5197 2904 5203 2936
rect 5229 2924 5235 2976
rect 5261 2964 5267 3036
rect 5261 2944 5267 2956
rect 5149 2704 5155 2836
rect 5197 2744 5203 2896
rect 5213 2724 5219 2916
rect 5309 2904 5315 2936
rect 5341 2924 5347 2936
rect 5389 2924 5395 3016
rect 5421 2984 5427 3076
rect 5437 3064 5443 3096
rect 5277 2724 5283 2836
rect 5293 2784 5299 2796
rect 5325 2704 5331 2816
rect 5341 2784 5347 2916
rect 5357 2704 5363 2836
rect 5421 2804 5427 2896
rect 5485 2784 5491 3296
rect 5549 3184 5555 3316
rect 5581 3304 5587 3516
rect 5613 3464 5619 3556
rect 5661 3544 5667 4117
rect 5709 4084 5715 4096
rect 5757 4084 5763 4096
rect 5677 3984 5683 4076
rect 5757 3944 5763 4076
rect 5837 3984 5843 4296
rect 5997 4284 6003 4496
rect 6029 4484 6035 4516
rect 6125 4464 6131 4536
rect 6141 4524 6147 4636
rect 6173 4624 6179 4716
rect 6221 4704 6227 4836
rect 6349 4724 6355 4836
rect 6205 4664 6211 4676
rect 6221 4624 6227 4676
rect 6317 4664 6323 4676
rect 6317 4524 6323 4616
rect 6333 4544 6339 4696
rect 6205 4504 6211 4516
rect 6317 4484 6323 4516
rect 6301 4324 6307 4376
rect 6093 4304 6099 4316
rect 5949 4164 5955 4256
rect 5869 4124 5875 4156
rect 5981 4144 5987 4176
rect 6045 4062 6051 4100
rect 6061 3984 6067 4076
rect 6077 4004 6083 4236
rect 6205 4223 6211 4276
rect 6189 4217 6211 4223
rect 6189 4184 6195 4217
rect 6125 4144 6131 4156
rect 6077 3944 6083 3996
rect 6093 3944 6099 4116
rect 6237 4104 6243 4136
rect 6269 4104 6275 4136
rect 5693 3864 5699 3936
rect 5693 3764 5699 3856
rect 5720 3806 5726 3814
rect 5734 3806 5740 3814
rect 5748 3806 5754 3814
rect 5762 3806 5768 3814
rect 5805 3784 5811 3916
rect 5837 3844 5843 3896
rect 5853 3824 5859 3876
rect 5885 3864 5891 3876
rect 5709 3743 5715 3776
rect 5700 3737 5715 3743
rect 5725 3723 5731 3756
rect 5821 3744 5827 3756
rect 5901 3744 5907 3756
rect 5789 3724 5795 3736
rect 5917 3724 5923 3736
rect 5709 3717 5731 3723
rect 5668 3537 5683 3543
rect 5661 3444 5667 3476
rect 5597 3384 5603 3436
rect 5565 3164 5571 3236
rect 5581 3124 5587 3296
rect 5613 3124 5619 3136
rect 5629 3124 5635 3276
rect 5677 3164 5683 3537
rect 5693 3344 5699 3716
rect 5709 3684 5715 3717
rect 5725 3684 5731 3696
rect 5725 3524 5731 3676
rect 5773 3584 5779 3716
rect 5789 3524 5795 3556
rect 5789 3504 5795 3516
rect 5805 3504 5811 3536
rect 5741 3464 5747 3496
rect 5821 3484 5827 3716
rect 5853 3524 5859 3696
rect 5885 3684 5891 3716
rect 5901 3504 5907 3596
rect 5720 3406 5726 3414
rect 5734 3406 5740 3414
rect 5748 3406 5754 3414
rect 5762 3406 5768 3414
rect 5821 3344 5827 3476
rect 5837 3464 5843 3496
rect 5885 3444 5891 3496
rect 5853 3324 5859 3436
rect 5885 3324 5891 3436
rect 5901 3364 5907 3496
rect 5933 3364 5939 3676
rect 5965 3484 5971 3876
rect 6045 3784 6051 3816
rect 5981 3424 5987 3656
rect 5908 3357 5923 3363
rect 5901 3303 5907 3336
rect 5892 3297 5907 3303
rect 5677 3104 5683 3156
rect 5821 3124 5827 3236
rect 5197 2664 5203 2676
rect 4813 2604 4819 2656
rect 4893 2584 4899 2656
rect 4701 2564 4707 2576
rect 4973 2564 4979 2636
rect 5053 2564 5059 2656
rect 5213 2624 5219 2636
rect 5341 2604 5347 2676
rect 5421 2664 5427 2676
rect 5277 2564 5283 2596
rect 5469 2584 5475 2736
rect 5501 2644 5507 2956
rect 5517 2924 5523 3056
rect 5533 2964 5539 3096
rect 5565 3084 5571 3096
rect 5581 3063 5587 3096
rect 5565 3057 5587 3063
rect 5565 2844 5571 3057
rect 5597 2984 5603 3076
rect 5693 3024 5699 3076
rect 5709 3044 5715 3056
rect 5720 3006 5726 3014
rect 5734 3006 5740 3014
rect 5748 3006 5754 3014
rect 5762 3006 5768 3014
rect 5789 2944 5795 3076
rect 5805 2944 5811 2976
rect 5693 2924 5699 2936
rect 5821 2924 5827 3116
rect 5837 3004 5843 3096
rect 5885 2924 5891 3036
rect 5917 2924 5923 3357
rect 5933 3324 5939 3356
rect 5949 3264 5955 3336
rect 5981 3324 5987 3416
rect 5956 3257 5971 3263
rect 5965 3084 5971 3257
rect 5981 3144 5987 3296
rect 5997 3284 6003 3396
rect 6029 3324 6035 3716
rect 6061 3524 6067 3756
rect 6077 3744 6083 3936
rect 6109 3904 6115 3916
rect 6093 3864 6099 3896
rect 6125 3884 6131 3956
rect 6141 3884 6147 3896
rect 6109 3764 6115 3856
rect 6157 3784 6163 3836
rect 6077 3724 6083 3736
rect 6077 3404 6083 3716
rect 6125 3664 6131 3756
rect 6205 3744 6211 3956
rect 6221 3884 6227 3956
rect 6237 3844 6243 3896
rect 6269 3864 6275 4096
rect 6285 4004 6291 4136
rect 6093 3444 6099 3456
rect 6125 3444 6131 3496
rect 6173 3464 6179 3516
rect 6013 3124 6019 3136
rect 6013 3104 6019 3116
rect 6029 3084 6035 3316
rect 6077 3264 6083 3336
rect 6061 3084 6067 3096
rect 6077 3084 6083 3256
rect 6093 3104 6099 3196
rect 5965 3024 5971 3076
rect 5981 3044 5987 3076
rect 5933 2924 5939 2936
rect 5981 2924 5987 3036
rect 4717 2544 4723 2556
rect 4605 2504 4611 2516
rect 4285 2304 4291 2376
rect 4573 2304 4579 2316
rect 3933 1884 3939 1916
rect 3949 1843 3955 2216
rect 3988 2117 4003 2123
rect 3965 1984 3971 2056
rect 3965 1864 3971 1896
rect 3949 1837 3971 1843
rect 3949 1724 3955 1736
rect 3965 1724 3971 1837
rect 3789 1524 3795 1576
rect 3805 1504 3811 1716
rect 3869 1644 3875 1700
rect 3981 1583 3987 1636
rect 3997 1584 4003 2117
rect 4013 2104 4019 2196
rect 4109 2124 4115 2296
rect 4317 2284 4323 2296
rect 4237 2164 4243 2256
rect 4013 2084 4019 2096
rect 4029 1984 4035 2036
rect 4061 1764 4067 2116
rect 4141 2062 4147 2100
rect 4152 2006 4158 2014
rect 4166 2006 4172 2014
rect 4180 2006 4186 2014
rect 4194 2006 4200 2014
rect 4173 1904 4179 1976
rect 4365 1924 4371 2256
rect 4397 2084 4403 2276
rect 4509 2164 4515 2236
rect 4397 2024 4403 2036
rect 4461 1984 4467 2036
rect 4541 1920 4547 1958
rect 4077 1824 4083 1876
rect 4077 1784 4083 1816
rect 4093 1804 4099 1836
rect 4125 1784 4131 1836
rect 4173 1784 4179 1896
rect 4333 1764 4339 1856
rect 4477 1824 4483 1876
rect 4525 1784 4531 1816
rect 4013 1684 4019 1716
rect 4045 1664 4051 1716
rect 4253 1683 4259 1716
rect 4237 1677 4259 1683
rect 4152 1606 4158 1614
rect 4166 1606 4172 1614
rect 4180 1606 4186 1614
rect 4194 1606 4200 1614
rect 4221 1584 4227 1676
rect 3965 1577 3987 1583
rect 3901 1520 3907 1558
rect 3965 1484 3971 1577
rect 3469 1364 3475 1456
rect 3997 1424 4003 1456
rect 3677 1364 3683 1416
rect 4109 1364 4115 1416
rect 4141 1344 4147 1396
rect 3341 1262 3347 1300
rect 3085 720 3091 758
rect 3149 744 3155 1056
rect 3165 924 3171 1016
rect 3245 964 3251 1056
rect 3341 862 3347 900
rect 3069 603 3075 676
rect 3149 664 3155 676
rect 3069 597 3091 603
rect 3069 524 3075 576
rect 3085 544 3091 597
rect 3101 544 3107 556
rect 3021 304 3027 336
rect 3117 324 3123 436
rect 2573 264 2579 296
rect 2605 164 2611 236
rect 2632 206 2638 214
rect 2646 206 2652 214
rect 2660 206 2666 214
rect 2674 206 2680 214
rect 2717 184 2723 296
rect 3021 284 3027 296
rect 3133 284 3139 476
rect 2765 164 2771 276
rect 2365 144 2371 156
rect 2509 144 2515 156
rect 2397 124 2403 136
rect 2605 124 2611 156
rect 2733 144 2739 156
rect 2765 144 2771 156
rect 2733 124 2739 136
rect 1117 104 1123 116
rect 2029 104 2035 116
rect 2861 104 2867 236
rect 2909 184 2915 236
rect 2925 124 2931 256
rect 3181 184 3187 656
rect 3357 644 3363 1256
rect 3373 1104 3379 1316
rect 3421 1264 3427 1316
rect 3501 1263 3507 1316
rect 3501 1257 3523 1263
rect 3581 1262 3587 1300
rect 3421 1204 3427 1236
rect 3501 1184 3507 1236
rect 3517 1204 3523 1257
rect 3645 1224 3651 1336
rect 3917 1324 3923 1336
rect 4237 1324 4243 1677
rect 4285 1504 4291 1576
rect 4253 1364 4259 1456
rect 4205 1262 4211 1300
rect 4237 1264 4243 1316
rect 3885 1204 3891 1236
rect 3645 1184 3651 1196
rect 3581 1124 3587 1176
rect 3901 1120 3907 1158
rect 3373 924 3379 1096
rect 3581 944 3587 996
rect 3613 964 3619 1056
rect 3645 1004 3651 1036
rect 3517 844 3523 900
rect 3405 724 3411 776
rect 3437 724 3443 836
rect 3613 744 3619 956
rect 3693 924 3699 1096
rect 3693 803 3699 916
rect 3677 797 3699 803
rect 3357 544 3363 636
rect 3437 524 3443 696
rect 3501 684 3507 716
rect 3533 664 3539 736
rect 3421 462 3427 500
rect 3405 320 3411 358
rect 3437 304 3443 516
rect 3485 344 3491 616
rect 3677 524 3683 797
rect 3773 744 3779 836
rect 3837 784 3843 1056
rect 3917 944 3923 1196
rect 3933 924 3939 1176
rect 3997 1104 4003 1196
rect 4013 1144 4019 1236
rect 4093 1184 4099 1216
rect 4152 1206 4158 1214
rect 4166 1206 4172 1214
rect 4180 1206 4186 1214
rect 4194 1206 4200 1214
rect 4045 1104 4051 1176
rect 4125 1144 4131 1156
rect 4109 1124 4115 1136
rect 4157 1104 4163 1176
rect 4269 1104 4275 1476
rect 4285 1184 4291 1496
rect 4317 1384 4323 1516
rect 4333 1424 4339 1756
rect 4365 1744 4371 1776
rect 4557 1764 4563 1916
rect 4509 1744 4515 1756
rect 4573 1724 4579 1896
rect 4589 1824 4595 2436
rect 4605 2320 4611 2358
rect 4781 2304 4787 2496
rect 4701 2184 4707 2256
rect 4701 2144 4707 2156
rect 4701 2064 4707 2116
rect 4669 1964 4675 1976
rect 4653 1924 4659 1956
rect 4621 1904 4627 1916
rect 4669 1884 4675 1956
rect 4765 1904 4771 2136
rect 4813 1944 4819 2536
rect 4685 1884 4691 1896
rect 4813 1884 4819 1936
rect 4829 1904 4835 2336
rect 4861 2244 4867 2256
rect 4845 2237 4860 2243
rect 4845 2164 4851 2237
rect 4845 1904 4851 1916
rect 4621 1744 4627 1836
rect 4589 1704 4595 1736
rect 4653 1724 4659 1876
rect 4429 1644 4435 1700
rect 4541 1644 4547 1696
rect 4573 1604 4579 1636
rect 4365 1524 4371 1536
rect 4445 1520 4451 1558
rect 4349 1404 4355 1436
rect 4413 1324 4419 1496
rect 4541 1424 4547 1456
rect 4573 1364 4579 1416
rect 3997 1064 4003 1096
rect 4061 1084 4067 1096
rect 4125 944 4131 1036
rect 4253 964 4259 1056
rect 4285 984 4291 1176
rect 4301 1084 4307 1236
rect 4333 1104 4339 1256
rect 4477 1244 4483 1300
rect 4397 1184 4403 1236
rect 4541 1124 4547 1176
rect 4301 1004 4307 1076
rect 4445 984 4451 1076
rect 4509 984 4515 1076
rect 4573 1064 4579 1356
rect 4653 1184 4659 1636
rect 4669 1484 4675 1636
rect 4621 1117 4636 1123
rect 4589 1084 4595 1096
rect 4285 944 4291 956
rect 4509 924 4515 976
rect 4525 944 4531 996
rect 4573 924 4579 956
rect 4605 944 4611 996
rect 3949 903 3955 916
rect 4013 904 4019 916
rect 3908 897 3955 903
rect 3901 684 3907 736
rect 3965 724 3971 736
rect 3981 724 3987 876
rect 4349 844 4355 900
rect 4381 884 4387 916
rect 3997 704 4003 836
rect 4152 806 4158 814
rect 4166 806 4172 814
rect 4180 806 4186 814
rect 4194 806 4200 814
rect 4381 720 4387 758
rect 4397 704 4403 876
rect 4461 824 4467 896
rect 4461 724 4467 816
rect 4317 684 4323 696
rect 3725 624 3731 676
rect 3757 443 3763 556
rect 3789 544 3795 596
rect 3869 584 3875 656
rect 3885 544 3891 676
rect 3901 544 3907 676
rect 3949 604 3955 636
rect 4013 544 4019 676
rect 3757 437 3779 443
rect 3005 164 3011 176
rect 3037 144 3043 156
rect 3213 124 3219 236
rect 3229 223 3235 296
rect 3485 284 3491 336
rect 3597 304 3603 436
rect 3709 324 3715 396
rect 3757 324 3763 376
rect 3341 264 3347 276
rect 3229 217 3251 223
rect 3245 184 3251 217
rect 3309 184 3315 256
rect 3373 184 3379 216
rect 3597 204 3603 236
rect 3629 224 3635 256
rect 781 44 787 96
rect 1133 44 1139 96
rect 1965 44 1971 96
rect 2077 62 2083 100
rect 3101 62 3107 100
rect 1112 6 1118 14
rect 1126 6 1132 14
rect 1140 6 1146 14
rect 1154 6 1160 14
rect 397 -23 419 -17
rect 429 -23 451 -17
rect 2157 -23 2163 16
rect 2429 -17 2435 36
rect 2413 -23 2435 -17
rect 2557 -17 2563 36
rect 2685 -17 2691 36
rect 3181 -17 3187 36
rect 2557 -23 2579 -17
rect 2685 -23 2707 -17
rect 3181 -23 3203 -17
rect 3229 -23 3235 136
rect 3245 124 3251 176
rect 3533 164 3539 196
rect 3693 144 3699 276
rect 3709 124 3715 296
rect 3757 124 3763 236
rect 3773 204 3779 437
rect 3789 304 3795 516
rect 3885 444 3891 496
rect 3949 404 3955 436
rect 3789 124 3795 296
rect 3853 284 3859 336
rect 4013 284 4019 536
rect 4077 364 4083 636
rect 4189 544 4195 596
rect 4285 564 4291 656
rect 4397 524 4403 696
rect 4461 604 4467 636
rect 4477 584 4483 876
rect 4493 684 4499 916
rect 4548 897 4563 903
rect 4516 717 4531 723
rect 4509 624 4515 636
rect 4525 584 4531 717
rect 4557 584 4563 897
rect 4589 683 4595 936
rect 4621 784 4627 1117
rect 4637 1104 4643 1116
rect 4669 1084 4675 1096
rect 4685 1083 4691 1876
rect 4749 1724 4755 1836
rect 4829 1724 4835 1896
rect 4717 1703 4723 1716
rect 4829 1703 4835 1716
rect 4717 1697 4739 1703
rect 4829 1697 4844 1703
rect 4733 1584 4739 1697
rect 4861 1644 4867 2036
rect 4877 1924 4883 2516
rect 5005 2484 5011 2516
rect 5149 2504 5155 2516
rect 4893 2304 4899 2336
rect 4909 2304 4915 2476
rect 5181 2462 5187 2500
rect 5501 2384 5507 2616
rect 5085 2320 5091 2358
rect 4925 2264 4931 2276
rect 5069 2224 5075 2296
rect 5037 2164 5043 2176
rect 4893 2104 4899 2116
rect 4941 2062 4947 2100
rect 4941 1864 4947 2016
rect 4957 1884 4963 1936
rect 4948 1857 4963 1863
rect 4893 1724 4899 1816
rect 4957 1764 4963 1857
rect 4733 1384 4739 1556
rect 4765 1344 4771 1636
rect 4797 1524 4803 1576
rect 4893 1484 4899 1636
rect 4941 1604 4947 1756
rect 5005 1744 5011 2116
rect 5037 2024 5043 2156
rect 5117 2124 5123 2216
rect 5181 2184 5187 2256
rect 5293 2184 5299 2276
rect 5389 2264 5395 2316
rect 5533 2304 5539 2576
rect 5549 2544 5555 2836
rect 5613 2784 5619 2796
rect 5629 2704 5635 2876
rect 5645 2864 5651 2916
rect 5693 2664 5699 2916
rect 5837 2904 5843 2916
rect 5725 2704 5731 2776
rect 5869 2704 5875 2796
rect 5885 2724 5891 2916
rect 5917 2804 5923 2916
rect 5924 2717 5948 2723
rect 5597 2564 5603 2656
rect 5661 2544 5667 2596
rect 5677 2524 5683 2636
rect 5693 2564 5699 2656
rect 5709 2644 5715 2696
rect 5853 2684 5859 2696
rect 5720 2606 5726 2614
rect 5734 2606 5740 2614
rect 5748 2606 5754 2614
rect 5762 2606 5768 2614
rect 5757 2524 5763 2536
rect 5789 2503 5795 2636
rect 5805 2524 5811 2596
rect 5885 2584 5891 2716
rect 5965 2703 5971 2836
rect 5981 2704 5987 2876
rect 5997 2824 6003 3076
rect 6077 3064 6083 3076
rect 6125 3064 6131 3076
rect 6013 2944 6019 3056
rect 6029 3004 6035 3036
rect 5997 2704 6003 2816
rect 6045 2744 6051 2976
rect 6077 2944 6083 3016
rect 6125 2944 6131 2996
rect 6141 2984 6147 3316
rect 6157 3224 6163 3316
rect 6189 3244 6195 3696
rect 6205 3524 6211 3716
rect 6237 3703 6243 3836
rect 6237 3697 6252 3703
rect 6269 3644 6275 3716
rect 6285 3704 6291 3716
rect 6269 3544 6275 3636
rect 6205 3504 6211 3516
rect 6237 3504 6243 3536
rect 6205 3364 6211 3496
rect 6253 3464 6259 3496
rect 6205 3344 6211 3356
rect 6221 3344 6227 3356
rect 6189 3104 6195 3216
rect 6237 3164 6243 3316
rect 6269 3124 6275 3336
rect 6301 3303 6307 4296
rect 6317 4284 6323 4296
rect 6333 4244 6339 4496
rect 6349 4123 6355 4636
rect 6365 4584 6371 4656
rect 6365 4384 6371 4476
rect 6381 4344 6387 4937
rect 6477 4744 6483 4836
rect 6605 4823 6611 4916
rect 6605 4817 6627 4823
rect 6397 4664 6403 4696
rect 6413 4664 6419 4676
rect 6429 4644 6435 4696
rect 6445 4684 6451 4696
rect 6493 4664 6499 4696
rect 6477 4604 6483 4636
rect 6525 4584 6531 4636
rect 6413 4156 6419 4536
rect 6445 4524 6451 4576
rect 6525 4484 6531 4556
rect 6557 4544 6563 4596
rect 6621 4524 6627 4817
rect 6653 4444 6659 4496
rect 6477 4284 6483 4336
rect 6445 4184 6451 4216
rect 6477 4144 6483 4236
rect 6340 4117 6355 4123
rect 6333 3743 6339 4036
rect 6349 3784 6355 4117
rect 6381 4024 6387 4136
rect 6477 4084 6483 4136
rect 6436 3917 6451 3923
rect 6365 3784 6371 3894
rect 6397 3804 6403 3876
rect 6429 3784 6435 3836
rect 6317 3737 6339 3743
rect 6317 3564 6323 3737
rect 6349 3724 6355 3736
rect 6333 3584 6339 3716
rect 6365 3684 6371 3696
rect 6333 3504 6339 3576
rect 6381 3544 6387 3776
rect 6413 3744 6419 3756
rect 6445 3704 6451 3917
rect 6477 3864 6483 3876
rect 6477 3744 6483 3756
rect 6349 3504 6355 3516
rect 6317 3324 6323 3416
rect 6333 3324 6339 3456
rect 6349 3404 6355 3496
rect 6365 3423 6371 3536
rect 6381 3443 6387 3516
rect 6397 3463 6403 3696
rect 6397 3457 6419 3463
rect 6381 3437 6403 3443
rect 6365 3417 6380 3423
rect 6365 3364 6371 3376
rect 6381 3324 6387 3416
rect 6397 3324 6403 3437
rect 6301 3297 6323 3303
rect 6317 3284 6323 3297
rect 6285 3124 6291 3236
rect 6365 3184 6371 3316
rect 6381 3204 6387 3316
rect 6397 3304 6403 3316
rect 6077 2904 6083 2936
rect 6109 2924 6115 2936
rect 6157 2904 6163 3096
rect 6221 2944 6227 3036
rect 6141 2864 6147 2896
rect 6189 2883 6195 2936
rect 6237 2924 6243 3096
rect 6253 3024 6259 3076
rect 6253 2944 6259 2956
rect 6253 2904 6259 2916
rect 6285 2903 6291 3116
rect 6349 3084 6355 3096
rect 6276 2897 6291 2903
rect 6189 2877 6211 2883
rect 6093 2704 6099 2836
rect 6205 2784 6211 2877
rect 6253 2784 6259 2856
rect 5956 2697 5971 2703
rect 5933 2684 5939 2696
rect 5933 2544 5939 2676
rect 5949 2524 5955 2636
rect 5965 2604 5971 2697
rect 6077 2684 6083 2696
rect 6125 2664 6131 2716
rect 6173 2704 6179 2756
rect 6269 2724 6275 2896
rect 6285 2784 6291 2836
rect 6285 2704 6291 2776
rect 6301 2764 6307 2936
rect 6349 2924 6355 2976
rect 6365 2924 6371 2956
rect 6349 2844 6355 2916
rect 6381 2744 6387 3156
rect 6397 3084 6403 3276
rect 6413 3244 6419 3457
rect 6429 3384 6435 3496
rect 6429 3184 6435 3356
rect 6445 3344 6451 3636
rect 6461 3524 6467 3696
rect 6477 3624 6483 3736
rect 6493 3684 6499 4416
rect 6509 3724 6515 4076
rect 6525 3924 6531 3976
rect 6541 3904 6547 3936
rect 6509 3684 6515 3716
rect 6461 3504 6467 3516
rect 6445 3164 6451 3316
rect 6461 3264 6467 3476
rect 6493 3464 6499 3616
rect 6509 3604 6515 3636
rect 6541 3624 6547 3636
rect 6557 3584 6563 4336
rect 6589 4284 6595 4296
rect 6589 4124 6595 4276
rect 6669 4264 6675 4736
rect 6685 4484 6691 4956
rect 6717 4944 6723 4976
rect 6813 4844 6819 4896
rect 6701 4504 6707 4536
rect 6765 4320 6771 4358
rect 6669 4164 6675 4256
rect 6701 4224 6707 4276
rect 6669 3983 6675 4156
rect 6765 4062 6771 4100
rect 6781 3984 6787 4696
rect 6877 4684 6883 4696
rect 6813 4584 6819 4676
rect 6653 3977 6675 3983
rect 6653 3864 6659 3977
rect 6781 3924 6787 3976
rect 6701 3764 6707 3796
rect 6477 3344 6483 3456
rect 6413 3064 6419 3076
rect 6445 3064 6451 3116
rect 6397 2984 6403 3056
rect 6461 3044 6467 3096
rect 6477 3004 6483 3336
rect 6493 3324 6499 3396
rect 6509 3304 6515 3436
rect 6525 3304 6531 3376
rect 6541 3324 6547 3336
rect 6573 3284 6579 3316
rect 6493 2984 6499 3236
rect 6525 3104 6531 3116
rect 6557 3103 6563 3136
rect 6548 3097 6563 3103
rect 6509 3064 6515 3076
rect 6541 2984 6547 3096
rect 6557 3004 6563 3076
rect 6509 2964 6515 2976
rect 6573 2944 6579 3096
rect 6349 2704 6355 2736
rect 6397 2724 6403 2936
rect 6413 2884 6419 2916
rect 6397 2704 6403 2716
rect 6013 2584 6019 2636
rect 6125 2584 6131 2656
rect 6269 2644 6275 2676
rect 6301 2664 6307 2696
rect 6141 2524 6147 2636
rect 6301 2544 6307 2656
rect 5780 2497 5795 2503
rect 6061 2324 6067 2376
rect 5421 2264 5427 2296
rect 5405 2257 5420 2263
rect 5373 2183 5379 2236
rect 5373 2177 5395 2183
rect 5069 1984 5075 2016
rect 5101 1904 5107 1976
rect 5069 1784 5075 1836
rect 5005 1724 5011 1736
rect 4973 1624 4979 1636
rect 4925 1424 4931 1456
rect 5005 1324 5011 1716
rect 5037 1684 5043 1716
rect 5069 1364 5075 1776
rect 5085 1644 5091 1696
rect 5101 1664 5107 1896
rect 5181 1884 5187 1956
rect 5197 1884 5203 2036
rect 5229 1964 5235 2136
rect 5373 2124 5379 2156
rect 5389 2144 5395 2177
rect 5405 2164 5411 2257
rect 5453 2144 5459 2236
rect 5485 2164 5491 2236
rect 5165 1864 5171 1876
rect 5229 1864 5235 1956
rect 5245 1864 5251 2116
rect 5293 2084 5299 2096
rect 5341 2064 5347 2096
rect 5261 1984 5267 2056
rect 5261 1864 5267 1896
rect 5133 1804 5139 1836
rect 5181 1744 5187 1836
rect 5213 1824 5219 1836
rect 5213 1764 5219 1776
rect 5085 1584 5091 1596
rect 5181 1584 5187 1656
rect 5085 1384 5091 1476
rect 5117 1384 5123 1576
rect 5309 1524 5315 1816
rect 5133 1517 5148 1523
rect 4797 1244 4803 1296
rect 4717 1144 4723 1156
rect 4676 1077 4691 1083
rect 4653 1004 4659 1076
rect 4717 984 4723 1076
rect 4733 984 4739 1236
rect 4749 1124 4755 1176
rect 4797 1124 4803 1136
rect 5085 1120 5091 1158
rect 4749 964 4755 1036
rect 4845 964 4851 1056
rect 4909 1004 4915 1096
rect 4877 944 4883 956
rect 4957 924 4963 996
rect 5069 984 5075 1016
rect 5101 984 5107 1296
rect 5133 984 5139 1517
rect 5197 1484 5203 1496
rect 5213 1484 5219 1516
rect 5197 1364 5203 1476
rect 5229 1463 5235 1496
rect 5277 1484 5283 1516
rect 5309 1504 5315 1516
rect 5325 1484 5331 1836
rect 5341 1704 5347 1870
rect 5373 1844 5379 1876
rect 5405 1784 5411 1876
rect 5453 1724 5459 1876
rect 5501 1784 5507 2296
rect 5549 2264 5555 2316
rect 5565 2304 5571 2316
rect 5581 2304 5587 2316
rect 5565 2164 5571 2276
rect 5613 2264 5619 2276
rect 5517 2124 5523 2136
rect 5549 2124 5555 2136
rect 5565 2104 5571 2156
rect 5629 2123 5635 2236
rect 5620 2117 5635 2123
rect 5549 2084 5555 2096
rect 5549 1824 5555 2076
rect 5565 1883 5571 2096
rect 5645 2084 5651 2156
rect 5661 2144 5667 2316
rect 5725 2304 5731 2316
rect 6189 2304 6195 2536
rect 6285 2524 6291 2536
rect 6301 2384 6307 2536
rect 6317 2504 6323 2636
rect 6349 2564 6355 2696
rect 6365 2684 6371 2696
rect 6413 2604 6419 2676
rect 6429 2644 6435 2716
rect 6445 2704 6451 2936
rect 6461 2924 6467 2936
rect 6461 2704 6467 2716
rect 6493 2704 6499 2716
rect 6445 2684 6451 2696
rect 6429 2584 6435 2636
rect 6445 2543 6451 2676
rect 6445 2537 6460 2543
rect 6413 2504 6419 2536
rect 6333 2324 6339 2376
rect 6461 2324 6467 2516
rect 6477 2484 6483 2496
rect 6509 2404 6515 2816
rect 6525 2704 6531 2876
rect 6589 2824 6595 3736
rect 6701 3604 6707 3756
rect 6797 3743 6803 4116
rect 6813 4004 6819 4436
rect 6797 3737 6819 3743
rect 6813 3724 6819 3737
rect 6797 3644 6803 3700
rect 6605 3144 6611 3496
rect 6621 3484 6627 3496
rect 6669 3484 6675 3596
rect 6669 3344 6675 3476
rect 6701 3443 6707 3496
rect 6733 3464 6739 3496
rect 6797 3464 6803 3616
rect 6685 3437 6707 3443
rect 6685 3344 6691 3437
rect 6717 3364 6723 3436
rect 6765 3424 6771 3436
rect 6621 3304 6627 3316
rect 6637 3284 6643 3296
rect 6685 3264 6691 3336
rect 6749 3284 6755 3318
rect 6621 2924 6627 3176
rect 6653 3084 6659 3096
rect 6669 3084 6675 3256
rect 6765 3084 6771 3196
rect 6765 3024 6771 3076
rect 6669 2944 6675 3016
rect 6573 2704 6579 2756
rect 6589 2704 6595 2796
rect 6605 2724 6611 2736
rect 6637 2704 6643 2716
rect 6733 2704 6739 3016
rect 6765 2704 6771 2736
rect 6525 2544 6531 2676
rect 6589 2564 6595 2696
rect 6557 2524 6563 2556
rect 6525 2504 6531 2516
rect 6237 2302 6243 2316
rect 5684 2277 5692 2283
rect 5661 2124 5667 2136
rect 5597 1904 5603 1936
rect 5645 1904 5651 1916
rect 5629 1897 5644 1903
rect 5565 1877 5580 1883
rect 5581 1864 5587 1876
rect 5453 1644 5459 1716
rect 5469 1684 5475 1716
rect 5325 1464 5331 1476
rect 5341 1464 5347 1596
rect 5373 1564 5379 1636
rect 5405 1584 5411 1616
rect 5421 1524 5427 1636
rect 5229 1457 5251 1463
rect 5165 1344 5171 1356
rect 5165 1084 5171 1096
rect 5181 964 5187 976
rect 5037 924 5043 956
rect 5197 943 5203 1356
rect 5229 1124 5235 1156
rect 5213 1104 5219 1116
rect 5245 1044 5251 1457
rect 5373 1463 5379 1516
rect 5437 1483 5443 1596
rect 5469 1524 5475 1616
rect 5501 1484 5507 1556
rect 5428 1477 5443 1483
rect 5373 1457 5388 1463
rect 5364 1437 5379 1443
rect 5261 1344 5267 1436
rect 5341 1304 5347 1336
rect 5373 1324 5379 1437
rect 5373 1244 5379 1316
rect 5261 1104 5267 1116
rect 5277 984 5283 1076
rect 5293 1064 5299 1076
rect 5188 937 5212 943
rect 4765 884 4771 916
rect 4653 744 4659 876
rect 4941 862 4947 900
rect 4685 724 4691 776
rect 4580 677 4595 683
rect 4253 444 4259 500
rect 4152 406 4158 414
rect 4166 406 4172 414
rect 4180 406 4186 414
rect 4194 406 4200 414
rect 4333 384 4339 476
rect 4221 324 4227 356
rect 4269 284 4275 376
rect 4349 324 4355 516
rect 4429 404 4435 556
rect 4573 544 4579 676
rect 4685 664 4691 696
rect 4781 684 4787 716
rect 5021 664 5027 736
rect 4580 537 4595 543
rect 4381 320 4387 358
rect 4445 304 4451 536
rect 4477 324 4483 436
rect 4541 424 4547 476
rect 4557 304 4563 516
rect 4573 384 4579 476
rect 3885 204 3891 256
rect 3965 164 3971 196
rect 4173 164 4179 236
rect 3933 144 3939 156
rect 4189 124 4195 136
rect 4285 124 4291 296
rect 4301 144 4307 256
rect 4477 204 4483 256
rect 4413 164 4419 196
rect 4589 164 4595 537
rect 4621 524 4627 656
rect 4813 604 4819 656
rect 4749 564 4755 596
rect 4653 444 4659 500
rect 4621 164 4627 316
rect 4669 304 4675 316
rect 4653 184 4659 276
rect 4669 264 4675 296
rect 4685 184 4691 416
rect 4733 324 4739 376
rect 4749 204 4755 556
rect 4989 544 4995 656
rect 5021 584 5027 656
rect 5069 584 5075 896
rect 5005 524 5011 536
rect 4941 504 4947 516
rect 4989 504 4995 516
rect 5021 503 5027 576
rect 5053 544 5059 556
rect 5012 497 5027 503
rect 4781 344 4787 396
rect 4781 284 4787 336
rect 4797 324 4803 416
rect 4973 384 4979 476
rect 4845 284 4851 336
rect 4845 164 4851 196
rect 3661 44 3667 96
rect 3837 44 3843 96
rect 4285 44 4291 96
rect 3309 -17 3315 36
rect 3741 -17 3747 36
rect 3789 -17 3795 36
rect 3309 -23 3331 -17
rect 3725 -23 3747 -17
rect 3773 -23 3795 -17
rect 4125 -17 4131 36
rect 4152 6 4158 14
rect 4166 6 4172 14
rect 4180 6 4186 14
rect 4194 6 4200 14
rect 4125 -23 4211 -17
rect 4637 -23 4643 156
rect 4877 144 4883 276
rect 4893 264 4899 296
rect 4989 264 4995 496
rect 5037 304 5043 516
rect 5053 344 5059 536
rect 5085 504 5091 696
rect 5101 544 5107 936
rect 5309 924 5315 1196
rect 5373 1104 5379 1156
rect 5117 723 5123 876
rect 5133 744 5139 876
rect 5117 717 5132 723
rect 5117 664 5123 717
rect 5165 523 5171 696
rect 5181 684 5187 716
rect 5181 564 5187 676
rect 5156 517 5171 523
rect 5117 484 5123 496
rect 5149 464 5155 516
rect 4941 144 4947 256
rect 5037 184 5043 276
rect 4941 62 4947 100
rect 4925 -23 4931 16
rect 5021 -23 5027 156
rect 5053 124 5059 296
rect 5133 264 5139 396
rect 5149 384 5155 436
rect 5213 404 5219 636
rect 5261 584 5267 896
rect 5277 884 5283 896
rect 5325 684 5331 1076
rect 5357 904 5363 916
rect 5373 904 5379 1096
rect 5389 724 5395 1456
rect 5469 1384 5475 1436
rect 5405 723 5411 1296
rect 5421 1104 5427 1116
rect 5453 1084 5459 1316
rect 5469 1044 5475 1096
rect 5485 1084 5491 1396
rect 5501 1324 5507 1476
rect 5501 1284 5507 1296
rect 5501 1144 5507 1276
rect 5517 1204 5523 1436
rect 5533 1404 5539 1636
rect 5581 1584 5587 1856
rect 5629 1844 5635 1897
rect 5629 1744 5635 1836
rect 5613 1604 5619 1736
rect 5661 1724 5667 2116
rect 5677 2104 5683 2276
rect 5933 2244 5939 2256
rect 5965 2224 5971 2276
rect 5720 2206 5726 2214
rect 5734 2206 5740 2214
rect 5748 2206 5754 2214
rect 5762 2206 5768 2214
rect 5869 2184 5875 2216
rect 5789 2124 5795 2156
rect 5805 2144 5811 2176
rect 6077 2124 6083 2136
rect 6205 2124 6211 2296
rect 6269 2244 6275 2276
rect 6285 2164 6291 2236
rect 6429 2224 6435 2276
rect 6461 2244 6467 2256
rect 6493 2184 6499 2216
rect 6557 2144 6563 2156
rect 6589 2124 6595 2536
rect 6605 2524 6611 2576
rect 6621 2524 6627 2556
rect 6637 2544 6643 2676
rect 6637 2264 6643 2496
rect 6669 2384 6675 2696
rect 6717 2483 6723 2536
rect 6701 2477 6723 2483
rect 6701 2243 6707 2477
rect 6692 2237 6707 2243
rect 6621 2164 6627 2236
rect 6685 2184 6691 2236
rect 5789 2104 5795 2116
rect 5757 1904 5763 1916
rect 5821 1904 5827 1956
rect 5533 1324 5539 1356
rect 5549 1344 5555 1456
rect 5565 1364 5571 1476
rect 5565 1284 5571 1356
rect 5581 1263 5587 1556
rect 5629 1524 5635 1696
rect 5645 1524 5651 1636
rect 5613 1384 5619 1496
rect 5565 1257 5587 1263
rect 5501 1084 5507 1136
rect 5565 1104 5571 1257
rect 5581 1164 5587 1236
rect 5581 1124 5587 1156
rect 5421 764 5427 936
rect 5469 924 5475 1036
rect 5437 724 5443 896
rect 5405 717 5427 723
rect 5357 584 5363 696
rect 5405 564 5411 696
rect 5421 684 5427 717
rect 5293 544 5299 556
rect 5405 544 5411 556
rect 5245 324 5251 536
rect 5389 524 5395 536
rect 5421 524 5427 636
rect 5485 524 5491 1016
rect 5517 924 5523 956
rect 5533 784 5539 876
rect 5549 744 5555 1076
rect 5565 1024 5571 1096
rect 5597 1084 5603 1316
rect 5613 1104 5619 1136
rect 5629 1104 5635 1116
rect 5645 1104 5651 1236
rect 5661 1164 5667 1696
rect 5677 1504 5683 1896
rect 5693 1484 5699 1876
rect 5821 1844 5827 1896
rect 5853 1864 5859 1876
rect 5720 1806 5726 1814
rect 5734 1806 5740 1814
rect 5748 1806 5754 1814
rect 5762 1806 5768 1814
rect 5869 1784 5875 1896
rect 5901 1864 5907 2116
rect 5933 2104 5939 2116
rect 5917 1844 5923 1916
rect 5789 1724 5795 1756
rect 5677 1444 5683 1476
rect 5709 1443 5715 1716
rect 5741 1564 5747 1716
rect 5805 1664 5811 1716
rect 5773 1504 5779 1616
rect 5773 1463 5779 1496
rect 5789 1484 5795 1556
rect 5821 1504 5827 1636
rect 5853 1624 5859 1716
rect 5917 1704 5923 1776
rect 5933 1604 5939 2096
rect 6013 2084 6019 2116
rect 6029 2104 6035 2116
rect 6413 2044 6419 2096
rect 6221 1924 6227 1936
rect 5949 1724 5955 1896
rect 5981 1864 5987 1916
rect 6205 1904 6211 1916
rect 5981 1764 5987 1836
rect 6077 1744 6083 1876
rect 6125 1764 6131 1816
rect 6141 1744 6147 1756
rect 6157 1724 6163 1836
rect 6173 1764 6179 1876
rect 6189 1844 6195 1896
rect 6221 1824 6227 1916
rect 6301 1904 6307 1916
rect 6317 1904 6323 1936
rect 6365 1904 6371 1956
rect 6237 1884 6243 1896
rect 6253 1884 6259 1896
rect 6237 1803 6243 1876
rect 6237 1797 6259 1803
rect 5949 1644 5955 1716
rect 6045 1684 6051 1718
rect 5837 1537 5852 1543
rect 5773 1457 5795 1463
rect 5693 1437 5715 1443
rect 5565 824 5571 836
rect 5581 804 5587 936
rect 5565 704 5571 776
rect 5517 544 5523 576
rect 5405 504 5411 516
rect 5261 324 5267 376
rect 5277 344 5283 476
rect 5485 464 5491 516
rect 5309 324 5315 376
rect 5165 284 5171 296
rect 5341 264 5347 296
rect 5357 264 5363 276
rect 5133 204 5139 256
rect 5213 164 5219 196
rect 5389 164 5395 336
rect 5437 324 5443 336
rect 5469 304 5475 456
rect 5501 364 5507 516
rect 5517 343 5523 536
rect 5533 524 5539 696
rect 5581 664 5587 716
rect 5613 704 5619 936
rect 5629 924 5635 1036
rect 5645 944 5651 956
rect 5677 944 5683 1036
rect 5629 683 5635 896
rect 5645 724 5651 916
rect 5677 864 5683 916
rect 5613 677 5635 683
rect 5597 643 5603 676
rect 5581 637 5603 643
rect 5581 584 5587 637
rect 5501 337 5523 343
rect 5405 184 5411 256
rect 5469 184 5475 296
rect 5501 284 5507 337
rect 5533 324 5539 516
rect 5549 504 5555 516
rect 5581 503 5587 536
rect 5572 497 5587 503
rect 5565 344 5571 496
rect 5597 384 5603 616
rect 5613 584 5619 677
rect 5677 664 5683 856
rect 5693 824 5699 1437
rect 5720 1406 5726 1414
rect 5734 1406 5740 1414
rect 5748 1406 5754 1414
rect 5762 1406 5768 1414
rect 5789 1323 5795 1457
rect 5837 1384 5843 1537
rect 5853 1524 5859 1536
rect 5853 1384 5859 1496
rect 5869 1324 5875 1436
rect 5885 1404 5891 1596
rect 5933 1504 5939 1516
rect 5949 1504 5955 1536
rect 5997 1504 6003 1576
rect 5901 1444 5907 1496
rect 5885 1344 5891 1376
rect 5773 1317 5795 1323
rect 5725 1304 5731 1316
rect 5725 1224 5731 1296
rect 5773 1184 5779 1317
rect 5917 1303 5923 1456
rect 5949 1304 5955 1496
rect 5997 1404 6003 1496
rect 5965 1384 5971 1396
rect 6013 1364 6019 1496
rect 5981 1337 6012 1343
rect 5917 1297 5939 1303
rect 5720 1006 5726 1014
rect 5734 1006 5740 1014
rect 5748 1006 5754 1014
rect 5762 1006 5768 1014
rect 5709 704 5715 836
rect 5725 824 5731 916
rect 5773 724 5779 736
rect 5789 703 5795 1196
rect 5805 964 5811 1116
rect 5821 1064 5827 1276
rect 5853 1164 5859 1296
rect 5837 1104 5843 1116
rect 5901 1104 5907 1136
rect 5917 1104 5923 1116
rect 5821 784 5827 1056
rect 5821 764 5827 776
rect 5853 744 5859 1076
rect 5885 1064 5891 1076
rect 5901 1044 5907 1076
rect 5901 784 5907 816
rect 5869 704 5875 756
rect 5789 697 5804 703
rect 5709 643 5715 676
rect 5677 637 5715 643
rect 5677 564 5683 637
rect 5720 606 5726 614
rect 5734 606 5740 614
rect 5748 606 5754 614
rect 5762 606 5768 614
rect 5677 544 5683 556
rect 5693 544 5699 596
rect 5805 584 5811 596
rect 5821 584 5827 676
rect 5837 544 5843 616
rect 5853 584 5859 696
rect 5885 584 5891 716
rect 5933 604 5939 1297
rect 5981 1284 5987 1337
rect 5997 1304 6003 1316
rect 5949 1264 5955 1276
rect 5949 1084 5955 1256
rect 5997 1204 6003 1296
rect 5965 1124 5971 1156
rect 6013 1124 6019 1316
rect 5997 944 6003 956
rect 6029 924 6035 1656
rect 6109 1523 6115 1636
rect 6173 1584 6179 1756
rect 6237 1724 6243 1756
rect 6253 1744 6259 1797
rect 6269 1664 6275 1716
rect 6285 1704 6291 1716
rect 6141 1524 6147 1536
rect 6093 1517 6115 1523
rect 6093 1484 6099 1517
rect 6061 1444 6067 1476
rect 6045 1324 6051 1376
rect 6061 1344 6067 1436
rect 6093 1324 6099 1396
rect 6109 1304 6115 1496
rect 6141 1424 6147 1436
rect 6173 1363 6179 1436
rect 6173 1357 6195 1363
rect 6189 1344 6195 1357
rect 6045 924 6051 976
rect 5965 904 5971 918
rect 6077 743 6083 1136
rect 6109 1024 6115 1296
rect 6237 1264 6243 1536
rect 6269 1524 6275 1596
rect 6317 1584 6323 1876
rect 6365 1824 6371 1896
rect 6381 1803 6387 1896
rect 6365 1797 6387 1803
rect 6365 1784 6371 1797
rect 6413 1764 6419 1796
rect 6429 1724 6435 2116
rect 6461 1724 6467 1776
rect 6333 1584 6339 1716
rect 6461 1704 6467 1716
rect 6381 1584 6387 1676
rect 6253 1464 6259 1496
rect 6301 1403 6307 1516
rect 6285 1397 6307 1403
rect 6173 1102 6179 1136
rect 6205 1084 6211 1216
rect 6269 1103 6275 1176
rect 6260 1097 6275 1103
rect 6237 1064 6243 1076
rect 6125 984 6131 1056
rect 6109 924 6115 936
rect 6157 924 6163 1016
rect 6061 737 6083 743
rect 6013 704 6019 716
rect 6061 684 6067 737
rect 5613 504 5619 536
rect 5645 517 5660 523
rect 5645 384 5651 517
rect 5853 504 5859 536
rect 5885 484 5891 536
rect 5517 304 5523 316
rect 5565 304 5571 316
rect 5597 304 5603 376
rect 5661 304 5667 436
rect 5677 304 5683 336
rect 5693 304 5699 476
rect 5917 464 5923 516
rect 5933 344 5939 436
rect 5949 384 5955 556
rect 5981 524 5987 536
rect 5549 203 5555 236
rect 5720 206 5726 214
rect 5734 206 5740 214
rect 5748 206 5754 214
rect 5762 206 5768 214
rect 5549 197 5571 203
rect 5085 44 5091 96
rect 5421 -17 5427 156
rect 5565 144 5571 197
rect 5821 164 5827 276
rect 5965 184 5971 516
rect 5997 504 6003 576
rect 6029 524 6035 656
rect 6093 644 6099 916
rect 6125 784 6131 896
rect 6125 704 6131 756
rect 6093 384 6099 636
rect 6141 624 6147 716
rect 6157 704 6163 916
rect 6173 884 6179 936
rect 6173 784 6179 796
rect 6125 564 6131 596
rect 6125 484 6131 518
rect 6157 444 6163 676
rect 6189 524 6195 536
rect 6205 504 6211 516
rect 6221 343 6227 996
rect 6237 944 6243 1056
rect 6253 904 6259 976
rect 6253 704 6259 756
rect 6285 704 6291 1397
rect 6317 1263 6323 1436
rect 6333 1324 6339 1336
rect 6317 1257 6339 1263
rect 6301 1124 6307 1156
rect 6301 1044 6307 1076
rect 6317 924 6323 1236
rect 6333 1083 6339 1257
rect 6349 1244 6355 1496
rect 6349 1104 6355 1196
rect 6365 1104 6371 1396
rect 6381 1324 6387 1436
rect 6397 1424 6403 1676
rect 6445 1504 6451 1636
rect 6461 1544 6467 1636
rect 6477 1564 6483 1956
rect 6493 1684 6499 1916
rect 6509 1904 6515 1936
rect 6525 1884 6531 1976
rect 6509 1784 6515 1836
rect 6525 1744 6531 1876
rect 6557 1843 6563 2116
rect 6621 1904 6627 2156
rect 6621 1864 6627 1896
rect 6557 1837 6579 1843
rect 6557 1784 6563 1796
rect 6445 1404 6451 1496
rect 6461 1464 6467 1496
rect 6461 1344 6467 1356
rect 6381 1204 6387 1316
rect 6413 1304 6419 1336
rect 6477 1324 6483 1416
rect 6493 1324 6499 1576
rect 6557 1544 6563 1596
rect 6541 1504 6547 1536
rect 6557 1504 6563 1536
rect 6413 1224 6419 1296
rect 6381 1104 6387 1156
rect 6477 1104 6483 1316
rect 6333 1077 6348 1083
rect 6349 963 6355 1076
rect 6349 957 6371 963
rect 6365 944 6371 957
rect 6349 923 6355 936
rect 6349 917 6364 923
rect 6301 704 6307 716
rect 6269 544 6275 556
rect 6285 544 6291 696
rect 6333 524 6339 776
rect 6349 684 6355 696
rect 6365 644 6371 696
rect 6381 684 6387 1056
rect 6429 1004 6435 1096
rect 6509 984 6515 1336
rect 6525 1324 6531 1476
rect 6573 1384 6579 1837
rect 6589 1804 6595 1856
rect 6541 1324 6547 1336
rect 6573 1324 6579 1356
rect 6525 1164 6531 1236
rect 6573 1144 6579 1316
rect 6525 1104 6531 1136
rect 6573 1104 6579 1136
rect 6468 917 6483 923
rect 6413 723 6419 916
rect 6429 744 6435 896
rect 6461 724 6467 836
rect 6413 717 6428 723
rect 6365 544 6371 616
rect 6349 524 6355 536
rect 6365 524 6371 536
rect 6253 384 6259 516
rect 6221 337 6243 343
rect 5981 304 5987 336
rect 6045 144 6051 276
rect 6077 144 6083 156
rect 6093 124 6099 336
rect 6109 302 6115 336
rect 6196 317 6211 323
rect 6189 304 6195 316
rect 6141 224 6147 276
rect 6013 104 6019 118
rect 6141 104 6147 176
rect 6189 144 6195 276
rect 6205 124 6211 317
rect 5501 62 5507 100
rect 6237 84 6243 337
rect 6285 284 6291 416
rect 6301 304 6307 436
rect 6317 304 6323 316
rect 6301 284 6307 296
rect 6253 104 6259 196
rect 6285 164 6291 276
rect 6333 184 6339 436
rect 6365 384 6371 436
rect 6381 424 6387 676
rect 6397 463 6403 636
rect 6397 457 6419 463
rect 6349 164 6355 336
rect 6365 304 6371 376
rect 6381 364 6387 376
rect 6381 304 6387 356
rect 6365 184 6371 256
rect 6397 164 6403 436
rect 6413 304 6419 457
rect 6429 204 6435 536
rect 6461 484 6467 536
rect 6477 524 6483 917
rect 6541 664 6547 1036
rect 6589 964 6595 1756
rect 6605 1504 6611 1816
rect 6621 1503 6627 1816
rect 6637 1524 6643 1956
rect 6653 1904 6659 2136
rect 6717 2124 6723 2136
rect 6717 1924 6723 1936
rect 6660 1897 6668 1903
rect 6653 1824 6659 1896
rect 6717 1784 6723 1836
rect 6733 1824 6739 2436
rect 6749 1804 6755 2276
rect 6781 1944 6787 3456
rect 6797 2004 6803 3436
rect 6813 3204 6819 3316
rect 6877 3304 6883 3376
rect 6861 3124 6867 3136
rect 6813 2984 6819 3016
rect 6861 2064 6867 2236
rect 6829 1984 6835 2036
rect 6765 1904 6771 1916
rect 6877 1884 6883 1896
rect 6781 1844 6787 1876
rect 6717 1744 6723 1756
rect 6813 1744 6819 1836
rect 6685 1524 6691 1556
rect 6717 1524 6723 1736
rect 6813 1662 6819 1700
rect 6829 1684 6835 1816
rect 6621 1497 6643 1503
rect 6637 1484 6643 1497
rect 6637 1344 6643 1476
rect 6701 1384 6707 1456
rect 6605 1184 6611 1296
rect 6573 924 6579 936
rect 6573 684 6579 916
rect 6541 583 6547 656
rect 6541 577 6563 583
rect 6477 304 6483 336
rect 6493 304 6499 536
rect 6541 524 6547 556
rect 6557 544 6563 577
rect 6605 544 6611 1096
rect 6637 784 6643 918
rect 6669 803 6675 1116
rect 6717 1084 6723 1376
rect 6749 1104 6755 1196
rect 6653 797 6675 803
rect 6653 524 6659 797
rect 6701 784 6707 876
rect 6685 664 6691 676
rect 6685 544 6691 656
rect 6669 524 6675 536
rect 6509 484 6515 496
rect 6589 444 6595 516
rect 6541 324 6547 336
rect 6605 324 6611 516
rect 6637 464 6643 516
rect 6621 324 6627 436
rect 6637 364 6643 456
rect 6669 384 6675 516
rect 6685 504 6691 516
rect 6669 324 6675 356
rect 6509 304 6515 316
rect 6493 284 6499 296
rect 6429 184 6435 196
rect 6285 144 6291 156
rect 6301 124 6307 156
rect 6413 144 6419 176
rect 6493 144 6499 216
rect 6541 184 6547 316
rect 6605 304 6611 316
rect 6589 284 6595 296
rect 6621 284 6627 296
rect 6557 124 6563 236
rect 6701 144 6707 756
rect 6717 684 6723 1076
rect 6765 844 6771 1636
rect 6845 1624 6851 1796
rect 6781 1504 6787 1516
rect 6813 1244 6819 1616
rect 6829 1364 6835 1456
rect 6781 1104 6787 1116
rect 6797 1104 6803 1116
rect 6813 1044 6819 1096
rect 6717 504 6723 656
rect 6781 584 6787 1036
rect 6829 1004 6835 1036
rect 6733 544 6739 556
rect 6717 384 6723 476
rect 6717 304 6723 316
rect 6749 304 6755 536
rect 6765 504 6771 516
rect 6797 444 6803 916
rect 6829 584 6835 836
rect 6845 764 6851 1236
rect 6861 984 6867 1096
rect 6877 984 6883 1096
rect 6845 464 6851 736
rect 6861 524 6867 556
rect 6813 384 6819 456
rect 6845 284 6851 336
rect 6733 264 6739 276
rect 6877 264 6883 536
rect 6813 184 6819 236
rect 6877 144 6883 256
rect 6701 124 6707 136
rect 6541 104 6547 116
rect 6365 84 6371 96
rect 5869 -17 5875 36
rect 5405 -23 5427 -17
rect 5853 -23 5875 -17
<< m3contact >>
rect 2638 5006 2646 5014
rect 2652 5006 2660 5014
rect 2666 5006 2674 5014
rect 2236 4996 2244 5004
rect 4844 4996 4852 5004
rect 4844 4976 4852 4984
rect 4876 4976 4884 4984
rect 860 4956 868 4964
rect 1612 4956 1620 4964
rect 1836 4956 1844 4964
rect 2220 4956 2228 4964
rect 2396 4956 2404 4964
rect 3148 4956 3156 4964
rect 3628 4956 3636 4964
rect 3868 4956 3876 4964
rect 4300 4956 4308 4964
rect 4620 4956 4628 4964
rect 5084 4956 5092 4964
rect 5116 4956 5124 4964
rect 5324 4956 5332 4964
rect 140 4936 148 4944
rect 348 4936 356 4944
rect 588 4936 596 4944
rect 252 4916 260 4924
rect 492 4916 500 4924
rect 364 4896 372 4904
rect 396 4896 404 4904
rect 412 4896 420 4904
rect 108 4816 116 4824
rect 140 4816 148 4824
rect 28 4476 36 4484
rect 12 4436 20 4444
rect 12 4316 20 4324
rect 76 4116 84 4124
rect 12 3896 20 3904
rect 76 3716 84 3724
rect 76 3476 84 3484
rect 76 3316 84 3324
rect 396 4756 404 4764
rect 332 4716 340 4724
rect 364 4716 372 4724
rect 876 4936 884 4944
rect 1100 4936 1108 4944
rect 1484 4936 1492 4944
rect 1612 4936 1620 4944
rect 860 4896 868 4904
rect 876 4876 884 4884
rect 700 4856 708 4864
rect 780 4836 788 4844
rect 716 4736 724 4744
rect 780 4736 788 4744
rect 844 4736 852 4744
rect 428 4716 436 4724
rect 684 4716 692 4724
rect 220 4676 228 4684
rect 380 4676 388 4684
rect 188 4596 196 4604
rect 348 4536 356 4544
rect 140 4496 148 4504
rect 140 4302 148 4304
rect 140 4296 148 4302
rect 220 4496 228 4504
rect 204 4456 212 4464
rect 300 4516 308 4524
rect 268 4436 276 4444
rect 236 4416 244 4424
rect 268 4316 276 4324
rect 732 4696 740 4704
rect 828 4696 836 4704
rect 460 4676 468 4684
rect 428 4556 436 4564
rect 716 4656 724 4664
rect 588 4636 596 4644
rect 556 4596 564 4604
rect 460 4536 468 4544
rect 444 4516 452 4524
rect 316 4496 324 4504
rect 412 4496 420 4504
rect 428 4496 436 4504
rect 236 4296 244 4304
rect 396 4476 404 4484
rect 396 4436 404 4444
rect 364 4416 372 4424
rect 412 4376 420 4384
rect 428 4356 436 4364
rect 444 4336 452 4344
rect 348 4296 356 4304
rect 428 4296 436 4304
rect 348 4176 356 4184
rect 220 4156 228 4164
rect 316 4156 324 4164
rect 220 4136 228 4144
rect 268 4136 276 4144
rect 188 4096 196 4104
rect 236 4116 244 4124
rect 268 4096 276 4104
rect 252 4076 260 4084
rect 204 4016 212 4024
rect 236 3976 244 3984
rect 140 3936 148 3944
rect 204 3916 212 3924
rect 252 3916 260 3924
rect 284 4076 292 4084
rect 252 3896 260 3904
rect 332 3896 340 3904
rect 236 3816 244 3824
rect 220 3796 228 3804
rect 188 3736 196 3744
rect 188 3596 196 3604
rect 300 3876 308 3884
rect 300 3816 308 3824
rect 332 3756 340 3764
rect 284 3736 292 3744
rect 428 4156 436 4164
rect 492 4496 500 4504
rect 684 4636 692 4644
rect 668 4516 676 4524
rect 556 4456 564 4464
rect 556 4356 564 4364
rect 572 4296 580 4304
rect 460 4236 468 4244
rect 508 4156 516 4164
rect 508 4136 516 4144
rect 524 4116 532 4124
rect 396 4076 404 4084
rect 476 4056 484 4064
rect 636 4496 644 4504
rect 700 4496 708 4504
rect 732 4516 740 4524
rect 716 4456 724 4464
rect 652 4376 660 4384
rect 700 4376 708 4384
rect 668 4316 676 4324
rect 652 4296 660 4304
rect 556 4176 564 4184
rect 540 4036 548 4044
rect 636 4256 644 4264
rect 652 4196 660 4204
rect 588 4116 596 4124
rect 620 4116 628 4124
rect 684 4116 692 4124
rect 572 4096 580 4104
rect 636 4096 644 4104
rect 652 4096 660 4104
rect 620 4056 628 4064
rect 508 4016 516 4024
rect 556 4016 564 4024
rect 428 3976 436 3984
rect 364 3956 372 3964
rect 476 3936 484 3944
rect 428 3916 436 3924
rect 492 3916 500 3924
rect 396 3896 404 3904
rect 476 3896 484 3904
rect 380 3876 388 3884
rect 636 3996 644 4004
rect 524 3896 532 3904
rect 588 3896 596 3904
rect 572 3876 580 3884
rect 604 3876 612 3884
rect 492 3836 500 3844
rect 476 3776 484 3784
rect 540 3776 548 3784
rect 460 3756 468 3764
rect 300 3716 308 3724
rect 252 3556 260 3564
rect 348 3556 356 3564
rect 236 3516 244 3524
rect 236 3496 244 3504
rect 300 3536 308 3544
rect 268 3516 276 3524
rect 348 3496 356 3504
rect 268 3476 276 3484
rect 348 3476 356 3484
rect 252 3456 260 3464
rect 332 3456 340 3464
rect 316 3436 324 3444
rect 524 3736 532 3744
rect 572 3756 580 3764
rect 444 3716 452 3724
rect 428 3696 436 3704
rect 380 3576 388 3584
rect 428 3596 436 3604
rect 460 3576 468 3584
rect 396 3536 404 3544
rect 380 3516 388 3524
rect 556 3696 564 3704
rect 588 3556 596 3564
rect 428 3496 436 3504
rect 476 3496 484 3504
rect 524 3496 532 3504
rect 556 3496 564 3504
rect 364 3436 372 3444
rect 444 3436 452 3444
rect 556 3396 564 3404
rect 412 3376 420 3384
rect 540 3376 548 3384
rect 396 3336 404 3344
rect 492 3356 500 3364
rect 476 3336 484 3344
rect 252 3316 260 3324
rect 300 3316 308 3324
rect 332 3316 340 3324
rect 396 3316 404 3324
rect 76 3296 84 3304
rect 108 3296 116 3304
rect 124 3296 132 3304
rect 204 3296 212 3304
rect 236 3276 244 3284
rect 268 3276 276 3284
rect 284 3096 292 3104
rect 140 3076 148 3084
rect 172 3056 180 3064
rect 236 3016 244 3024
rect 156 2956 164 2964
rect 204 2936 212 2944
rect 28 2916 36 2924
rect 140 2916 148 2924
rect 12 2896 20 2904
rect 60 2896 68 2904
rect 108 2876 116 2884
rect 172 2876 180 2884
rect 172 2776 180 2784
rect 396 3296 404 3304
rect 348 3276 356 3284
rect 332 3116 340 3124
rect 380 3156 388 3164
rect 460 3156 468 3164
rect 364 3096 372 3104
rect 316 3016 324 3024
rect 284 2956 292 2964
rect 268 2936 276 2944
rect 412 3116 420 3124
rect 428 3076 436 3084
rect 540 3336 548 3344
rect 668 3996 676 4004
rect 732 4436 740 4444
rect 764 4656 772 4664
rect 828 4656 836 4664
rect 812 4636 820 4644
rect 940 4896 948 4904
rect 892 4836 900 4844
rect 956 4876 964 4884
rect 1228 4836 1236 4844
rect 940 4756 948 4764
rect 1118 4806 1126 4814
rect 1132 4806 1140 4814
rect 1146 4806 1154 4814
rect 988 4736 996 4744
rect 1052 4696 1060 4704
rect 924 4676 932 4684
rect 860 4616 868 4624
rect 844 4596 852 4604
rect 780 4556 788 4564
rect 876 4556 884 4564
rect 860 4536 868 4544
rect 764 4336 772 4344
rect 844 4496 852 4504
rect 860 4456 868 4464
rect 844 4316 852 4324
rect 748 4276 756 4284
rect 780 4276 788 4284
rect 844 4296 852 4304
rect 796 4256 804 4264
rect 876 4256 884 4264
rect 732 4216 740 4224
rect 1116 4656 1124 4664
rect 988 4636 996 4644
rect 1004 4616 1012 4624
rect 988 4556 996 4564
rect 1100 4536 1108 4544
rect 1068 4516 1076 4524
rect 972 4436 980 4444
rect 908 4196 916 4204
rect 988 4316 996 4324
rect 908 4176 916 4184
rect 972 4176 980 4184
rect 796 4136 804 4144
rect 844 4136 852 4144
rect 1036 4436 1044 4444
rect 1004 4196 1012 4204
rect 988 4136 996 4144
rect 1036 4136 1044 4144
rect 924 4116 932 4124
rect 940 4076 948 4084
rect 796 4056 804 4064
rect 780 4036 788 4044
rect 780 3916 788 3924
rect 668 3856 676 3864
rect 652 3776 660 3784
rect 636 3756 644 3764
rect 668 3756 676 3764
rect 652 3736 660 3744
rect 892 3956 900 3964
rect 812 3936 820 3944
rect 844 3916 852 3924
rect 988 4016 996 4024
rect 1020 3996 1028 4004
rect 956 3956 964 3964
rect 700 3876 708 3884
rect 796 3836 804 3844
rect 700 3756 708 3764
rect 700 3736 708 3744
rect 748 3816 756 3824
rect 828 3896 836 3904
rect 876 3876 884 3884
rect 1036 3956 1044 3964
rect 972 3856 980 3864
rect 828 3756 836 3764
rect 812 3736 820 3744
rect 684 3716 692 3724
rect 796 3716 804 3724
rect 620 3696 628 3704
rect 732 3696 740 3704
rect 620 3676 628 3684
rect 668 3656 676 3664
rect 700 3556 708 3564
rect 684 3536 692 3544
rect 652 3516 660 3524
rect 636 3496 644 3504
rect 620 3476 628 3484
rect 604 3396 612 3404
rect 700 3516 708 3524
rect 716 3516 724 3524
rect 780 3656 788 3664
rect 748 3516 756 3524
rect 780 3496 788 3504
rect 732 3476 740 3484
rect 716 3456 724 3464
rect 668 3416 676 3424
rect 764 3436 772 3444
rect 700 3356 708 3364
rect 716 3336 724 3344
rect 796 3336 804 3344
rect 620 3316 628 3324
rect 588 3296 596 3304
rect 652 3296 660 3304
rect 860 3496 868 3504
rect 956 3796 964 3804
rect 908 3716 916 3724
rect 956 3716 964 3724
rect 940 3656 948 3664
rect 940 3636 948 3644
rect 892 3516 900 3524
rect 876 3456 884 3464
rect 828 3416 836 3424
rect 828 3376 836 3384
rect 844 3296 852 3304
rect 700 3276 708 3284
rect 604 3136 612 3144
rect 748 3176 756 3184
rect 668 3156 676 3164
rect 508 3116 516 3124
rect 924 3576 932 3584
rect 908 3396 916 3404
rect 1036 3696 1044 3704
rect 1004 3676 1012 3684
rect 972 3636 980 3644
rect 1036 3636 1044 3644
rect 956 3556 964 3564
rect 1004 3516 1012 3524
rect 940 3416 948 3424
rect 908 3376 916 3384
rect 924 3376 932 3384
rect 924 3336 932 3344
rect 940 3236 948 3244
rect 908 3116 916 3124
rect 876 3096 884 3104
rect 556 3076 564 3084
rect 604 3076 612 3084
rect 556 3056 564 3064
rect 444 2936 452 2944
rect 540 2936 548 2944
rect 300 2916 308 2924
rect 348 2916 356 2924
rect 428 2916 436 2924
rect 476 2916 484 2924
rect 60 2676 68 2684
rect 140 2676 148 2684
rect 172 2656 180 2664
rect 204 2616 212 2624
rect 380 2896 388 2904
rect 332 2876 340 2884
rect 428 2876 436 2884
rect 332 2776 340 2784
rect 524 2876 532 2884
rect 476 2776 484 2784
rect 380 2696 388 2704
rect 364 2656 372 2664
rect 316 2636 324 2644
rect 124 2596 132 2604
rect 108 2556 116 2564
rect 140 2556 148 2564
rect 60 2536 68 2544
rect 12 2496 20 2504
rect 44 2496 52 2504
rect 268 2616 276 2624
rect 348 2536 356 2544
rect 444 2516 452 2524
rect 188 2296 196 2304
rect 428 2276 436 2284
rect 28 2176 36 2184
rect 188 2256 196 2264
rect 236 2256 244 2264
rect 268 2176 276 2184
rect 396 2176 404 2184
rect 140 2156 148 2164
rect 92 2136 100 2144
rect 236 2136 244 2144
rect 12 2096 20 2104
rect 108 2036 116 2044
rect 92 2016 100 2024
rect 140 2016 148 2024
rect 92 1916 100 1924
rect 12 1896 20 1904
rect 60 1896 68 1904
rect 76 1896 84 1904
rect 60 1736 68 1744
rect 28 1516 36 1524
rect 92 1856 100 1864
rect 156 1876 164 1884
rect 140 1836 148 1844
rect 300 1856 308 1864
rect 332 1856 340 1864
rect 172 1756 180 1764
rect 140 1736 148 1744
rect 508 2656 516 2664
rect 1276 4916 1284 4924
rect 1356 4916 1364 4924
rect 1340 4836 1348 4844
rect 1372 4836 1380 4844
rect 1324 4716 1332 4724
rect 1484 4816 1492 4824
rect 1260 4696 1268 4704
rect 1308 4696 1316 4704
rect 1388 4696 1396 4704
rect 1244 4656 1252 4664
rect 1196 4616 1204 4624
rect 1180 4556 1188 4564
rect 1292 4656 1300 4664
rect 1276 4636 1284 4644
rect 1340 4636 1348 4644
rect 1292 4616 1300 4624
rect 1292 4556 1300 4564
rect 1244 4536 1252 4544
rect 1116 4456 1124 4464
rect 1164 4436 1172 4444
rect 1118 4406 1126 4414
rect 1132 4406 1140 4414
rect 1146 4406 1154 4414
rect 1276 4516 1284 4524
rect 1276 4456 1284 4464
rect 1212 4296 1220 4304
rect 1228 4296 1236 4304
rect 1164 4136 1172 4144
rect 1148 4096 1156 4104
rect 1148 4056 1156 4064
rect 1118 4006 1126 4014
rect 1132 4006 1140 4014
rect 1146 4006 1154 4014
rect 1196 4216 1204 4224
rect 1244 4136 1252 4144
rect 1404 4636 1412 4644
rect 1468 4636 1476 4644
rect 1660 4916 1668 4924
rect 1516 4896 1524 4904
rect 1564 4896 1572 4904
rect 1644 4896 1652 4904
rect 1548 4876 1556 4884
rect 1676 4876 1684 4884
rect 1756 4856 1764 4864
rect 1596 4836 1604 4844
rect 1500 4616 1508 4624
rect 1644 4736 1652 4744
rect 1676 4736 1684 4744
rect 1724 4716 1732 4724
rect 1804 4716 1812 4724
rect 1628 4696 1636 4704
rect 1692 4696 1700 4704
rect 1596 4676 1604 4684
rect 1644 4656 1652 4664
rect 1564 4636 1572 4644
rect 1628 4536 1636 4544
rect 1340 4296 1348 4304
rect 1308 4156 1316 4164
rect 1292 4116 1300 4124
rect 1276 4076 1284 4084
rect 1228 3956 1236 3964
rect 1260 3956 1268 3964
rect 1084 3936 1092 3944
rect 1132 3936 1140 3944
rect 1180 3936 1188 3944
rect 1196 3936 1204 3944
rect 1084 3896 1092 3904
rect 1084 3716 1092 3724
rect 1212 3916 1220 3924
rect 1180 3896 1188 3904
rect 1164 3836 1172 3844
rect 1148 3816 1156 3824
rect 1116 3696 1124 3704
rect 1196 3876 1204 3884
rect 1196 3716 1204 3724
rect 1148 3676 1156 3684
rect 1164 3676 1172 3684
rect 1180 3676 1188 3684
rect 1084 3656 1092 3664
rect 1068 3576 1076 3584
rect 1068 3536 1076 3544
rect 1052 3476 1060 3484
rect 972 3436 980 3444
rect 1020 3436 1028 3444
rect 1036 3436 1044 3444
rect 1118 3606 1126 3614
rect 1132 3606 1140 3614
rect 1146 3606 1154 3614
rect 1244 3936 1252 3944
rect 1292 3956 1300 3964
rect 1292 3916 1300 3924
rect 1276 3896 1284 3904
rect 1276 3876 1284 3884
rect 1340 4216 1348 4224
rect 1372 4396 1380 4404
rect 1452 4516 1460 4524
rect 1420 4496 1428 4504
rect 1388 4356 1396 4364
rect 1356 4156 1364 4164
rect 1372 4136 1380 4144
rect 1324 4036 1332 4044
rect 1324 3956 1332 3964
rect 1372 4096 1380 4104
rect 1356 3936 1364 3944
rect 1340 3896 1348 3904
rect 1292 3856 1300 3864
rect 1276 3836 1284 3844
rect 1292 3836 1300 3844
rect 1356 3816 1364 3824
rect 1404 4196 1412 4204
rect 1788 4696 1796 4704
rect 1772 4676 1780 4684
rect 1804 4676 1812 4684
rect 2012 4936 2020 4944
rect 2044 4936 2052 4944
rect 2252 4936 2260 4944
rect 2492 4936 2500 4944
rect 2748 4936 2756 4944
rect 2924 4936 2932 4944
rect 3036 4936 3044 4944
rect 3340 4936 3348 4944
rect 3452 4936 3460 4944
rect 1868 4916 1876 4924
rect 1980 4916 1988 4924
rect 2140 4916 2148 4924
rect 2364 4916 2372 4924
rect 2060 4836 2068 4844
rect 1948 4696 1956 4704
rect 2156 4696 2164 4704
rect 2412 4696 2420 4704
rect 1740 4656 1748 4664
rect 1836 4656 1844 4664
rect 1820 4636 1828 4644
rect 1724 4576 1732 4584
rect 1756 4576 1764 4584
rect 1708 4536 1716 4544
rect 1500 4516 1508 4524
rect 1548 4516 1556 4524
rect 1628 4516 1636 4524
rect 1644 4516 1652 4524
rect 1484 4396 1492 4404
rect 1516 4336 1524 4344
rect 1468 4316 1476 4324
rect 1612 4496 1620 4504
rect 1564 4476 1572 4484
rect 1548 4376 1556 4384
rect 1532 4296 1540 4304
rect 1532 4276 1540 4284
rect 1548 4176 1556 4184
rect 1516 4136 1524 4144
rect 1500 4116 1508 4124
rect 1388 3996 1396 4004
rect 1484 4076 1492 4084
rect 1548 4096 1556 4104
rect 1404 3976 1412 3984
rect 1388 3956 1396 3964
rect 1436 3936 1444 3944
rect 1436 3916 1444 3924
rect 1404 3896 1412 3904
rect 1340 3756 1348 3764
rect 1372 3756 1380 3764
rect 1228 3736 1236 3744
rect 1260 3736 1268 3744
rect 1228 3696 1236 3704
rect 1228 3656 1236 3664
rect 1164 3576 1172 3584
rect 1212 3576 1220 3584
rect 1148 3536 1156 3544
rect 1148 3496 1156 3504
rect 1196 3536 1204 3544
rect 1276 3616 1284 3624
rect 1260 3516 1268 3524
rect 1340 3676 1348 3684
rect 1388 3736 1396 3744
rect 1484 3896 1492 3904
rect 1452 3876 1460 3884
rect 1484 3876 1492 3884
rect 1436 3856 1444 3864
rect 1500 3856 1508 3864
rect 1516 3816 1524 3824
rect 1452 3796 1460 3804
rect 1500 3796 1508 3804
rect 1484 3776 1492 3784
rect 1372 3716 1380 3724
rect 1324 3556 1332 3564
rect 1308 3516 1316 3524
rect 1180 3496 1188 3504
rect 1212 3496 1220 3504
rect 1260 3496 1268 3504
rect 1132 3456 1140 3464
rect 988 3356 996 3364
rect 1036 3356 1044 3364
rect 1084 3356 1092 3364
rect 1292 3456 1300 3464
rect 1228 3436 1236 3444
rect 1324 3496 1332 3504
rect 1324 3456 1332 3464
rect 1212 3376 1220 3384
rect 1276 3376 1284 3384
rect 1116 3316 1124 3324
rect 1148 3318 1156 3324
rect 1148 3316 1156 3318
rect 972 3276 980 3284
rect 1020 3276 1028 3284
rect 972 3216 980 3224
rect 1036 3236 1044 3244
rect 1004 3116 1012 3124
rect 1020 3096 1028 3104
rect 956 3076 964 3084
rect 860 3056 868 3064
rect 604 2936 612 2944
rect 748 2936 756 2944
rect 604 2916 612 2924
rect 956 2936 964 2944
rect 972 2936 980 2944
rect 940 2896 948 2904
rect 780 2856 788 2864
rect 684 2776 692 2784
rect 588 2716 596 2724
rect 652 2716 660 2724
rect 876 2696 884 2704
rect 556 2676 564 2684
rect 572 2676 580 2684
rect 604 2676 612 2684
rect 540 2596 548 2604
rect 508 2536 516 2544
rect 668 2636 676 2644
rect 652 2596 660 2604
rect 700 2596 708 2604
rect 844 2636 852 2644
rect 892 2596 900 2604
rect 1356 3556 1364 3564
rect 1388 3516 1396 3524
rect 1500 3576 1508 3584
rect 1420 3476 1428 3484
rect 1356 3436 1364 3444
rect 1340 3336 1348 3344
rect 1180 3296 1188 3304
rect 1118 3206 1126 3214
rect 1132 3206 1140 3214
rect 1146 3206 1154 3214
rect 1100 3076 1108 3084
rect 1132 3056 1140 3064
rect 1116 2976 1124 2984
rect 1084 2936 1092 2944
rect 1020 2916 1028 2924
rect 1052 2916 1060 2924
rect 1004 2896 1012 2904
rect 1068 2896 1076 2904
rect 1052 2876 1060 2884
rect 1118 2806 1126 2814
rect 1132 2806 1140 2814
rect 1146 2806 1154 2814
rect 1004 2736 1012 2744
rect 1084 2716 1092 2724
rect 1116 2696 1124 2704
rect 1116 2676 1124 2684
rect 1084 2656 1092 2664
rect 1340 3236 1348 3244
rect 1404 3456 1412 3464
rect 1420 3436 1428 3444
rect 1468 3416 1476 3424
rect 1500 3376 1508 3384
rect 1420 3356 1428 3364
rect 1708 4516 1716 4524
rect 1692 4396 1700 4404
rect 1612 4356 1620 4364
rect 1692 4336 1700 4344
rect 1596 4316 1604 4324
rect 1692 4316 1700 4324
rect 1596 4296 1604 4304
rect 1628 4296 1636 4304
rect 1596 4236 1604 4244
rect 1580 3916 1588 3924
rect 1580 3796 1588 3804
rect 1564 3536 1572 3544
rect 1548 3516 1556 3524
rect 1644 4276 1652 4284
rect 2300 4676 2308 4684
rect 2316 4676 2324 4684
rect 1980 4616 1988 4624
rect 1852 4536 1860 4544
rect 2620 4916 2628 4924
rect 2908 4916 2916 4924
rect 2524 4816 2532 4824
rect 2812 4816 2820 4824
rect 2764 4716 2772 4724
rect 2732 4696 2740 4704
rect 2764 4696 2772 4704
rect 2524 4676 2532 4684
rect 2204 4616 2212 4624
rect 2028 4576 2036 4584
rect 1996 4536 2004 4544
rect 1740 4516 1748 4524
rect 1804 4518 1812 4524
rect 1804 4516 1812 4518
rect 1964 4516 1972 4524
rect 2092 4516 2100 4524
rect 2140 4516 2148 4524
rect 2188 4516 2196 4524
rect 1740 4496 1748 4504
rect 1852 4496 1860 4504
rect 1820 4476 1828 4484
rect 1788 4356 1796 4364
rect 1772 4316 1780 4324
rect 1932 4476 1940 4484
rect 1804 4296 1812 4304
rect 1676 4196 1684 4204
rect 1644 4116 1652 4124
rect 1692 4156 1700 4164
rect 1708 4136 1716 4144
rect 1788 4276 1796 4284
rect 1740 4196 1748 4204
rect 1804 4256 1812 4264
rect 1740 4096 1748 4104
rect 1724 4056 1732 4064
rect 1980 4396 1988 4404
rect 1900 4296 1908 4304
rect 2012 4296 2020 4304
rect 2108 4296 2116 4304
rect 1868 4276 1876 4284
rect 1916 4276 1924 4284
rect 1852 4256 1860 4264
rect 1884 4256 1892 4264
rect 1932 4256 1940 4264
rect 1852 4236 1860 4244
rect 2188 4376 2196 4384
rect 2172 4316 2180 4324
rect 2444 4576 2452 4584
rect 2220 4476 2228 4484
rect 2268 4476 2276 4484
rect 2156 4276 2164 4284
rect 2140 4256 2148 4264
rect 2172 4256 2180 4264
rect 2316 4376 2324 4384
rect 2252 4336 2260 4344
rect 2284 4316 2292 4324
rect 2252 4296 2260 4304
rect 2060 4236 2068 4244
rect 1820 4176 1828 4184
rect 2092 4216 2100 4224
rect 2124 4196 2132 4204
rect 2156 4196 2164 4204
rect 1836 4136 1844 4144
rect 1948 4136 1956 4144
rect 1804 4116 1812 4124
rect 1788 3996 1796 4004
rect 1772 3956 1780 3964
rect 1724 3916 1732 3924
rect 1756 3916 1764 3924
rect 1884 4096 1892 4104
rect 1884 3936 1892 3944
rect 1868 3916 1876 3924
rect 1676 3876 1684 3884
rect 1772 3876 1780 3884
rect 1660 3836 1668 3844
rect 1628 3816 1636 3824
rect 1660 3816 1668 3824
rect 1612 3716 1620 3724
rect 1628 3696 1636 3704
rect 1692 3796 1700 3804
rect 1804 3816 1812 3824
rect 1884 3876 1892 3884
rect 1868 3856 1876 3864
rect 1932 4036 1940 4044
rect 2012 4016 2020 4024
rect 2044 4016 2052 4024
rect 1932 3916 1940 3924
rect 2012 3916 2020 3924
rect 1948 3896 1956 3904
rect 1996 3896 2004 3904
rect 1996 3876 2004 3884
rect 1964 3856 1972 3864
rect 1900 3836 1908 3844
rect 1948 3836 1956 3844
rect 1852 3776 1860 3784
rect 1868 3776 1876 3784
rect 1964 3776 1972 3784
rect 1772 3756 1780 3764
rect 1740 3736 1748 3744
rect 1788 3736 1796 3744
rect 1708 3716 1716 3724
rect 1756 3716 1764 3724
rect 1836 3716 1844 3724
rect 1660 3616 1668 3624
rect 1628 3536 1636 3544
rect 1580 3516 1588 3524
rect 1596 3516 1604 3524
rect 1644 3516 1652 3524
rect 1692 3556 1700 3564
rect 1676 3496 1684 3504
rect 1932 3756 1940 3764
rect 2204 4136 2212 4144
rect 2348 4316 2356 4324
rect 2268 4136 2276 4144
rect 2236 4116 2244 4124
rect 2638 4606 2646 4614
rect 2652 4606 2660 4614
rect 2666 4606 2674 4614
rect 2796 4656 2804 4664
rect 2812 4596 2820 4604
rect 2828 4556 2836 4564
rect 2796 4536 2804 4544
rect 3020 4916 3028 4924
rect 3660 4936 3668 4944
rect 4060 4936 4068 4944
rect 4332 4936 4340 4944
rect 4396 4936 4404 4944
rect 4652 4936 4660 4944
rect 4764 4936 4772 4944
rect 3228 4916 3236 4924
rect 3548 4916 3556 4924
rect 3628 4916 3636 4924
rect 4028 4916 4036 4924
rect 3308 4836 3316 4844
rect 3340 4836 3348 4844
rect 4012 4836 4020 4844
rect 3324 4816 3332 4824
rect 3260 4736 3268 4744
rect 3164 4716 3172 4724
rect 3196 4716 3204 4724
rect 3308 4716 3316 4724
rect 3004 4696 3012 4704
rect 3276 4696 3284 4704
rect 2940 4656 2948 4664
rect 2988 4656 2996 4664
rect 2924 4556 2932 4564
rect 2572 4516 2580 4524
rect 2604 4516 2612 4524
rect 2716 4516 2724 4524
rect 2796 4516 2804 4524
rect 2476 4336 2484 4344
rect 2460 4276 2468 4284
rect 2348 4256 2356 4264
rect 2412 4256 2420 4264
rect 2444 4256 2452 4264
rect 2364 4156 2372 4164
rect 2444 4216 2452 4224
rect 2380 4136 2388 4144
rect 2268 3936 2276 3944
rect 2204 3916 2212 3924
rect 2332 3936 2340 3944
rect 2348 3916 2356 3924
rect 2108 3876 2116 3884
rect 2172 3836 2180 3844
rect 2060 3756 2068 3764
rect 1868 3696 1876 3704
rect 2044 3696 2052 3704
rect 1532 3476 1540 3484
rect 1612 3476 1620 3484
rect 1628 3456 1636 3464
rect 1580 3416 1588 3424
rect 1596 3416 1604 3424
rect 1532 3336 1540 3344
rect 1612 3336 1620 3344
rect 2044 3556 2052 3564
rect 1836 3436 1844 3444
rect 1884 3416 1892 3424
rect 1676 3376 1684 3384
rect 1676 3356 1684 3364
rect 1404 3316 1412 3324
rect 1516 3316 1524 3324
rect 1596 3316 1604 3324
rect 1660 3316 1668 3324
rect 1372 3136 1380 3144
rect 2140 3736 2148 3744
rect 2124 3596 2132 3604
rect 2252 3816 2260 3824
rect 2284 3816 2292 3824
rect 2204 3736 2212 3744
rect 2268 3716 2276 3724
rect 2204 3656 2212 3664
rect 2220 3516 2228 3524
rect 2236 3496 2244 3504
rect 2252 3476 2260 3484
rect 2204 3456 2212 3464
rect 2092 3436 2100 3444
rect 2060 3396 2068 3404
rect 1596 3296 1604 3304
rect 1548 3276 1556 3284
rect 1980 3296 1988 3304
rect 1452 3176 1460 3184
rect 1564 3176 1572 3184
rect 1468 3116 1476 3124
rect 1532 3116 1540 3124
rect 1404 3096 1412 3104
rect 1500 3096 1508 3104
rect 1244 3076 1252 3084
rect 1612 3096 1620 3104
rect 1548 3076 1556 3084
rect 1356 3056 1364 3064
rect 1276 3016 1284 3024
rect 1340 3016 1348 3024
rect 1468 2976 1476 2984
rect 1420 2956 1428 2964
rect 1308 2936 1316 2944
rect 1196 2856 1204 2864
rect 1532 2936 1540 2944
rect 1516 2896 1524 2904
rect 1500 2876 1508 2884
rect 1340 2856 1348 2864
rect 1532 2856 1540 2864
rect 1324 2836 1332 2844
rect 1372 2716 1380 2724
rect 1180 2636 1188 2644
rect 1292 2636 1300 2644
rect 1068 2616 1076 2624
rect 988 2596 996 2604
rect 1036 2596 1044 2604
rect 1244 2596 1252 2604
rect 972 2576 980 2584
rect 1052 2556 1060 2564
rect 1196 2556 1204 2564
rect 828 2536 836 2544
rect 1084 2536 1092 2544
rect 588 2516 596 2524
rect 780 2516 788 2524
rect 508 2496 516 2504
rect 572 2496 580 2504
rect 764 2456 772 2464
rect 652 2316 660 2324
rect 780 2316 788 2324
rect 1118 2406 1126 2414
rect 1132 2406 1140 2414
rect 1146 2406 1154 2414
rect 1004 2316 1012 2324
rect 588 2296 596 2304
rect 764 2296 772 2304
rect 796 2296 804 2304
rect 572 2276 580 2284
rect 620 2256 628 2264
rect 524 2236 532 2244
rect 492 2156 500 2164
rect 588 2156 596 2164
rect 428 2036 436 2044
rect 492 1956 500 1964
rect 572 1936 580 1944
rect 508 1916 516 1924
rect 556 1876 564 1884
rect 476 1856 484 1864
rect 524 1776 532 1784
rect 332 1756 340 1764
rect 380 1756 388 1764
rect 252 1716 260 1724
rect 332 1676 340 1684
rect 92 1616 100 1624
rect 140 1616 148 1624
rect 76 1376 84 1384
rect 28 1116 36 1124
rect 60 1116 68 1124
rect 12 1036 20 1044
rect 12 916 20 924
rect 60 1036 68 1044
rect 284 1576 292 1584
rect 108 1516 116 1524
rect 332 1516 340 1524
rect 348 1516 356 1524
rect 140 1496 148 1504
rect 188 1476 196 1484
rect 124 1316 132 1324
rect 188 1236 196 1244
rect 236 1476 244 1484
rect 300 1476 308 1484
rect 316 1476 324 1484
rect 348 1476 356 1484
rect 316 1456 324 1464
rect 268 1376 276 1384
rect 412 1616 420 1624
rect 444 1556 452 1564
rect 412 1516 420 1524
rect 396 1476 404 1484
rect 428 1476 436 1484
rect 412 1456 420 1464
rect 268 1336 276 1344
rect 348 1336 356 1344
rect 380 1316 388 1324
rect 396 1316 404 1324
rect 236 1296 244 1304
rect 268 1296 276 1304
rect 284 1236 292 1244
rect 220 1116 228 1124
rect 252 1116 260 1124
rect 380 1276 388 1284
rect 364 1116 372 1124
rect 156 1096 164 1104
rect 268 1096 276 1104
rect 332 1096 340 1104
rect 60 676 68 684
rect 92 936 100 944
rect 252 1076 260 1084
rect 172 916 180 924
rect 140 896 148 904
rect 172 896 180 904
rect 316 996 324 1004
rect 268 976 276 984
rect 220 956 228 964
rect 236 936 244 944
rect 204 916 212 924
rect 188 716 196 724
rect 204 696 212 704
rect 300 936 308 944
rect 236 876 244 884
rect 268 856 276 864
rect 252 716 260 724
rect 348 1056 356 1064
rect 428 1076 436 1084
rect 380 976 388 984
rect 364 956 372 964
rect 428 1016 436 1024
rect 428 976 436 984
rect 380 916 388 924
rect 412 916 420 924
rect 348 716 356 724
rect 300 696 308 704
rect 316 676 324 684
rect 396 876 404 884
rect 380 716 388 724
rect 380 696 388 704
rect 92 656 100 664
rect 268 656 276 664
rect 204 636 212 644
rect 92 536 100 544
rect 220 556 228 564
rect 300 556 308 564
rect 268 536 276 544
rect 412 836 420 844
rect 428 716 436 724
rect 604 1876 612 1884
rect 700 2276 708 2284
rect 748 2276 756 2284
rect 668 2256 676 2264
rect 700 2236 708 2244
rect 732 2196 740 2204
rect 812 2196 820 2204
rect 780 2176 788 2184
rect 876 2176 884 2184
rect 684 2036 692 2044
rect 636 1976 644 1984
rect 796 1936 804 1944
rect 716 1916 724 1924
rect 764 1916 772 1924
rect 828 1916 836 1924
rect 636 1896 644 1904
rect 700 1896 708 1904
rect 732 1896 740 1904
rect 620 1856 628 1864
rect 1116 2296 1124 2304
rect 1180 2296 1188 2304
rect 1196 2256 1204 2264
rect 1036 2236 1044 2244
rect 1084 2156 1092 2164
rect 1564 2876 1572 2884
rect 1548 2796 1556 2804
rect 1692 3156 1700 3164
rect 2220 3396 2228 3404
rect 2172 3336 2180 3344
rect 2092 3316 2100 3324
rect 1660 3096 1668 3104
rect 1628 3076 1636 3084
rect 1884 3076 1892 3084
rect 2060 3076 2068 3084
rect 1628 3056 1636 3064
rect 1708 3056 1716 3064
rect 1772 3056 1780 3064
rect 1852 3056 1860 3064
rect 1884 3056 1892 3064
rect 1628 2996 1636 3004
rect 1612 2916 1620 2924
rect 1612 2836 1620 2844
rect 1580 2776 1588 2784
rect 1564 2756 1572 2764
rect 1772 3036 1780 3044
rect 1708 2956 1716 2964
rect 1804 3016 1812 3024
rect 1804 2936 1812 2944
rect 1804 2896 1812 2904
rect 1788 2836 1796 2844
rect 1708 2796 1716 2804
rect 1740 2716 1748 2724
rect 1852 2796 1860 2804
rect 1564 2676 1572 2684
rect 1708 2676 1716 2684
rect 1532 2656 1540 2664
rect 1308 2596 1316 2604
rect 1276 2276 1284 2284
rect 1420 2596 1428 2604
rect 1836 2596 1844 2604
rect 1564 2556 1572 2564
rect 1404 2536 1412 2544
rect 1692 2536 1700 2544
rect 1836 2536 1844 2544
rect 1372 2416 1380 2424
rect 1564 2496 1572 2504
rect 1532 2396 1540 2404
rect 1564 2396 1572 2404
rect 1404 2376 1412 2384
rect 1484 2296 1492 2304
rect 1356 2276 1364 2284
rect 1308 2256 1316 2264
rect 1340 2256 1348 2264
rect 1356 2216 1364 2224
rect 1340 2196 1348 2204
rect 1388 2196 1396 2204
rect 1356 2156 1364 2164
rect 956 2136 964 2144
rect 1244 2136 1252 2144
rect 1676 2516 1684 2524
rect 1804 2516 1812 2524
rect 1676 2416 1684 2424
rect 1676 2376 1684 2384
rect 1596 2316 1604 2324
rect 1676 2336 1684 2344
rect 1596 2276 1604 2284
rect 1756 2276 1764 2284
rect 1740 2256 1748 2264
rect 1564 2236 1572 2244
rect 1740 2236 1748 2244
rect 1548 2176 1556 2184
rect 1580 2216 1588 2224
rect 1500 2156 1508 2164
rect 1564 2156 1572 2164
rect 1052 1956 1060 1964
rect 908 1902 916 1904
rect 908 1896 916 1902
rect 652 1876 660 1884
rect 780 1876 788 1884
rect 844 1876 852 1884
rect 588 1816 596 1824
rect 636 1756 644 1764
rect 700 1856 708 1864
rect 924 1856 932 1864
rect 700 1756 708 1764
rect 588 1736 596 1744
rect 652 1736 660 1744
rect 684 1736 692 1744
rect 556 1696 564 1704
rect 620 1696 628 1704
rect 652 1696 660 1704
rect 556 1676 564 1684
rect 540 1616 548 1624
rect 796 1776 804 1784
rect 892 1736 900 1744
rect 796 1716 804 1724
rect 748 1696 756 1704
rect 908 1636 916 1644
rect 876 1616 884 1624
rect 732 1556 740 1564
rect 796 1556 804 1564
rect 492 1516 500 1524
rect 524 1516 532 1524
rect 588 1516 596 1524
rect 684 1516 692 1524
rect 860 1516 868 1524
rect 556 1496 564 1504
rect 636 1496 644 1504
rect 668 1496 676 1504
rect 540 1436 548 1444
rect 524 1416 532 1424
rect 508 1396 516 1404
rect 492 1376 500 1384
rect 620 1456 628 1464
rect 604 1356 612 1364
rect 540 1336 548 1344
rect 508 1296 516 1304
rect 460 1196 468 1204
rect 588 1316 596 1324
rect 572 1296 580 1304
rect 524 1196 532 1204
rect 556 1116 564 1124
rect 716 1436 724 1444
rect 748 1456 756 1464
rect 732 1416 740 1424
rect 684 1396 692 1404
rect 668 1376 676 1384
rect 636 1336 644 1344
rect 668 1316 676 1324
rect 668 1136 676 1144
rect 716 1376 724 1384
rect 764 1356 772 1364
rect 748 1336 756 1344
rect 716 1296 724 1304
rect 764 1296 772 1304
rect 780 1136 788 1144
rect 764 1116 772 1124
rect 604 1096 612 1104
rect 668 1096 676 1104
rect 716 1096 724 1104
rect 476 1076 484 1084
rect 508 1076 516 1084
rect 460 976 468 984
rect 524 976 532 984
rect 588 976 596 984
rect 476 956 484 964
rect 652 956 660 964
rect 540 936 548 944
rect 636 936 644 944
rect 540 916 548 924
rect 524 876 532 884
rect 508 856 516 864
rect 460 716 468 724
rect 412 556 420 564
rect 508 696 516 704
rect 476 676 484 684
rect 524 636 532 644
rect 508 596 516 604
rect 492 576 500 584
rect 364 536 372 544
rect 444 536 452 544
rect 220 516 228 524
rect 188 496 196 504
rect 252 496 260 504
rect 124 436 132 444
rect 172 436 180 444
rect 28 296 36 304
rect 28 136 36 144
rect 140 276 148 284
rect 332 316 340 324
rect 572 856 580 864
rect 588 856 596 864
rect 556 836 564 844
rect 604 696 612 704
rect 572 616 580 624
rect 540 556 548 564
rect 492 496 500 504
rect 508 496 516 504
rect 412 336 420 344
rect 492 336 500 344
rect 460 316 468 324
rect 412 296 420 304
rect 428 276 436 284
rect 460 276 468 284
rect 380 256 388 264
rect 172 156 180 164
rect 204 156 212 164
rect 172 136 180 144
rect 284 116 292 124
rect 540 516 548 524
rect 700 1076 708 1084
rect 828 1436 836 1444
rect 812 1416 820 1424
rect 860 1416 868 1424
rect 940 1536 948 1544
rect 1036 1516 1044 1524
rect 1052 1496 1060 1504
rect 1118 2006 1126 2014
rect 1132 2006 1140 2014
rect 1146 2006 1154 2014
rect 1404 1916 1412 1924
rect 1500 1896 1508 1904
rect 1084 1876 1092 1884
rect 1196 1876 1204 1884
rect 1084 1696 1092 1704
rect 1116 1656 1124 1664
rect 1180 1776 1188 1784
rect 1228 1856 1236 1864
rect 1420 1876 1428 1884
rect 1340 1756 1348 1764
rect 1372 1736 1380 1744
rect 1196 1716 1204 1724
rect 1228 1716 1236 1724
rect 1180 1696 1188 1704
rect 1212 1676 1220 1684
rect 1148 1636 1156 1644
rect 1118 1606 1126 1614
rect 1132 1606 1140 1614
rect 1146 1606 1154 1614
rect 1244 1696 1252 1704
rect 1404 1756 1412 1764
rect 1500 1756 1508 1764
rect 1468 1716 1476 1724
rect 1244 1636 1252 1644
rect 1228 1576 1236 1584
rect 1196 1516 1204 1524
rect 908 1476 916 1484
rect 924 1456 932 1464
rect 1180 1456 1188 1464
rect 908 1336 916 1344
rect 924 1316 932 1324
rect 988 1316 996 1324
rect 812 1136 820 1144
rect 876 1116 884 1124
rect 1052 1416 1060 1424
rect 1020 1236 1028 1244
rect 988 1176 996 1184
rect 988 1156 996 1164
rect 956 1096 964 1104
rect 876 1076 884 1084
rect 700 1056 708 1064
rect 796 1056 804 1064
rect 796 996 804 1004
rect 716 956 724 964
rect 1020 1116 1028 1124
rect 1020 1096 1028 1104
rect 1020 1056 1028 1064
rect 940 1016 948 1024
rect 988 1016 996 1024
rect 1004 1016 1012 1024
rect 908 956 916 964
rect 684 916 692 924
rect 828 876 836 884
rect 860 836 868 844
rect 972 936 980 944
rect 924 916 932 924
rect 1084 1356 1092 1364
rect 1116 1336 1124 1344
rect 1212 1476 1220 1484
rect 1068 1176 1076 1184
rect 1052 1116 1060 1124
rect 1068 1096 1076 1104
rect 1118 1206 1126 1214
rect 1132 1206 1140 1214
rect 1146 1206 1154 1214
rect 1180 1176 1188 1184
rect 1116 1116 1124 1124
rect 1148 1116 1156 1124
rect 1276 1536 1284 1544
rect 1548 1796 1556 1804
rect 1708 2156 1716 2164
rect 1644 1896 1652 1904
rect 1580 1756 1588 1764
rect 1612 1756 1620 1764
rect 1564 1716 1572 1724
rect 1484 1696 1492 1704
rect 1532 1696 1540 1704
rect 1516 1676 1524 1684
rect 1548 1676 1556 1684
rect 1436 1636 1444 1644
rect 1500 1636 1508 1644
rect 1420 1596 1428 1604
rect 1324 1576 1332 1584
rect 1388 1576 1396 1584
rect 1340 1556 1348 1564
rect 1292 1456 1300 1464
rect 1276 1416 1284 1424
rect 1260 1316 1268 1324
rect 1244 1276 1252 1284
rect 1228 1176 1236 1184
rect 1260 1176 1268 1184
rect 1212 1136 1220 1144
rect 1212 1116 1220 1124
rect 1276 1116 1284 1124
rect 1244 1096 1252 1104
rect 1212 1016 1220 1024
rect 1100 976 1108 984
rect 1180 956 1188 964
rect 1036 916 1044 924
rect 1004 896 1012 904
rect 1260 1036 1268 1044
rect 1276 996 1284 1004
rect 1116 896 1124 904
rect 1228 896 1236 904
rect 924 876 932 884
rect 972 876 980 884
rect 908 836 916 844
rect 876 816 884 824
rect 860 756 868 764
rect 732 716 740 724
rect 636 676 644 684
rect 588 596 596 604
rect 668 636 676 644
rect 652 616 660 624
rect 828 616 836 624
rect 876 616 884 624
rect 892 616 900 624
rect 844 576 852 584
rect 1468 1496 1476 1504
rect 1388 1476 1396 1484
rect 1388 1376 1396 1384
rect 1324 1256 1332 1264
rect 1340 1256 1348 1264
rect 1340 1056 1348 1064
rect 1308 976 1316 984
rect 1340 936 1348 944
rect 1388 1096 1396 1104
rect 1548 1596 1556 1604
rect 1612 1596 1620 1604
rect 1596 1536 1604 1544
rect 1516 1496 1524 1504
rect 1548 1496 1556 1504
rect 1500 1476 1508 1484
rect 1580 1476 1588 1484
rect 1484 1456 1492 1464
rect 1564 1456 1572 1464
rect 1516 1436 1524 1444
rect 1532 1416 1540 1424
rect 1548 1356 1556 1364
rect 1436 1316 1444 1324
rect 1484 1316 1492 1324
rect 1564 1316 1572 1324
rect 1420 1236 1428 1244
rect 1468 1276 1476 1284
rect 1484 1236 1492 1244
rect 1436 1196 1444 1204
rect 1628 1556 1636 1564
rect 1996 2996 2004 3004
rect 1900 2976 1908 2984
rect 2124 3296 2132 3304
rect 2156 3276 2164 3284
rect 2156 3256 2164 3264
rect 2108 3156 2116 3164
rect 2204 3176 2212 3184
rect 2236 3356 2244 3364
rect 2444 4116 2452 4124
rect 2412 4096 2420 4104
rect 2380 3916 2388 3924
rect 2812 4436 2820 4444
rect 2604 4276 2612 4284
rect 2572 4256 2580 4264
rect 2638 4206 2646 4214
rect 2652 4206 2660 4214
rect 2666 4206 2674 4214
rect 2572 4156 2580 4164
rect 2476 4136 2484 4144
rect 2588 4136 2596 4144
rect 2476 4096 2484 4104
rect 2428 3936 2436 3944
rect 2508 3936 2516 3944
rect 2396 3876 2404 3884
rect 2316 3836 2324 3844
rect 2364 3836 2372 3844
rect 2476 3876 2484 3884
rect 2412 3816 2420 3824
rect 2540 4056 2548 4064
rect 2684 4056 2692 4064
rect 2828 4276 2836 4284
rect 2812 4256 2820 4264
rect 2796 4196 2804 4204
rect 2812 4196 2820 4204
rect 2860 4196 2868 4204
rect 2780 4156 2788 4164
rect 3100 4676 3108 4684
rect 3100 4656 3108 4664
rect 3052 4556 3060 4564
rect 3004 4536 3012 4544
rect 3084 4556 3092 4564
rect 3068 4456 3076 4464
rect 2988 4316 2996 4324
rect 3036 4316 3044 4324
rect 2956 4296 2964 4304
rect 3004 4296 3012 4304
rect 2972 4276 2980 4284
rect 2924 4256 2932 4264
rect 2988 4256 2996 4264
rect 2844 4016 2852 4024
rect 2908 4016 2916 4024
rect 2748 3996 2756 4004
rect 2780 3976 2788 3984
rect 2716 3956 2724 3964
rect 2588 3936 2596 3944
rect 2764 3896 2772 3904
rect 2524 3856 2532 3864
rect 2540 3836 2548 3844
rect 2508 3796 2516 3804
rect 2572 3816 2580 3824
rect 2638 3806 2646 3814
rect 2652 3806 2660 3814
rect 2666 3806 2674 3814
rect 2540 3776 2548 3784
rect 2300 3756 2308 3764
rect 2348 3756 2356 3764
rect 2508 3756 2516 3764
rect 2828 3756 2836 3764
rect 2300 3736 2308 3744
rect 2364 3736 2372 3744
rect 2412 3696 2420 3704
rect 2332 3676 2340 3684
rect 2396 3636 2404 3644
rect 2284 3536 2292 3544
rect 2284 3516 2292 3524
rect 2268 3396 2276 3404
rect 2268 3376 2276 3384
rect 2364 3536 2372 3544
rect 2316 3496 2324 3504
rect 2300 3476 2308 3484
rect 2380 3476 2388 3484
rect 2284 3356 2292 3364
rect 3052 4296 3060 4304
rect 3036 4156 3044 4164
rect 3036 4096 3044 4104
rect 2972 4036 2980 4044
rect 3004 3996 3012 4004
rect 3068 4256 3076 4264
rect 3084 4236 3092 4244
rect 3244 4676 3252 4684
rect 3324 4676 3332 4684
rect 3212 4656 3220 4664
rect 3196 4616 3204 4624
rect 3116 4536 3124 4544
rect 3148 4476 3156 4484
rect 3196 4536 3204 4544
rect 3228 4516 3236 4524
rect 3212 4476 3220 4484
rect 3180 4416 3188 4424
rect 3228 4356 3236 4364
rect 3196 4336 3204 4344
rect 3132 4296 3140 4304
rect 3180 4296 3188 4304
rect 3132 4276 3140 4284
rect 3052 3936 3060 3944
rect 3036 3896 3044 3904
rect 2924 3876 2932 3884
rect 2924 3836 2932 3844
rect 2956 3836 2964 3844
rect 3036 3836 3044 3844
rect 2908 3816 2916 3824
rect 2876 3756 2884 3764
rect 2716 3736 2724 3744
rect 2844 3736 2852 3744
rect 2844 3716 2852 3724
rect 2812 3656 2820 3664
rect 2780 3616 2788 3624
rect 2988 3756 2996 3764
rect 2940 3736 2948 3744
rect 2812 3556 2820 3564
rect 2908 3556 2916 3564
rect 2732 3536 2740 3544
rect 2412 3496 2420 3504
rect 2444 3496 2452 3504
rect 2540 3496 2548 3504
rect 2572 3496 2580 3504
rect 2540 3476 2548 3484
rect 2638 3406 2646 3414
rect 2652 3406 2660 3414
rect 2666 3406 2674 3414
rect 2348 3316 2356 3324
rect 2252 3256 2260 3264
rect 2252 3196 2260 3204
rect 2300 3136 2308 3144
rect 2092 3096 2100 3104
rect 2076 3056 2084 3064
rect 2172 3076 2180 3084
rect 2268 3076 2276 3084
rect 2044 3036 2052 3044
rect 2156 3036 2164 3044
rect 2268 3036 2276 3044
rect 2172 2996 2180 3004
rect 2220 3016 2228 3024
rect 2188 2956 2196 2964
rect 2188 2936 2196 2944
rect 1964 2896 1972 2904
rect 2044 2896 2052 2904
rect 2012 2836 2020 2844
rect 2188 2896 2196 2904
rect 2236 2836 2244 2844
rect 2044 2816 2052 2824
rect 2396 3316 2404 3324
rect 2508 3336 2516 3344
rect 2828 3336 2836 3344
rect 2572 3296 2580 3304
rect 2444 3196 2452 3204
rect 2476 3196 2484 3204
rect 2428 3096 2436 3104
rect 2364 3076 2372 3084
rect 2412 3056 2420 3064
rect 2460 3056 2468 3064
rect 2428 3036 2436 3044
rect 2524 3136 2532 3144
rect 2828 3216 2836 3224
rect 2700 3196 2708 3204
rect 2668 3096 2676 3104
rect 2476 3016 2484 3024
rect 2700 3016 2708 3024
rect 2748 3016 2756 3024
rect 2638 3006 2646 3014
rect 2652 3006 2660 3014
rect 2666 3006 2674 3014
rect 2476 2976 2484 2984
rect 2412 2936 2420 2944
rect 2444 2936 2452 2944
rect 2508 2956 2516 2964
rect 2716 2936 2724 2944
rect 2380 2896 2388 2904
rect 2524 2896 2532 2904
rect 2332 2736 2340 2744
rect 1900 2696 1908 2704
rect 2188 2696 2196 2704
rect 2316 2696 2324 2704
rect 1868 2576 1876 2584
rect 1804 2396 1812 2404
rect 1852 2396 1860 2404
rect 1804 2236 1812 2244
rect 2060 2656 2068 2664
rect 2092 2576 2100 2584
rect 2172 2576 2180 2584
rect 1980 2536 1988 2544
rect 2204 2616 2212 2624
rect 2252 2616 2260 2624
rect 2300 2616 2308 2624
rect 2236 2576 2244 2584
rect 2284 2576 2292 2584
rect 2268 2536 2276 2544
rect 2092 2516 2100 2524
rect 2188 2516 2196 2524
rect 2012 2496 2020 2504
rect 2172 2356 2180 2364
rect 2428 2856 2436 2864
rect 2428 2796 2436 2804
rect 2972 3516 2980 3524
rect 3004 3656 3012 3664
rect 2972 3476 2980 3484
rect 2988 3236 2996 3244
rect 2908 3216 2916 3224
rect 2940 3216 2948 3224
rect 2860 3196 2868 3204
rect 2956 3176 2964 3184
rect 3020 3636 3028 3644
rect 3116 4076 3124 4084
rect 3132 4056 3140 4064
rect 3164 4156 3172 4164
rect 3308 4576 3316 4584
rect 3308 4536 3316 4544
rect 3324 4516 3332 4524
rect 3276 4476 3284 4484
rect 3260 4456 3268 4464
rect 3292 4436 3300 4444
rect 3308 4356 3316 4364
rect 3276 4336 3284 4344
rect 3196 4256 3204 4264
rect 3212 4256 3220 4264
rect 3228 4236 3236 4244
rect 3212 4216 3220 4224
rect 3228 4076 3236 4084
rect 3180 3996 3188 4004
rect 3212 3996 3220 4004
rect 3180 3976 3188 3984
rect 3148 3956 3156 3964
rect 3148 3916 3156 3924
rect 3196 3956 3204 3964
rect 3260 4256 3268 4264
rect 3292 4256 3300 4264
rect 3324 4316 3332 4324
rect 3324 4276 3332 4284
rect 3468 4816 3476 4824
rect 3596 4816 3604 4824
rect 3580 4716 3588 4724
rect 3356 4696 3364 4704
rect 3468 4696 3476 4704
rect 3484 4696 3492 4704
rect 3532 4696 3540 4704
rect 3436 4676 3444 4684
rect 3404 4656 3412 4664
rect 3468 4656 3476 4664
rect 3532 4656 3540 4664
rect 3388 4636 3396 4644
rect 3436 4636 3444 4644
rect 3356 4556 3364 4564
rect 3500 4616 3508 4624
rect 3500 4596 3508 4604
rect 3484 4576 3492 4584
rect 3452 4556 3460 4564
rect 3388 4536 3396 4544
rect 3356 4436 3364 4444
rect 3420 4436 3428 4444
rect 3404 4416 3412 4424
rect 3420 4376 3428 4384
rect 3404 4296 3412 4304
rect 3356 4256 3364 4264
rect 3372 4256 3380 4264
rect 3404 4216 3412 4224
rect 3260 4136 3268 4144
rect 3276 4116 3284 4124
rect 3260 3936 3268 3944
rect 3132 3876 3140 3884
rect 3084 3836 3092 3844
rect 3116 3836 3124 3844
rect 3132 3836 3140 3844
rect 3068 3756 3076 3764
rect 3100 3756 3108 3764
rect 3196 3796 3204 3804
rect 3292 3876 3300 3884
rect 3244 3856 3252 3864
rect 3244 3796 3252 3804
rect 3164 3756 3172 3764
rect 3212 3756 3220 3764
rect 3260 3756 3268 3764
rect 3020 3516 3028 3524
rect 3052 3516 3060 3524
rect 3036 3476 3044 3484
rect 3036 3336 3044 3344
rect 3020 3236 3028 3244
rect 2972 3156 2980 3164
rect 3004 3156 3012 3164
rect 2860 3136 2868 3144
rect 2956 3136 2964 3144
rect 2892 3076 2900 3084
rect 2908 3056 2916 3064
rect 2940 2976 2948 2984
rect 2988 3136 2996 3144
rect 3004 3116 3012 3124
rect 3004 3096 3012 3104
rect 2972 2956 2980 2964
rect 2892 2896 2900 2904
rect 2780 2816 2788 2824
rect 2476 2776 2484 2784
rect 2748 2776 2756 2784
rect 2764 2736 2772 2744
rect 2748 2716 2756 2724
rect 2828 2796 2836 2804
rect 2812 2716 2820 2724
rect 2588 2696 2596 2704
rect 2604 2696 2612 2704
rect 2716 2696 2724 2704
rect 2492 2656 2500 2664
rect 2588 2616 2596 2624
rect 2412 2596 2420 2604
rect 2460 2596 2468 2604
rect 2412 2556 2420 2564
rect 2332 2516 2340 2524
rect 2300 2396 2308 2404
rect 2396 2356 2404 2364
rect 2364 2316 2372 2324
rect 2076 2296 2084 2304
rect 2284 2276 2292 2284
rect 1884 2256 1892 2264
rect 2044 2256 2052 2264
rect 1884 2216 1892 2224
rect 2332 2296 2340 2304
rect 2332 2276 2340 2284
rect 2316 2176 2324 2184
rect 1836 2156 1844 2164
rect 2156 2156 2164 2164
rect 1836 2136 1844 2144
rect 1900 2136 1908 2144
rect 2012 2136 2020 2144
rect 2092 1976 2100 1984
rect 1804 1956 1812 1964
rect 1708 1856 1716 1864
rect 1996 1856 2004 1864
rect 2028 1856 2036 1864
rect 1836 1836 1844 1844
rect 1692 1816 1700 1824
rect 1692 1756 1700 1764
rect 1660 1736 1668 1744
rect 1676 1716 1684 1724
rect 1740 1676 1748 1684
rect 1660 1596 1668 1604
rect 1708 1556 1716 1564
rect 1676 1502 1684 1504
rect 1676 1496 1684 1502
rect 1596 1436 1604 1444
rect 1628 1436 1636 1444
rect 1612 1416 1620 1424
rect 1596 1376 1604 1384
rect 1676 1416 1684 1424
rect 1612 1336 1620 1344
rect 1580 1296 1588 1304
rect 1484 1116 1492 1124
rect 1468 1096 1476 1104
rect 1372 1036 1380 1044
rect 1372 956 1380 964
rect 1356 916 1364 924
rect 1308 876 1316 884
rect 1340 896 1348 904
rect 1292 856 1300 864
rect 1324 856 1332 864
rect 1100 836 1108 844
rect 1276 836 1284 844
rect 1292 836 1300 844
rect 972 816 980 824
rect 940 716 948 724
rect 1118 806 1126 814
rect 1132 806 1140 814
rect 1146 806 1154 814
rect 1276 796 1284 804
rect 1324 716 1332 724
rect 1020 696 1028 704
rect 1148 696 1156 704
rect 1068 676 1076 684
rect 940 576 948 584
rect 940 556 948 564
rect 924 536 932 544
rect 604 516 612 524
rect 700 518 708 524
rect 700 516 708 518
rect 876 496 884 504
rect 796 456 804 464
rect 572 336 580 344
rect 588 316 596 324
rect 636 316 644 324
rect 604 296 612 304
rect 588 276 596 284
rect 636 196 644 204
rect 684 196 692 204
rect 652 156 660 164
rect 908 436 916 444
rect 908 416 916 424
rect 956 516 964 524
rect 940 496 948 504
rect 940 436 948 444
rect 1132 656 1140 664
rect 1276 696 1284 704
rect 1228 676 1236 684
rect 1116 636 1124 644
rect 1196 636 1204 644
rect 1228 636 1236 644
rect 1100 596 1108 604
rect 1132 596 1140 604
rect 1132 556 1140 564
rect 1228 556 1236 564
rect 1180 536 1188 544
rect 1052 516 1060 524
rect 1196 516 1204 524
rect 972 416 980 424
rect 1180 416 1188 424
rect 1118 406 1126 414
rect 1132 406 1140 414
rect 1146 406 1154 414
rect 1004 376 1012 384
rect 1036 356 1044 364
rect 1068 356 1076 364
rect 1036 336 1044 344
rect 1260 616 1268 624
rect 1324 656 1332 664
rect 1308 576 1316 584
rect 1260 556 1268 564
rect 1308 536 1316 544
rect 1324 516 1332 524
rect 1388 876 1396 884
rect 1388 836 1396 844
rect 1436 1036 1444 1044
rect 1452 1016 1460 1024
rect 1500 1096 1508 1104
rect 1564 1102 1572 1104
rect 1564 1096 1572 1102
rect 1532 1076 1540 1084
rect 1436 936 1444 944
rect 1468 936 1476 944
rect 1452 916 1460 924
rect 1436 896 1444 904
rect 1436 816 1444 824
rect 1420 776 1428 784
rect 1404 756 1412 764
rect 1420 736 1428 744
rect 1484 876 1492 884
rect 1564 896 1572 904
rect 1500 816 1508 824
rect 1548 796 1556 804
rect 1468 716 1476 724
rect 1532 716 1540 724
rect 1372 696 1380 704
rect 1404 696 1412 704
rect 1436 676 1444 684
rect 1564 736 1572 744
rect 1532 656 1540 664
rect 1500 576 1508 584
rect 1404 556 1412 564
rect 1196 336 1204 344
rect 1100 316 1108 324
rect 1228 316 1236 324
rect 988 296 996 304
rect 1100 296 1108 304
rect 924 276 932 284
rect 988 276 996 284
rect 1052 276 1060 284
rect 972 256 980 264
rect 1116 256 1124 264
rect 940 196 948 204
rect 1036 196 1044 204
rect 908 156 916 164
rect 1004 156 1012 164
rect 1260 256 1268 264
rect 1244 156 1252 164
rect 444 136 452 144
rect 508 136 516 144
rect 844 136 850 144
rect 850 136 852 144
rect 892 136 900 144
rect 1292 476 1300 484
rect 1324 476 1332 484
rect 1388 516 1396 524
rect 1372 496 1380 504
rect 1452 496 1460 504
rect 1356 476 1364 484
rect 1404 476 1412 484
rect 1436 476 1444 484
rect 1356 376 1364 384
rect 1340 296 1348 304
rect 1372 296 1380 304
rect 1372 276 1380 284
rect 1596 1276 1604 1284
rect 1692 1236 1700 1244
rect 1676 1176 1684 1184
rect 1628 1156 1636 1164
rect 1628 916 1636 924
rect 1628 796 1636 804
rect 1596 716 1604 724
rect 1660 716 1668 724
rect 1692 836 1700 844
rect 1692 736 1700 744
rect 1884 1816 1892 1824
rect 2060 1816 2068 1824
rect 2108 1916 2116 1924
rect 2140 1896 2148 1904
rect 2124 1856 2132 1864
rect 1980 1756 1988 1764
rect 2092 1756 2100 1764
rect 1948 1736 1956 1744
rect 1788 1696 1796 1704
rect 1804 1696 1812 1704
rect 1820 1676 1828 1684
rect 1852 1716 1860 1724
rect 1884 1716 1892 1724
rect 1868 1696 1876 1704
rect 1772 1636 1780 1644
rect 1836 1636 1844 1644
rect 1740 1496 1748 1504
rect 1900 1696 1908 1704
rect 1932 1556 1940 1564
rect 1916 1496 1924 1504
rect 1852 1476 1860 1484
rect 1820 1456 1828 1464
rect 1756 1396 1764 1404
rect 1724 1296 1732 1304
rect 1868 1396 1876 1404
rect 1868 1356 1876 1364
rect 2044 1736 2052 1744
rect 2092 1736 2100 1744
rect 2140 1736 2148 1744
rect 2028 1676 2036 1684
rect 1964 1556 1972 1564
rect 1948 1536 1956 1544
rect 2012 1516 2020 1524
rect 1964 1496 1972 1504
rect 1948 1416 1956 1424
rect 2268 2136 2276 2144
rect 2316 2136 2324 2144
rect 2348 2236 2356 2244
rect 2348 2216 2356 2224
rect 2444 2536 2452 2544
rect 2684 2676 2692 2684
rect 2700 2656 2708 2664
rect 2638 2606 2646 2614
rect 2652 2606 2660 2614
rect 2666 2606 2674 2614
rect 2748 2576 2756 2584
rect 2684 2436 2692 2444
rect 2428 2336 2436 2344
rect 2716 2396 2724 2404
rect 2700 2296 2702 2304
rect 2702 2296 2708 2304
rect 2412 2256 2420 2264
rect 2428 2236 2436 2244
rect 2364 2196 2372 2204
rect 2396 2196 2404 2204
rect 2364 2176 2372 2184
rect 2380 2136 2388 2144
rect 2508 2176 2516 2184
rect 2172 1896 2180 1904
rect 2172 1796 2180 1804
rect 2268 2116 2276 2124
rect 2492 2116 2500 2124
rect 2380 2096 2388 2104
rect 2732 2236 2740 2244
rect 2638 2206 2646 2214
rect 2652 2206 2660 2214
rect 2666 2206 2674 2214
rect 3196 3736 3204 3744
rect 3244 3736 3252 3744
rect 3260 3716 3268 3724
rect 3292 3716 3300 3724
rect 3196 3696 3204 3704
rect 3100 3596 3108 3604
rect 3084 3456 3092 3464
rect 3084 3396 3092 3404
rect 3068 3316 3076 3324
rect 3084 3296 3092 3304
rect 3036 3096 3044 3104
rect 3068 3096 3076 3104
rect 3084 3016 3092 3024
rect 3068 2956 3076 2964
rect 2924 2716 2932 2724
rect 2860 2676 2868 2684
rect 2876 2636 2884 2644
rect 2844 2616 2852 2624
rect 3164 3676 3172 3684
rect 3148 3576 3156 3584
rect 3116 3556 3124 3564
rect 3164 3536 3172 3544
rect 3132 3496 3140 3504
rect 3276 3656 3284 3664
rect 3260 3616 3268 3624
rect 3228 3516 3236 3524
rect 3212 3496 3220 3504
rect 3244 3496 3252 3504
rect 3116 3476 3124 3484
rect 3132 3476 3140 3484
rect 3196 3476 3204 3484
rect 3212 3476 3220 3484
rect 3244 3476 3252 3484
rect 3196 3456 3204 3464
rect 3180 3416 3188 3424
rect 3228 3436 3236 3444
rect 3180 3376 3188 3384
rect 3164 3356 3172 3364
rect 3148 3316 3156 3324
rect 3196 3336 3204 3344
rect 3148 3156 3156 3164
rect 3116 3136 3124 3144
rect 3180 3136 3188 3144
rect 3260 3396 3268 3404
rect 3340 4156 3348 4164
rect 3324 4096 3332 4104
rect 3356 4096 3364 4104
rect 3372 4076 3380 4084
rect 3340 4056 3348 4064
rect 3340 3996 3348 4004
rect 3340 3936 3348 3944
rect 3372 3916 3380 3924
rect 3404 4056 3412 4064
rect 3404 3996 3412 4004
rect 3356 3856 3364 3864
rect 3468 4536 3476 4544
rect 3516 4556 3524 4564
rect 3484 4516 3492 4524
rect 3500 4416 3508 4424
rect 3452 4356 3460 4364
rect 3484 4356 3492 4364
rect 3452 4316 3460 4324
rect 3484 4276 3492 4284
rect 3772 4736 3780 4744
rect 3660 4716 3668 4724
rect 3724 4716 3732 4724
rect 3756 4716 3764 4724
rect 3612 4676 3620 4684
rect 3564 4556 3572 4564
rect 3548 4536 3556 4544
rect 3596 4616 3604 4624
rect 3564 4516 3572 4524
rect 3580 4516 3588 4524
rect 3548 4416 3556 4424
rect 3564 4316 3572 4324
rect 3660 4536 3668 4544
rect 3676 4496 3684 4504
rect 3628 4456 3636 4464
rect 3628 4396 3636 4404
rect 3708 4656 3716 4664
rect 3708 4596 3716 4604
rect 3900 4676 3908 4684
rect 3868 4616 3876 4624
rect 3932 4616 3940 4624
rect 3756 4556 3764 4564
rect 3788 4536 3796 4544
rect 3820 4536 3828 4544
rect 3724 4516 3732 4524
rect 3740 4516 3748 4524
rect 3772 4496 3780 4504
rect 3804 4496 3812 4504
rect 3692 4416 3700 4424
rect 3660 4376 3668 4384
rect 3660 4356 3668 4364
rect 3436 4256 3444 4264
rect 3468 4256 3476 4264
rect 3484 4236 3492 4244
rect 3452 4216 3460 4224
rect 3468 4216 3476 4224
rect 3436 4196 3444 4204
rect 3436 4076 3444 4084
rect 3500 4196 3508 4204
rect 3468 4156 3476 4164
rect 3484 4156 3492 4164
rect 3468 4016 3476 4024
rect 3436 3936 3444 3944
rect 3452 3936 3460 3944
rect 3436 3916 3444 3924
rect 3596 4276 3604 4284
rect 3548 4256 3556 4264
rect 3532 4196 3540 4204
rect 3532 4116 3540 4124
rect 3516 4096 3524 4104
rect 3516 4076 3524 4084
rect 3500 4016 3508 4024
rect 3500 3956 3508 3964
rect 3436 3856 3444 3864
rect 3372 3816 3380 3824
rect 3420 3816 3428 3824
rect 3324 3776 3332 3784
rect 3388 3776 3396 3784
rect 3420 3756 3428 3764
rect 3340 3616 3348 3624
rect 3372 3696 3380 3704
rect 3404 3676 3412 3684
rect 3468 3776 3476 3784
rect 3468 3716 3476 3724
rect 3564 4236 3572 4244
rect 3612 4256 3620 4264
rect 3580 4176 3588 4184
rect 3564 4116 3572 4124
rect 3644 4336 3652 4344
rect 3724 4436 3732 4444
rect 3708 4336 3716 4344
rect 3900 4596 3908 4604
rect 3932 4596 3940 4604
rect 3884 4516 3892 4524
rect 3820 4476 3828 4484
rect 3676 4316 3684 4324
rect 3740 4316 3748 4324
rect 3676 4296 3684 4304
rect 3660 4236 3668 4244
rect 3628 4176 3636 4184
rect 3612 4156 3620 4164
rect 3628 4136 3636 4144
rect 3612 4096 3620 4104
rect 3596 4076 3604 4084
rect 3644 4076 3652 4084
rect 3660 4076 3668 4084
rect 3548 3996 3556 4004
rect 3516 3816 3524 3824
rect 3532 3756 3540 3764
rect 3580 4016 3588 4024
rect 3612 4016 3620 4024
rect 3580 3956 3588 3964
rect 3612 3956 3620 3964
rect 3628 3916 3636 3924
rect 3596 3856 3604 3864
rect 3580 3796 3588 3804
rect 3628 3816 3636 3824
rect 3628 3796 3636 3804
rect 3612 3756 3620 3764
rect 3500 3696 3508 3704
rect 3612 3716 3620 3724
rect 3580 3696 3588 3704
rect 3484 3676 3492 3684
rect 3436 3656 3444 3664
rect 3484 3656 3492 3664
rect 3324 3596 3332 3604
rect 3356 3596 3364 3604
rect 3420 3596 3428 3604
rect 3292 3576 3300 3584
rect 3308 3576 3316 3584
rect 3436 3556 3444 3564
rect 3484 3556 3492 3564
rect 3564 3556 3572 3564
rect 3324 3536 3332 3544
rect 3388 3516 3396 3524
rect 3660 4036 3668 4044
rect 3660 3916 3668 3924
rect 3708 4236 3716 4244
rect 3708 4196 3716 4204
rect 3724 4116 3732 4124
rect 3692 4096 3700 4104
rect 3692 4076 3700 4084
rect 3724 4076 3732 4084
rect 3756 4276 3764 4284
rect 3836 4396 3844 4404
rect 3820 4356 3828 4364
rect 3804 4316 3812 4324
rect 3788 4256 3796 4264
rect 3788 4176 3796 4184
rect 3772 4156 3780 4164
rect 3756 4116 3764 4124
rect 3884 4476 3892 4484
rect 3900 4436 3908 4444
rect 3836 4316 3844 4324
rect 3868 4316 3876 4324
rect 3884 4316 3892 4324
rect 3980 4536 3988 4544
rect 3948 4436 3956 4444
rect 3996 4456 4004 4464
rect 4060 4836 4068 4844
rect 4158 4806 4166 4814
rect 4172 4806 4180 4814
rect 4186 4806 4194 4814
rect 4364 4916 4372 4924
rect 4092 4776 4100 4784
rect 4220 4776 4228 4784
rect 4268 4776 4276 4784
rect 4332 4776 4340 4784
rect 4204 4716 4212 4724
rect 4284 4716 4292 4724
rect 4204 4696 4212 4704
rect 4236 4696 4244 4704
rect 4300 4696 4308 4704
rect 4460 4696 4466 4704
rect 4466 4696 4468 4704
rect 4156 4676 4164 4684
rect 4236 4656 4244 4664
rect 4028 4556 4036 4564
rect 4108 4556 4116 4564
rect 4140 4536 4148 4544
rect 4012 4416 4020 4424
rect 4076 4416 4084 4424
rect 4060 4356 4068 4364
rect 3900 4296 3908 4304
rect 3916 4276 3924 4284
rect 3836 4216 3844 4224
rect 3852 4196 3860 4204
rect 3836 4176 3844 4184
rect 3900 4156 3908 4164
rect 3964 4276 3972 4284
rect 3948 4256 3956 4264
rect 3996 4176 4004 4184
rect 3948 4156 3956 4164
rect 4012 4156 4020 4164
rect 3868 4136 3876 4144
rect 3932 4136 3940 4144
rect 4158 4406 4166 4414
rect 4172 4406 4180 4414
rect 4186 4406 4194 4414
rect 4364 4676 4372 4684
rect 4348 4636 4356 4644
rect 4348 4596 4356 4604
rect 4364 4456 4372 4464
rect 4652 4676 4660 4684
rect 4540 4656 4548 4664
rect 4748 4656 4756 4664
rect 4540 4616 4548 4624
rect 4620 4616 4628 4624
rect 4860 4916 4868 4924
rect 4924 4916 4930 4924
rect 4930 4916 4932 4924
rect 4508 4556 4516 4564
rect 4780 4556 4788 4564
rect 4812 4556 4820 4564
rect 4428 4536 4436 4544
rect 4380 4416 4388 4424
rect 4460 4416 4468 4424
rect 4268 4396 4276 4404
rect 4380 4396 4388 4404
rect 4492 4316 4500 4324
rect 4732 4536 4740 4544
rect 5004 4816 5012 4824
rect 5036 4816 5044 4824
rect 4924 4676 4932 4684
rect 4844 4656 4852 4664
rect 4924 4656 4932 4664
rect 4956 4656 4964 4664
rect 4892 4616 4900 4624
rect 4972 4556 4980 4564
rect 4764 4496 4772 4504
rect 4508 4296 4516 4304
rect 4684 4296 4692 4304
rect 4428 4256 4436 4264
rect 4252 4216 4260 4224
rect 4300 4216 4308 4224
rect 4220 4156 4228 4164
rect 3820 4116 3828 4124
rect 4028 4116 4036 4124
rect 3804 4096 3812 4104
rect 3772 4076 3780 4084
rect 3788 4076 3796 4084
rect 3820 4056 3828 4064
rect 3868 4056 3876 4064
rect 3740 4036 3748 4044
rect 3756 3996 3764 4004
rect 3772 3996 3780 4004
rect 3740 3976 3748 3984
rect 4364 4196 4372 4204
rect 4412 4196 4420 4204
rect 4492 4196 4500 4204
rect 4332 4156 4340 4164
rect 4476 4116 4484 4124
rect 4092 4096 4100 4104
rect 3932 4076 3940 4084
rect 3964 4056 3972 4064
rect 3916 4036 3924 4044
rect 3900 4016 3908 4024
rect 3692 3936 3700 3944
rect 3740 3936 3748 3944
rect 3756 3916 3764 3924
rect 3676 3796 3684 3804
rect 3676 3756 3684 3764
rect 3660 3696 3668 3704
rect 3724 3876 3732 3884
rect 3868 3916 3876 3924
rect 3836 3876 3844 3884
rect 3772 3776 3780 3784
rect 3756 3716 3764 3724
rect 3708 3696 3716 3704
rect 3724 3696 3732 3704
rect 3692 3656 3700 3664
rect 3756 3656 3764 3664
rect 3724 3616 3732 3624
rect 3884 3896 3892 3904
rect 3788 3696 3796 3704
rect 3804 3696 3812 3704
rect 3852 3696 3860 3704
rect 3884 3696 3892 3704
rect 3804 3656 3812 3664
rect 3820 3656 3828 3664
rect 3772 3596 3780 3604
rect 3804 3596 3812 3604
rect 3740 3536 3748 3544
rect 3756 3536 3764 3544
rect 3820 3536 3828 3544
rect 3340 3496 3348 3504
rect 3436 3496 3444 3504
rect 3292 3456 3300 3464
rect 3372 3476 3380 3484
rect 3308 3436 3316 3444
rect 3404 3456 3412 3464
rect 3420 3456 3428 3464
rect 3292 3416 3300 3424
rect 3244 3336 3252 3344
rect 3228 3316 3236 3324
rect 3228 3296 3236 3304
rect 3212 3276 3220 3284
rect 3212 3156 3220 3164
rect 3116 3116 3124 3124
rect 3132 3116 3140 3124
rect 3164 3116 3172 3124
rect 3244 3276 3252 3284
rect 3324 3376 3332 3384
rect 3324 3336 3332 3344
rect 3388 3416 3396 3424
rect 3372 3396 3380 3404
rect 3404 3356 3412 3364
rect 3532 3496 3540 3504
rect 3452 3396 3460 3404
rect 3484 3456 3492 3464
rect 3580 3436 3588 3444
rect 3548 3376 3556 3384
rect 3516 3356 3524 3364
rect 3468 3336 3476 3344
rect 3484 3336 3492 3344
rect 3276 3316 3284 3324
rect 3356 3316 3364 3324
rect 3276 3116 3284 3124
rect 3132 2956 3140 2964
rect 3180 2956 3188 2964
rect 3148 2936 3156 2944
rect 3084 2816 3092 2824
rect 3004 2796 3012 2804
rect 3148 2796 3156 2804
rect 3100 2776 3108 2784
rect 2972 2736 2980 2744
rect 2972 2696 2980 2704
rect 3100 2696 3108 2704
rect 3068 2656 3076 2664
rect 3132 2616 3140 2624
rect 2956 2596 2964 2604
rect 2972 2596 2980 2604
rect 3020 2596 3028 2604
rect 2908 2556 2916 2564
rect 2940 2556 2948 2564
rect 3100 2516 3108 2524
rect 2908 2496 2916 2504
rect 2908 2456 2916 2464
rect 3116 2476 3124 2484
rect 2844 2416 2852 2424
rect 2956 2416 2964 2424
rect 2940 2316 2948 2324
rect 2876 2296 2884 2304
rect 2908 2296 2916 2304
rect 3164 2516 3172 2524
rect 3244 3056 3252 3064
rect 3244 2976 3252 2984
rect 3276 2976 3284 2984
rect 3228 2936 3236 2944
rect 3212 2916 3220 2924
rect 3276 2936 3284 2944
rect 3372 3296 3380 3304
rect 3596 3336 3604 3344
rect 3708 3496 3716 3504
rect 3660 3476 3668 3484
rect 3676 3476 3684 3484
rect 3644 3456 3652 3464
rect 3660 3436 3668 3444
rect 3644 3396 3652 3404
rect 3692 3436 3700 3444
rect 3756 3476 3764 3484
rect 3740 3396 3748 3404
rect 3724 3356 3732 3364
rect 3820 3496 3828 3504
rect 3772 3376 3780 3384
rect 3804 3336 3812 3344
rect 3452 3316 3460 3324
rect 3564 3316 3572 3324
rect 3628 3316 3636 3324
rect 3388 3216 3396 3224
rect 3308 3196 3316 3204
rect 3340 3156 3348 3164
rect 3308 3116 3316 3124
rect 3308 2976 3316 2984
rect 3308 2956 3316 2964
rect 3212 2896 3220 2904
rect 3244 2896 3252 2904
rect 3292 2896 3300 2904
rect 3228 2876 3236 2884
rect 3196 2756 3204 2764
rect 3180 2476 3188 2484
rect 3180 2416 3188 2424
rect 3004 2296 3012 2304
rect 3068 2296 3076 2304
rect 3132 2296 3140 2304
rect 3164 2296 3172 2304
rect 2860 2256 2868 2264
rect 2940 2256 2948 2264
rect 2588 2156 2596 2164
rect 2812 2156 2820 2164
rect 2940 2156 2948 2164
rect 2556 2116 2564 2124
rect 2572 2096 2580 2104
rect 2540 2076 2548 2084
rect 2780 2096 2788 2104
rect 2988 2156 2996 2164
rect 2956 2136 2964 2144
rect 2988 2116 2996 2124
rect 3020 2236 3028 2244
rect 3084 2236 3092 2244
rect 3020 2176 3028 2184
rect 3052 2156 3060 2164
rect 3036 2136 3044 2144
rect 3036 2096 3044 2104
rect 3068 2096 3076 2104
rect 3004 2056 3012 2064
rect 3036 2056 3044 2064
rect 2524 1996 2532 2004
rect 2556 1996 2564 2004
rect 2700 1996 2708 2004
rect 2780 1996 2788 2004
rect 2812 1996 2820 2004
rect 2268 1956 2276 1964
rect 2380 1916 2388 1924
rect 2252 1896 2260 1904
rect 3004 1896 3012 1904
rect 2204 1876 2212 1884
rect 2300 1876 2306 1884
rect 2306 1876 2308 1884
rect 2604 1876 2612 1884
rect 2892 1876 2900 1884
rect 2236 1856 2244 1864
rect 2492 1856 2500 1864
rect 2460 1836 2468 1844
rect 2588 1776 2596 1784
rect 3052 1856 3060 1864
rect 2638 1806 2646 1814
rect 2652 1806 2660 1814
rect 2666 1806 2674 1814
rect 2700 1776 2708 1784
rect 2652 1756 2660 1764
rect 2156 1636 2164 1644
rect 2060 1536 2068 1544
rect 2092 1536 2100 1544
rect 2172 1536 2180 1544
rect 2156 1516 2164 1524
rect 2092 1496 2100 1504
rect 2124 1496 2132 1504
rect 2028 1476 2036 1484
rect 2140 1476 2148 1484
rect 2188 1456 2196 1464
rect 2092 1396 2100 1404
rect 1964 1356 1972 1364
rect 1788 1336 1796 1344
rect 1948 1336 1956 1344
rect 1916 1316 1924 1324
rect 1772 1296 1780 1304
rect 1740 1256 1748 1264
rect 1740 1236 1748 1244
rect 1756 1196 1764 1204
rect 1740 1116 1748 1124
rect 1724 1076 1732 1084
rect 1772 1156 1780 1164
rect 1756 1096 1764 1104
rect 1788 1116 1796 1124
rect 1820 1156 1828 1164
rect 1804 1056 1812 1064
rect 1788 976 1796 984
rect 1756 956 1764 964
rect 1724 936 1732 944
rect 1740 876 1748 884
rect 1756 816 1764 824
rect 1724 756 1732 764
rect 1756 756 1764 764
rect 1724 716 1732 724
rect 1756 716 1764 724
rect 1628 696 1636 704
rect 1708 696 1716 704
rect 1740 696 1748 704
rect 1724 676 1732 684
rect 1612 656 1620 664
rect 1596 636 1604 644
rect 1708 656 1716 664
rect 1644 576 1652 584
rect 1516 516 1524 524
rect 1580 516 1588 524
rect 1564 496 1572 504
rect 1468 376 1476 384
rect 1420 316 1428 324
rect 1436 296 1444 304
rect 1420 276 1428 284
rect 1420 256 1428 264
rect 572 116 580 124
rect 780 116 788 124
rect 924 116 932 124
rect 1852 1276 1860 1284
rect 1996 1276 2004 1284
rect 1964 1256 1972 1264
rect 1900 1236 1908 1244
rect 2028 1236 2036 1244
rect 1996 1196 2004 1204
rect 1900 1116 1908 1124
rect 1932 1116 1940 1124
rect 1964 1116 1972 1124
rect 2076 1116 2084 1124
rect 1996 1096 2004 1104
rect 2028 1096 2036 1104
rect 1884 1076 1892 1084
rect 1932 1076 1940 1084
rect 2012 1076 2020 1084
rect 1836 876 1844 884
rect 1820 856 1828 864
rect 1868 1056 1876 1064
rect 1948 1056 1956 1064
rect 1964 936 1972 944
rect 2044 936 2052 944
rect 1932 916 1940 924
rect 1868 816 1876 824
rect 1852 716 1860 724
rect 1932 716 1940 724
rect 1836 696 1844 704
rect 1932 696 1940 704
rect 1804 656 1812 664
rect 1628 516 1636 524
rect 1644 516 1652 524
rect 1596 476 1604 484
rect 1564 316 1572 324
rect 1484 296 1492 304
rect 1500 296 1508 304
rect 1596 302 1604 304
rect 1596 296 1604 302
rect 1532 276 1540 284
rect 1452 196 1460 204
rect 1692 496 1700 504
rect 1676 476 1684 484
rect 1708 476 1716 484
rect 1724 476 1732 484
rect 1756 476 1764 484
rect 1756 416 1764 424
rect 1692 376 1700 384
rect 1724 376 1732 384
rect 1820 516 1828 524
rect 2028 676 2036 684
rect 2044 676 2052 684
rect 1916 656 1924 664
rect 2060 656 2068 664
rect 1932 556 1940 564
rect 2284 1496 2292 1504
rect 2204 1436 2212 1444
rect 2124 1216 2132 1224
rect 2556 1736 2564 1744
rect 2636 1736 2644 1744
rect 2332 1616 2340 1624
rect 2380 1616 2388 1624
rect 2844 1736 2852 1744
rect 2508 1716 2516 1724
rect 2748 1716 2756 1724
rect 2556 1696 2564 1704
rect 2460 1516 2468 1524
rect 2380 1496 2388 1504
rect 2476 1496 2484 1504
rect 2332 1456 2340 1464
rect 2428 1476 2436 1484
rect 2492 1476 2500 1484
rect 2412 1436 2420 1444
rect 2524 1436 2532 1444
rect 2396 1416 2404 1424
rect 2364 1396 2372 1404
rect 2300 1236 2308 1244
rect 2364 1236 2372 1244
rect 2220 1196 2228 1204
rect 2236 1196 2244 1204
rect 2188 1176 2196 1184
rect 2108 956 2116 964
rect 2220 1116 2228 1124
rect 2172 1096 2180 1104
rect 2188 1096 2196 1104
rect 2268 1096 2276 1104
rect 2364 1176 2372 1184
rect 2380 1176 2388 1184
rect 2428 1396 2436 1404
rect 2604 1496 2612 1504
rect 2732 1456 2740 1464
rect 2652 1436 2660 1444
rect 2638 1406 2646 1414
rect 2652 1406 2660 1414
rect 2666 1406 2674 1414
rect 2556 1376 2564 1384
rect 2684 1376 2692 1384
rect 2460 1356 2468 1364
rect 2524 1356 2532 1364
rect 2652 1336 2660 1344
rect 2556 1316 2564 1324
rect 2444 1276 2452 1284
rect 2412 1236 2420 1244
rect 2444 1236 2452 1244
rect 2412 1196 2420 1204
rect 2396 1136 2404 1144
rect 2396 1116 2404 1124
rect 2428 1176 2436 1184
rect 2604 1296 2612 1304
rect 2508 1236 2516 1244
rect 2492 1196 2500 1204
rect 2524 1196 2532 1204
rect 2492 1116 2500 1124
rect 2604 1156 2612 1164
rect 2572 1136 2580 1144
rect 2588 1136 2596 1144
rect 2380 1076 2388 1084
rect 2172 1056 2180 1064
rect 2204 1056 2212 1064
rect 2252 1056 2260 1064
rect 2172 956 2180 964
rect 2252 1016 2260 1024
rect 2236 996 2244 1004
rect 2316 1036 2324 1044
rect 2300 1016 2308 1024
rect 2332 1016 2340 1024
rect 2428 1036 2436 1044
rect 2396 996 2404 1004
rect 2316 956 2324 964
rect 2476 936 2484 944
rect 2492 936 2500 944
rect 2556 1056 2564 1064
rect 2380 836 2388 844
rect 2492 836 2500 844
rect 2316 736 2324 744
rect 2236 696 2244 704
rect 2300 696 2308 704
rect 2124 676 2132 684
rect 2268 656 2276 664
rect 2140 556 2148 564
rect 2156 556 2164 564
rect 2092 516 2100 524
rect 2060 496 2068 504
rect 2124 456 2132 464
rect 2716 1316 2724 1324
rect 2796 1416 2804 1424
rect 2956 1636 2964 1644
rect 2876 1456 2884 1464
rect 2748 1376 2756 1384
rect 2748 1356 2756 1364
rect 2796 1336 2804 1344
rect 2684 1136 2692 1144
rect 2668 1076 2676 1084
rect 2652 1036 2660 1044
rect 2638 1006 2646 1014
rect 2652 1006 2660 1014
rect 2666 1006 2674 1014
rect 2796 1276 2804 1284
rect 2892 1416 2900 1424
rect 2844 1396 2852 1404
rect 3068 1516 3076 1524
rect 3036 1476 3038 1484
rect 3038 1476 3044 1484
rect 3036 1456 3044 1464
rect 3020 1396 3028 1404
rect 3052 1416 3060 1424
rect 2892 1356 2900 1364
rect 2956 1356 2964 1364
rect 3052 1356 3060 1364
rect 2876 1316 2884 1324
rect 2956 1316 2964 1324
rect 2908 1296 2916 1304
rect 2940 1296 2948 1304
rect 2940 1276 2948 1284
rect 2828 1216 2836 1224
rect 2972 1296 2980 1304
rect 3004 1296 3012 1304
rect 3020 1256 3028 1264
rect 3100 2176 3108 2184
rect 3100 2116 3108 2124
rect 3100 1896 3108 1904
rect 3132 2256 3140 2264
rect 3212 2576 3220 2584
rect 3260 2836 3268 2844
rect 3356 3016 3364 3024
rect 3324 2936 3332 2944
rect 3356 2936 3364 2944
rect 3324 2896 3332 2904
rect 3372 2896 3380 2904
rect 3532 3276 3540 3284
rect 3788 3316 3796 3324
rect 3868 3476 3876 3484
rect 3852 3456 3860 3464
rect 3836 3396 3844 3404
rect 4060 4016 4068 4024
rect 3916 3996 3924 4004
rect 3948 3996 3956 4004
rect 3980 3836 3988 3844
rect 3996 3816 4004 3824
rect 3932 3696 3940 3704
rect 3948 3676 3956 3684
rect 3932 3656 3940 3664
rect 4076 3816 4084 3824
rect 4028 3776 4036 3784
rect 4028 3736 4036 3744
rect 4158 4006 4166 4014
rect 4172 4006 4180 4014
rect 4186 4006 4194 4014
rect 4172 3936 4180 3944
rect 4316 3996 4324 4004
rect 4636 4276 4644 4284
rect 4780 4396 4788 4404
rect 4860 4436 4868 4444
rect 4844 4396 4852 4404
rect 4828 4376 4836 4384
rect 4812 4256 4820 4264
rect 4700 4216 4708 4224
rect 4844 4216 4852 4224
rect 4636 4176 4644 4184
rect 4524 4156 4532 4164
rect 4668 4156 4676 4164
rect 4508 4116 4516 4124
rect 4540 4116 4548 4124
rect 4396 3896 4404 3904
rect 4492 3896 4500 3904
rect 4252 3816 4260 3824
rect 4284 3876 4292 3884
rect 4364 3876 4372 3884
rect 4412 3876 4420 3884
rect 4268 3796 4276 3804
rect 4332 3756 4340 3764
rect 4028 3716 4036 3724
rect 4124 3716 4132 3724
rect 4172 3656 4180 3664
rect 4220 3656 4228 3664
rect 4028 3636 4036 3644
rect 3980 3616 3988 3624
rect 4012 3576 4020 3584
rect 4158 3606 4166 3614
rect 4172 3606 4180 3614
rect 4186 3606 4194 3614
rect 4236 3576 4244 3584
rect 4156 3496 4164 3504
rect 4060 3476 4068 3484
rect 4140 3476 4148 3484
rect 4060 3456 4068 3464
rect 3980 3376 3988 3384
rect 3964 3336 3972 3344
rect 3996 3356 4004 3364
rect 4012 3336 4020 3344
rect 3900 3316 3908 3324
rect 4028 3316 4036 3324
rect 3612 3296 3620 3304
rect 3676 3296 3684 3304
rect 3756 3296 3764 3304
rect 3820 3296 3828 3304
rect 3756 3276 3764 3284
rect 3916 3296 3924 3304
rect 4220 3376 4228 3384
rect 4076 3356 4084 3364
rect 4124 3356 4132 3364
rect 4108 3336 4116 3344
rect 4220 3336 4228 3344
rect 4332 3636 4340 3644
rect 4332 3616 4340 3624
rect 4364 3616 4372 3624
rect 4476 3876 4484 3884
rect 4460 3716 4468 3724
rect 4524 3756 4532 3764
rect 4492 3676 4500 3684
rect 4284 3576 4292 3584
rect 4428 3576 4436 3584
rect 4748 4076 4756 4084
rect 4636 3816 4644 3824
rect 4684 3836 4692 3844
rect 4668 3756 4676 3764
rect 4572 3716 4580 3724
rect 4348 3516 4356 3524
rect 4252 3496 4260 3504
rect 4268 3456 4276 3464
rect 4268 3356 4276 3364
rect 4300 3476 4308 3484
rect 4828 4036 4836 4044
rect 4924 4176 4932 4184
rect 4860 4136 4868 4144
rect 4892 4136 4900 4144
rect 4876 4116 4884 4124
rect 4876 4036 4884 4044
rect 4876 3956 4884 3964
rect 4860 3936 4868 3944
rect 4860 3896 4868 3904
rect 4828 3876 4836 3884
rect 4844 3876 4852 3884
rect 4780 3856 4788 3864
rect 4844 3836 4852 3844
rect 4828 3696 4836 3704
rect 4812 3576 4820 3584
rect 4668 3496 4676 3504
rect 4780 3496 4788 3504
rect 4316 3456 4324 3464
rect 4572 3456 4580 3464
rect 4332 3436 4340 3444
rect 4380 3436 4388 3444
rect 4284 3336 4292 3344
rect 4092 3316 4100 3324
rect 4236 3316 4244 3324
rect 4300 3316 4308 3324
rect 4556 3376 4564 3384
rect 4348 3336 4356 3344
rect 4268 3296 4276 3304
rect 4364 3296 4372 3304
rect 4044 3276 4052 3284
rect 3468 3256 3476 3264
rect 3548 3256 3556 3264
rect 3660 3256 3668 3264
rect 3692 3256 3700 3264
rect 3452 3196 3460 3204
rect 3404 3136 3412 3144
rect 3436 3116 3444 3124
rect 3532 3176 3540 3184
rect 3692 3176 3700 3184
rect 3468 3156 3476 3164
rect 3484 3096 3492 3104
rect 3420 3056 3428 3064
rect 3452 3056 3460 3064
rect 3340 2756 3348 2764
rect 3260 2676 3262 2684
rect 3262 2676 3268 2684
rect 3356 2676 3364 2684
rect 3276 2576 3284 2584
rect 3292 2556 3300 2564
rect 3260 2536 3268 2544
rect 3260 2516 3268 2524
rect 3340 2536 3348 2544
rect 3292 2516 3300 2524
rect 3276 2476 3284 2484
rect 3436 3016 3444 3024
rect 3452 2956 3460 2964
rect 3452 2936 3460 2944
rect 3436 2876 3444 2884
rect 3404 2816 3412 2824
rect 3420 2816 3428 2824
rect 3436 2776 3444 2784
rect 3420 2756 3428 2764
rect 3404 2736 3412 2744
rect 3404 2716 3412 2724
rect 3580 3116 3588 3124
rect 3628 3116 3636 3124
rect 3612 3096 3620 3104
rect 3596 3076 3604 3084
rect 3580 3056 3588 3064
rect 3516 3036 3524 3044
rect 3548 3036 3556 3044
rect 3628 3016 3636 3024
rect 3692 3016 3700 3024
rect 3708 2976 3716 2984
rect 3564 2956 3572 2964
rect 3644 2956 3652 2964
rect 3596 2936 3604 2944
rect 3468 2896 3476 2904
rect 3516 2876 3524 2884
rect 3612 2856 3620 2864
rect 3468 2836 3476 2844
rect 3484 2836 3492 2844
rect 3468 2796 3476 2804
rect 3452 2756 3460 2764
rect 3500 2796 3508 2804
rect 3580 2776 3588 2784
rect 3628 2776 3636 2784
rect 3404 2696 3412 2704
rect 3420 2696 3428 2704
rect 3436 2656 3444 2664
rect 3484 2656 3492 2664
rect 3468 2556 3476 2564
rect 3388 2536 3396 2544
rect 3372 2476 3380 2484
rect 3420 2476 3428 2484
rect 3356 2456 3364 2464
rect 3228 2416 3236 2424
rect 3372 2396 3380 2404
rect 3308 2316 3316 2324
rect 3196 2276 3204 2284
rect 3212 2216 3220 2224
rect 3180 2196 3188 2204
rect 3308 2176 3316 2184
rect 3340 2156 3348 2164
rect 3276 2116 3284 2124
rect 3324 2116 3332 2124
rect 3132 2096 3140 2104
rect 3628 2736 3636 2744
rect 3612 2716 3620 2724
rect 3548 2656 3556 2664
rect 3948 3096 3956 3104
rect 3884 3056 3892 3064
rect 3852 2956 3860 2964
rect 3884 2936 3892 2944
rect 3756 2916 3764 2924
rect 4044 2916 4052 2924
rect 3756 2836 3764 2844
rect 3980 2816 3988 2824
rect 3788 2776 3796 2784
rect 3772 2716 3780 2724
rect 3708 2656 3716 2664
rect 3500 2616 3508 2624
rect 3516 2476 3524 2484
rect 3500 2276 3508 2284
rect 3484 2236 3492 2244
rect 3372 2156 3380 2164
rect 3420 2156 3428 2164
rect 3676 2616 3684 2624
rect 3644 2596 3652 2604
rect 3692 2576 3700 2584
rect 3724 2556 3732 2564
rect 3548 2476 3556 2484
rect 3676 2516 3684 2524
rect 3660 2436 3668 2444
rect 3612 2416 3620 2424
rect 3548 2396 3556 2404
rect 3548 2376 3556 2384
rect 3452 2136 3460 2144
rect 3372 2116 3380 2124
rect 3420 2116 3428 2124
rect 3468 2096 3476 2104
rect 3500 2096 3508 2104
rect 3356 2076 3364 2084
rect 3340 2056 3348 2064
rect 3228 1996 3236 2004
rect 3196 1896 3204 1904
rect 3244 1976 3252 1984
rect 3308 1916 3316 1924
rect 3228 1856 3236 1864
rect 3388 2036 3396 2044
rect 3404 1916 3412 1924
rect 3468 1916 3476 1924
rect 3404 1896 3412 1904
rect 3452 1896 3460 1904
rect 3388 1876 3390 1884
rect 3390 1876 3396 1884
rect 3356 1796 3364 1804
rect 3404 1796 3412 1804
rect 3148 1756 3156 1764
rect 3372 1756 3380 1764
rect 3132 1736 3140 1744
rect 3180 1736 3188 1744
rect 3164 1716 3172 1724
rect 3212 1716 3220 1724
rect 3132 1696 3140 1704
rect 3116 1536 3124 1544
rect 3116 1356 3124 1364
rect 3084 1296 3092 1304
rect 2956 1196 2964 1204
rect 2972 1196 2980 1204
rect 3068 1196 3076 1204
rect 2876 1076 2884 1084
rect 2844 1056 2852 1064
rect 2924 1016 2932 1024
rect 2956 1016 2964 1024
rect 2956 956 2964 964
rect 2588 796 2596 804
rect 2748 936 2756 944
rect 3228 1696 3236 1704
rect 3292 1636 3300 1644
rect 3196 1516 3204 1524
rect 3260 1456 3268 1464
rect 3292 1456 3300 1464
rect 3180 1196 3188 1204
rect 3228 1136 3236 1144
rect 3020 1096 3028 1104
rect 3084 1096 3092 1104
rect 3116 1076 3124 1084
rect 3164 1076 3172 1084
rect 3036 1036 3044 1044
rect 2716 796 2724 804
rect 2780 796 2788 804
rect 2684 776 2692 784
rect 2604 756 2612 764
rect 2636 756 2644 764
rect 2908 736 2916 744
rect 3020 896 3028 904
rect 3004 736 3012 744
rect 2892 696 2900 704
rect 2940 696 2948 704
rect 2988 696 2996 704
rect 2396 656 2404 664
rect 2492 656 2500 664
rect 2524 656 2532 664
rect 2348 616 2356 624
rect 2156 516 2164 524
rect 2188 496 2196 504
rect 1772 296 1780 304
rect 1868 296 1876 304
rect 1644 196 1652 204
rect 1468 156 1476 164
rect 1596 156 1604 164
rect 1564 136 1572 144
rect 1804 276 1812 284
rect 1852 276 1860 284
rect 1964 276 1972 284
rect 1980 276 1988 284
rect 1740 256 1748 264
rect 1820 256 1828 264
rect 1660 176 1668 184
rect 1788 196 1796 204
rect 1836 176 1844 184
rect 2524 616 2532 624
rect 2556 576 2564 584
rect 2572 556 2580 564
rect 2892 676 2900 684
rect 2956 676 2964 684
rect 2876 636 2884 644
rect 2638 606 2646 614
rect 2652 606 2660 614
rect 2666 606 2674 614
rect 2764 536 2772 544
rect 2604 516 2612 524
rect 2668 516 2676 524
rect 2524 396 2532 404
rect 2780 396 2788 404
rect 2332 376 2340 384
rect 2492 376 2500 384
rect 2460 296 2468 304
rect 2188 276 2196 284
rect 2172 176 2180 184
rect 1676 156 1684 164
rect 1740 156 1748 164
rect 1964 156 1972 164
rect 2076 156 2084 164
rect 2140 156 2148 164
rect 1868 136 1876 144
rect 2876 496 2884 504
rect 2796 376 2804 384
rect 2924 656 2932 664
rect 2988 616 2996 624
rect 2972 576 2980 584
rect 2956 556 2964 564
rect 2972 536 2980 544
rect 3020 556 3028 564
rect 3052 936 3060 944
rect 3052 816 3060 824
rect 3500 1876 3508 1884
rect 3452 1536 3460 1544
rect 3612 2336 3620 2344
rect 3628 2316 3636 2324
rect 3644 2296 3652 2304
rect 3564 2276 3572 2284
rect 3660 2276 3668 2284
rect 3788 2696 3796 2704
rect 4156 3236 4164 3244
rect 4158 3206 4166 3214
rect 4172 3206 4180 3214
rect 4186 3206 4194 3214
rect 4716 3476 4724 3484
rect 4764 3476 4772 3484
rect 4908 3976 4916 3984
rect 4956 4476 4964 4484
rect 4956 4376 4964 4384
rect 5260 4916 5268 4924
rect 5116 4856 5124 4864
rect 5228 4876 5236 4884
rect 5292 4936 5300 4944
rect 5388 4936 5396 4944
rect 5292 4896 5300 4904
rect 5388 4896 5396 4904
rect 5356 4856 5364 4864
rect 5276 4776 5284 4784
rect 5260 4716 5268 4724
rect 5308 4716 5316 4724
rect 5084 4656 5092 4664
rect 5132 4656 5140 4664
rect 5180 4656 5188 4664
rect 5180 4636 5188 4644
rect 5148 4596 5156 4604
rect 5100 4556 5108 4564
rect 4988 4436 4996 4444
rect 5148 4436 5156 4444
rect 5132 4376 5140 4384
rect 5068 4336 5076 4344
rect 5020 4296 5028 4304
rect 5036 4296 5044 4304
rect 4972 4136 4980 4144
rect 4956 4116 4964 4124
rect 5084 4296 5092 4304
rect 5068 4276 5076 4284
rect 5020 4236 5028 4244
rect 5052 4216 5060 4224
rect 5020 4136 5028 4144
rect 5036 4116 5044 4124
rect 5004 4096 5012 4104
rect 5036 4096 5044 4104
rect 4940 4036 4948 4044
rect 5068 4136 5076 4144
rect 5068 4016 5076 4024
rect 5052 3996 5060 4004
rect 5036 3956 5044 3964
rect 4988 3936 4996 3944
rect 4924 3916 4932 3924
rect 4908 3876 4916 3884
rect 4892 3816 4900 3824
rect 4892 3756 4900 3764
rect 4876 3576 4884 3584
rect 4764 3456 4772 3464
rect 4860 3456 4868 3464
rect 4716 3376 4724 3384
rect 4700 3356 4708 3364
rect 4396 3176 4404 3184
rect 4524 3156 4532 3164
rect 4828 3436 4836 3444
rect 4780 3376 4788 3384
rect 4764 3356 4772 3364
rect 4748 3336 4756 3344
rect 4780 3276 4788 3284
rect 4652 3116 4660 3124
rect 4748 3116 4756 3124
rect 4940 3856 4948 3864
rect 4924 3776 4932 3784
rect 4940 3776 4948 3784
rect 4908 3716 4916 3724
rect 4908 3476 4916 3484
rect 4956 3476 4964 3484
rect 4908 3456 4916 3464
rect 4940 3456 4948 3464
rect 4972 3416 4980 3424
rect 4812 3316 4820 3324
rect 4828 3276 4836 3284
rect 4796 3176 4804 3184
rect 4828 3156 4836 3164
rect 4796 3116 4804 3124
rect 4108 3096 4116 3104
rect 4684 3096 4692 3104
rect 4780 3096 4788 3104
rect 4076 3076 4084 3084
rect 4204 3076 4212 3084
rect 4140 3036 4148 3044
rect 4444 3076 4452 3084
rect 4700 3076 4708 3084
rect 4716 3076 4724 3084
rect 4860 3176 4868 3184
rect 4844 3116 4852 3124
rect 4396 3036 4404 3044
rect 4412 3016 4420 3024
rect 4268 2996 4276 3004
rect 4316 2996 4324 3004
rect 4236 2956 4244 2964
rect 4524 2976 4532 2984
rect 4636 2976 4644 2984
rect 4364 2956 4372 2964
rect 4476 2956 4484 2964
rect 4652 2956 4660 2964
rect 4732 2956 4740 2964
rect 4332 2936 4340 2944
rect 4540 2936 4548 2944
rect 4652 2936 4660 2944
rect 4684 2936 4692 2944
rect 4060 2876 4068 2884
rect 4158 2806 4166 2814
rect 4172 2806 4180 2814
rect 4186 2806 4194 2814
rect 4028 2776 4036 2784
rect 4092 2776 4100 2784
rect 4060 2736 4068 2744
rect 4556 2776 4564 2784
rect 3868 2696 3876 2704
rect 4508 2696 4516 2704
rect 3836 2676 3844 2684
rect 3804 2556 3812 2564
rect 3804 2536 3812 2544
rect 3948 2636 3956 2644
rect 3868 2556 3876 2564
rect 4396 2676 4404 2684
rect 4108 2656 4116 2664
rect 4252 2656 4260 2664
rect 4028 2596 4036 2604
rect 3980 2536 3988 2544
rect 4012 2556 4020 2564
rect 3852 2516 3860 2524
rect 3836 2496 3844 2504
rect 3884 2496 3892 2504
rect 3916 2496 3924 2504
rect 3772 2456 3780 2464
rect 3788 2456 3796 2464
rect 3852 2456 3860 2464
rect 3900 2456 3908 2464
rect 3884 2436 3892 2444
rect 3836 2416 3844 2424
rect 3788 2376 3796 2384
rect 3852 2376 3860 2384
rect 3756 2356 3764 2364
rect 3756 2336 3764 2344
rect 3724 2296 3732 2304
rect 3708 2276 3716 2284
rect 3676 2216 3684 2224
rect 3804 2356 3812 2364
rect 3820 2336 3828 2344
rect 3852 2296 3860 2304
rect 3836 2276 3844 2284
rect 3804 2236 3812 2244
rect 3756 2196 3764 2204
rect 3772 2196 3780 2204
rect 3596 2136 3604 2144
rect 3580 1976 3588 1984
rect 3564 1856 3572 1864
rect 3548 1816 3556 1824
rect 3532 1776 3540 1784
rect 3564 1696 3572 1704
rect 3452 1516 3460 1524
rect 3516 1516 3524 1524
rect 3404 1456 3412 1464
rect 3708 1956 3716 1964
rect 3756 2136 3764 2144
rect 3804 1976 3812 1984
rect 3724 1936 3732 1944
rect 3756 1916 3764 1924
rect 3820 1916 3828 1924
rect 3836 1896 3844 1904
rect 3612 1876 3620 1884
rect 3692 1876 3700 1884
rect 3724 1876 3732 1884
rect 3692 1836 3700 1844
rect 3836 1836 3844 1844
rect 3676 1816 3684 1824
rect 3660 1796 3668 1804
rect 3772 1796 3780 1804
rect 3932 2416 3940 2424
rect 4060 2616 4068 2624
rect 4108 2576 4116 2584
rect 4108 2556 4116 2564
rect 4044 2536 4052 2544
rect 4428 2596 4436 2604
rect 4508 2596 4516 2604
rect 4396 2556 4404 2564
rect 4140 2536 4148 2544
rect 4364 2536 4372 2544
rect 4140 2516 4148 2524
rect 4156 2496 4164 2504
rect 4236 2456 4244 2464
rect 4012 2376 4020 2384
rect 4158 2406 4166 2414
rect 4172 2406 4180 2414
rect 4186 2406 4194 2414
rect 4236 2336 4244 2344
rect 3932 2316 3940 2324
rect 4028 2316 4036 2324
rect 4108 2316 4116 2324
rect 3900 2296 3908 2304
rect 3900 2176 3908 2184
rect 3916 2136 3924 2144
rect 3900 1936 3908 1944
rect 4284 2496 4292 2504
rect 4556 2576 4564 2584
rect 4572 2516 4580 2524
rect 4700 2896 4708 2904
rect 4812 3076 4820 3084
rect 4796 3056 4804 3064
rect 4780 3016 4788 3024
rect 4812 2996 4820 3004
rect 4860 3056 4868 3064
rect 4876 3056 4884 3064
rect 4844 2996 4852 3004
rect 4876 2956 4884 2964
rect 4796 2936 4804 2944
rect 4828 2936 4836 2944
rect 4860 2936 4868 2944
rect 4764 2916 4772 2924
rect 4748 2896 4756 2904
rect 4716 2876 4724 2884
rect 4828 2916 4836 2924
rect 4860 2916 4868 2924
rect 4812 2796 4820 2804
rect 4684 2696 4692 2704
rect 4972 3316 4980 3324
rect 4940 3176 4948 3184
rect 4972 3256 4980 3264
rect 4956 3156 4964 3164
rect 4908 3136 4916 3144
rect 5068 3916 5076 3924
rect 5100 4076 5108 4084
rect 5100 3976 5108 3984
rect 5726 5006 5734 5014
rect 5740 5006 5748 5014
rect 5754 5006 5762 5014
rect 5516 4996 5524 5004
rect 6316 4976 6324 4984
rect 6716 4976 6724 4984
rect 5676 4956 5684 4964
rect 5788 4956 5796 4964
rect 6060 4956 6068 4964
rect 6684 4956 6692 4964
rect 5452 4936 5460 4944
rect 5420 4916 5428 4924
rect 5708 4916 5716 4924
rect 5596 4876 5604 4884
rect 5516 4836 5524 4844
rect 5852 4936 5860 4944
rect 6252 4936 6260 4944
rect 5836 4716 5844 4724
rect 5868 4916 5876 4924
rect 6028 4916 6036 4924
rect 5500 4696 5508 4704
rect 5788 4696 5796 4704
rect 5420 4676 5428 4684
rect 5596 4656 5604 4664
rect 5500 4636 5508 4644
rect 5532 4636 5540 4644
rect 5420 4596 5428 4604
rect 5308 4556 5316 4564
rect 5532 4616 5540 4624
rect 5516 4596 5524 4604
rect 5260 4536 5268 4544
rect 5468 4536 5476 4544
rect 5180 4376 5188 4384
rect 5212 4376 5220 4384
rect 5420 4496 5428 4504
rect 5500 4496 5508 4504
rect 5324 4316 5332 4324
rect 5292 4296 5300 4304
rect 5228 4276 5236 4284
rect 5196 4256 5204 4264
rect 5260 4256 5268 4264
rect 5180 4236 5188 4244
rect 5196 4236 5204 4244
rect 5260 4236 5268 4244
rect 5340 4276 5348 4284
rect 5292 4236 5300 4244
rect 5356 4236 5364 4244
rect 5276 4216 5284 4224
rect 5292 4136 5300 4144
rect 5404 4196 5412 4204
rect 5404 4156 5412 4164
rect 5388 4116 5396 4124
rect 5180 4076 5188 4084
rect 5148 3936 5156 3944
rect 5292 4036 5300 4044
rect 5308 4036 5316 4044
rect 5212 4016 5220 4024
rect 5228 3956 5236 3964
rect 5084 3896 5092 3904
rect 5036 3876 5044 3884
rect 5052 3876 5060 3884
rect 5100 3876 5108 3884
rect 5148 3896 5156 3904
rect 5212 3896 5220 3904
rect 5356 3956 5364 3964
rect 5276 3896 5284 3904
rect 5164 3876 5172 3884
rect 5228 3876 5236 3884
rect 5164 3856 5172 3864
rect 5212 3856 5220 3864
rect 5036 3816 5044 3824
rect 5116 3816 5124 3824
rect 5004 3756 5012 3764
rect 5004 3716 5012 3724
rect 5180 3816 5188 3824
rect 5116 3736 5124 3744
rect 5228 3796 5236 3804
rect 5340 3876 5348 3884
rect 5308 3836 5316 3844
rect 5260 3776 5268 3784
rect 5308 3776 5316 3784
rect 5260 3756 5268 3764
rect 5036 3696 5044 3704
rect 5116 3716 5124 3724
rect 5164 3716 5172 3724
rect 5036 3476 5044 3484
rect 5020 3316 5028 3324
rect 5036 3296 5044 3304
rect 5068 3316 5076 3324
rect 5052 3276 5060 3284
rect 5004 3216 5012 3224
rect 4988 3176 4996 3184
rect 5052 3196 5060 3204
rect 5100 3676 5108 3684
rect 5196 3616 5204 3624
rect 5196 3556 5204 3564
rect 5100 3496 5108 3504
rect 5404 3816 5412 3824
rect 5372 3796 5380 3804
rect 5404 3756 5412 3764
rect 5340 3736 5348 3744
rect 5372 3736 5380 3744
rect 5292 3696 5300 3704
rect 5324 3696 5332 3704
rect 5100 3456 5108 3464
rect 5116 3456 5124 3464
rect 5212 3456 5220 3464
rect 5228 3456 5236 3464
rect 5116 3436 5124 3444
rect 5228 3436 5236 3444
rect 5164 3336 5172 3344
rect 5148 3316 5156 3324
rect 5116 3296 5124 3304
rect 5260 3496 5268 3504
rect 5308 3636 5316 3644
rect 5356 3656 5364 3664
rect 5324 3556 5332 3564
rect 5308 3536 5316 3544
rect 5276 3476 5284 3484
rect 5308 3456 5316 3464
rect 5212 3336 5220 3344
rect 5228 3336 5236 3344
rect 5180 3256 5188 3264
rect 5148 3216 5156 3224
rect 5036 3136 5044 3144
rect 5052 3136 5060 3144
rect 5084 3136 5092 3144
rect 5180 3136 5188 3144
rect 4940 3116 4948 3124
rect 5004 3116 5012 3124
rect 4956 3076 4964 3084
rect 5020 3076 5028 3084
rect 4972 3056 4980 3064
rect 4956 2956 4964 2964
rect 4972 2936 4980 2944
rect 5196 3116 5204 3124
rect 4988 2916 4996 2924
rect 4636 2676 4644 2684
rect 4892 2676 4900 2684
rect 5020 2836 5028 2844
rect 5068 2956 5076 2964
rect 5132 3096 5140 3104
rect 5164 3096 5172 3104
rect 5116 2976 5124 2984
rect 5228 3316 5236 3324
rect 5308 3316 5316 3324
rect 5260 3296 5268 3304
rect 5340 3476 5348 3484
rect 5356 3316 5364 3324
rect 5324 3296 5332 3304
rect 5276 3216 5284 3224
rect 5308 3196 5316 3204
rect 5276 3136 5284 3144
rect 5324 3136 5332 3144
rect 5500 4456 5508 4464
rect 5468 4436 5476 4444
rect 5436 4376 5444 4384
rect 5516 4376 5524 4384
rect 5468 4316 5476 4324
rect 5500 4296 5508 4304
rect 5516 4216 5524 4224
rect 5516 4116 5524 4124
rect 5484 4096 5492 4104
rect 5500 4096 5508 4104
rect 5452 3956 5460 3964
rect 5468 3936 5476 3944
rect 5452 3916 5460 3924
rect 5436 3776 5444 3784
rect 5452 3696 5460 3704
rect 5468 3676 5476 3684
rect 5436 3616 5444 3624
rect 5420 3596 5428 3604
rect 5420 3536 5428 3544
rect 5388 3516 5396 3524
rect 5388 3456 5396 3464
rect 5404 3436 5412 3444
rect 5388 3416 5396 3424
rect 5388 3396 5396 3404
rect 5372 3276 5380 3284
rect 5404 3336 5412 3344
rect 5484 3596 5492 3604
rect 5468 3576 5476 3584
rect 5692 4676 5700 4684
rect 5676 4656 5684 4664
rect 5772 4676 5780 4684
rect 5756 4656 5764 4664
rect 5772 4656 5780 4664
rect 5726 4606 5734 4614
rect 5740 4606 5748 4614
rect 5754 4606 5762 4614
rect 5692 4596 5700 4604
rect 5852 4676 5860 4684
rect 5900 4656 5908 4664
rect 5932 4616 5940 4624
rect 6348 4836 6356 4844
rect 6012 4716 6020 4724
rect 6092 4716 6100 4724
rect 6172 4716 6180 4724
rect 5996 4696 6004 4704
rect 6060 4696 6068 4704
rect 6124 4696 6132 4704
rect 5964 4676 5972 4684
rect 6012 4676 6020 4684
rect 6092 4676 6100 4684
rect 5916 4536 5924 4544
rect 5948 4536 5956 4544
rect 6060 4576 6068 4584
rect 6108 4656 6116 4664
rect 6108 4616 6116 4624
rect 6124 4556 6132 4564
rect 6060 4536 6068 4544
rect 6092 4536 6100 4544
rect 5628 4516 5636 4524
rect 5708 4516 5716 4524
rect 5820 4516 5828 4524
rect 5548 4496 5556 4504
rect 5548 4316 5556 4324
rect 5964 4496 5972 4504
rect 5996 4496 6004 4504
rect 5932 4476 5940 4484
rect 5836 4316 5844 4324
rect 5964 4316 5972 4324
rect 5836 4296 5844 4304
rect 5740 4276 5748 4284
rect 5612 4256 5620 4264
rect 5708 4256 5716 4264
rect 5628 4236 5636 4244
rect 5548 4196 5556 4204
rect 5548 4176 5556 4184
rect 5548 4116 5556 4124
rect 5564 4096 5572 4104
rect 5692 4216 5700 4224
rect 5726 4206 5734 4214
rect 5740 4206 5748 4214
rect 5754 4206 5762 4214
rect 5644 4136 5652 4144
rect 5660 4136 5668 4144
rect 5596 4116 5604 4124
rect 5596 4096 5604 4104
rect 5644 3956 5652 3964
rect 5548 3916 5556 3924
rect 5628 3916 5636 3924
rect 5564 3856 5572 3864
rect 5644 3816 5652 3824
rect 5564 3716 5572 3724
rect 5628 3676 5636 3684
rect 5532 3616 5540 3624
rect 5500 3556 5508 3564
rect 5612 3556 5620 3564
rect 5452 3516 5460 3524
rect 5484 3516 5492 3524
rect 5516 3516 5524 3524
rect 5580 3516 5588 3524
rect 5484 3496 5492 3504
rect 5516 3496 5524 3504
rect 5564 3496 5572 3504
rect 5532 3476 5540 3484
rect 5436 3436 5444 3444
rect 5564 3416 5572 3424
rect 5564 3356 5572 3364
rect 5452 3336 5460 3344
rect 5532 3336 5540 3344
rect 5484 3316 5492 3324
rect 5388 3236 5396 3244
rect 5436 3296 5444 3304
rect 5452 3296 5460 3304
rect 5516 3296 5524 3304
rect 5420 3136 5428 3144
rect 5340 3116 5348 3124
rect 5420 3116 5428 3124
rect 5468 3256 5476 3264
rect 5388 3076 5396 3084
rect 5420 3076 5428 3084
rect 5292 3056 5300 3064
rect 5228 2976 5236 2984
rect 5212 2956 5220 2964
rect 5164 2936 5172 2944
rect 5196 2936 5204 2944
rect 5180 2916 5188 2924
rect 5388 3016 5396 3024
rect 5260 2956 5268 2964
rect 5308 2936 5316 2944
rect 5340 2936 5348 2944
rect 5116 2876 5124 2884
rect 5100 2816 5108 2824
rect 5196 2736 5204 2744
rect 5436 3056 5444 3064
rect 5324 2916 5332 2924
rect 5452 2916 5460 2924
rect 5324 2816 5332 2824
rect 5292 2796 5300 2804
rect 5276 2716 5284 2724
rect 5340 2776 5348 2784
rect 5420 2796 5428 2804
rect 5500 3276 5508 3284
rect 5676 4116 5684 4124
rect 5756 4096 5764 4104
rect 5676 4076 5684 4084
rect 5708 4076 5716 4084
rect 6028 4476 6036 4484
rect 6348 4716 6356 4724
rect 6220 4696 6228 4704
rect 6268 4696 6276 4704
rect 6348 4696 6356 4704
rect 6204 4656 6212 4664
rect 6316 4656 6324 4664
rect 6172 4616 6180 4624
rect 6220 4616 6228 4624
rect 6316 4616 6324 4624
rect 6156 4556 6164 4564
rect 6252 4556 6260 4564
rect 6364 4656 6372 4664
rect 6348 4636 6356 4644
rect 6332 4536 6340 4544
rect 6220 4516 6228 4524
rect 6172 4496 6180 4504
rect 6204 4496 6212 4504
rect 6268 4476 6276 4484
rect 6300 4476 6308 4484
rect 6316 4476 6324 4484
rect 6124 4456 6132 4464
rect 6284 4456 6292 4464
rect 6092 4316 6100 4324
rect 6300 4296 6308 4304
rect 5996 4276 6004 4284
rect 5948 4256 5956 4264
rect 6172 4256 6180 4264
rect 6012 4236 6020 4244
rect 6076 4236 6084 4244
rect 5980 4176 5988 4184
rect 5868 4156 5876 4164
rect 6060 4076 6068 4084
rect 6124 4156 6132 4164
rect 6220 4136 6228 4144
rect 6236 4136 6244 4144
rect 6220 4116 6228 4124
rect 6076 3996 6084 4004
rect 6268 4096 6276 4104
rect 6124 3956 6132 3964
rect 6204 3956 6212 3964
rect 6220 3956 6228 3964
rect 5692 3936 5700 3944
rect 6044 3936 6052 3944
rect 6092 3936 6100 3944
rect 5788 3876 5796 3884
rect 5708 3836 5716 3844
rect 5726 3806 5734 3814
rect 5740 3806 5748 3814
rect 5754 3806 5762 3814
rect 5916 3902 5924 3904
rect 5916 3896 5924 3902
rect 5836 3836 5844 3844
rect 5884 3856 5892 3864
rect 5852 3816 5860 3824
rect 5708 3776 5716 3784
rect 5772 3776 5780 3784
rect 5804 3776 5812 3784
rect 5692 3756 5700 3764
rect 5724 3756 5732 3764
rect 5820 3756 5828 3764
rect 5900 3756 5908 3764
rect 5692 3716 5700 3724
rect 5660 3536 5668 3544
rect 5628 3516 5636 3524
rect 5628 3476 5636 3484
rect 5596 3436 5604 3444
rect 5660 3436 5668 3444
rect 5580 3296 5588 3304
rect 5564 3236 5572 3244
rect 5532 3176 5540 3184
rect 5548 3176 5556 3184
rect 5564 3156 5572 3164
rect 5628 3276 5636 3284
rect 5612 3136 5620 3144
rect 5788 3716 5796 3724
rect 5820 3716 5828 3724
rect 5916 3716 5924 3724
rect 5708 3676 5716 3684
rect 5724 3676 5732 3684
rect 5788 3556 5796 3564
rect 5804 3536 5812 3544
rect 5724 3516 5732 3524
rect 5788 3516 5796 3524
rect 5884 3676 5892 3684
rect 5932 3676 5940 3684
rect 5900 3596 5908 3604
rect 5852 3516 5860 3524
rect 5820 3476 5828 3484
rect 5740 3456 5748 3464
rect 5726 3406 5734 3414
rect 5740 3406 5748 3414
rect 5754 3406 5762 3414
rect 5836 3456 5844 3464
rect 5884 3436 5892 3444
rect 6044 3816 6052 3824
rect 5996 3756 6004 3764
rect 5980 3716 5988 3724
rect 6028 3716 6036 3724
rect 5980 3656 5988 3664
rect 5996 3496 6004 3504
rect 5980 3416 5988 3424
rect 5900 3356 5908 3364
rect 5724 3318 5732 3324
rect 5724 3316 5732 3318
rect 5868 3316 5876 3324
rect 5820 3236 5828 3244
rect 5676 3156 5684 3164
rect 5500 3116 5508 3124
rect 5580 3116 5588 3124
rect 5820 3116 5828 3124
rect 5564 3096 5572 3104
rect 5516 3056 5524 3064
rect 5484 2776 5492 2784
rect 5468 2736 5476 2744
rect 5388 2716 5396 2724
rect 5148 2696 5156 2704
rect 5244 2696 5252 2704
rect 5388 2696 5396 2704
rect 5452 2702 5460 2704
rect 5452 2696 5460 2702
rect 5068 2676 5076 2684
rect 5292 2676 5300 2684
rect 5340 2676 5348 2684
rect 4780 2656 4788 2664
rect 4892 2656 4900 2664
rect 5004 2656 5012 2664
rect 5196 2656 5204 2664
rect 4812 2596 4820 2604
rect 4620 2576 4628 2584
rect 4700 2576 4708 2584
rect 5212 2616 5220 2624
rect 5420 2656 5428 2664
rect 5276 2596 5284 2604
rect 5340 2596 5348 2604
rect 5548 3076 5556 3084
rect 5628 3076 5636 3084
rect 5692 3076 5700 3084
rect 5532 2956 5540 2964
rect 5708 3036 5716 3044
rect 5692 3016 5700 3024
rect 5726 3006 5734 3014
rect 5740 3006 5748 3014
rect 5754 3006 5762 3014
rect 5596 2976 5604 2984
rect 5692 2936 5700 2944
rect 5788 2936 5796 2944
rect 5804 2936 5812 2944
rect 5884 3036 5892 3044
rect 5836 2996 5844 3004
rect 5932 3356 5940 3364
rect 5996 3396 6004 3404
rect 5964 3276 5972 3284
rect 5948 3256 5956 3264
rect 5948 3136 5956 3144
rect 6108 3896 6116 3904
rect 6188 3916 6196 3924
rect 6140 3876 6148 3884
rect 6188 3876 6196 3884
rect 6092 3856 6100 3864
rect 6108 3856 6116 3864
rect 6156 3836 6164 3844
rect 6076 3736 6084 3744
rect 6092 3696 6100 3704
rect 6236 3896 6244 3904
rect 6284 3996 6292 4004
rect 6268 3856 6276 3864
rect 6188 3736 6196 3744
rect 6188 3696 6196 3704
rect 6124 3656 6132 3664
rect 6140 3496 6148 3504
rect 6108 3476 6116 3484
rect 6092 3456 6100 3464
rect 6172 3456 6180 3464
rect 6124 3436 6132 3444
rect 6076 3396 6084 3404
rect 6092 3376 6100 3384
rect 6140 3336 6148 3344
rect 5996 3276 6004 3284
rect 5980 3136 5988 3144
rect 6012 3136 6020 3144
rect 5980 3096 5988 3104
rect 6012 3096 6020 3104
rect 6092 3296 6100 3304
rect 6076 3256 6084 3264
rect 6092 3196 6100 3204
rect 6108 3096 6116 3104
rect 5980 3076 5988 3084
rect 5996 3076 6004 3084
rect 6028 3076 6036 3084
rect 6060 3076 6068 3084
rect 6124 3076 6132 3084
rect 5980 3036 5988 3044
rect 5964 3016 5972 3024
rect 5932 2936 5940 2944
rect 5628 2876 5636 2884
rect 5564 2836 5572 2844
rect 5500 2636 5508 2644
rect 5500 2616 5508 2624
rect 4716 2556 4724 2564
rect 5052 2556 5060 2564
rect 5100 2556 5108 2564
rect 5436 2556 5444 2564
rect 4812 2536 4820 2544
rect 4844 2536 4852 2544
rect 5068 2536 5076 2544
rect 5244 2536 5252 2544
rect 4604 2496 4612 2504
rect 4780 2496 4788 2504
rect 4588 2436 4596 2444
rect 4284 2376 4292 2384
rect 4268 2316 4276 2324
rect 4572 2316 4580 2324
rect 3996 2276 4004 2284
rect 4028 2256 4036 2264
rect 3948 2216 3956 2224
rect 3932 1916 3940 1924
rect 4012 2196 4020 2204
rect 3964 2136 3972 2144
rect 3964 2116 3972 2124
rect 3964 2056 3972 2064
rect 3980 1936 3988 1944
rect 3964 1856 3972 1864
rect 3868 1736 3876 1744
rect 3948 1736 3956 1744
rect 4316 2276 4324 2284
rect 4236 2256 4244 2264
rect 4252 2256 4260 2264
rect 4364 2256 4372 2264
rect 4236 2156 4244 2164
rect 4204 2136 4212 2144
rect 4012 2076 4020 2084
rect 4028 2036 4036 2044
rect 4044 1936 4052 1944
rect 4012 1916 4020 1924
rect 4028 1896 4036 1904
rect 4158 2006 4166 2014
rect 4172 2006 4180 2014
rect 4186 2006 4194 2014
rect 4172 1976 4180 1984
rect 4284 1976 4292 1984
rect 4508 2156 4516 2164
rect 4428 2116 4436 2124
rect 4508 2116 4514 2124
rect 4514 2116 4516 2124
rect 4396 2076 4404 2084
rect 4396 2016 4404 2024
rect 4460 1976 4468 1984
rect 4364 1916 4372 1924
rect 4556 1916 4564 1924
rect 4172 1896 4180 1904
rect 4076 1876 4084 1884
rect 4124 1836 4132 1844
rect 4076 1816 4084 1824
rect 4092 1796 4100 1804
rect 4204 1876 4212 1884
rect 4332 1856 4340 1864
rect 4444 1856 4452 1864
rect 4124 1776 4132 1784
rect 4476 1816 4484 1824
rect 4524 1816 4532 1824
rect 4364 1776 4372 1784
rect 4060 1756 4068 1764
rect 4012 1676 4020 1684
rect 4220 1676 4228 1684
rect 4044 1656 4052 1664
rect 4158 1606 4166 1614
rect 4172 1606 4180 1614
rect 4186 1606 4194 1614
rect 3804 1496 3812 1504
rect 3868 1496 3876 1504
rect 3996 1576 4004 1584
rect 4076 1496 4084 1504
rect 4156 1456 4164 1464
rect 3676 1416 3684 1424
rect 3996 1416 4004 1424
rect 4108 1416 4116 1424
rect 3948 1376 3956 1384
rect 4140 1396 4148 1404
rect 3916 1336 3924 1344
rect 3276 1276 3284 1284
rect 3356 1256 3364 1264
rect 3292 1136 3300 1144
rect 3260 1116 3268 1124
rect 3276 1076 3284 1084
rect 3244 1056 3252 1064
rect 3116 956 3124 964
rect 3084 896 3092 904
rect 3164 1016 3172 1024
rect 3276 936 3284 944
rect 3148 736 3156 744
rect 3340 736 3348 744
rect 3068 676 3076 684
rect 3052 636 3060 644
rect 3148 656 3156 664
rect 3068 576 3076 584
rect 3036 536 3044 544
rect 3100 556 3108 564
rect 2956 496 2964 504
rect 3020 496 3028 504
rect 2908 376 2916 384
rect 3020 336 3028 344
rect 3084 316 3092 324
rect 3116 316 3124 324
rect 2764 296 2772 304
rect 2892 296 2900 304
rect 3020 296 3028 304
rect 3052 296 3060 304
rect 3084 296 3092 304
rect 2572 256 2580 264
rect 2604 236 2612 244
rect 2652 236 2660 244
rect 2638 206 2646 214
rect 2652 206 2660 214
rect 2666 206 2674 214
rect 2732 276 2740 284
rect 2764 276 2772 284
rect 2844 276 2852 284
rect 3036 276 3044 284
rect 3132 276 3140 284
rect 2668 176 2676 184
rect 2716 176 2724 184
rect 2924 256 2932 264
rect 3084 256 3092 264
rect 2444 156 2452 164
rect 2508 156 2516 164
rect 2764 156 2772 164
rect 2828 156 2836 164
rect 2364 136 2372 144
rect 2396 136 2404 144
rect 2732 136 2740 144
rect 2828 136 2836 144
rect 2252 116 2260 124
rect 2348 116 2356 124
rect 2380 116 2388 124
rect 2476 116 2484 124
rect 1116 96 1124 104
rect 2028 96 2036 104
rect 2908 176 2916 184
rect 3148 236 3156 244
rect 3420 1256 3428 1264
rect 3420 1196 3428 1204
rect 4284 1576 4292 1584
rect 4252 1456 4260 1464
rect 4252 1356 4260 1364
rect 3756 1316 3764 1324
rect 4028 1316 4036 1324
rect 4236 1256 4244 1264
rect 3836 1236 3844 1244
rect 4012 1236 4020 1244
rect 3644 1216 3652 1224
rect 3516 1196 3524 1204
rect 3644 1196 3652 1204
rect 3884 1196 3892 1204
rect 3916 1196 3924 1204
rect 3996 1196 4004 1204
rect 3500 1176 3508 1184
rect 3692 1096 3700 1104
rect 3724 1096 3732 1104
rect 3484 1076 3492 1084
rect 3452 1056 3460 1064
rect 3612 1056 3620 1064
rect 3580 996 3588 1004
rect 3420 956 3428 964
rect 3644 996 3652 1004
rect 3836 1076 3844 1084
rect 3804 1056 3812 1064
rect 3836 1056 3844 1064
rect 3804 936 3812 944
rect 3820 916 3828 924
rect 3532 736 3540 744
rect 3612 736 3620 744
rect 3436 716 3444 724
rect 3500 716 3508 724
rect 3356 636 3364 644
rect 3324 556 3332 564
rect 3484 616 3492 624
rect 3596 576 3604 584
rect 3564 536 3572 544
rect 3900 956 3908 964
rect 3932 1176 3940 1184
rect 3916 936 3924 944
rect 4092 1216 4100 1224
rect 4158 1206 4166 1214
rect 4172 1206 4180 1214
rect 4186 1206 4194 1214
rect 4044 1176 4052 1184
rect 4156 1176 4164 1184
rect 4124 1156 4132 1164
rect 4108 1136 4116 1144
rect 4252 1156 4260 1164
rect 4508 1756 4516 1764
rect 4668 2276 4676 2284
rect 4700 2176 4708 2184
rect 4668 2156 4676 2164
rect 4700 2156 4708 2164
rect 4764 2136 4772 2144
rect 4668 1976 4676 1984
rect 4652 1956 4660 1964
rect 4668 1956 4676 1964
rect 4652 1916 4660 1924
rect 4620 1896 4628 1904
rect 4652 1896 4660 1904
rect 4796 2096 4804 2104
rect 4860 2516 4868 2524
rect 4988 2516 4996 2524
rect 4828 2336 4836 2344
rect 4812 1936 4820 1944
rect 4684 1896 4692 1904
rect 4764 1896 4772 1904
rect 4860 2256 4868 2264
rect 4844 1916 4852 1924
rect 4652 1876 4660 1884
rect 4684 1876 4692 1884
rect 4588 1816 4596 1824
rect 4588 1776 4596 1784
rect 4588 1736 4596 1744
rect 4476 1716 4484 1724
rect 4572 1716 4580 1724
rect 4636 1716 4644 1724
rect 4540 1636 4548 1644
rect 4652 1636 4660 1644
rect 4572 1596 4580 1604
rect 4364 1536 4372 1544
rect 4412 1496 4420 1504
rect 4620 1496 4628 1504
rect 4332 1416 4340 1424
rect 4348 1396 4356 1404
rect 4316 1376 4324 1384
rect 4380 1356 4388 1364
rect 4508 1476 4516 1484
rect 4540 1416 4548 1424
rect 4572 1416 4580 1424
rect 4540 1336 4548 1344
rect 4364 1316 4372 1324
rect 4412 1316 4420 1324
rect 4444 1316 4452 1324
rect 4332 1256 4340 1264
rect 4284 1176 4292 1184
rect 3996 1096 4004 1104
rect 4060 1096 4068 1104
rect 4268 1096 4276 1104
rect 3980 1076 3988 1084
rect 4028 1076 4036 1084
rect 4076 1076 4084 1084
rect 4172 1076 4180 1084
rect 4252 1056 4260 1064
rect 4396 1176 4404 1184
rect 4540 1096 4548 1104
rect 4300 1076 4308 1084
rect 4508 1076 4516 1084
rect 4412 1056 4420 1064
rect 4300 996 4308 1004
rect 4668 1476 4676 1484
rect 4652 1176 4660 1184
rect 4588 1096 4596 1104
rect 4572 1056 4580 1064
rect 4524 996 4532 1004
rect 4604 996 4612 1004
rect 4284 976 4292 984
rect 4508 976 4516 984
rect 4284 956 4292 964
rect 4124 936 4132 944
rect 4428 936 4436 944
rect 4572 956 4580 964
rect 4588 936 4596 944
rect 3932 916 3940 924
rect 3948 916 3956 924
rect 4012 916 4020 924
rect 4508 916 4516 924
rect 3868 896 3876 904
rect 4092 896 4100 904
rect 3772 736 3780 744
rect 3900 736 3908 744
rect 3964 736 3972 744
rect 4380 876 4388 884
rect 4396 876 4404 884
rect 3980 716 3988 724
rect 4158 806 4166 814
rect 4172 806 4180 814
rect 4186 806 4194 814
rect 4044 716 4052 724
rect 4460 816 4468 824
rect 3996 696 4004 704
rect 4316 696 4324 704
rect 3884 676 3892 684
rect 3692 636 3700 644
rect 3724 616 3732 624
rect 3788 596 3796 604
rect 3756 556 3764 564
rect 3580 516 3588 524
rect 3676 516 3684 524
rect 3868 576 3876 584
rect 3948 596 3956 604
rect 3996 576 4004 584
rect 3884 536 3892 544
rect 3900 536 3908 544
rect 3932 536 3940 544
rect 4012 536 4020 544
rect 3484 336 3492 344
rect 3212 236 3220 244
rect 3004 176 3012 184
rect 3180 176 3188 184
rect 3036 156 3044 164
rect 3708 396 3716 404
rect 3596 296 3604 304
rect 3708 296 3716 304
rect 3660 276 3668 284
rect 3340 256 3348 264
rect 3372 216 3380 224
rect 3628 216 3636 224
rect 3532 196 3540 204
rect 3596 196 3604 204
rect 3308 176 3316 184
rect 3228 136 3236 144
rect 3132 116 3140 124
rect 2444 96 2452 104
rect 2508 96 2516 104
rect 2540 96 2548 104
rect 2812 96 2820 104
rect 2860 96 2868 104
rect 2156 16 2164 24
rect 1118 6 1126 14
rect 1132 6 1140 14
rect 1146 6 1154 14
rect 3292 136 3300 144
rect 3564 136 3572 144
rect 3692 136 3700 144
rect 3756 236 3764 244
rect 3948 396 3956 404
rect 3852 336 3860 344
rect 3772 196 3780 204
rect 4188 596 4196 604
rect 4156 556 4164 564
rect 4284 556 4292 564
rect 4460 596 4468 604
rect 4508 616 4516 624
rect 4540 696 4548 704
rect 4572 836 4580 844
rect 4604 916 4612 924
rect 4636 1116 4644 1124
rect 4668 1076 4676 1084
rect 4700 1856 4708 1864
rect 4748 1836 4756 1844
rect 4844 1756 4852 1764
rect 4732 1716 4740 1724
rect 4828 1716 4836 1724
rect 5148 2496 5156 2504
rect 4908 2476 4916 2484
rect 5004 2476 5012 2484
rect 4892 2336 4900 2344
rect 5532 2576 5540 2584
rect 5388 2316 5396 2324
rect 4924 2276 4932 2284
rect 5004 2256 5012 2264
rect 5148 2276 5156 2284
rect 5292 2276 5300 2284
rect 5068 2216 5076 2224
rect 5116 2216 5124 2224
rect 5036 2176 5044 2184
rect 5004 2136 5012 2144
rect 4892 2096 4900 2104
rect 4940 2016 4948 2024
rect 4876 1916 4884 1924
rect 4876 1896 4884 1904
rect 4956 1936 4964 1944
rect 4892 1816 4900 1824
rect 4860 1636 4868 1644
rect 4732 1556 4740 1564
rect 4700 1456 4708 1464
rect 4748 1456 4756 1464
rect 4796 1496 4804 1504
rect 5612 2796 5620 2804
rect 5580 2776 5588 2784
rect 5596 2716 5604 2724
rect 5644 2856 5652 2864
rect 5628 2696 5636 2704
rect 5628 2676 5636 2684
rect 5836 2896 5844 2904
rect 5868 2876 5876 2884
rect 5868 2796 5876 2804
rect 5724 2776 5732 2784
rect 5836 2756 5844 2764
rect 5980 2876 5988 2884
rect 5964 2836 5972 2844
rect 5916 2796 5924 2804
rect 5804 2696 5812 2704
rect 5596 2656 5604 2664
rect 5692 2656 5700 2664
rect 5660 2596 5668 2604
rect 5548 2536 5556 2544
rect 5852 2676 5860 2684
rect 5708 2636 5716 2644
rect 5788 2636 5796 2644
rect 5726 2606 5734 2614
rect 5740 2606 5748 2614
rect 5754 2606 5762 2614
rect 5692 2556 5700 2564
rect 5580 2516 5588 2524
rect 5756 2516 5764 2524
rect 5804 2596 5812 2604
rect 5932 2696 5940 2704
rect 6012 3056 6020 3064
rect 6076 3056 6084 3064
rect 6076 3016 6084 3024
rect 6028 2996 6036 3004
rect 6044 2976 6052 2984
rect 6028 2856 6036 2864
rect 5996 2816 6004 2824
rect 6124 2996 6132 3004
rect 6252 3696 6260 3704
rect 6220 3676 6228 3684
rect 6284 3696 6292 3704
rect 6268 3636 6276 3644
rect 6236 3536 6244 3544
rect 6268 3536 6276 3544
rect 6204 3516 6212 3524
rect 6236 3496 6244 3504
rect 6220 3476 6228 3484
rect 6252 3456 6260 3464
rect 6268 3436 6276 3444
rect 6204 3356 6212 3364
rect 6220 3356 6228 3364
rect 6252 3336 6260 3344
rect 6268 3336 6276 3344
rect 6188 3236 6196 3244
rect 6156 3216 6164 3224
rect 6188 3216 6196 3224
rect 6236 3156 6244 3164
rect 6316 4276 6324 4284
rect 6332 4236 6340 4244
rect 6316 4136 6324 4144
rect 6364 4476 6372 4484
rect 6524 4836 6532 4844
rect 6476 4736 6484 4744
rect 6524 4716 6532 4724
rect 6556 4696 6564 4704
rect 6396 4656 6404 4664
rect 6412 4656 6420 4664
rect 6444 4676 6452 4684
rect 6572 4676 6580 4684
rect 6492 4656 6500 4664
rect 6428 4636 6436 4644
rect 6588 4636 6596 4644
rect 6476 4596 6484 4604
rect 6556 4596 6564 4604
rect 6444 4576 6452 4584
rect 6524 4576 6532 4584
rect 6412 4536 6420 4544
rect 6380 4336 6388 4344
rect 6668 4736 6676 4744
rect 6524 4476 6532 4484
rect 6492 4416 6500 4424
rect 6476 4336 6484 4344
rect 6476 4236 6484 4244
rect 6444 4216 6452 4224
rect 6364 4096 6372 4104
rect 6476 4076 6484 4084
rect 6380 4016 6388 4024
rect 6396 3796 6404 3804
rect 6348 3776 6356 3784
rect 6380 3776 6388 3784
rect 6428 3776 6436 3784
rect 6348 3716 6356 3724
rect 6364 3676 6372 3684
rect 6332 3576 6340 3584
rect 6316 3556 6324 3564
rect 6412 3756 6420 3764
rect 6428 3736 6436 3744
rect 6396 3716 6404 3724
rect 6460 3896 6468 3904
rect 6476 3856 6484 3864
rect 6476 3736 6484 3744
rect 6396 3696 6404 3704
rect 6444 3696 6452 3704
rect 6364 3536 6372 3544
rect 6380 3536 6388 3544
rect 6348 3516 6356 3524
rect 6332 3476 6340 3484
rect 6332 3456 6340 3464
rect 6316 3416 6324 3424
rect 6412 3476 6420 3484
rect 6380 3416 6388 3424
rect 6348 3396 6356 3404
rect 6364 3376 6372 3384
rect 6348 3356 6356 3364
rect 6332 3316 6340 3324
rect 6364 3316 6372 3324
rect 6332 3296 6340 3304
rect 6300 3276 6308 3284
rect 6316 3276 6324 3284
rect 6284 3236 6292 3244
rect 6396 3296 6404 3304
rect 6396 3276 6404 3284
rect 6380 3196 6388 3204
rect 6332 3176 6340 3184
rect 6380 3156 6388 3164
rect 6268 3116 6276 3124
rect 6236 3096 6244 3104
rect 6076 2936 6084 2944
rect 6108 2936 6116 2944
rect 6204 2956 6212 2964
rect 6220 2936 6228 2944
rect 6172 2916 6180 2924
rect 6156 2896 6164 2904
rect 6252 3016 6260 3024
rect 6252 2956 6260 2964
rect 6236 2916 6244 2924
rect 6204 2896 6212 2904
rect 6252 2896 6260 2904
rect 6332 3096 6340 3104
rect 6348 3096 6356 3104
rect 6348 2976 6356 2984
rect 6316 2956 6324 2964
rect 6332 2956 6340 2964
rect 6140 2856 6148 2864
rect 6092 2836 6100 2844
rect 6044 2736 6052 2744
rect 6252 2856 6260 2864
rect 6172 2756 6180 2764
rect 5884 2576 5892 2584
rect 5884 2556 5892 2564
rect 5820 2536 5828 2544
rect 5932 2536 5940 2544
rect 6076 2696 6084 2704
rect 5996 2676 6004 2684
rect 6044 2676 6052 2684
rect 6284 2836 6292 2844
rect 6284 2776 6292 2784
rect 6236 2716 6244 2724
rect 6268 2716 6276 2724
rect 6364 2956 6372 2964
rect 6348 2836 6356 2844
rect 6300 2756 6308 2764
rect 6428 3356 6436 3364
rect 6412 3236 6420 3244
rect 6556 4336 6564 4344
rect 6508 4236 6516 4244
rect 6508 4096 6516 4104
rect 6508 4076 6516 4084
rect 6540 3936 6548 3944
rect 6492 3676 6500 3684
rect 6508 3676 6516 3684
rect 6476 3616 6484 3624
rect 6492 3616 6500 3624
rect 6460 3516 6468 3524
rect 6476 3496 6484 3504
rect 6444 3336 6452 3344
rect 6444 3316 6452 3324
rect 6428 3176 6436 3184
rect 6540 3616 6548 3624
rect 6508 3596 6516 3604
rect 6588 4276 6596 4284
rect 6700 4696 6708 4704
rect 6876 4696 6884 4704
rect 6748 4676 6756 4684
rect 6700 4496 6708 4504
rect 6684 4476 6692 4484
rect 6668 4256 6676 4264
rect 6700 4216 6708 4224
rect 6700 4136 6708 4144
rect 6812 4676 6820 4684
rect 6620 3876 6628 3884
rect 6780 3976 6788 3984
rect 6780 3916 6788 3924
rect 6700 3796 6708 3804
rect 6588 3736 6596 3744
rect 6556 3576 6564 3584
rect 6476 3456 6484 3464
rect 6492 3396 6500 3404
rect 6460 3256 6468 3264
rect 6444 3156 6452 3164
rect 6444 3116 6452 3124
rect 6428 3096 6436 3104
rect 6412 3076 6420 3084
rect 6396 3056 6404 3064
rect 6460 3036 6468 3044
rect 6524 3376 6532 3384
rect 6540 3336 6548 3344
rect 6556 3316 6564 3324
rect 6572 3316 6580 3324
rect 6508 3296 6516 3304
rect 6524 3296 6532 3304
rect 6492 3276 6500 3284
rect 6492 3236 6500 3244
rect 6476 2996 6484 3004
rect 6556 3136 6564 3144
rect 6524 3116 6532 3124
rect 6508 3076 6516 3084
rect 6556 2996 6564 3004
rect 6540 2976 6548 2984
rect 6508 2956 6516 2964
rect 6396 2936 6404 2944
rect 6460 2936 6468 2944
rect 6572 2936 6580 2944
rect 6348 2736 6356 2744
rect 6380 2736 6388 2744
rect 6412 2876 6420 2884
rect 6396 2716 6404 2724
rect 6364 2696 6372 2704
rect 6188 2676 6196 2684
rect 6124 2656 6132 2664
rect 6220 2656 6228 2664
rect 6012 2636 6020 2644
rect 5964 2596 5972 2604
rect 6300 2656 6308 2664
rect 6268 2636 6276 2644
rect 6028 2576 6036 2584
rect 6124 2576 6132 2584
rect 6220 2576 6228 2584
rect 6188 2536 6196 2544
rect 6284 2536 6292 2544
rect 6300 2536 6308 2544
rect 5884 2518 5892 2524
rect 5884 2516 5892 2518
rect 5948 2516 5956 2524
rect 6124 2516 6132 2524
rect 6140 2516 6148 2524
rect 6108 2376 6116 2384
rect 5564 2316 5572 2324
rect 5580 2316 5588 2324
rect 5660 2316 5668 2324
rect 5724 2316 5732 2324
rect 5500 2296 5508 2304
rect 5404 2276 5412 2284
rect 5340 2256 5348 2264
rect 5180 2176 5188 2184
rect 5276 2176 5284 2184
rect 5372 2156 5380 2164
rect 5036 2016 5044 2024
rect 5068 2016 5076 2024
rect 5100 1976 5108 1984
rect 5180 1956 5188 1964
rect 5068 1776 5076 1784
rect 5004 1716 5012 1724
rect 4972 1616 4980 1624
rect 4940 1596 4948 1604
rect 4924 1416 4932 1424
rect 4924 1356 4932 1364
rect 4764 1336 4772 1344
rect 4892 1336 4900 1344
rect 5036 1676 5044 1684
rect 5084 1716 5092 1724
rect 5420 2256 5428 2264
rect 5468 2256 5476 2264
rect 5484 2156 5492 2164
rect 5436 2136 5444 2144
rect 5452 2136 5460 2144
rect 5484 2136 5492 2144
rect 5452 2116 5460 2124
rect 5228 1956 5236 1964
rect 5164 1876 5172 1884
rect 5196 1876 5204 1884
rect 5276 2096 5284 2104
rect 5292 2076 5300 2084
rect 5260 2056 5268 2064
rect 5340 2056 5348 2064
rect 5452 1896 5460 1904
rect 5452 1876 5460 1884
rect 5164 1856 5172 1864
rect 5244 1856 5252 1864
rect 5260 1856 5268 1864
rect 5180 1836 5188 1844
rect 5308 1836 5316 1844
rect 5324 1836 5332 1844
rect 5132 1796 5140 1804
rect 5212 1816 5220 1824
rect 5308 1816 5316 1824
rect 5212 1776 5220 1784
rect 5100 1656 5108 1664
rect 5180 1656 5188 1664
rect 5084 1596 5092 1604
rect 5116 1576 5124 1584
rect 5084 1476 5092 1484
rect 5100 1456 5108 1464
rect 5068 1356 5076 1364
rect 4716 1156 4724 1164
rect 4700 1076 4708 1084
rect 4652 996 4660 1004
rect 4748 1176 4756 1184
rect 4828 1156 4836 1164
rect 4796 1136 4804 1144
rect 4764 1076 4772 1084
rect 4812 1076 4820 1084
rect 4844 1056 4852 1064
rect 4652 976 4660 984
rect 4716 976 4724 984
rect 4732 976 4740 984
rect 5020 1076 5028 1084
rect 4988 1056 4996 1064
rect 5068 1016 5076 1024
rect 4908 996 4916 1004
rect 4956 996 4964 1004
rect 4748 956 4756 964
rect 4876 956 4884 964
rect 5116 1096 5124 1104
rect 5212 1516 5220 1524
rect 5308 1516 5316 1524
rect 5148 1496 5156 1504
rect 5180 1496 5188 1504
rect 5196 1496 5204 1504
rect 5372 1836 5380 1844
rect 5404 1776 5412 1784
rect 5420 1756 5428 1764
rect 5564 2276 5572 2284
rect 5596 2276 5604 2284
rect 5548 2256 5556 2264
rect 5612 2256 5620 2264
rect 5516 2136 5524 2144
rect 5548 2136 5556 2144
rect 5644 2156 5652 2164
rect 5564 2096 5572 2104
rect 5516 2076 5524 2084
rect 5548 2076 5556 2084
rect 6524 2876 6532 2884
rect 6508 2816 6516 2824
rect 6460 2736 6468 2744
rect 6460 2716 6468 2724
rect 6444 2696 6452 2704
rect 6492 2696 6500 2704
rect 6428 2636 6436 2644
rect 6412 2596 6420 2604
rect 6428 2576 6436 2584
rect 6348 2556 6356 2564
rect 6412 2536 6420 2544
rect 6332 2516 6340 2524
rect 6444 2516 6452 2524
rect 6316 2496 6324 2504
rect 6444 2476 6452 2484
rect 6300 2376 6308 2384
rect 6476 2476 6484 2484
rect 6732 3736 6740 3744
rect 6812 3996 6820 4004
rect 6812 3976 6820 3984
rect 6796 3616 6804 3624
rect 6668 3596 6676 3604
rect 6700 3596 6708 3604
rect 6604 3496 6612 3504
rect 6620 3476 6628 3484
rect 6732 3456 6740 3464
rect 6764 3416 6772 3424
rect 6716 3356 6724 3364
rect 6668 3336 6676 3344
rect 6716 3336 6724 3344
rect 6668 3316 6676 3324
rect 6620 3296 6628 3304
rect 6636 3276 6644 3284
rect 6668 3276 6676 3284
rect 6748 3276 6756 3284
rect 6668 3256 6676 3264
rect 6684 3256 6692 3264
rect 6620 3176 6628 3184
rect 6604 3136 6612 3144
rect 6604 3116 6612 3124
rect 6636 3096 6644 3104
rect 6764 3196 6772 3204
rect 6732 3102 6740 3104
rect 6732 3096 6740 3102
rect 6652 3076 6660 3084
rect 6668 3016 6676 3024
rect 6732 3016 6740 3024
rect 6764 3016 6772 3024
rect 6700 2936 6708 2944
rect 6588 2816 6596 2824
rect 6588 2796 6596 2804
rect 6572 2756 6580 2764
rect 6540 2716 6548 2724
rect 6668 2756 6676 2764
rect 6604 2736 6612 2744
rect 6636 2736 6644 2744
rect 6636 2716 6644 2724
rect 6764 2736 6772 2744
rect 6572 2696 6580 2704
rect 6668 2696 6676 2704
rect 6524 2676 6532 2684
rect 6636 2676 6644 2684
rect 6652 2676 6660 2684
rect 6604 2576 6612 2584
rect 6556 2556 6564 2564
rect 6588 2556 6596 2564
rect 6588 2536 6596 2544
rect 6572 2516 6580 2524
rect 6524 2496 6532 2504
rect 6508 2396 6516 2404
rect 6236 2316 6244 2324
rect 6460 2316 6468 2324
rect 5852 2296 5860 2304
rect 6076 2296 6084 2304
rect 6204 2296 6212 2304
rect 5676 2276 5684 2284
rect 5660 2136 5668 2144
rect 5596 1936 5604 1944
rect 5612 1896 5620 1904
rect 5580 1856 5588 1864
rect 5564 1836 5572 1844
rect 5548 1816 5556 1824
rect 5548 1756 5556 1764
rect 5548 1736 5556 1744
rect 5340 1696 5348 1704
rect 5564 1696 5572 1704
rect 5468 1676 5476 1684
rect 5452 1636 5460 1644
rect 5340 1596 5348 1604
rect 5276 1476 5284 1484
rect 5404 1616 5412 1624
rect 5372 1556 5380 1564
rect 5468 1616 5476 1624
rect 5436 1596 5444 1604
rect 5372 1516 5380 1524
rect 5420 1516 5428 1524
rect 5164 1356 5172 1364
rect 5196 1356 5204 1364
rect 5148 1316 5156 1324
rect 5180 1276 5188 1284
rect 5164 1096 5172 1104
rect 5180 976 5188 984
rect 5036 956 5044 964
rect 5020 936 5028 944
rect 5084 936 5092 944
rect 5100 936 5108 944
rect 5180 936 5188 944
rect 5228 1156 5236 1164
rect 5212 1116 5220 1124
rect 5324 1456 5332 1464
rect 5388 1496 5396 1504
rect 5420 1496 5428 1504
rect 5500 1556 5508 1564
rect 5484 1456 5492 1464
rect 5260 1336 5268 1344
rect 5308 1318 5316 1324
rect 5308 1316 5316 1318
rect 5340 1296 5348 1304
rect 5372 1236 5380 1244
rect 5308 1196 5316 1204
rect 5260 1136 5268 1144
rect 5260 1116 5268 1124
rect 5244 1036 5252 1044
rect 5292 1056 5300 1064
rect 4764 876 4772 884
rect 4652 736 4660 744
rect 5020 736 5028 744
rect 4780 716 4788 724
rect 4636 676 4644 684
rect 4476 576 4484 584
rect 4412 536 4420 544
rect 4284 516 4292 524
rect 4396 516 4404 524
rect 4158 406 4166 414
rect 4172 406 4180 414
rect 4186 406 4194 414
rect 4268 376 4276 384
rect 4332 376 4340 384
rect 4076 356 4084 364
rect 4220 356 4228 364
rect 4140 336 4148 344
rect 4108 316 4116 324
rect 4108 296 4116 304
rect 4140 296 4148 304
rect 4620 656 4628 664
rect 4684 656 4692 664
rect 4972 656 4980 664
rect 5036 656 5044 664
rect 4492 536 4500 544
rect 4540 536 4548 544
rect 4572 536 4580 544
rect 4428 396 4436 404
rect 4348 316 4356 324
rect 4556 516 4564 524
rect 4540 416 4548 424
rect 4476 316 4484 324
rect 4572 376 4580 384
rect 4284 296 4292 304
rect 4348 296 4356 304
rect 4444 296 4452 304
rect 4012 276 4020 284
rect 4156 276 4164 284
rect 4268 276 4276 284
rect 4044 236 4052 244
rect 3884 196 3892 204
rect 3964 196 3972 204
rect 3932 156 3940 164
rect 4172 156 4180 164
rect 4124 136 4126 144
rect 4126 136 4132 144
rect 4188 136 4196 144
rect 4444 276 4452 284
rect 4412 196 4420 204
rect 4476 196 4484 204
rect 4748 596 4756 604
rect 4812 596 4820 604
rect 4908 576 4916 584
rect 4716 536 4724 544
rect 4620 516 4628 524
rect 4684 416 4692 424
rect 4636 376 4644 384
rect 4620 316 4628 324
rect 4668 316 4676 324
rect 4668 256 4676 264
rect 4732 376 4740 384
rect 4700 276 4708 284
rect 5084 716 5092 724
rect 5020 576 5028 584
rect 4924 536 4932 544
rect 4940 516 4948 524
rect 5004 516 5012 524
rect 4988 496 4996 504
rect 5052 556 5060 564
rect 5036 516 5044 524
rect 4972 476 4980 484
rect 4796 416 4804 424
rect 4780 396 4788 404
rect 4780 336 4788 344
rect 4764 296 4772 304
rect 4844 336 4852 344
rect 4828 316 4836 324
rect 4828 296 4836 304
rect 4860 316 4868 324
rect 4748 196 4756 204
rect 4844 196 4852 204
rect 4300 136 4308 144
rect 4380 136 4388 144
rect 4588 136 4596 144
rect 3244 116 3252 124
rect 3660 116 3668 124
rect 3788 116 3796 124
rect 3836 116 3844 124
rect 4044 116 4052 124
rect 4284 116 4292 124
rect 4492 116 4500 124
rect 4124 36 4132 44
rect 4156 36 4164 44
rect 4158 6 4166 14
rect 4172 6 4180 14
rect 4186 6 4194 14
rect 5372 1156 5380 1164
rect 5372 1096 5380 1104
rect 5324 1076 5332 1084
rect 5228 856 5236 864
rect 5132 736 5140 744
rect 5180 716 5188 724
rect 5116 656 5124 664
rect 5100 536 5108 544
rect 5148 516 5156 524
rect 5180 556 5188 564
rect 5196 556 5204 564
rect 5084 496 5092 504
rect 5068 476 5076 484
rect 5116 476 5124 484
rect 5148 456 5156 464
rect 5132 396 5140 404
rect 5052 336 5060 344
rect 5036 296 5044 304
rect 5036 276 5044 284
rect 4892 256 4900 264
rect 4988 256 4996 264
rect 4940 136 4948 144
rect 4764 116 4772 124
rect 4988 116 4996 124
rect 4924 16 4932 24
rect 5276 876 5284 884
rect 5356 956 5364 964
rect 5356 896 5364 904
rect 5372 896 5380 904
rect 5484 1396 5492 1404
rect 5468 1376 5476 1384
rect 5404 1356 5412 1364
rect 5436 1336 5444 1344
rect 5468 1316 5476 1324
rect 5404 1296 5412 1304
rect 5388 716 5396 724
rect 5420 1116 5428 1124
rect 5436 1116 5444 1124
rect 5420 1076 5428 1084
rect 5452 1076 5460 1084
rect 5500 1316 5508 1324
rect 5500 1276 5508 1284
rect 5644 1896 5652 1904
rect 5628 1836 5636 1844
rect 5596 1716 5604 1724
rect 5932 2236 5940 2244
rect 5868 2216 5876 2224
rect 5964 2216 5972 2224
rect 5726 2206 5734 2214
rect 5740 2206 5748 2214
rect 5754 2206 5762 2214
rect 5804 2176 5812 2184
rect 5772 2136 5780 2144
rect 5900 2136 5908 2144
rect 5996 2136 6004 2144
rect 6076 2136 6084 2144
rect 6108 2136 6116 2144
rect 6332 2296 6340 2304
rect 6268 2236 6276 2244
rect 6284 2236 6292 2244
rect 6460 2236 6468 2244
rect 6428 2216 6436 2224
rect 6492 2216 6500 2224
rect 6556 2156 6564 2164
rect 6316 2136 6324 2144
rect 6460 2136 6468 2144
rect 6620 2556 6628 2564
rect 6652 2516 6660 2524
rect 6636 2496 6644 2504
rect 6684 2516 6692 2524
rect 6684 2496 6692 2504
rect 6748 2518 6756 2524
rect 6748 2516 6756 2518
rect 6684 2236 6692 2244
rect 6732 2436 6740 2444
rect 6620 2156 6628 2164
rect 5692 2116 5700 2124
rect 5788 2116 5796 2124
rect 5980 2116 5988 2124
rect 6124 2116 6130 2124
rect 6130 2116 6132 2124
rect 6556 2116 6564 2124
rect 6588 2116 6596 2124
rect 5676 2096 5684 2104
rect 5788 2096 5796 2104
rect 5820 1956 5828 1964
rect 5788 1936 5796 1944
rect 5756 1916 5764 1924
rect 5772 1896 5780 1904
rect 5884 1896 5892 1904
rect 5628 1696 5636 1704
rect 5612 1596 5620 1604
rect 5580 1556 5588 1564
rect 5564 1476 5572 1484
rect 5548 1456 5556 1464
rect 5532 1396 5540 1404
rect 5532 1356 5540 1364
rect 5564 1276 5572 1284
rect 5644 1516 5652 1524
rect 5628 1496 5636 1504
rect 5612 1376 5620 1384
rect 5596 1316 5604 1324
rect 5516 1196 5524 1204
rect 5500 1136 5508 1144
rect 5516 1116 5524 1124
rect 5532 1116 5540 1124
rect 5580 1156 5588 1164
rect 5580 1116 5588 1124
rect 5532 1076 5540 1084
rect 5548 1076 5556 1084
rect 5468 1036 5476 1044
rect 5484 1016 5492 1024
rect 5420 756 5428 764
rect 5356 696 5364 704
rect 5388 702 5396 704
rect 5388 696 5396 702
rect 5404 696 5412 704
rect 5324 676 5332 684
rect 5436 716 5444 724
rect 5420 636 5428 644
rect 5292 556 5300 564
rect 5404 556 5412 564
rect 5244 536 5252 544
rect 5388 536 5396 544
rect 5228 516 5236 524
rect 5212 396 5220 404
rect 5148 376 5156 384
rect 5436 536 5444 544
rect 5516 916 5524 924
rect 5532 896 5540 904
rect 5532 876 5540 884
rect 5644 1236 5652 1244
rect 5612 1136 5620 1144
rect 5628 1116 5636 1124
rect 5692 1876 5700 1884
rect 5676 1496 5684 1504
rect 5852 1856 5860 1864
rect 5820 1836 5828 1844
rect 5726 1806 5734 1814
rect 5740 1806 5748 1814
rect 5754 1806 5762 1814
rect 5932 2096 5940 2104
rect 5900 1856 5908 1864
rect 5916 1836 5924 1844
rect 5772 1776 5780 1784
rect 5868 1776 5876 1784
rect 5788 1756 5796 1764
rect 5820 1716 5828 1724
rect 5692 1476 5700 1484
rect 5676 1436 5684 1444
rect 5820 1696 5828 1704
rect 5804 1656 5812 1664
rect 5820 1636 5828 1644
rect 5772 1616 5780 1624
rect 5740 1556 5748 1564
rect 5740 1516 5748 1524
rect 5788 1556 5796 1564
rect 5916 1696 5924 1704
rect 5852 1616 5860 1624
rect 6028 2096 6036 2104
rect 6012 2076 6020 2084
rect 6364 1956 6372 1964
rect 6220 1936 6228 1944
rect 6316 1936 6324 1944
rect 5980 1916 5988 1924
rect 6204 1916 6212 1924
rect 6284 1916 6292 1924
rect 6300 1916 6308 1924
rect 5964 1876 5972 1884
rect 6092 1896 6100 1904
rect 6172 1876 6180 1884
rect 5980 1856 5988 1864
rect 5980 1836 5988 1844
rect 5980 1756 5988 1764
rect 6156 1836 6164 1844
rect 6124 1816 6132 1824
rect 6140 1756 6148 1764
rect 6076 1736 6084 1744
rect 5948 1716 5956 1724
rect 6188 1836 6196 1844
rect 6396 1936 6404 1944
rect 6236 1896 6244 1904
rect 6252 1876 6260 1884
rect 6300 1876 6308 1884
rect 6316 1876 6324 1884
rect 6220 1816 6228 1824
rect 6172 1756 6180 1764
rect 6236 1756 6244 1764
rect 6156 1716 6164 1724
rect 6044 1676 6052 1684
rect 6028 1656 6036 1664
rect 5948 1636 5956 1644
rect 5884 1596 5892 1604
rect 5932 1596 5940 1604
rect 5820 1496 5828 1504
rect 5804 1476 5812 1484
rect 5676 1316 5684 1324
rect 5660 1156 5668 1164
rect 5596 1076 5604 1084
rect 5628 1036 5636 1044
rect 5564 1016 5572 1024
rect 5612 936 5620 944
rect 5564 816 5572 824
rect 5596 896 5604 904
rect 5580 796 5588 804
rect 5564 776 5572 784
rect 5532 696 5540 704
rect 5516 636 5524 644
rect 5516 576 5524 584
rect 5308 516 5316 524
rect 5340 496 5348 504
rect 5404 496 5412 504
rect 5468 456 5476 464
rect 5484 456 5492 464
rect 5308 376 5316 384
rect 5276 336 5284 344
rect 5388 336 5396 344
rect 5436 336 5444 344
rect 5244 316 5252 324
rect 5164 296 5172 304
rect 5308 296 5316 304
rect 5372 276 5380 284
rect 5340 256 5348 264
rect 5356 256 5364 264
rect 5132 196 5140 204
rect 5212 196 5220 204
rect 5500 356 5508 364
rect 5644 956 5652 964
rect 5676 936 5684 944
rect 5644 916 5652 924
rect 5628 896 5636 904
rect 5612 696 5620 704
rect 5676 856 5684 864
rect 5580 656 5588 664
rect 5596 616 5604 624
rect 5580 576 5588 584
rect 5532 516 5540 524
rect 5468 296 5476 304
rect 5404 276 5412 284
rect 5404 256 5412 264
rect 5548 496 5556 504
rect 5726 1406 5734 1414
rect 5740 1406 5748 1414
rect 5754 1406 5762 1414
rect 5852 1536 5860 1544
rect 5852 1496 5860 1504
rect 5996 1576 6004 1584
rect 5948 1536 5956 1544
rect 5932 1516 5940 1524
rect 5916 1476 5924 1484
rect 5916 1456 5924 1464
rect 5900 1436 5908 1444
rect 5884 1396 5892 1404
rect 5884 1376 5892 1384
rect 5724 1296 5732 1304
rect 5724 1216 5732 1224
rect 5868 1316 5876 1324
rect 5900 1296 5908 1304
rect 5932 1316 5940 1324
rect 5964 1436 5972 1444
rect 5964 1396 5972 1404
rect 5996 1396 6004 1404
rect 6012 1356 6020 1364
rect 5820 1276 5828 1284
rect 5788 1196 5796 1204
rect 5740 1076 5748 1084
rect 5772 1036 5780 1044
rect 5726 1006 5734 1014
rect 5740 1006 5748 1014
rect 5754 1006 5762 1014
rect 5756 956 5764 964
rect 5724 916 5732 924
rect 5740 916 5748 924
rect 5692 816 5700 824
rect 5692 716 5700 724
rect 5724 816 5732 824
rect 5772 736 5780 744
rect 5804 1116 5812 1124
rect 5868 1176 5876 1184
rect 5852 1156 5860 1164
rect 5900 1136 5908 1144
rect 5836 1096 5844 1104
rect 5868 1096 5876 1104
rect 5916 1096 5924 1104
rect 5852 1076 5860 1084
rect 5804 956 5812 964
rect 5836 976 5844 984
rect 5820 776 5828 784
rect 5804 756 5812 764
rect 5820 756 5828 764
rect 5884 1056 5892 1064
rect 5900 1036 5908 1044
rect 5900 816 5908 824
rect 5868 756 5876 764
rect 5836 736 5844 744
rect 5852 736 5860 744
rect 5852 696 5860 704
rect 5676 656 5684 664
rect 5726 606 5734 614
rect 5740 606 5748 614
rect 5754 606 5762 614
rect 5692 596 5700 604
rect 5804 596 5812 604
rect 5676 556 5684 564
rect 5836 616 5844 624
rect 5820 576 5828 584
rect 5964 1296 5972 1304
rect 6012 1316 6020 1324
rect 5996 1296 6004 1304
rect 5980 1276 5988 1284
rect 5948 1256 5956 1264
rect 5996 1196 6004 1204
rect 5964 1156 5972 1164
rect 6012 1116 6020 1124
rect 5948 1076 5956 1084
rect 5996 1076 6004 1084
rect 6012 1036 6020 1044
rect 5996 956 6004 964
rect 6300 1756 6308 1764
rect 6268 1716 6276 1724
rect 6188 1696 6196 1704
rect 6236 1676 6244 1684
rect 6284 1696 6292 1704
rect 6268 1656 6276 1664
rect 6268 1596 6276 1604
rect 6140 1536 6148 1544
rect 6220 1536 6228 1544
rect 6204 1496 6212 1504
rect 6060 1476 6068 1484
rect 6044 1376 6052 1384
rect 6092 1396 6100 1404
rect 6060 1336 6068 1344
rect 6140 1416 6148 1424
rect 6124 1336 6132 1344
rect 6172 1336 6180 1344
rect 6204 1316 6212 1324
rect 6108 1296 6116 1304
rect 6172 1296 6180 1304
rect 6204 1296 6212 1304
rect 6044 1156 6052 1164
rect 6044 976 6052 984
rect 6028 916 6036 924
rect 5964 896 5972 904
rect 6364 1816 6372 1824
rect 6412 1796 6420 1804
rect 6524 1976 6532 1984
rect 6476 1956 6484 1964
rect 6460 1776 6468 1784
rect 6396 1716 6404 1724
rect 6428 1716 6436 1724
rect 6364 1696 6372 1704
rect 6460 1696 6468 1704
rect 6380 1676 6388 1684
rect 6332 1576 6340 1584
rect 6300 1516 6308 1524
rect 6284 1496 6292 1504
rect 6252 1456 6260 1464
rect 6252 1376 6260 1384
rect 6236 1256 6244 1264
rect 6204 1216 6212 1224
rect 6172 1136 6180 1144
rect 6268 1176 6276 1184
rect 6252 1136 6260 1144
rect 6124 1056 6132 1064
rect 6236 1056 6244 1064
rect 6108 1016 6116 1024
rect 6156 1016 6164 1024
rect 6220 996 6228 1004
rect 6188 936 6196 944
rect 6108 916 6116 924
rect 6012 716 6020 724
rect 6028 656 6036 664
rect 5932 596 5940 604
rect 5884 576 5892 584
rect 5996 576 6004 584
rect 5948 556 5956 564
rect 5612 536 5620 544
rect 5852 536 5860 544
rect 5628 496 5636 504
rect 5692 476 5700 484
rect 5884 476 5892 484
rect 5596 376 5604 384
rect 5564 336 5572 344
rect 5516 316 5524 324
rect 5532 316 5540 324
rect 5676 336 5684 344
rect 5916 456 5924 464
rect 5980 536 5988 544
rect 5964 516 5972 524
rect 5724 336 5732 344
rect 5932 336 5940 344
rect 5564 296 5572 304
rect 5660 296 5668 304
rect 5836 296 5844 304
rect 5500 276 5508 284
rect 5596 276 5604 284
rect 5916 276 5924 284
rect 5726 206 5734 214
rect 5740 206 5748 214
rect 5754 206 5762 214
rect 5468 176 5476 184
rect 5180 136 5188 144
rect 5052 116 5060 124
rect 5084 116 5092 124
rect 5292 116 5300 124
rect 5756 176 5764 184
rect 6124 756 6132 764
rect 6108 736 6116 744
rect 6092 636 6100 644
rect 6028 516 6036 524
rect 5996 496 6004 504
rect 6204 916 6212 924
rect 6204 896 6212 904
rect 6172 876 6180 884
rect 6172 796 6180 804
rect 6140 616 6148 624
rect 6124 596 6132 604
rect 6124 476 6132 484
rect 6188 536 6196 544
rect 6204 496 6212 504
rect 6156 436 6164 444
rect 6092 376 6100 384
rect 6092 336 6100 344
rect 6108 336 6116 344
rect 6252 976 6260 984
rect 6236 936 6244 944
rect 6252 756 6260 764
rect 6236 736 6244 744
rect 6268 716 6276 724
rect 6332 1336 6340 1344
rect 6316 1236 6324 1244
rect 6300 1156 6308 1164
rect 6300 1076 6308 1084
rect 6300 1036 6308 1044
rect 6300 936 6308 944
rect 6364 1396 6372 1404
rect 6348 1236 6356 1244
rect 6348 1196 6356 1204
rect 6412 1556 6420 1564
rect 6508 1936 6516 1944
rect 6492 1916 6500 1924
rect 6508 1836 6516 1844
rect 6652 2136 6660 2144
rect 6636 1956 6644 1964
rect 6604 1856 6612 1864
rect 6556 1796 6564 1804
rect 6524 1736 6532 1744
rect 6492 1676 6500 1684
rect 6556 1596 6564 1604
rect 6492 1576 6500 1584
rect 6476 1556 6484 1564
rect 6460 1536 6468 1544
rect 6428 1456 6436 1464
rect 6396 1416 6404 1424
rect 6460 1456 6468 1464
rect 6476 1416 6484 1424
rect 6444 1396 6452 1404
rect 6460 1336 6468 1344
rect 6380 1316 6388 1324
rect 6540 1536 6548 1544
rect 6556 1536 6564 1544
rect 6508 1496 6516 1504
rect 6508 1336 6516 1344
rect 6412 1296 6420 1304
rect 6444 1276 6452 1284
rect 6412 1216 6420 1224
rect 6380 1196 6388 1204
rect 6396 1176 6404 1184
rect 6380 1156 6388 1164
rect 6348 1096 6356 1104
rect 6476 1096 6484 1104
rect 6348 1076 6356 1084
rect 6380 1056 6388 1064
rect 6364 936 6372 944
rect 6300 916 6308 924
rect 6364 916 6372 924
rect 6332 776 6340 784
rect 6300 716 6308 724
rect 6268 556 6276 564
rect 6284 536 6292 544
rect 6348 696 6356 704
rect 6476 1056 6484 1064
rect 6428 996 6436 1004
rect 6604 1816 6612 1824
rect 6620 1816 6628 1824
rect 6588 1796 6596 1804
rect 6588 1756 6596 1764
rect 6572 1376 6580 1384
rect 6572 1356 6580 1364
rect 6540 1336 6548 1344
rect 6524 1316 6532 1324
rect 6524 1156 6532 1164
rect 6524 1136 6532 1144
rect 6572 1136 6580 1144
rect 6444 936 6452 944
rect 6460 916 6468 924
rect 6428 736 6436 744
rect 6444 736 6452 744
rect 6460 716 6468 724
rect 6396 696 6404 704
rect 6428 696 6436 704
rect 6364 636 6372 644
rect 6364 616 6372 624
rect 6348 536 6356 544
rect 6364 536 6372 544
rect 6252 516 6260 524
rect 6332 436 6340 444
rect 6364 436 6372 444
rect 6284 416 6292 424
rect 6252 376 6260 384
rect 5980 296 5988 304
rect 6044 276 6052 284
rect 5884 176 5892 184
rect 5964 176 5972 184
rect 5596 156 5604 164
rect 5820 156 5828 164
rect 6076 156 6084 164
rect 5468 116 5476 124
rect 6188 316 6196 324
rect 6172 276 6180 284
rect 6188 276 6196 284
rect 6140 216 6148 224
rect 6140 176 6148 184
rect 6220 316 6228 324
rect 6012 96 6020 104
rect 6092 96 6100 104
rect 6268 336 6276 344
rect 6316 316 6324 324
rect 6300 296 6308 304
rect 6300 276 6308 284
rect 6252 196 6260 204
rect 6396 636 6404 644
rect 6428 536 6436 544
rect 6460 536 6468 544
rect 6412 516 6420 524
rect 6380 416 6388 424
rect 6364 376 6372 384
rect 6380 376 6388 384
rect 6348 336 6356 344
rect 6380 356 6388 364
rect 6364 256 6372 264
rect 6444 496 6452 504
rect 6524 696 6532 704
rect 6604 1496 6612 1504
rect 6716 2116 6724 2124
rect 6716 1936 6724 1944
rect 6652 1896 6660 1904
rect 6716 1896 6724 1904
rect 6668 1856 6676 1864
rect 6700 1856 6708 1864
rect 6652 1816 6660 1824
rect 6748 2296 6756 2304
rect 6732 1816 6740 1824
rect 6796 3436 6804 3444
rect 6876 3296 6884 3304
rect 6812 3196 6820 3204
rect 6860 3116 6868 3124
rect 6812 3016 6820 3024
rect 6876 2576 6884 2584
rect 6860 2056 6868 2064
rect 6796 1996 6804 2004
rect 6828 1976 6836 1984
rect 6780 1936 6788 1944
rect 6764 1916 6772 1924
rect 6876 1896 6884 1904
rect 6764 1876 6772 1884
rect 6780 1836 6788 1844
rect 6748 1796 6756 1804
rect 6716 1776 6724 1784
rect 6828 1816 6836 1824
rect 6716 1736 6724 1744
rect 6748 1736 6756 1744
rect 6812 1736 6820 1744
rect 6684 1556 6692 1564
rect 6700 1536 6708 1544
rect 6748 1716 6756 1724
rect 6844 1796 6852 1804
rect 6828 1676 6836 1684
rect 6764 1636 6772 1644
rect 6636 1516 6644 1524
rect 6716 1516 6724 1524
rect 6684 1496 6692 1504
rect 6700 1456 6708 1464
rect 6716 1376 6724 1384
rect 6652 1316 6660 1324
rect 6684 1316 6692 1324
rect 6604 1296 6612 1304
rect 6684 1296 6692 1304
rect 6668 1116 6676 1124
rect 6604 1096 6612 1104
rect 6588 956 6596 964
rect 6572 936 6580 944
rect 6540 656 6548 664
rect 6540 556 6548 564
rect 6508 536 6516 544
rect 6460 476 6468 484
rect 6476 476 6484 484
rect 6476 336 6484 344
rect 6748 1196 6756 1204
rect 6732 1076 6740 1084
rect 6700 876 6708 884
rect 6636 776 6644 784
rect 6636 716 6644 724
rect 6604 536 6612 544
rect 6668 776 6676 784
rect 6700 756 6708 764
rect 6668 696 6676 704
rect 6684 656 6692 664
rect 6668 536 6676 544
rect 6684 536 6692 544
rect 6508 516 6516 524
rect 6604 516 6612 524
rect 6508 476 6516 484
rect 6588 436 6596 444
rect 6540 336 6548 344
rect 6636 456 6644 464
rect 6684 496 6692 504
rect 6668 376 6676 384
rect 6636 356 6644 364
rect 6668 356 6676 364
rect 6508 316 6516 324
rect 6604 316 6612 324
rect 6620 316 6628 324
rect 6492 296 6500 304
rect 6476 276 6484 284
rect 6492 216 6500 224
rect 6428 196 6436 204
rect 6412 176 6420 184
rect 6284 156 6292 164
rect 6300 156 6308 164
rect 6396 156 6404 164
rect 6284 136 6292 144
rect 6620 296 6628 304
rect 6588 276 6596 284
rect 6604 276 6612 284
rect 6540 176 6548 184
rect 6316 136 6324 144
rect 6620 176 6628 184
rect 6812 1616 6820 1624
rect 6844 1616 6852 1624
rect 6780 1516 6788 1524
rect 6796 1496 6804 1504
rect 6796 1316 6804 1324
rect 6812 1236 6820 1244
rect 6844 1236 6852 1244
rect 6796 1116 6804 1124
rect 6780 1096 6788 1104
rect 6812 1096 6820 1104
rect 6812 1036 6820 1044
rect 6764 836 6772 844
rect 6716 676 6724 684
rect 6732 676 6740 684
rect 6716 656 6724 664
rect 6828 996 6836 1004
rect 6780 576 6788 584
rect 6732 556 6740 564
rect 6716 496 6724 504
rect 6716 476 6724 484
rect 6716 316 6724 324
rect 6780 516 6788 524
rect 6764 496 6772 504
rect 6828 836 6836 844
rect 6876 1096 6884 1104
rect 6860 976 6868 984
rect 6844 756 6852 764
rect 6844 736 6852 744
rect 6812 496 6820 504
rect 6860 556 6868 564
rect 6876 536 6884 544
rect 6812 456 6820 464
rect 6844 456 6852 464
rect 6796 436 6804 444
rect 6844 336 6852 344
rect 6748 296 6756 304
rect 6732 276 6740 284
rect 6748 276 6756 284
rect 6732 256 6740 264
rect 6876 256 6884 264
rect 6812 236 6820 244
rect 6588 136 6596 144
rect 6700 136 6708 144
rect 6396 116 6404 124
rect 6556 116 6564 124
rect 6732 116 6740 124
rect 6844 116 6852 124
rect 6300 96 6308 104
rect 6540 96 6548 104
rect 6812 96 6820 104
rect 6236 76 6244 84
rect 6364 76 6372 84
<< metal3 >>
rect 2632 5014 2680 5016
rect 2632 5006 2636 5014
rect 2646 5006 2652 5014
rect 2660 5006 2666 5014
rect 2676 5006 2680 5014
rect 2632 5004 2680 5006
rect 5720 5014 5768 5016
rect 5720 5006 5724 5014
rect 5734 5006 5740 5014
rect 5748 5006 5754 5014
rect 5764 5006 5768 5014
rect 5720 5004 5768 5006
rect 2244 4997 2252 5003
rect 4852 4977 4876 4983
rect 6324 4977 6716 4983
rect 868 4957 1612 4963
rect 1844 4957 2220 4963
rect 2228 4957 2396 4963
rect 2925 4957 3148 4963
rect 2925 4944 2931 4957
rect 3156 4957 3628 4963
rect 3876 4957 4300 4963
rect 4628 4957 5084 4963
rect 5124 4957 5324 4963
rect 5684 4957 5788 4963
rect 5796 4957 6060 4963
rect 6068 4957 6684 4963
rect 148 4937 348 4943
rect 596 4937 876 4943
rect 1108 4937 1484 4943
rect 1620 4937 2012 4943
rect 2052 4937 2252 4943
rect 2500 4937 2748 4943
rect 2756 4937 2924 4943
rect 3044 4937 3340 4943
rect 3460 4937 3660 4943
rect 4340 4937 4396 4943
rect 4660 4937 4764 4943
rect 5300 4937 5388 4943
rect 5396 4937 5452 4943
rect 5860 4937 6252 4943
rect 260 4917 492 4923
rect 1284 4917 1356 4923
rect 1668 4917 1868 4923
rect 1988 4917 2140 4923
rect 2372 4917 2620 4923
rect 2916 4917 3020 4923
rect 3236 4917 3548 4923
rect 3636 4917 4028 4923
rect 4061 4923 4067 4936
rect 4061 4917 4364 4923
rect 4868 4917 4924 4923
rect 4932 4917 5260 4923
rect 5428 4917 5708 4923
rect 5876 4917 6028 4923
rect 372 4897 396 4903
rect 420 4897 460 4903
rect 468 4897 860 4903
rect 948 4897 1516 4903
rect 1572 4897 1644 4903
rect 5300 4897 5388 4903
rect 884 4877 956 4883
rect 1556 4877 1676 4883
rect 5236 4877 5596 4883
rect 708 4857 1756 4863
rect 5124 4857 5356 4863
rect 788 4837 892 4843
rect 1236 4837 1340 4843
rect 1348 4837 1372 4843
rect 1604 4837 2060 4843
rect 3316 4837 3340 4843
rect 4020 4837 4060 4843
rect 5492 4837 5516 4843
rect 6356 4837 6524 4843
rect 116 4817 140 4823
rect 1492 4817 2524 4823
rect 2532 4817 2812 4823
rect 3332 4817 3468 4823
rect 3476 4817 3596 4823
rect 5012 4817 5036 4823
rect 1112 4814 1160 4816
rect 1112 4806 1116 4814
rect 1126 4806 1132 4814
rect 1140 4806 1146 4814
rect 1156 4806 1160 4814
rect 1112 4804 1160 4806
rect 4152 4814 4200 4816
rect 4152 4806 4156 4814
rect 4166 4806 4172 4814
rect 4180 4806 4186 4814
rect 4196 4806 4200 4814
rect 4152 4804 4200 4806
rect 4100 4777 4220 4783
rect 4276 4777 4332 4783
rect 4340 4777 5276 4783
rect 404 4757 940 4763
rect 724 4737 780 4743
rect 852 4737 988 4743
rect 1652 4737 1676 4743
rect 3268 4737 3772 4743
rect 6484 4737 6668 4743
rect 340 4717 364 4723
rect 372 4717 428 4723
rect 692 4717 1324 4723
rect 1732 4717 1804 4723
rect 3172 4717 3196 4723
rect 3316 4717 3580 4723
rect 3668 4717 3724 4723
rect 3764 4717 3980 4723
rect 4212 4717 4284 4723
rect 5268 4717 5308 4723
rect 5844 4717 6012 4723
rect 6100 4717 6172 4723
rect 6180 4717 6348 4723
rect 6532 4717 6540 4723
rect 740 4697 828 4703
rect 1060 4697 1260 4703
rect 1316 4697 1388 4703
rect 1396 4697 1628 4703
rect 1700 4697 1788 4703
rect 1796 4697 1948 4703
rect 2164 4697 2412 4703
rect 2740 4697 2764 4703
rect 3012 4697 3276 4703
rect 3284 4697 3356 4703
rect 3364 4697 3468 4703
rect 3492 4697 3532 4703
rect 4212 4697 4236 4703
rect 4308 4697 4460 4703
rect 5508 4697 5788 4703
rect 6004 4697 6060 4703
rect 6068 4697 6124 4703
rect 6132 4697 6220 4703
rect 6276 4697 6348 4703
rect 6452 4697 6556 4703
rect 6884 4697 6915 4703
rect 228 4677 380 4683
rect 468 4677 924 4683
rect 932 4677 940 4683
rect 948 4677 1596 4683
rect 1780 4677 1804 4683
rect 1812 4677 2300 4683
rect 2324 4677 2524 4683
rect 3108 4677 3219 4683
rect 3213 4664 3219 4677
rect 3252 4677 3324 4683
rect 3444 4677 3612 4683
rect 3908 4677 4156 4683
rect 4372 4677 4652 4683
rect 4932 4677 5420 4683
rect 5700 4677 5772 4683
rect 5860 4677 5964 4683
rect 6020 4677 6092 4683
rect 6349 4683 6355 4696
rect 6349 4677 6444 4683
rect 6516 4677 6572 4683
rect 6756 4677 6812 4683
rect 724 4657 764 4663
rect 836 4657 1116 4663
rect 1252 4657 1292 4663
rect 1652 4657 1740 4663
rect 1748 4657 1836 4663
rect 2804 4657 2940 4663
rect 2996 4657 3100 4663
rect 3220 4657 3404 4663
rect 3412 4657 3436 4663
rect 3476 4657 3532 4663
rect 3540 4657 3708 4663
rect 3716 4657 3820 4663
rect 4244 4657 4540 4663
rect 4756 4657 4844 4663
rect 4852 4657 4924 4663
rect 4964 4657 5084 4663
rect 5092 4657 5132 4663
rect 5188 4657 5596 4663
rect 5604 4657 5676 4663
rect 5684 4657 5756 4663
rect 5780 4657 5900 4663
rect 6116 4657 6204 4663
rect 6212 4657 6316 4663
rect 6324 4657 6364 4663
rect 6372 4657 6396 4663
rect 6420 4657 6492 4663
rect 596 4637 684 4643
rect 820 4637 988 4643
rect 1284 4637 1340 4643
rect 1412 4637 1468 4643
rect 1572 4637 1612 4643
rect 1620 4637 1820 4643
rect 3396 4637 3436 4643
rect 4356 4637 5180 4643
rect 5508 4637 5532 4643
rect 5901 4643 5907 4656
rect 5901 4637 6348 4643
rect 6356 4637 6428 4643
rect 6596 4637 6732 4643
rect 868 4617 1004 4623
rect 1012 4617 1196 4623
rect 1300 4617 1500 4623
rect 1988 4617 2204 4623
rect 3204 4617 3500 4623
rect 3604 4617 3868 4623
rect 3940 4617 4540 4623
rect 4548 4617 4620 4623
rect 4852 4617 4892 4623
rect 5524 4617 5532 4623
rect 5940 4617 6108 4623
rect 6180 4617 6220 4623
rect 6228 4617 6316 4623
rect 2632 4614 2680 4616
rect 2632 4606 2636 4614
rect 2646 4606 2652 4614
rect 2660 4606 2666 4614
rect 2676 4606 2680 4614
rect 2632 4604 2680 4606
rect 5720 4614 5768 4616
rect 5720 4606 5724 4614
rect 5734 4606 5740 4614
rect 5748 4606 5754 4614
rect 5764 4606 5768 4614
rect 5720 4604 5768 4606
rect 196 4597 556 4603
rect 564 4597 844 4603
rect 2820 4597 2956 4603
rect 3508 4597 3708 4603
rect 3716 4597 3900 4603
rect 3940 4597 4348 4603
rect 5156 4597 5420 4603
rect 5524 4597 5692 4603
rect 6484 4597 6556 4603
rect 1732 4577 1756 4583
rect 2036 4577 2444 4583
rect 3316 4577 3484 4583
rect 6068 4577 6444 4583
rect 6532 4577 6572 4583
rect 788 4557 876 4563
rect 884 4557 988 4563
rect 996 4557 1180 4563
rect 1188 4557 1292 4563
rect 2836 4557 2924 4563
rect 3060 4557 3084 4563
rect 3364 4557 3452 4563
rect 3460 4557 3516 4563
rect 3572 4557 3756 4563
rect 4036 4557 4108 4563
rect 4516 4557 4780 4563
rect 4820 4557 4972 4563
rect 5108 4557 5308 4563
rect 6132 4557 6156 4563
rect 6164 4557 6252 4563
rect 356 4537 460 4543
rect 868 4537 1100 4543
rect 1108 4537 1244 4543
rect 1636 4537 1644 4543
rect 1860 4537 1996 4543
rect 2804 4537 3004 4543
rect 3124 4537 3196 4543
rect 3316 4537 3388 4543
rect 3396 4537 3468 4543
rect 3556 4537 3660 4543
rect 3796 4537 3820 4543
rect 3988 4537 4140 4543
rect 4436 4537 4732 4543
rect 5268 4537 5468 4543
rect 5924 4537 5948 4543
rect 5956 4537 6060 4543
rect 6100 4537 6332 4543
rect 6340 4537 6412 4543
rect 308 4517 444 4523
rect 676 4517 732 4523
rect 1076 4517 1276 4523
rect 1460 4517 1500 4523
rect 1556 4517 1628 4523
rect 1652 4517 1708 4523
rect 1748 4517 1804 4523
rect 1972 4517 2092 4523
rect 2148 4517 2188 4523
rect 2580 4517 2604 4523
rect 2724 4517 2796 4523
rect 3236 4517 3324 4523
rect 3492 4517 3564 4523
rect 3588 4517 3692 4523
rect 3700 4517 3724 4523
rect 3748 4517 3884 4523
rect 5636 4517 5708 4523
rect 5828 4517 6220 4523
rect 148 4497 220 4503
rect 324 4497 412 4503
rect 420 4497 428 4503
rect 500 4497 636 4503
rect 644 4497 652 4503
rect 708 4497 844 4503
rect 1428 4497 1612 4503
rect 1748 4497 1852 4503
rect 3684 4497 3772 4503
rect 3780 4497 3804 4503
rect 4772 4497 4780 4503
rect 5428 4497 5500 4503
rect 5556 4497 5964 4503
rect 6004 4497 6172 4503
rect 6212 4497 6284 4503
rect 6644 4497 6700 4503
rect 36 4477 396 4483
rect 1572 4477 1820 4483
rect 1828 4477 1932 4483
rect 2228 4477 2268 4483
rect 3156 4477 3212 4483
rect 3220 4477 3276 4483
rect 3828 4477 3884 4483
rect 4964 4477 5932 4483
rect 5940 4477 6028 4483
rect 6276 4477 6300 4483
rect 6372 4477 6524 4483
rect 6532 4477 6684 4483
rect 212 4457 556 4463
rect 724 4457 860 4463
rect 1124 4457 1276 4463
rect 3076 4457 3260 4463
rect 3268 4457 3628 4463
rect 4004 4457 4364 4463
rect 4372 4457 5500 4463
rect 6132 4457 6284 4463
rect 20 4437 268 4443
rect 276 4437 396 4443
rect 740 4437 972 4443
rect 1044 4437 1164 4443
rect 2772 4437 2812 4443
rect 3300 4437 3356 4443
rect 3364 4437 3420 4443
rect 3428 4437 3724 4443
rect 3908 4437 3948 4443
rect 4868 4437 4988 4443
rect 5156 4437 5468 4443
rect 244 4417 364 4423
rect 3188 4417 3404 4423
rect 3508 4417 3548 4423
rect 3556 4417 3692 4423
rect 4020 4417 4076 4423
rect 4388 4417 4460 4423
rect 6500 4417 6508 4423
rect 1112 4414 1160 4416
rect 1112 4406 1116 4414
rect 1126 4406 1132 4414
rect 1140 4406 1146 4414
rect 1156 4406 1160 4414
rect 1112 4404 1160 4406
rect 4152 4414 4200 4416
rect 4152 4406 4156 4414
rect 4166 4406 4172 4414
rect 4180 4406 4186 4414
rect 4196 4406 4200 4414
rect 4152 4404 4200 4406
rect 1380 4397 1484 4403
rect 1492 4397 1692 4403
rect 1700 4397 1980 4403
rect 3636 4397 3836 4403
rect 4276 4397 4380 4403
rect 4788 4397 4844 4403
rect 420 4377 652 4383
rect 660 4377 700 4383
rect 708 4377 1548 4383
rect 2196 4377 2316 4383
rect 3428 4377 3468 4383
rect 4836 4377 4956 4383
rect 5140 4377 5180 4383
rect 5220 4377 5436 4383
rect 5444 4377 5516 4383
rect 564 4357 1388 4363
rect 1620 4357 1788 4363
rect 3236 4357 3308 4363
rect 3460 4357 3484 4363
rect 3668 4357 3692 4363
rect 3828 4357 4060 4363
rect 452 4337 764 4343
rect 1524 4337 1692 4343
rect 2260 4337 2476 4343
rect 3204 4337 3276 4343
rect 3284 4337 3644 4343
rect 3652 4337 3708 4343
rect 3716 4337 3724 4343
rect 5076 4337 6380 4343
rect 6388 4337 6476 4343
rect 6484 4337 6556 4343
rect 20 4317 268 4323
rect 276 4317 332 4323
rect 573 4317 668 4323
rect 573 4304 579 4317
rect 852 4317 988 4323
rect 1476 4317 1596 4323
rect 1700 4317 1772 4323
rect 2180 4317 2284 4323
rect 2292 4317 2348 4323
rect 2996 4317 3036 4323
rect 3332 4317 3452 4323
rect 3460 4317 3564 4323
rect 3661 4317 3676 4323
rect 148 4297 236 4303
rect 356 4297 364 4303
rect 372 4297 428 4303
rect 436 4297 572 4303
rect 660 4297 844 4303
rect 1220 4297 1228 4303
rect 1236 4297 1340 4303
rect 1540 4297 1596 4303
rect 1636 4297 1804 4303
rect 1908 4297 2012 4303
rect 2116 4297 2252 4303
rect 2964 4297 3004 4303
rect 3012 4297 3052 4303
rect 3060 4297 3132 4303
rect 3188 4297 3340 4303
rect 3348 4297 3404 4303
rect 3661 4303 3667 4317
rect 3684 4317 3740 4323
rect 3812 4317 3836 4323
rect 3844 4317 3868 4323
rect 3892 4317 4492 4323
rect 5476 4317 5548 4323
rect 5556 4317 5580 4323
rect 5844 4317 5964 4323
rect 5972 4317 6092 4323
rect 3469 4297 3667 4303
rect 756 4277 780 4283
rect 1540 4277 1612 4283
rect 1652 4277 1788 4283
rect 1796 4277 1868 4283
rect 1876 4277 1916 4283
rect 2164 4277 2355 4283
rect 2349 4264 2355 4277
rect 2468 4277 2604 4283
rect 2740 4277 2828 4283
rect 2964 4277 2972 4283
rect 3060 4277 3132 4283
rect 3469 4283 3475 4297
rect 3684 4297 3900 4303
rect 4516 4297 4684 4303
rect 4692 4297 5020 4303
rect 5044 4297 5084 4303
rect 5092 4297 5292 4303
rect 5508 4297 5836 4303
rect 6308 4297 6316 4303
rect 3332 4277 3475 4283
rect 3492 4277 3596 4283
rect 3764 4277 3852 4283
rect 3924 4277 3964 4283
rect 4644 4277 5068 4283
rect 5236 4277 5340 4283
rect 5348 4277 5356 4283
rect 5364 4277 5612 4283
rect 5748 4277 5996 4283
rect 6324 4277 6588 4283
rect 644 4257 796 4263
rect 804 4257 876 4263
rect 1812 4257 1852 4263
rect 1892 4257 1932 4263
rect 2148 4257 2172 4263
rect 2356 4257 2412 4263
rect 2452 4257 2572 4263
rect 2580 4257 2812 4263
rect 2932 4257 2988 4263
rect 3076 4257 3196 4263
rect 3220 4257 3260 4263
rect 3300 4257 3356 4263
rect 3380 4257 3436 4263
rect 3476 4257 3548 4263
rect 3620 4257 3788 4263
rect 3956 4257 3980 4263
rect 3988 4257 4428 4263
rect 4820 4257 5196 4263
rect 5268 4257 5420 4263
rect 5428 4257 5612 4263
rect 5716 4257 5948 4263
rect 5956 4257 6172 4263
rect 6180 4257 6668 4263
rect 468 4237 876 4243
rect 1604 4237 1644 4243
rect 1860 4237 2060 4243
rect 3092 4237 3228 4243
rect 3476 4237 3484 4243
rect 3572 4237 3660 4243
rect 3716 4237 3884 4243
rect 5028 4237 5180 4243
rect 5204 4237 5260 4243
rect 5300 4237 5356 4243
rect 5364 4237 5628 4243
rect 6020 4237 6076 4243
rect 6164 4237 6332 4243
rect 6484 4237 6508 4243
rect 740 4217 780 4223
rect 788 4217 1196 4223
rect 1204 4217 1340 4223
rect 1348 4217 1708 4223
rect 2100 4217 2444 4223
rect 3220 4217 3404 4223
rect 3444 4217 3452 4223
rect 3476 4217 3836 4223
rect 4260 4217 4300 4223
rect 4708 4217 4844 4223
rect 5060 4217 5276 4223
rect 5524 4217 5692 4223
rect 6452 4217 6700 4223
rect 2632 4214 2680 4216
rect 2632 4206 2636 4214
rect 2646 4206 2652 4214
rect 2660 4206 2666 4214
rect 2676 4206 2680 4214
rect 2632 4204 2680 4206
rect 5720 4214 5768 4216
rect 5720 4206 5724 4214
rect 5734 4206 5740 4214
rect 5748 4206 5754 4214
rect 5764 4206 5768 4214
rect 5720 4204 5768 4206
rect 1012 4197 1036 4203
rect 1412 4197 1676 4203
rect 1684 4197 1740 4203
rect 2132 4197 2156 4203
rect 2708 4197 2796 4203
rect 2820 4197 2860 4203
rect 3348 4197 3436 4203
rect 3508 4197 3532 4203
rect 3540 4197 3708 4203
rect 3716 4197 3852 4203
rect 4372 4197 4412 4203
rect 4500 4197 5404 4203
rect 5412 4197 5548 4203
rect 356 4177 556 4183
rect 564 4177 588 4183
rect 916 4177 972 4183
rect 1556 4177 1820 4183
rect 2932 4177 3580 4183
rect 3588 4177 3628 4183
rect 3636 4177 3788 4183
rect 3844 4177 3996 4183
rect 4644 4177 4924 4183
rect 5556 4177 5980 4183
rect 228 4157 300 4163
rect 324 4157 428 4163
rect 436 4157 508 4163
rect 1316 4157 1356 4163
rect 1700 4157 1708 4163
rect 2372 4157 2572 4163
rect 2580 4157 2780 4163
rect 3044 4157 3164 4163
rect 3252 4157 3340 4163
rect 3348 4157 3468 4163
rect 3492 4157 3612 4163
rect 3780 4157 3900 4163
rect 3908 4157 3916 4163
rect 3956 4157 4012 4163
rect 4228 4157 4332 4163
rect 4340 4157 4524 4163
rect 4532 4157 4668 4163
rect 5412 4157 5868 4163
rect 5972 4157 6124 4163
rect 6708 4157 6764 4163
rect 228 4137 268 4143
rect 516 4137 796 4143
rect 852 4137 988 4143
rect 1044 4137 1164 4143
rect 1252 4137 1372 4143
rect 1524 4137 1708 4143
rect 1716 4137 1836 4143
rect 1844 4137 1948 4143
rect 2212 4137 2268 4143
rect 2276 4137 2380 4143
rect 2484 4137 2588 4143
rect 3268 4137 3628 4143
rect 3636 4137 3868 4143
rect 3940 4137 3980 4143
rect 4868 4137 4892 4143
rect 4980 4137 5020 4143
rect 5076 4137 5292 4143
rect 5620 4137 5644 4143
rect 5668 4137 5676 4143
rect 6228 4137 6236 4143
rect 6244 4137 6316 4143
rect 6708 4137 6828 4143
rect 84 4117 236 4123
rect 532 4117 588 4123
rect 628 4117 684 4123
rect 932 4117 1292 4123
rect 1300 4117 1500 4123
rect 1652 4117 1772 4123
rect 1780 4117 1804 4123
rect 2244 4117 2444 4123
rect 3284 4117 3532 4123
rect 3572 4117 3596 4123
rect 3732 4117 3756 4123
rect 3764 4117 3820 4123
rect 3892 4117 4028 4123
rect 4484 4117 4508 4123
rect 4516 4117 4540 4123
rect 4884 4117 4956 4123
rect 4964 4117 5036 4123
rect 5044 4117 5388 4123
rect 5396 4117 5516 4123
rect 5556 4117 5596 4123
rect 5684 4117 6220 4123
rect 196 4097 268 4103
rect 580 4097 620 4103
rect 644 4097 652 4103
rect 660 4097 1148 4103
rect 1380 4097 1548 4103
rect 1748 4097 1884 4103
rect 2420 4097 2476 4103
rect 3044 4097 3324 4103
rect 3332 4097 3356 4103
rect 3524 4097 3612 4103
rect 3700 4097 3804 4103
rect 3812 4097 4092 4103
rect 5012 4097 5036 4103
rect 5428 4097 5484 4103
rect 5508 4097 5564 4103
rect 5604 4097 5756 4103
rect 6276 4097 6364 4103
rect 6372 4097 6508 4103
rect 260 4077 284 4083
rect 404 4077 652 4083
rect 948 4077 1276 4083
rect 1284 4077 1484 4083
rect 3124 4077 3228 4083
rect 3236 4077 3372 4083
rect 3444 4077 3516 4083
rect 3604 4077 3644 4083
rect 3668 4077 3692 4083
rect 3732 4077 3772 4083
rect 3796 4077 3852 4083
rect 3860 4077 3932 4083
rect 4756 4077 5100 4083
rect 5108 4077 5180 4083
rect 5492 4077 5516 4083
rect 5716 4077 6060 4083
rect 6484 4077 6508 4083
rect 484 4057 620 4063
rect 628 4057 796 4063
rect 1156 4057 1260 4063
rect 1268 4057 1724 4063
rect 2548 4057 2684 4063
rect 3140 4057 3148 4063
rect 3348 4057 3404 4063
rect 3412 4057 3820 4063
rect 3876 4057 3964 4063
rect 548 4037 780 4043
rect 788 4037 1324 4043
rect 1332 4037 1932 4043
rect 2868 4037 2972 4043
rect 3412 4037 3660 4043
rect 3748 4037 3916 4043
rect 4836 4037 4876 4043
rect 4948 4037 5292 4043
rect 5316 4037 5324 4043
rect 212 4017 508 4023
rect 516 4017 556 4023
rect 564 4017 988 4023
rect 2020 4017 2044 4023
rect 2852 4017 2908 4023
rect 3476 4017 3500 4023
rect 3508 4017 3580 4023
rect 3620 4017 3900 4023
rect 3908 4017 4060 4023
rect 5076 4017 5212 4023
rect 1112 4014 1160 4016
rect 1112 4006 1116 4014
rect 1126 4006 1132 4014
rect 1140 4006 1146 4014
rect 1156 4006 1160 4014
rect 1112 4004 1160 4006
rect 4152 4014 4200 4016
rect 4152 4006 4156 4014
rect 4166 4006 4172 4014
rect 4180 4006 4186 4014
rect 4196 4006 4200 4014
rect 4152 4004 4200 4006
rect 308 3997 636 4003
rect 676 3997 1020 4003
rect 1396 3997 1788 4003
rect 2756 3997 3004 4003
rect 3188 3997 3212 4003
rect 3348 3997 3404 4003
rect 3556 3997 3756 4003
rect 3780 3997 3916 4003
rect 3924 3997 3948 4003
rect 4324 3997 5052 4003
rect 6084 3997 6284 4003
rect 6516 3997 6812 4003
rect 244 3977 428 3983
rect 692 3977 1404 3983
rect 2788 3977 3180 3983
rect 3188 3977 3740 3983
rect 4916 3977 5100 3983
rect 6788 3977 6812 3983
rect 372 3957 716 3963
rect 900 3957 956 3963
rect 1044 3957 1228 3963
rect 1268 3957 1292 3963
rect 1332 3957 1388 3963
rect 1780 3957 2716 3963
rect 3156 3957 3196 3963
rect 3204 3957 3500 3963
rect 3588 3957 3612 3963
rect 4788 3957 4812 3963
rect 4884 3957 5036 3963
rect 5236 3957 5356 3963
rect 5364 3957 5452 3963
rect 5652 3957 5900 3963
rect 5908 3957 6124 3963
rect 6132 3957 6204 3963
rect 6212 3957 6220 3963
rect 148 3937 476 3943
rect 820 3937 1084 3943
rect 1140 3937 1180 3943
rect 1204 3937 1244 3943
rect 1252 3937 1356 3943
rect 1428 3937 1436 3943
rect 1773 3937 1884 3943
rect 1773 3924 1779 3937
rect 2276 3937 2332 3943
rect 2340 3937 2428 3943
rect 2516 3937 2588 3943
rect 3060 3937 3260 3943
rect 3348 3937 3436 3943
rect 3460 3937 3628 3943
rect 3636 3937 3692 3943
rect 3748 3937 4172 3943
rect 4868 3937 4988 3943
rect 4996 3937 5148 3943
rect 5204 3937 5468 3943
rect 5700 3937 6044 3943
rect 6100 3937 6540 3943
rect 212 3917 252 3923
rect 436 3917 492 3923
rect 788 3917 844 3923
rect 1044 3917 1212 3923
rect 1300 3917 1436 3923
rect 1588 3917 1724 3923
rect 1764 3917 1772 3923
rect 1876 3917 1932 3923
rect 1940 3917 2012 3923
rect 2212 3917 2348 3923
rect 2356 3917 2380 3923
rect 3156 3917 3372 3923
rect 3444 3917 3628 3923
rect 3668 3917 3756 3923
rect 3764 3917 3868 3923
rect 4932 3917 5068 3923
rect 5460 3917 5548 3923
rect 5636 3917 6188 3923
rect 6196 3917 6780 3923
rect -19 3897 12 3903
rect 260 3897 332 3903
rect 340 3897 396 3903
rect 484 3897 524 3903
rect 836 3897 1084 3903
rect 1188 3897 1276 3903
rect 1284 3897 1340 3903
rect 1412 3897 1484 3903
rect 1956 3897 1996 3903
rect 2036 3897 2764 3903
rect 3044 3897 3884 3903
rect 4404 3897 4492 3903
rect 4868 3897 5068 3903
rect 5092 3897 5148 3903
rect 5156 3897 5212 3903
rect 5284 3897 5916 3903
rect 6116 3897 6236 3903
rect 6420 3897 6460 3903
rect 308 3877 380 3883
rect 580 3877 604 3883
rect 660 3877 700 3883
rect 884 3877 1196 3883
rect 1284 3877 1388 3883
rect 1396 3877 1452 3883
rect 1492 3877 1676 3883
rect 1780 3877 1884 3883
rect 2004 3877 2108 3883
rect 2404 3877 2476 3883
rect 2932 3877 3020 3883
rect 3028 3877 3132 3883
rect 3300 3877 3596 3883
rect 3604 3877 3724 3883
rect 3844 3877 4284 3883
rect 4308 3877 4364 3883
rect 4372 3877 4412 3883
rect 4484 3877 4828 3883
rect 4852 3877 4908 3883
rect 4916 3877 5036 3883
rect 5060 3877 5100 3883
rect 5108 3877 5164 3883
rect 5172 3877 5228 3883
rect 5348 3877 5788 3883
rect 5796 3877 6140 3883
rect 6196 3877 6620 3883
rect 340 3857 668 3863
rect 980 3857 1292 3863
rect 1428 3857 1436 3863
rect 1508 3857 1516 3863
rect 1876 3857 1964 3863
rect 2420 3857 2524 3863
rect 3252 3857 3356 3863
rect 3444 3857 3468 3863
rect 3476 3857 3596 3863
rect 4788 3857 4940 3863
rect 5172 3857 5196 3863
rect 5220 3857 5356 3863
rect 5572 3857 5884 3863
rect 6100 3857 6108 3863
rect 6116 3857 6268 3863
rect 6356 3857 6476 3863
rect 500 3837 796 3843
rect 1172 3837 1276 3843
rect 1300 3837 1660 3843
rect 1668 3837 1900 3843
rect 1908 3837 1948 3843
rect 1956 3837 2172 3843
rect 2180 3837 2316 3843
rect 2324 3837 2364 3843
rect 2548 3837 2924 3843
rect 2932 3837 2956 3843
rect 3044 3837 3084 3843
rect 3092 3837 3116 3843
rect 3140 3837 3980 3843
rect 4692 3837 4844 3843
rect 4948 3837 5308 3843
rect 5620 3837 5708 3843
rect 5844 3837 5868 3843
rect 5876 3837 6156 3843
rect 244 3817 300 3823
rect 308 3817 748 3823
rect 1156 3817 1356 3823
rect 1364 3817 1516 3823
rect 1636 3817 1660 3823
rect 1668 3817 1804 3823
rect 2292 3817 2412 3823
rect 2916 3817 2956 3823
rect 3188 3817 3372 3823
rect 3428 3817 3516 3823
rect 3524 3817 3628 3823
rect 3988 3817 3996 3823
rect 4084 3817 4252 3823
rect 4644 3817 4892 3823
rect 5044 3817 5116 3823
rect 5188 3817 5404 3823
rect 5412 3817 5644 3823
rect 5652 3817 5676 3823
rect 5860 3817 6044 3823
rect 2632 3814 2680 3816
rect 2632 3806 2636 3814
rect 2646 3806 2652 3814
rect 2660 3806 2666 3814
rect 2676 3806 2680 3814
rect 2632 3804 2680 3806
rect 5720 3814 5768 3816
rect 5720 3806 5724 3814
rect 5734 3806 5740 3814
rect 5748 3806 5754 3814
rect 5764 3806 5768 3814
rect 5720 3804 5768 3806
rect 228 3797 956 3803
rect 1460 3797 1500 3803
rect 1508 3797 1580 3803
rect 1700 3797 2124 3803
rect 2132 3797 2508 3803
rect 3204 3797 3244 3803
rect 3588 3797 3628 3803
rect 3668 3797 3676 3803
rect 4276 3797 4908 3803
rect 5236 3797 5372 3803
rect 6404 3797 6700 3803
rect 372 3777 476 3783
rect 548 3777 652 3783
rect 1492 3777 1852 3783
rect 1876 3777 1964 3783
rect 1972 3777 2540 3783
rect 3220 3777 3324 3783
rect 3396 3777 3468 3783
rect 3476 3777 3772 3783
rect 4036 3777 4924 3783
rect 4948 3777 5260 3783
rect 5316 3777 5436 3783
rect 5684 3777 5708 3783
rect 5780 3777 5804 3783
rect 6196 3777 6348 3783
rect 6388 3777 6428 3783
rect 340 3757 460 3763
rect 580 3757 636 3763
rect 676 3757 700 3763
rect 724 3757 828 3763
rect 836 3757 1340 3763
rect 1348 3757 1372 3763
rect 1780 3757 1932 3763
rect 2068 3757 2300 3763
rect 2356 3757 2508 3763
rect 2836 3757 2876 3763
rect 2884 3757 2924 3763
rect 2996 3757 3068 3763
rect 3108 3757 3164 3763
rect 3220 3757 3260 3763
rect 3428 3757 3532 3763
rect 3620 3757 3676 3763
rect 4340 3757 4524 3763
rect 4532 3757 4668 3763
rect 4900 3757 5004 3763
rect 5268 3757 5404 3763
rect 5412 3757 5692 3763
rect 5732 3757 5820 3763
rect 6004 3757 6380 3763
rect 6388 3757 6412 3763
rect 196 3737 284 3743
rect 292 3737 524 3743
rect 532 3737 652 3743
rect 708 3737 812 3743
rect 1236 3737 1260 3743
rect 1396 3737 1740 3743
rect 1796 3737 2140 3743
rect 2212 3737 2300 3743
rect 2372 3737 2716 3743
rect 2852 3737 2940 3743
rect 3204 3737 3244 3743
rect 3444 3737 4028 3743
rect 5124 3737 5340 3743
rect 5380 3737 6076 3743
rect 6084 3737 6188 3743
rect 6292 3737 6316 3743
rect 6436 3737 6476 3743
rect 6580 3737 6588 3743
rect 6740 3737 6796 3743
rect 84 3717 300 3723
rect 452 3717 684 3723
rect 804 3717 908 3723
rect 948 3717 956 3723
rect 1092 3717 1196 3723
rect 1204 3717 1372 3723
rect 1620 3717 1708 3723
rect 1764 3717 1836 3723
rect 2276 3717 2844 3723
rect 2852 3717 2860 3723
rect 3268 3717 3292 3723
rect 3412 3717 3468 3723
rect 3620 3717 3628 3723
rect 3636 3717 3756 3723
rect 4036 3717 4124 3723
rect 4468 3717 4572 3723
rect 4916 3717 5004 3723
rect 5012 3717 5116 3723
rect 5172 3717 5564 3723
rect 5572 3717 5692 3723
rect 5796 3717 5820 3723
rect 5828 3717 5916 3723
rect 5988 3717 6028 3723
rect 6356 3717 6396 3723
rect 436 3697 556 3703
rect 628 3697 732 3703
rect 989 3697 1036 3703
rect 989 3683 995 3697
rect 1124 3697 1228 3703
rect 1636 3697 1868 3703
rect 2052 3697 2412 3703
rect 3204 3697 3372 3703
rect 3389 3697 3500 3703
rect 628 3677 995 3683
rect 1012 3677 1148 3683
rect 1172 3677 1180 3683
rect 1188 3677 1340 3683
rect 2189 3677 2332 3683
rect 676 3657 780 3663
rect 948 3657 1084 3663
rect 2189 3663 2195 3677
rect 3389 3683 3395 3697
rect 3588 3697 3660 3703
rect 3668 3697 3708 3703
rect 3732 3697 3788 3703
rect 3812 3697 3852 3703
rect 3892 3697 3932 3703
rect 4836 3697 5036 3703
rect 5300 3697 5324 3703
rect 5332 3697 5452 3703
rect 5789 3703 5795 3716
rect 5460 3697 5795 3703
rect 5805 3697 6092 3703
rect 3172 3677 3395 3683
rect 3412 3677 3484 3683
rect 3492 3677 3948 3683
rect 4116 3677 4492 3683
rect 5108 3677 5468 3683
rect 5636 3677 5708 3683
rect 5805 3683 5811 3697
rect 6100 3697 6188 3703
rect 6260 3697 6284 3703
rect 6404 3697 6444 3703
rect 5732 3677 5811 3683
rect 5892 3677 5932 3683
rect 6228 3677 6364 3683
rect 6484 3677 6492 3683
rect 6516 3677 6572 3683
rect 1236 3657 2195 3663
rect 2212 3657 2812 3663
rect 3012 3657 3244 3663
rect 3284 3657 3436 3663
rect 3492 3657 3692 3663
rect 3764 3657 3804 3663
rect 3828 3657 3932 3663
rect 4180 3657 4220 3663
rect 5364 3657 5980 3663
rect 5988 3657 6124 3663
rect 948 3637 972 3643
rect 1044 3637 2396 3643
rect 3028 3637 4028 3643
rect 4036 3637 4332 3643
rect 5316 3637 6268 3643
rect 1284 3617 1660 3623
rect 2788 3617 3260 3623
rect 3348 3617 3724 3623
rect 3764 3617 3980 3623
rect 4340 3617 4364 3623
rect 5204 3617 5436 3623
rect 5540 3617 5548 3623
rect 6484 3617 6492 3623
rect 6500 3617 6540 3623
rect 6548 3617 6796 3623
rect 1112 3614 1160 3616
rect 1112 3606 1116 3614
rect 1126 3606 1132 3614
rect 1140 3606 1146 3614
rect 1156 3606 1160 3614
rect 1112 3604 1160 3606
rect 4152 3614 4200 3616
rect 4152 3606 4156 3614
rect 4166 3606 4172 3614
rect 4180 3606 4186 3614
rect 4196 3606 4200 3614
rect 4152 3604 4200 3606
rect 196 3597 428 3603
rect 2132 3597 3100 3603
rect 3108 3597 3324 3603
rect 3364 3597 3420 3603
rect 3780 3597 3804 3603
rect 5396 3597 5420 3603
rect 5492 3597 5644 3603
rect 5908 3597 6508 3603
rect 6676 3597 6700 3603
rect 388 3577 460 3583
rect 468 3577 924 3583
rect 932 3577 1068 3583
rect 1172 3577 1212 3583
rect 1508 3577 1516 3583
rect 3156 3577 3292 3583
rect 3316 3577 3340 3583
rect 3508 3577 3660 3583
rect 4020 3577 4236 3583
rect 4244 3577 4284 3583
rect 4292 3577 4428 3583
rect 4820 3577 4876 3583
rect 5476 3577 6332 3583
rect 6564 3577 6700 3583
rect 260 3557 348 3563
rect 596 3557 700 3563
rect 964 3557 1324 3563
rect 1332 3557 1356 3563
rect 1364 3557 1692 3563
rect 2052 3557 2812 3563
rect 2820 3557 2908 3563
rect 3124 3557 3148 3563
rect 3156 3557 3436 3563
rect 3444 3557 3468 3563
rect 3492 3557 3564 3563
rect 5204 3557 5324 3563
rect 5508 3557 5612 3563
rect 5620 3557 5788 3563
rect 6068 3557 6316 3563
rect 308 3537 396 3543
rect 692 3537 780 3543
rect 1076 3537 1148 3543
rect 1204 3537 1260 3543
rect 1572 3537 1628 3543
rect 1636 3537 2284 3543
rect 2372 3537 2732 3543
rect 3124 3537 3164 3543
rect 3172 3537 3276 3543
rect 3284 3537 3308 3543
rect 3332 3537 3740 3543
rect 3764 3537 3820 3543
rect 5236 3537 5308 3543
rect 5428 3537 5660 3543
rect 5812 3537 6236 3543
rect 6276 3537 6364 3543
rect 244 3517 268 3523
rect 388 3517 531 3523
rect 525 3504 531 3517
rect 660 3517 700 3523
rect 724 3517 748 3523
rect 900 3517 908 3523
rect 1012 3517 1260 3523
rect 1316 3517 1388 3523
rect 1556 3517 1580 3523
rect 1604 3517 1644 3523
rect 2228 3517 2284 3523
rect 2980 3517 3020 3523
rect 3060 3517 3180 3523
rect 3236 3517 3363 3523
rect 244 3497 348 3503
rect 436 3497 476 3503
rect 532 3497 556 3503
rect 644 3497 780 3503
rect 868 3497 1148 3503
rect 1188 3497 1212 3503
rect 1268 3497 1324 3503
rect 2244 3497 2316 3503
rect 2420 3497 2444 3503
rect 2548 3497 2572 3503
rect 3140 3497 3212 3503
rect 3252 3497 3340 3503
rect 3357 3503 3363 3517
rect 3396 3517 3571 3523
rect 3565 3504 3571 3517
rect 4356 3517 5283 3523
rect 3357 3497 3436 3503
rect 3444 3497 3532 3503
rect 3572 3497 3708 3503
rect 3716 3497 3820 3503
rect 4164 3497 4252 3503
rect 4676 3497 4780 3503
rect 5108 3497 5260 3503
rect 5277 3503 5283 3517
rect 5396 3517 5452 3523
rect 5469 3517 5484 3523
rect 5469 3503 5475 3517
rect 5524 3517 5580 3523
rect 5636 3517 5724 3523
rect 5796 3517 5852 3523
rect 6212 3517 6348 3523
rect 6468 3517 6604 3523
rect 5277 3497 5475 3503
rect 5492 3497 5516 3503
rect 5572 3497 5868 3503
rect 6004 3497 6140 3503
rect 6244 3497 6476 3503
rect 6484 3497 6604 3503
rect 84 3477 268 3483
rect 356 3477 620 3483
rect 740 3477 1052 3483
rect 1060 3477 1420 3483
rect 1428 3477 1532 3483
rect 1540 3477 1612 3483
rect 2260 3477 2300 3483
rect 2388 3477 2540 3483
rect 2980 3477 3036 3483
rect 3044 3477 3116 3483
rect 3140 3477 3196 3483
rect 3220 3477 3244 3483
rect 3252 3477 3372 3483
rect 3380 3477 3660 3483
rect 3668 3477 3676 3483
rect 3684 3477 3756 3483
rect 3764 3477 3868 3483
rect 4068 3477 4140 3483
rect 4724 3477 4764 3483
rect 4772 3477 4780 3483
rect 4788 3477 4908 3483
rect 4964 3477 5036 3483
rect 5284 3477 5340 3483
rect 5540 3477 5628 3483
rect 5828 3477 6108 3483
rect 6228 3477 6332 3483
rect 6340 3477 6355 3483
rect 260 3457 332 3463
rect 340 3457 716 3463
rect 884 3457 1132 3463
rect 1140 3457 1292 3463
rect 1332 3457 1388 3463
rect 1412 3457 1628 3463
rect 2212 3457 2700 3463
rect 3092 3457 3196 3463
rect 3300 3457 3404 3463
rect 3428 3457 3484 3463
rect 3652 3457 3660 3463
rect 3860 3457 4060 3463
rect 4276 3457 4316 3463
rect 4580 3457 4764 3463
rect 4868 3457 4908 3463
rect 4948 3457 5100 3463
rect 5124 3457 5212 3463
rect 5236 3457 5308 3463
rect 5396 3457 5740 3463
rect 5748 3457 5836 3463
rect 6100 3457 6172 3463
rect 6180 3457 6252 3463
rect 6324 3457 6332 3463
rect 6349 3463 6355 3477
rect 6420 3477 6620 3483
rect 6644 3477 6668 3483
rect 6349 3457 6476 3463
rect 6612 3457 6732 3463
rect 324 3437 364 3443
rect 372 3437 444 3443
rect 452 3437 764 3443
rect 772 3437 972 3443
rect 980 3437 1020 3443
rect 1044 3437 1228 3443
rect 1364 3437 1420 3443
rect 1844 3437 2092 3443
rect 3236 3437 3308 3443
rect 3348 3437 3468 3443
rect 3588 3437 3660 3443
rect 3700 3437 4332 3443
rect 4340 3437 4380 3443
rect 4836 3437 5116 3443
rect 5236 3437 5404 3443
rect 5444 3437 5580 3443
rect 5604 3437 5660 3443
rect 5668 3437 5884 3443
rect 6132 3437 6268 3443
rect 6548 3437 6796 3443
rect 676 3417 828 3423
rect 948 3417 1468 3423
rect 1476 3417 1580 3423
rect 1604 3417 1884 3423
rect 3188 3417 3292 3423
rect 3300 3417 3388 3423
rect 3693 3423 3699 3436
rect 3396 3417 3699 3423
rect 4980 3417 5388 3423
rect 5460 3417 5564 3423
rect 5988 3417 6316 3423
rect 6388 3417 6764 3423
rect 2632 3414 2680 3416
rect 2632 3406 2636 3414
rect 2646 3406 2652 3414
rect 2660 3406 2666 3414
rect 2676 3406 2680 3414
rect 2632 3404 2680 3406
rect 5720 3414 5768 3416
rect 5720 3406 5724 3414
rect 5734 3406 5740 3414
rect 5748 3406 5754 3414
rect 5764 3406 5768 3414
rect 5720 3404 5768 3406
rect 564 3397 604 3403
rect 916 3397 2060 3403
rect 2228 3397 2268 3403
rect 3092 3397 3212 3403
rect 3268 3397 3372 3403
rect 3380 3397 3452 3403
rect 3469 3397 3644 3403
rect 420 3377 540 3383
rect 836 3377 908 3383
rect 932 3377 940 3383
rect 1220 3377 1276 3383
rect 1508 3377 1548 3383
rect 1684 3377 2268 3383
rect 2276 3377 2412 3383
rect 3188 3377 3324 3383
rect 3469 3383 3475 3397
rect 3748 3397 3836 3403
rect 6004 3397 6076 3403
rect 6356 3397 6492 3403
rect 3341 3377 3475 3383
rect 500 3357 684 3363
rect 708 3357 988 3363
rect 1044 3357 1084 3363
rect 1092 3357 1420 3363
rect 1428 3357 1676 3363
rect 2244 3357 2284 3363
rect 3341 3363 3347 3377
rect 3556 3377 3772 3383
rect 3780 3377 3980 3383
rect 3988 3377 4220 3383
rect 4564 3377 4716 3383
rect 4788 3377 6092 3383
rect 6372 3377 6524 3383
rect 3172 3357 3347 3363
rect 3412 3357 3516 3363
rect 3524 3357 3724 3363
rect 3732 3357 3916 3363
rect 3924 3357 3996 3363
rect 4084 3357 4124 3363
rect 4276 3357 4700 3363
rect 4772 3357 4812 3363
rect 4820 3357 5564 3363
rect 5588 3357 5900 3363
rect 5940 3357 6204 3363
rect 6228 3357 6348 3363
rect 6388 3357 6428 3363
rect 6644 3357 6716 3363
rect 404 3337 476 3343
rect 548 3337 716 3343
rect 804 3337 924 3343
rect 1348 3337 1532 3343
rect 1556 3337 1612 3343
rect 2180 3337 2508 3343
rect 2836 3337 3036 3343
rect 3204 3337 3244 3343
rect 3316 3337 3324 3343
rect 3332 3337 3468 3343
rect 3476 3337 3484 3343
rect 3492 3337 3596 3343
rect 3604 3337 3804 3343
rect 3812 3337 3955 3343
rect 84 3317 252 3323
rect 308 3317 332 3323
rect 404 3317 620 3323
rect 1124 3317 1148 3323
rect 1412 3317 1516 3323
rect 1524 3317 1596 3323
rect 1604 3317 1660 3323
rect 2100 3317 2124 3323
rect 2356 3317 2396 3323
rect 3076 3317 3148 3323
rect 3213 3317 3228 3323
rect 84 3297 108 3303
rect 132 3297 172 3303
rect 212 3297 396 3303
rect 596 3297 652 3303
rect 852 3297 1180 3303
rect 1604 3297 1676 3303
rect 1988 3297 2124 3303
rect 2132 3297 2572 3303
rect 3213 3303 3219 3317
rect 3284 3317 3356 3323
rect 3364 3317 3452 3323
rect 3460 3317 3564 3323
rect 3572 3317 3628 3323
rect 3636 3317 3788 3323
rect 3796 3317 3900 3323
rect 3949 3323 3955 3337
rect 3972 3337 4012 3343
rect 4116 3337 4220 3343
rect 4228 3337 4284 3343
rect 4356 3337 4748 3343
rect 5172 3337 5212 3343
rect 5236 3337 5404 3343
rect 5460 3337 5532 3343
rect 6148 3337 6252 3343
rect 6276 3337 6444 3343
rect 6452 3337 6540 3343
rect 6676 3337 6716 3343
rect 3949 3317 4028 3323
rect 4100 3317 4236 3323
rect 4244 3317 4300 3323
rect 4820 3317 4972 3323
rect 5028 3317 5068 3323
rect 5156 3317 5228 3323
rect 5236 3317 5308 3323
rect 5364 3317 5484 3323
rect 5732 3317 5868 3323
rect 6340 3317 6364 3323
rect 6452 3317 6556 3323
rect 6580 3317 6668 3323
rect 3092 3297 3219 3303
rect 3236 3297 3372 3303
rect 3572 3297 3612 3303
rect 3684 3297 3756 3303
rect 3828 3297 3916 3303
rect 4276 3297 4364 3303
rect 4724 3297 4940 3303
rect 5044 3297 5116 3303
rect 5268 3297 5324 3303
rect 5428 3297 5436 3303
rect 5460 3297 5516 3303
rect 5588 3297 6092 3303
rect 6340 3297 6396 3303
rect 6404 3297 6508 3303
rect 6532 3297 6620 3303
rect 6628 3297 6876 3303
rect 244 3277 268 3283
rect 356 3277 700 3283
rect 980 3277 1020 3283
rect 1556 3277 2156 3283
rect 3220 3277 3244 3283
rect 3677 3283 3683 3296
rect 3540 3277 3683 3283
rect 3764 3277 4044 3283
rect 4788 3277 4828 3283
rect 5060 3277 5068 3283
rect 5380 3277 5500 3283
rect 5636 3277 5964 3283
rect 6004 3277 6300 3283
rect 6324 3277 6396 3283
rect 6500 3277 6636 3283
rect 6676 3277 6748 3283
rect 2164 3257 2252 3263
rect 3476 3257 3548 3263
rect 3668 3257 3692 3263
rect 4980 3257 5180 3263
rect 5476 3257 5948 3263
rect 6084 3257 6460 3263
rect 6468 3257 6668 3263
rect 6676 3257 6684 3263
rect 948 3237 1036 3243
rect 1044 3237 1340 3243
rect 2996 3237 3020 3243
rect 3028 3237 3852 3243
rect 4164 3237 5388 3243
rect 5572 3237 5644 3243
rect 5652 3237 5820 3243
rect 6196 3237 6284 3243
rect 6420 3237 6492 3243
rect 948 3217 972 3223
rect 2836 3217 2908 3223
rect 2916 3217 2940 3223
rect 3396 3217 3500 3223
rect 5012 3217 5148 3223
rect 5284 3217 6156 3223
rect 6164 3217 6188 3223
rect 1112 3214 1160 3216
rect 1112 3206 1116 3214
rect 1126 3206 1132 3214
rect 1140 3206 1146 3214
rect 1156 3206 1160 3214
rect 1112 3204 1160 3206
rect 4152 3214 4200 3216
rect 4152 3206 4156 3214
rect 4166 3206 4172 3214
rect 4180 3206 4186 3214
rect 4196 3206 4200 3214
rect 4152 3204 4200 3206
rect 2260 3197 2444 3203
rect 2484 3197 2700 3203
rect 2708 3197 2860 3203
rect 3316 3197 3452 3203
rect 5060 3197 5308 3203
rect 6100 3197 6380 3203
rect 6772 3197 6812 3203
rect 756 3177 1452 3183
rect 1572 3177 1900 3183
rect 1908 3177 2204 3183
rect 2964 3177 3372 3183
rect 3380 3177 3532 3183
rect 3700 3177 3756 3183
rect 4404 3177 4796 3183
rect 4813 3177 4860 3183
rect 388 3157 460 3163
rect 468 3157 668 3163
rect 685 3157 1692 3163
rect 685 3143 691 3157
rect 1700 3157 2108 3163
rect 2980 3157 3004 3163
rect 3156 3157 3212 3163
rect 3348 3157 3468 3163
rect 4813 3163 4819 3177
rect 4996 3177 5532 3183
rect 5556 3177 6332 3183
rect 6436 3177 6620 3183
rect 4532 3157 4819 3163
rect 4836 3157 4956 3163
rect 4964 3157 5564 3163
rect 5684 3157 6236 3163
rect 6388 3157 6444 3163
rect 612 3137 691 3143
rect 1380 3137 2300 3143
rect 2532 3137 2860 3143
rect 2868 3137 2956 3143
rect 2996 3137 3116 3143
rect 3188 3137 3404 3143
rect 4749 3137 4908 3143
rect 4749 3124 4755 3137
rect 4916 3137 5036 3143
rect 5060 3137 5084 3143
rect 5188 3137 5276 3143
rect 5332 3137 5420 3143
rect 5956 3137 5980 3143
rect 5988 3137 6012 3143
rect 6564 3137 6604 3143
rect 340 3117 412 3123
rect 420 3117 508 3123
rect 916 3117 1004 3123
rect 1476 3117 1532 3123
rect 2804 3117 3004 3123
rect 3140 3117 3164 3123
rect 3284 3117 3308 3123
rect 3316 3117 3436 3123
rect 3588 3117 3628 3123
rect 4660 3117 4748 3123
rect 4804 3117 4844 3123
rect 4948 3117 5004 3123
rect 5204 3117 5340 3123
rect 5428 3117 5500 3123
rect 5508 3117 5580 3123
rect 5828 3117 6268 3123
rect 6452 3117 6524 3123
rect 6532 3117 6604 3123
rect 6612 3117 6860 3123
rect 292 3097 364 3103
rect 372 3097 876 3103
rect 1028 3097 1404 3103
rect 1508 3097 1612 3103
rect 1668 3097 2092 3103
rect 2436 3097 2668 3103
rect 3012 3097 3036 3103
rect 3277 3103 3283 3116
rect 3076 3097 3283 3103
rect 3492 3097 3612 3103
rect 3956 3097 4108 3103
rect 4692 3097 4780 3103
rect 4788 3097 5132 3103
rect 5140 3097 5164 3103
rect 5172 3097 5564 3103
rect 5588 3097 5980 3103
rect 5988 3097 5996 3103
rect 6020 3097 6108 3103
rect 6244 3097 6332 3103
rect 6356 3097 6428 3103
rect 6644 3097 6732 3103
rect 148 3077 428 3083
rect 564 3077 604 3083
rect 612 3077 956 3083
rect 1108 3077 1244 3083
rect 1556 3077 1628 3083
rect 1892 3077 2060 3083
rect 2180 3077 2268 3083
rect 2372 3077 2572 3083
rect 2580 3077 2764 3083
rect 2772 3077 2892 3083
rect 2900 3077 3436 3083
rect 4084 3077 4204 3083
rect 4452 3077 4700 3083
rect 4724 3077 4812 3083
rect 4964 3077 5020 3083
rect 5396 3077 5420 3083
rect 5556 3077 5628 3083
rect 5700 3077 5980 3083
rect 6004 3077 6028 3083
rect 6068 3077 6124 3083
rect 6164 3077 6412 3083
rect 6516 3077 6652 3083
rect 564 3057 620 3063
rect 868 3057 1132 3063
rect 1364 3057 1628 3063
rect 1716 3057 1772 3063
rect 1860 3057 1868 3063
rect 1892 3057 2076 3063
rect 2420 3057 2460 3063
rect 2916 3057 3244 3063
rect 3252 3057 3420 3063
rect 3460 3057 3532 3063
rect 3588 3057 3884 3063
rect 4804 3057 4860 3063
rect 4884 3057 4972 3063
rect 5300 3057 5436 3063
rect 5444 3057 5516 3063
rect 6020 3057 6076 3063
rect 6404 3057 6412 3063
rect 6548 3057 6668 3063
rect 1780 3037 2044 3043
rect 2276 3037 2428 3043
rect 3524 3037 3548 3043
rect 4148 3037 4396 3043
rect 5716 3037 5884 3043
rect 5988 3037 6460 3043
rect 244 3017 316 3023
rect 1284 3017 1340 3023
rect 1812 3017 2220 3023
rect 2228 3017 2476 3023
rect 2708 3017 2748 3023
rect 3092 3017 3356 3023
rect 3444 3017 3628 3023
rect 3700 3017 4412 3023
rect 4788 3017 5388 3023
rect 5396 3017 5692 3023
rect 5972 3017 6067 3023
rect 2632 3014 2680 3016
rect 2632 3006 2636 3014
rect 2646 3006 2652 3014
rect 2660 3006 2666 3014
rect 2676 3006 2680 3014
rect 2632 3004 2680 3006
rect 5720 3014 5768 3016
rect 5720 3006 5724 3014
rect 5734 3006 5740 3014
rect 5748 3006 5754 3014
rect 5764 3006 5768 3014
rect 5720 3004 5768 3006
rect 1636 2997 1996 3003
rect 2004 2997 2172 3003
rect 4276 2997 4316 3003
rect 4820 2997 4844 3003
rect 5844 2997 6028 3003
rect 6061 3003 6067 3017
rect 6084 3017 6252 3023
rect 6676 3017 6732 3023
rect 6740 3017 6764 3023
rect 6772 3017 6812 3023
rect 6061 2997 6124 3003
rect 6132 2997 6476 3003
rect 6484 2997 6556 3003
rect 1124 2977 1468 2983
rect 2484 2977 2940 2983
rect 3252 2977 3276 2983
rect 3316 2977 3708 2983
rect 4532 2977 4636 2983
rect 4644 2977 5116 2983
rect 5236 2977 5580 2983
rect 5604 2977 6044 2983
rect 6356 2977 6540 2983
rect 164 2957 284 2963
rect 1428 2957 1708 2963
rect 1805 2957 2188 2963
rect 1805 2944 1811 2957
rect 2205 2957 2508 2963
rect 212 2937 268 2943
rect 276 2937 444 2943
rect 452 2937 540 2943
rect 548 2937 604 2943
rect 756 2937 956 2943
rect 980 2937 1084 2943
rect 1316 2937 1532 2943
rect 2205 2943 2211 2957
rect 2980 2957 3068 2963
rect 3076 2957 3132 2963
rect 3140 2957 3180 2963
rect 3188 2957 3308 2963
rect 3316 2957 3452 2963
rect 3572 2957 3644 2963
rect 3860 2957 4236 2963
rect 4244 2957 4364 2963
rect 4372 2957 4476 2963
rect 4564 2957 4652 2963
rect 4740 2957 4876 2963
rect 4964 2957 5068 2963
rect 5076 2957 5212 2963
rect 5220 2957 5260 2963
rect 5540 2957 6204 2963
rect 6260 2957 6316 2963
rect 6340 2957 6364 2963
rect 6372 2957 6508 2963
rect 2196 2937 2211 2943
rect 2420 2937 2444 2943
rect 2724 2937 2796 2943
rect 3156 2937 3228 2943
rect 3284 2937 3324 2943
rect 3364 2937 3452 2943
rect 3604 2937 3884 2943
rect 4340 2937 4540 2943
rect 4660 2937 4684 2943
rect 4804 2937 4828 2943
rect 4868 2937 4972 2943
rect 5172 2937 5196 2943
rect 5316 2937 5340 2943
rect 5700 2937 5788 2943
rect 5812 2937 5932 2943
rect 5940 2937 6076 2943
rect 6116 2937 6220 2943
rect 6228 2937 6396 2943
rect 6404 2937 6460 2943
rect 6468 2937 6572 2943
rect 36 2917 140 2923
rect 148 2917 300 2923
rect 308 2917 348 2923
rect 436 2917 476 2923
rect 612 2917 1020 2923
rect 1060 2917 1612 2923
rect 3220 2917 3756 2923
rect 3764 2917 3788 2923
rect 4772 2917 4828 2923
rect 4868 2917 4988 2923
rect 5188 2917 5228 2923
rect 5236 2917 5324 2923
rect 5460 2917 6028 2923
rect 6036 2917 6172 2923
rect 6180 2917 6236 2923
rect -19 2897 12 2903
rect 68 2897 380 2903
rect 948 2897 1004 2903
rect 1076 2897 1516 2903
rect 1524 2897 1804 2903
rect 1972 2897 2044 2903
rect 2196 2897 2380 2903
rect 2532 2897 2892 2903
rect 3220 2897 3244 2903
rect 3300 2897 3324 2903
rect 3380 2897 3468 2903
rect 4708 2897 4716 2903
rect 4756 2897 5836 2903
rect 5844 2897 6156 2903
rect 6212 2897 6252 2903
rect 6708 2897 6764 2903
rect 116 2877 172 2883
rect 340 2877 428 2883
rect 532 2877 1052 2883
rect 1508 2877 1564 2883
rect 3236 2877 3436 2883
rect 3524 2877 4060 2883
rect 4724 2877 5116 2883
rect 5124 2877 5628 2883
rect 5876 2877 5980 2883
rect 6157 2883 6163 2896
rect 6157 2877 6412 2883
rect 6420 2877 6524 2883
rect 788 2857 1196 2863
rect 1204 2857 1340 2863
rect 1348 2857 1532 2863
rect 2436 2857 3612 2863
rect 3620 2857 3724 2863
rect 5652 2857 6028 2863
rect 6148 2857 6252 2863
rect 884 2837 1324 2843
rect 1620 2837 1788 2843
rect 1796 2837 2012 2843
rect 2020 2837 2156 2843
rect 2164 2837 2236 2843
rect 3268 2837 3468 2843
rect 3492 2837 3756 2843
rect 5028 2837 5564 2843
rect 5972 2837 5996 2843
rect 6004 2837 6092 2843
rect 6292 2837 6348 2843
rect 2052 2817 2780 2823
rect 3092 2817 3404 2823
rect 3428 2817 3980 2823
rect 5108 2817 5324 2823
rect 5332 2817 5996 2823
rect 6516 2817 6588 2823
rect 1112 2814 1160 2816
rect 1112 2806 1116 2814
rect 1126 2806 1132 2814
rect 1140 2806 1146 2814
rect 1156 2806 1160 2814
rect 1112 2804 1160 2806
rect 4152 2814 4200 2816
rect 4152 2806 4156 2814
rect 4166 2806 4172 2814
rect 4180 2806 4186 2814
rect 4196 2806 4200 2814
rect 4152 2804 4200 2806
rect 1556 2797 1708 2803
rect 1860 2797 2428 2803
rect 2836 2797 3004 2803
rect 3156 2797 3468 2803
rect 4820 2797 5068 2803
rect 5076 2797 5292 2803
rect 5428 2797 5612 2803
rect 5876 2797 5916 2803
rect 5924 2797 6588 2803
rect 180 2777 332 2783
rect 484 2777 684 2783
rect 2388 2777 2476 2783
rect 2756 2777 3100 2783
rect 3444 2777 3580 2783
rect 3636 2777 3788 2783
rect 3796 2777 4028 2783
rect 4036 2777 4092 2783
rect 4100 2777 4556 2783
rect 5348 2777 5484 2783
rect 5492 2777 5580 2783
rect 5732 2777 6284 2783
rect 1572 2757 3148 2763
rect 3204 2757 3340 2763
rect 3348 2757 3420 2763
rect 3460 2757 3660 2763
rect 3668 2757 3820 2763
rect 5844 2757 6172 2763
rect 6308 2757 6572 2763
rect 6580 2757 6668 2763
rect 1012 2737 2332 2743
rect 2772 2737 2972 2743
rect 3412 2737 3628 2743
rect 4068 2737 4108 2743
rect 5204 2737 5468 2743
rect 6052 2737 6348 2743
rect 6356 2737 6380 2743
rect 6468 2737 6604 2743
rect 6644 2737 6764 2743
rect 596 2717 652 2723
rect 1092 2717 1372 2723
rect 1380 2717 1740 2723
rect 2756 2717 2812 2723
rect 3412 2717 3596 2723
rect 3620 2717 3772 2723
rect 5284 2717 5388 2723
rect 5604 2717 6236 2723
rect 6244 2717 6268 2723
rect 6404 2717 6412 2723
rect 6420 2717 6460 2723
rect 6548 2717 6636 2723
rect 388 2697 876 2703
rect 1124 2697 1900 2703
rect 2196 2697 2316 2703
rect 2596 2697 2604 2703
rect 2612 2697 2716 2703
rect 2724 2697 2972 2703
rect 3108 2697 3404 2703
rect 3428 2697 3756 2703
rect 3796 2697 3852 2703
rect 3860 2697 3868 2703
rect 4516 2697 4684 2703
rect 5156 2697 5244 2703
rect 5396 2697 5452 2703
rect 5636 2697 5804 2703
rect 5940 2697 6076 2703
rect 6084 2697 6364 2703
rect 6372 2697 6444 2703
rect 6500 2697 6572 2703
rect 6612 2697 6668 2703
rect 68 2677 140 2683
rect 564 2677 572 2683
rect 580 2677 604 2683
rect 612 2677 1116 2683
rect 1572 2677 1708 2683
rect 2692 2677 2732 2683
rect 3268 2677 3356 2683
rect 3444 2677 3836 2683
rect 4404 2677 4636 2683
rect 4900 2677 5068 2683
rect 5300 2677 5340 2683
rect 5636 2677 5852 2683
rect 6004 2677 6044 2683
rect 6052 2677 6188 2683
rect 6196 2677 6348 2683
rect 6356 2677 6524 2683
rect 6532 2677 6636 2683
rect 6644 2677 6652 2683
rect 180 2657 364 2663
rect 516 2657 1084 2663
rect 1540 2657 1868 2663
rect 1876 2657 2060 2663
rect 2500 2657 2700 2663
rect 3076 2657 3436 2663
rect 3492 2657 3532 2663
rect 3540 2657 3548 2663
rect 3572 2657 3708 2663
rect 3764 2657 4108 2663
rect 4260 2657 4556 2663
rect 4788 2657 4892 2663
rect 5012 2657 5196 2663
rect 5204 2657 5420 2663
rect 5428 2657 5596 2663
rect 5604 2657 5692 2663
rect 5853 2663 5859 2676
rect 5853 2657 6124 2663
rect 6228 2657 6300 2663
rect 324 2637 668 2643
rect 676 2637 844 2643
rect 852 2637 1180 2643
rect 1188 2637 1292 2643
rect 2884 2637 3948 2643
rect 5508 2637 5708 2643
rect 5716 2637 5788 2643
rect 5796 2637 6012 2643
rect 6276 2637 6428 2643
rect 212 2617 268 2623
rect 1076 2617 2204 2623
rect 2212 2617 2252 2623
rect 2308 2617 2588 2623
rect 2852 2617 3132 2623
rect 3140 2617 3500 2623
rect 3508 2617 3676 2623
rect 3684 2617 4060 2623
rect 5220 2617 5484 2623
rect 5508 2617 5548 2623
rect 2632 2614 2680 2616
rect 2632 2606 2636 2614
rect 2646 2606 2652 2614
rect 2660 2606 2666 2614
rect 2676 2606 2680 2614
rect 2632 2604 2680 2606
rect 5720 2614 5768 2616
rect 5720 2606 5724 2614
rect 5734 2606 5740 2614
rect 5748 2606 5754 2614
rect 5764 2606 5768 2614
rect 5720 2604 5768 2606
rect 132 2597 540 2603
rect 660 2597 700 2603
rect 900 2597 988 2603
rect 1044 2597 1228 2603
rect 1252 2597 1308 2603
rect 1316 2597 1420 2603
rect 1428 2597 1836 2603
rect 2420 2597 2460 2603
rect 2980 2597 3020 2603
rect 3652 2597 3692 2603
rect 3700 2597 4028 2603
rect 4436 2597 4508 2603
rect 4516 2597 4812 2603
rect 4820 2597 5276 2603
rect 5348 2597 5660 2603
rect 5812 2597 5964 2603
rect 6420 2597 6668 2603
rect 980 2577 1868 2583
rect 2100 2577 2172 2583
rect 2180 2577 2236 2583
rect 2292 2577 2748 2583
rect 2756 2577 3212 2583
rect 3284 2577 3404 2583
rect 3508 2577 3692 2583
rect 4116 2577 4460 2583
rect 4628 2577 4700 2583
rect 5524 2577 5532 2583
rect 5892 2577 6028 2583
rect 6132 2577 6220 2583
rect 6436 2577 6604 2583
rect 6612 2577 6876 2583
rect 116 2557 140 2563
rect 1060 2557 1068 2563
rect 1204 2557 1564 2563
rect 1572 2557 1580 2563
rect 2420 2557 2908 2563
rect 2948 2557 3292 2563
rect 3476 2557 3724 2563
rect 3812 2557 3868 2563
rect 4020 2557 4108 2563
rect 4372 2557 4396 2563
rect 4404 2557 4716 2563
rect 5060 2557 5100 2563
rect 5108 2557 5436 2563
rect 5700 2557 5884 2563
rect 6356 2557 6556 2563
rect 6596 2557 6620 2563
rect -19 2537 60 2543
rect 356 2537 508 2543
rect 836 2537 1084 2543
rect 1412 2537 1692 2543
rect 1844 2537 1980 2543
rect 2276 2537 2444 2543
rect 3268 2537 3308 2543
rect 3348 2537 3372 2543
rect 3396 2537 3804 2543
rect 3988 2537 4044 2543
rect 4148 2537 4364 2543
rect 4820 2537 4844 2543
rect 5076 2537 5244 2543
rect 5556 2537 5820 2543
rect 5828 2537 5932 2543
rect 6196 2537 6284 2543
rect 6308 2537 6412 2543
rect 6548 2537 6588 2543
rect 452 2517 588 2523
rect 788 2517 1676 2523
rect 1684 2517 1804 2523
rect 2100 2517 2188 2523
rect 2340 2517 3100 2523
rect 3156 2517 3164 2523
rect 3268 2517 3292 2523
rect 3684 2517 3852 2523
rect 3924 2517 4140 2523
rect 4580 2517 4860 2523
rect 4868 2517 4988 2523
rect 5492 2517 5580 2523
rect 5764 2517 5884 2523
rect 5956 2517 6124 2523
rect 6148 2517 6332 2523
rect 6420 2517 6444 2523
rect 6580 2517 6652 2523
rect 6692 2517 6748 2523
rect -19 2497 12 2503
rect 52 2497 508 2503
rect 516 2497 572 2503
rect 1572 2497 2012 2503
rect 2900 2497 2908 2503
rect 3101 2497 3827 2503
rect 3101 2483 3107 2497
rect 2909 2477 3107 2483
rect 2909 2464 2915 2477
rect 3124 2477 3180 2483
rect 3188 2477 3212 2483
rect 3252 2477 3276 2483
rect 3380 2477 3420 2483
rect 3524 2477 3548 2483
rect 3821 2483 3827 2497
rect 3844 2497 3884 2503
rect 3892 2497 3916 2503
rect 4164 2497 4268 2503
rect 4292 2497 4604 2503
rect 4788 2497 5148 2503
rect 6324 2497 6524 2503
rect 6580 2497 6636 2503
rect 6676 2497 6684 2503
rect 3821 2477 4908 2483
rect 4916 2477 5004 2483
rect 6452 2477 6476 2483
rect 772 2457 2908 2463
rect 2932 2457 3276 2463
rect 3284 2457 3356 2463
rect 3364 2457 3772 2463
rect 3780 2457 3788 2463
rect 3796 2457 3852 2463
rect 3908 2457 4236 2463
rect 2612 2437 2684 2443
rect 2692 2437 3372 2443
rect 3380 2437 3660 2443
rect 3668 2437 3884 2443
rect 3892 2437 4588 2443
rect 6740 2437 6796 2443
rect 1380 2417 1676 2423
rect 2852 2417 2860 2423
rect 3188 2417 3228 2423
rect 3412 2417 3612 2423
rect 3844 2417 3932 2423
rect 1112 2414 1160 2416
rect 1112 2406 1116 2414
rect 1126 2406 1132 2414
rect 1140 2406 1146 2414
rect 1156 2406 1160 2414
rect 1112 2404 1160 2406
rect 4152 2414 4200 2416
rect 4152 2406 4156 2414
rect 4166 2406 4172 2414
rect 4180 2406 4186 2414
rect 4196 2406 4200 2414
rect 4152 2404 4200 2406
rect 1540 2397 1564 2403
rect 1812 2397 1852 2403
rect 1860 2397 2300 2403
rect 2308 2397 2716 2403
rect 2724 2397 3372 2403
rect 3556 2397 4131 2403
rect 1236 2377 1404 2383
rect 1684 2377 3548 2383
rect 3796 2377 3852 2383
rect 3860 2377 4012 2383
rect 4125 2383 4131 2397
rect 6516 2397 6540 2403
rect 4125 2377 4284 2383
rect 6116 2377 6300 2383
rect 2180 2357 2396 2363
rect 3316 2357 3692 2363
rect 3764 2357 3804 2363
rect 6612 2357 6828 2363
rect 1684 2337 2428 2343
rect 3284 2337 3612 2343
rect 3764 2337 3820 2343
rect 4244 2337 4828 2343
rect 4836 2337 4892 2343
rect 660 2317 780 2323
rect 1012 2317 1596 2323
rect 2372 2317 2380 2323
rect 2388 2317 2940 2323
rect 3316 2317 3628 2323
rect 3940 2317 4028 2323
rect 4116 2317 4268 2323
rect 4276 2317 4572 2323
rect 5396 2317 5564 2323
rect 5588 2317 5660 2323
rect 5668 2317 5724 2323
rect 6244 2317 6460 2323
rect 196 2297 588 2303
rect 772 2297 796 2303
rect 1124 2297 1180 2303
rect 1188 2297 1484 2303
rect 2084 2297 2332 2303
rect 2708 2297 2876 2303
rect 2884 2297 2908 2303
rect 3012 2297 3068 2303
rect 3076 2297 3132 2303
rect 3172 2297 3644 2303
rect 3732 2297 3852 2303
rect 3860 2297 3900 2303
rect 5508 2297 5852 2303
rect 6084 2297 6204 2303
rect 6212 2297 6332 2303
rect 6756 2297 6860 2303
rect 436 2277 572 2283
rect 708 2277 748 2283
rect 756 2277 1276 2283
rect 1284 2277 1356 2283
rect 1604 2277 1756 2283
rect 2292 2277 2332 2283
rect 2340 2277 3196 2283
rect 3508 2277 3564 2283
rect 3668 2277 3708 2283
rect 3844 2277 3852 2283
rect 4004 2277 4316 2283
rect 4676 2277 4924 2283
rect 5156 2277 5292 2283
rect 5412 2277 5564 2283
rect 5604 2277 5676 2283
rect 196 2257 236 2263
rect 628 2257 668 2263
rect 1204 2257 1308 2263
rect 1348 2257 1580 2263
rect 1588 2257 1740 2263
rect 1892 2257 1932 2263
rect 2052 2257 2412 2263
rect 2948 2257 3132 2263
rect 3140 2257 3244 2263
rect 4036 2257 4236 2263
rect 4260 2257 4364 2263
rect 4868 2257 5004 2263
rect 5348 2257 5420 2263
rect 5428 2257 5468 2263
rect 5476 2257 5548 2263
rect 5556 2257 5612 2263
rect 532 2237 700 2243
rect 1044 2237 1564 2243
rect 1748 2237 1804 2243
rect 2356 2237 2428 2243
rect 2436 2237 2732 2243
rect 3028 2237 3084 2243
rect 3444 2237 3484 2243
rect 3764 2237 3804 2243
rect 5940 2237 6268 2243
rect 6276 2237 6284 2243
rect 6292 2237 6460 2243
rect 6468 2237 6684 2243
rect 1364 2217 1388 2223
rect 1588 2217 1884 2223
rect 1892 2217 2348 2223
rect 2740 2217 3212 2223
rect 3220 2217 3676 2223
rect 3732 2217 3948 2223
rect 5076 2217 5116 2223
rect 5876 2217 5964 2223
rect 6436 2217 6492 2223
rect 2632 2214 2680 2216
rect 2632 2206 2636 2214
rect 2646 2206 2652 2214
rect 2660 2206 2666 2214
rect 2676 2206 2680 2214
rect 2632 2204 2680 2206
rect 5720 2214 5768 2216
rect 5720 2206 5724 2214
rect 5734 2206 5740 2214
rect 5748 2206 5754 2214
rect 5764 2206 5768 2214
rect 5720 2204 5768 2206
rect 740 2197 812 2203
rect 1348 2197 1388 2203
rect 2372 2197 2396 2203
rect 3188 2197 3756 2203
rect 3780 2197 4012 2203
rect 4052 2197 4108 2203
rect 36 2177 268 2183
rect 276 2177 396 2183
rect 404 2177 780 2183
rect 788 2177 876 2183
rect 1556 2177 1580 2183
rect 2324 2177 2364 2183
rect 2516 2177 3020 2183
rect 3108 2177 3308 2183
rect 3757 2183 3763 2196
rect 3757 2177 3900 2183
rect 4708 2177 5036 2183
rect 5044 2177 5180 2183
rect 5284 2177 5804 2183
rect 148 2157 492 2163
rect 500 2157 588 2163
rect 596 2157 963 2163
rect 957 2144 963 2157
rect 1076 2157 1084 2163
rect 1092 2157 1356 2163
rect 1364 2157 1500 2163
rect 1572 2157 1708 2163
rect 1844 2157 2156 2163
rect 2596 2157 2604 2163
rect 2820 2157 2892 2163
rect 2948 2157 2988 2163
rect 3060 2157 3340 2163
rect 3380 2157 3420 2163
rect 4244 2157 4508 2163
rect 4516 2157 4668 2163
rect 4708 2157 5372 2163
rect 5492 2157 5644 2163
rect 6564 2157 6620 2163
rect 100 2137 236 2143
rect 964 2137 1244 2143
rect 1844 2137 1900 2143
rect 2020 2137 2268 2143
rect 2324 2137 2380 2143
rect 2964 2137 3036 2143
rect 3220 2137 3452 2143
rect 3604 2137 3756 2143
rect 3892 2137 3916 2143
rect 3924 2137 3964 2143
rect 4212 2137 4764 2143
rect 5012 2137 5436 2143
rect 5460 2137 5484 2143
rect 5524 2137 5548 2143
rect 5668 2137 5772 2143
rect 5780 2137 5900 2143
rect 6004 2137 6076 2143
rect 6116 2137 6316 2143
rect 6468 2137 6652 2143
rect 1396 2117 2268 2123
rect 2317 2123 2323 2136
rect 2276 2117 2323 2123
rect 2500 2117 2556 2123
rect 2564 2117 2732 2123
rect 2996 2117 3100 2123
rect 3108 2117 3276 2123
rect 3332 2117 3372 2123
rect 3428 2117 3916 2123
rect 3972 2117 4332 2123
rect 4340 2117 4428 2123
rect 4436 2117 4508 2123
rect 5460 2117 5692 2123
rect 5796 2117 5980 2123
rect 5988 2117 5996 2123
rect 6004 2117 6124 2123
rect 6564 2117 6588 2123
rect 6596 2117 6716 2123
rect -19 2097 12 2103
rect 2388 2097 2572 2103
rect 2580 2097 2780 2103
rect 3044 2097 3068 2103
rect 3140 2097 3468 2103
rect 3476 2097 3500 2103
rect 4804 2097 4892 2103
rect 5284 2097 5564 2103
rect 5684 2097 5788 2103
rect 5940 2097 6028 2103
rect 2548 2077 3356 2083
rect 4020 2077 4268 2083
rect 4372 2077 4396 2083
rect 5300 2077 5516 2083
rect 5556 2077 6012 2083
rect 3012 2057 3036 2063
rect 3348 2057 3964 2063
rect 5268 2057 5340 2063
rect 6804 2057 6860 2063
rect 116 2037 428 2043
rect 436 2037 684 2043
rect 3396 2037 4028 2043
rect 100 2017 140 2023
rect 4404 2017 4940 2023
rect 5044 2017 5068 2023
rect 1112 2014 1160 2016
rect 1112 2006 1116 2014
rect 1126 2006 1132 2014
rect 1140 2006 1146 2014
rect 1156 2006 1160 2014
rect 1112 2004 1160 2006
rect 4152 2014 4200 2016
rect 4152 2006 4156 2014
rect 4166 2006 4172 2014
rect 4180 2006 4186 2014
rect 4196 2006 4200 2014
rect 4152 2004 4200 2006
rect 2532 1997 2556 2003
rect 2564 1997 2700 2003
rect 2708 1997 2780 2003
rect 2820 1997 3228 2003
rect 6804 1997 6828 2003
rect 644 1977 2092 1983
rect 3252 1977 3580 1983
rect 3764 1977 3804 1983
rect 3828 1977 4172 1983
rect 4276 1977 4284 1983
rect 4468 1977 4668 1983
rect 4948 1977 5100 1983
rect 6196 1977 6348 1983
rect 6532 1977 6828 1983
rect 500 1957 1052 1963
rect 1812 1957 2268 1963
rect 2276 1957 3708 1963
rect 3716 1957 4652 1963
rect 4676 1957 5180 1963
rect 5188 1957 5228 1963
rect 5828 1957 6364 1963
rect 6484 1957 6540 1963
rect 580 1937 796 1943
rect 3732 1937 3756 1943
rect 3908 1937 3980 1943
rect 3988 1937 4044 1943
rect 4372 1937 4812 1943
rect 4820 1937 4956 1943
rect 5604 1937 5788 1943
rect 6228 1937 6316 1943
rect 6324 1937 6396 1943
rect 6429 1937 6508 1943
rect 100 1917 508 1923
rect 724 1917 764 1923
rect 836 1917 1404 1923
rect 2116 1917 2380 1923
rect 3316 1917 3404 1923
rect 3476 1917 3756 1923
rect 3764 1917 3820 1923
rect 3940 1917 4012 1923
rect 4372 1917 4556 1923
rect 4660 1917 4844 1923
rect 4852 1917 4876 1923
rect 5764 1917 5980 1923
rect 6212 1917 6284 1923
rect 6429 1923 6435 1937
rect 6580 1937 6716 1943
rect 6772 1937 6780 1943
rect 6308 1917 6435 1923
rect 6452 1917 6492 1923
rect 6500 1917 6764 1923
rect -19 1897 12 1903
rect 68 1897 76 1903
rect 84 1897 636 1903
rect 708 1897 732 1903
rect 1508 1897 1644 1903
rect 2148 1897 2172 1903
rect 2180 1897 2252 1903
rect 3012 1897 3100 1903
rect 3204 1897 3404 1903
rect 3460 1897 3836 1903
rect 4036 1897 4044 1903
rect 4180 1897 4620 1903
rect 4660 1897 4684 1903
rect 4772 1897 4876 1903
rect 5460 1897 5612 1903
rect 5652 1897 5772 1903
rect 5892 1897 6092 1903
rect 6244 1897 6652 1903
rect 6724 1897 6876 1903
rect 164 1877 172 1883
rect 564 1877 604 1883
rect 660 1877 780 1883
rect 788 1877 844 1883
rect 852 1877 1084 1883
rect 1092 1877 1196 1883
rect 1428 1877 2204 1883
rect 2212 1877 2300 1883
rect 2612 1877 2892 1883
rect 3396 1877 3500 1883
rect 3620 1877 3692 1883
rect 3700 1877 3724 1883
rect 4084 1877 4204 1883
rect 4212 1877 4364 1883
rect 4468 1877 4652 1883
rect 4692 1877 5164 1883
rect 5204 1877 5452 1883
rect 5700 1877 5964 1883
rect 5972 1877 6172 1883
rect 6260 1877 6300 1883
rect 6324 1877 6476 1883
rect 6484 1877 6764 1883
rect 100 1857 300 1863
rect 340 1857 476 1863
rect 628 1857 700 1863
rect 932 1857 1228 1863
rect 1716 1857 1996 1863
rect 2036 1857 2124 1863
rect 2244 1857 2492 1863
rect 3060 1857 3084 1863
rect 3236 1857 3564 1863
rect 3972 1857 4012 1863
rect 4340 1857 4444 1863
rect 4452 1857 4700 1863
rect 5172 1857 5244 1863
rect 5252 1857 5260 1863
rect 5588 1857 5852 1863
rect 5860 1857 5900 1863
rect 5988 1857 6124 1863
rect 6132 1857 6604 1863
rect 6644 1857 6668 1863
rect 6676 1857 6700 1863
rect 1748 1837 1836 1843
rect 1997 1843 2003 1856
rect 1844 1837 1987 1843
rect 1997 1837 2460 1843
rect 180 1817 588 1823
rect 1700 1817 1884 1823
rect 1981 1823 1987 1837
rect 3700 1837 3836 1843
rect 4116 1837 4124 1843
rect 4132 1837 4748 1843
rect 5188 1837 5308 1843
rect 5332 1837 5372 1843
rect 5572 1837 5628 1843
rect 5684 1837 5820 1843
rect 5924 1837 5980 1843
rect 6164 1837 6188 1843
rect 6516 1837 6780 1843
rect 1981 1817 2060 1823
rect 3556 1817 3676 1823
rect 3684 1817 4076 1823
rect 4484 1817 4524 1823
rect 4596 1817 4892 1823
rect 5220 1817 5308 1823
rect 5316 1817 5548 1823
rect 6132 1817 6220 1823
rect 6372 1817 6604 1823
rect 6628 1817 6652 1823
rect 6740 1817 6828 1823
rect 2632 1814 2680 1816
rect 2632 1806 2636 1814
rect 2646 1806 2652 1814
rect 2660 1806 2666 1814
rect 2676 1806 2680 1814
rect 2632 1804 2680 1806
rect 5720 1814 5768 1816
rect 5720 1806 5724 1814
rect 5734 1806 5740 1814
rect 5748 1806 5754 1814
rect 5764 1806 5768 1814
rect 5720 1804 5768 1806
rect 1556 1797 2172 1803
rect 3364 1797 3404 1803
rect 3412 1797 3660 1803
rect 3668 1797 3772 1803
rect 3780 1797 4092 1803
rect 5140 1797 5324 1803
rect 6420 1797 6556 1803
rect 6564 1797 6588 1803
rect 6756 1797 6844 1803
rect 532 1777 796 1783
rect 1188 1777 2588 1783
rect 2596 1777 2700 1783
rect 2717 1777 3532 1783
rect 180 1757 332 1763
rect 340 1757 380 1763
rect 644 1757 700 1763
rect 1348 1757 1404 1763
rect 1508 1757 1580 1763
rect 1620 1757 1692 1763
rect 1700 1757 1980 1763
rect 2100 1757 2652 1763
rect 2717 1763 2723 1777
rect 3540 1777 4124 1783
rect 4372 1777 4588 1783
rect 5076 1777 5212 1783
rect 5220 1777 5404 1783
rect 5780 1777 5868 1783
rect 6468 1777 6636 1783
rect 6676 1777 6716 1783
rect 2660 1757 2723 1763
rect 3156 1757 3372 1763
rect 4068 1757 4508 1763
rect 4916 1757 5420 1763
rect 5556 1757 5788 1763
rect 5796 1757 5980 1763
rect 6148 1757 6172 1763
rect 6244 1757 6300 1763
rect 6596 1757 6796 1763
rect 68 1737 140 1743
rect 308 1737 588 1743
rect 596 1737 652 1743
rect 692 1737 892 1743
rect 1380 1737 1587 1743
rect 1581 1724 1587 1737
rect 1668 1737 1948 1743
rect 1956 1737 2028 1743
rect 2036 1737 2044 1743
rect 2100 1737 2140 1743
rect 2148 1737 2556 1743
rect 2564 1737 2636 1743
rect 2804 1737 2844 1743
rect 3140 1737 3180 1743
rect 3188 1737 3468 1743
rect 3876 1737 3948 1743
rect 4596 1737 5548 1743
rect 6084 1737 6524 1743
rect 6532 1737 6716 1743
rect 6756 1737 6812 1743
rect 260 1717 796 1723
rect 1204 1717 1228 1723
rect 1236 1717 1468 1723
rect 1476 1717 1564 1723
rect 1588 1717 1676 1723
rect 1860 1717 1884 1723
rect 2516 1717 2748 1723
rect 3172 1717 3212 1723
rect 4484 1717 4572 1723
rect 4644 1717 4732 1723
rect 4740 1717 4828 1723
rect 5012 1717 5084 1723
rect 5604 1717 5820 1723
rect 5956 1717 6156 1723
rect 6276 1717 6396 1723
rect 6436 1717 6748 1723
rect 532 1697 556 1703
rect 564 1697 620 1703
rect 660 1697 748 1703
rect 756 1697 1084 1703
rect 1092 1697 1180 1703
rect 1252 1697 1484 1703
rect 1540 1697 1788 1703
rect 1812 1697 1868 1703
rect 1876 1697 1900 1703
rect 2564 1697 3132 1703
rect 3236 1697 3436 1703
rect 3444 1697 3564 1703
rect 5268 1697 5340 1703
rect 5348 1697 5564 1703
rect 5572 1697 5628 1703
rect 5828 1697 5836 1703
rect 5924 1697 6188 1703
rect 6196 1697 6284 1703
rect 6372 1697 6460 1703
rect 340 1677 556 1683
rect 1220 1677 1516 1683
rect 1556 1677 1740 1683
rect 1828 1677 2028 1683
rect 4020 1677 4220 1683
rect 5044 1677 5196 1683
rect 5204 1677 5468 1683
rect 6052 1677 6236 1683
rect 6388 1677 6492 1683
rect 6804 1677 6828 1683
rect 436 1657 1116 1663
rect 1940 1657 4044 1663
rect 4052 1657 5100 1663
rect 5188 1657 5676 1663
rect 5812 1657 6028 1663
rect 6036 1657 6268 1663
rect 1156 1637 1244 1643
rect 1252 1637 1436 1643
rect 1444 1637 1484 1643
rect 1508 1637 1772 1643
rect 1780 1637 1836 1643
rect 1844 1637 2156 1643
rect 2964 1637 3292 1643
rect 4548 1637 4652 1643
rect 4868 1637 5036 1643
rect 5300 1637 5452 1643
rect 5460 1637 5804 1643
rect 5828 1637 5948 1643
rect 6068 1637 6092 1643
rect 6708 1637 6764 1643
rect 100 1617 140 1623
rect 420 1617 540 1623
rect 548 1617 876 1623
rect 2340 1617 2380 1623
rect 4980 1617 5068 1623
rect 5412 1617 5468 1623
rect 5780 1617 5852 1623
rect 6820 1617 6844 1623
rect 1112 1614 1160 1616
rect 1112 1606 1116 1614
rect 1126 1606 1132 1614
rect 1140 1606 1146 1614
rect 1156 1606 1160 1614
rect 1112 1604 1160 1606
rect 4152 1614 4200 1616
rect 4152 1606 4156 1614
rect 4166 1606 4172 1614
rect 4180 1606 4186 1614
rect 4196 1606 4200 1614
rect 4152 1604 4200 1606
rect 1428 1597 1548 1603
rect 1620 1597 1660 1603
rect 4580 1597 4588 1603
rect 4948 1597 5084 1603
rect 5092 1597 5340 1603
rect 5348 1597 5436 1603
rect 5620 1597 5884 1603
rect 6276 1597 6556 1603
rect 292 1577 364 1583
rect 372 1577 1228 1583
rect 1332 1577 1388 1583
rect 4004 1577 4284 1583
rect 5124 1577 5996 1583
rect 6004 1577 6332 1583
rect 6340 1577 6492 1583
rect 452 1557 732 1563
rect 804 1557 1340 1563
rect 1348 1557 1628 1563
rect 1636 1557 1708 1563
rect 1940 1557 1964 1563
rect 4740 1557 4844 1563
rect 5380 1557 5500 1563
rect 5588 1557 5740 1563
rect 5796 1557 6412 1563
rect 6484 1557 6684 1563
rect 685 1537 940 1543
rect 685 1524 691 1537
rect 1284 1537 1596 1543
rect 1604 1537 1948 1543
rect 1956 1537 2060 1543
rect 2100 1537 2172 1543
rect 3124 1537 3452 1543
rect 3460 1537 3564 1543
rect 4372 1537 5452 1543
rect 5860 1537 5948 1543
rect 6148 1537 6220 1543
rect 6468 1537 6540 1543
rect 6564 1537 6700 1543
rect 6708 1537 6828 1543
rect 36 1517 108 1523
rect 116 1517 332 1523
rect 356 1517 412 1523
rect 500 1517 524 1523
rect 596 1517 684 1523
rect 868 1517 1036 1523
rect 1044 1517 1196 1523
rect 1917 1517 2012 1523
rect 1917 1504 1923 1517
rect 2164 1517 2460 1523
rect 3076 1517 3196 1523
rect 3460 1517 3516 1523
rect 5220 1517 5308 1523
rect 5380 1517 5420 1523
rect 5652 1517 5740 1523
rect 5812 1517 5891 1523
rect 148 1497 524 1503
rect 564 1497 636 1503
rect 676 1497 1052 1503
rect 1476 1497 1516 1503
rect 1556 1497 1676 1503
rect 1748 1497 1916 1503
rect 1972 1497 2092 1503
rect 2132 1497 2284 1503
rect 2388 1497 2476 1503
rect 2484 1497 2604 1503
rect 3812 1497 3868 1503
rect 4084 1497 4412 1503
rect 4628 1497 4796 1503
rect 5156 1497 5180 1503
rect 5204 1497 5388 1503
rect 5396 1497 5420 1503
rect 5460 1497 5628 1503
rect 5684 1497 5820 1503
rect 5844 1497 5852 1503
rect 5885 1503 5891 1517
rect 5940 1517 6300 1523
rect 6461 1523 6467 1536
rect 6308 1517 6467 1523
rect 6724 1517 6780 1523
rect 5885 1497 6204 1503
rect 6212 1497 6220 1503
rect 6228 1497 6284 1503
rect 6516 1497 6604 1503
rect 6692 1497 6796 1503
rect 180 1477 188 1483
rect 196 1477 236 1483
rect 244 1477 300 1483
rect 324 1477 348 1483
rect 404 1477 428 1483
rect 916 1477 1212 1483
rect 1396 1477 1500 1483
rect 1588 1477 1852 1483
rect 2036 1477 2140 1483
rect 2436 1477 2492 1483
rect 3044 1477 3052 1483
rect 4516 1477 4668 1483
rect 5092 1477 5276 1483
rect 5284 1477 5564 1483
rect 5700 1477 5804 1483
rect 5924 1477 6060 1483
rect 324 1457 412 1463
rect 420 1457 620 1463
rect 756 1457 924 1463
rect 1012 1457 1180 1463
rect 1188 1457 1292 1463
rect 1492 1457 1564 1463
rect 1572 1457 1820 1463
rect 2196 1457 2332 1463
rect 2340 1457 2732 1463
rect 2740 1457 2876 1463
rect 3044 1457 3260 1463
rect 3300 1457 3404 1463
rect 4164 1457 4252 1463
rect 4708 1457 4748 1463
rect 4756 1457 5100 1463
rect 5332 1457 5484 1463
rect 5693 1463 5699 1476
rect 5556 1457 5699 1463
rect 5924 1457 5932 1463
rect 5972 1457 6252 1463
rect 6436 1457 6460 1463
rect 6468 1457 6572 1463
rect 6580 1457 6700 1463
rect 548 1437 716 1443
rect 724 1437 828 1443
rect 1524 1437 1596 1443
rect 1636 1437 1740 1443
rect 2212 1437 2412 1443
rect 2420 1437 2524 1443
rect 2573 1437 2652 1443
rect 532 1417 732 1423
rect 740 1417 812 1423
rect 820 1417 860 1423
rect 868 1417 1052 1423
rect 1060 1417 1276 1423
rect 1540 1417 1612 1423
rect 1620 1417 1676 1423
rect 1780 1417 1948 1423
rect 2573 1423 2579 1437
rect 5684 1437 5795 1443
rect 2404 1417 2579 1423
rect 2900 1417 3052 1423
rect 3684 1417 3756 1423
rect 3764 1417 3996 1423
rect 4004 1417 4108 1423
rect 4116 1417 4332 1423
rect 4548 1417 4572 1423
rect 4580 1417 4924 1423
rect 5789 1423 5795 1437
rect 5908 1437 5964 1443
rect 5789 1417 6140 1423
rect 6404 1417 6476 1423
rect 2632 1414 2680 1416
rect 2632 1406 2636 1414
rect 2646 1406 2652 1414
rect 2660 1406 2666 1414
rect 2676 1406 2680 1414
rect 2632 1404 2680 1406
rect 5720 1414 5768 1416
rect 5720 1406 5724 1414
rect 5734 1406 5740 1414
rect 5748 1406 5754 1414
rect 5764 1406 5768 1414
rect 5720 1404 5768 1406
rect 516 1397 684 1403
rect 1764 1397 1868 1403
rect 1940 1397 2092 1403
rect 2372 1397 2428 1403
rect 2852 1397 2860 1403
rect 2868 1397 3020 1403
rect 4148 1397 4348 1403
rect 5492 1397 5532 1403
rect 5892 1397 5964 1403
rect 6004 1397 6092 1403
rect 6372 1397 6444 1403
rect 84 1377 268 1383
rect 500 1377 668 1383
rect 724 1377 1388 1383
rect 1604 1377 2556 1383
rect 2692 1377 2748 1383
rect 3796 1377 3948 1383
rect 3956 1377 4316 1383
rect 5476 1377 5612 1383
rect 5620 1377 5699 1383
rect 612 1357 764 1363
rect 1092 1357 1548 1363
rect 1876 1357 1964 1363
rect 2468 1357 2524 1363
rect 2532 1357 2748 1363
rect 2756 1357 2892 1363
rect 3060 1357 3116 1363
rect 4260 1357 4380 1363
rect 4932 1357 5068 1363
rect 5172 1357 5196 1363
rect 5412 1357 5532 1363
rect 5540 1357 5676 1363
rect 5693 1363 5699 1377
rect 5892 1377 6044 1383
rect 6052 1377 6252 1383
rect 6580 1377 6716 1383
rect 5693 1357 6012 1363
rect 6020 1357 6572 1363
rect 276 1337 348 1343
rect 356 1337 540 1343
rect 644 1337 748 1343
rect 916 1337 1116 1343
rect 1236 1337 1612 1343
rect 1796 1337 1948 1343
rect 2660 1337 2764 1343
rect 2804 1337 3052 1343
rect 3924 1337 4339 1343
rect 4333 1324 4339 1337
rect 4548 1337 4764 1343
rect 4900 1337 5260 1343
rect 5428 1337 5436 1343
rect 5444 1337 6060 1343
rect 6068 1337 6124 1343
rect 6180 1337 6332 1343
rect 6468 1337 6508 1343
rect 6516 1337 6540 1343
rect 132 1317 380 1323
rect 404 1317 588 1323
rect 676 1317 924 1323
rect 996 1317 1004 1323
rect 1268 1317 1436 1323
rect 1492 1317 1564 1323
rect 1924 1317 1932 1323
rect 2564 1317 2716 1323
rect 2724 1317 2732 1323
rect 2884 1317 2956 1323
rect 3764 1317 4028 1323
rect 4340 1317 4364 1323
rect 4420 1317 4444 1323
rect 5076 1317 5148 1323
rect 5316 1317 5468 1323
rect 5508 1317 5596 1323
rect 5684 1317 5868 1323
rect 5940 1317 5964 1323
rect 6020 1317 6124 1323
rect 6212 1317 6380 1323
rect 6532 1317 6652 1323
rect 6692 1317 6796 1323
rect 244 1297 268 1303
rect 516 1297 572 1303
rect 580 1297 716 1303
rect 772 1297 1580 1303
rect 1732 1297 1772 1303
rect 2612 1297 2908 1303
rect 2948 1297 2972 1303
rect 3012 1297 3084 1303
rect 5348 1297 5404 1303
rect 5412 1297 5724 1303
rect 5908 1297 5964 1303
rect 6004 1297 6108 1303
rect 6180 1297 6204 1303
rect 6420 1297 6604 1303
rect 6676 1297 6684 1303
rect 388 1277 1228 1283
rect 1252 1277 1468 1283
rect 1604 1277 1852 1283
rect 1860 1277 1996 1283
rect 2004 1277 2444 1283
rect 2772 1277 2796 1283
rect 2948 1277 3276 1283
rect 5188 1277 5500 1283
rect 5572 1277 5820 1283
rect 5828 1277 5932 1283
rect 5988 1277 6444 1283
rect 285 1257 1324 1263
rect 285 1244 291 1257
rect 1348 1257 1740 1263
rect 1972 1257 3020 1263
rect 3364 1257 3420 1263
rect 4244 1257 4332 1263
rect 5956 1257 6236 1263
rect 196 1237 284 1243
rect 1028 1237 1036 1243
rect 1341 1243 1347 1256
rect 1044 1237 1347 1243
rect 1428 1237 1484 1243
rect 1492 1237 1692 1243
rect 1748 1237 1900 1243
rect 1908 1237 2028 1243
rect 2308 1237 2364 1243
rect 2397 1237 2412 1243
rect 2397 1223 2403 1237
rect 2452 1237 2508 1243
rect 3844 1237 4012 1243
rect 5380 1237 5644 1243
rect 5652 1237 6316 1243
rect 6324 1237 6348 1243
rect 6820 1237 6844 1243
rect 2132 1217 2403 1223
rect 2413 1217 2828 1223
rect 1112 1214 1160 1216
rect 1112 1206 1116 1214
rect 1126 1206 1132 1214
rect 1140 1206 1146 1214
rect 1156 1206 1160 1214
rect 1112 1204 1160 1206
rect 2413 1204 2419 1217
rect 3652 1217 4092 1223
rect 5732 1217 6204 1223
rect 6212 1217 6412 1223
rect 4152 1214 4200 1216
rect 4152 1206 4156 1214
rect 4166 1206 4172 1214
rect 4180 1206 4186 1214
rect 4196 1206 4200 1214
rect 4152 1204 4200 1206
rect 468 1197 524 1203
rect 1444 1197 1756 1203
rect 2004 1197 2220 1203
rect 2244 1197 2412 1203
rect 2500 1197 2524 1203
rect 2532 1197 2956 1203
rect 2964 1197 2972 1203
rect 2980 1197 3068 1203
rect 3076 1197 3180 1203
rect 3188 1197 3420 1203
rect 3524 1197 3644 1203
rect 3892 1197 3916 1203
rect 3924 1197 3996 1203
rect 5316 1197 5516 1203
rect 5524 1197 5788 1203
rect 5796 1197 5996 1203
rect 6356 1197 6380 1203
rect 6388 1197 6748 1203
rect 996 1177 1068 1183
rect 1188 1177 1228 1183
rect 1268 1177 1676 1183
rect 2196 1177 2364 1183
rect 2388 1177 2428 1183
rect 3508 1177 3932 1183
rect 3940 1177 4044 1183
rect 4052 1177 4156 1183
rect 4164 1177 4284 1183
rect 4404 1177 4492 1183
rect 4660 1177 4748 1183
rect 4756 1177 5868 1183
rect 6276 1177 6396 1183
rect 996 1157 1628 1163
rect 1636 1157 1772 1163
rect 1828 1157 2604 1163
rect 3860 1157 4124 1163
rect 4132 1157 4252 1163
rect 4436 1157 4716 1163
rect 4724 1157 4828 1163
rect 5236 1157 5260 1163
rect 5268 1157 5372 1163
rect 5588 1157 5660 1163
rect 5668 1157 5804 1163
rect 5812 1157 5852 1163
rect 5860 1157 5964 1163
rect 6052 1157 6300 1163
rect 6308 1157 6380 1163
rect 6532 1157 6540 1163
rect 676 1137 780 1143
rect 788 1137 812 1143
rect 1220 1137 1283 1143
rect 1277 1124 1283 1137
rect 2388 1137 2396 1143
rect 2580 1137 2588 1143
rect 2596 1137 2684 1143
rect 3092 1137 3228 1143
rect 3236 1137 3292 1143
rect 4116 1137 4796 1143
rect 4804 1137 5260 1143
rect 5508 1137 5612 1143
rect 5844 1137 5900 1143
rect 6180 1137 6252 1143
rect 6292 1137 6348 1143
rect 6532 1137 6572 1143
rect 36 1117 60 1123
rect 228 1117 252 1123
rect 564 1117 764 1123
rect 884 1117 1020 1123
rect 1060 1117 1116 1123
rect 1156 1117 1212 1123
rect 1268 1117 1276 1123
rect 1284 1117 1484 1123
rect 1748 1117 1788 1123
rect 1940 1117 1964 1123
rect 2084 1117 2220 1123
rect 2404 1117 2492 1123
rect 3220 1117 3260 1123
rect 4644 1117 5196 1123
rect 5204 1117 5212 1123
rect 5268 1117 5420 1123
rect 5444 1117 5516 1123
rect 5540 1117 5580 1123
rect 5636 1117 5804 1123
rect 5812 1117 6012 1123
rect 6020 1117 6668 1123
rect 6676 1117 6796 1123
rect 164 1097 268 1103
rect 276 1097 332 1103
rect 340 1097 604 1103
rect 676 1097 716 1103
rect 964 1097 1020 1103
rect 1076 1097 1244 1103
rect 1396 1097 1468 1103
rect 1508 1097 1564 1103
rect 1764 1097 1932 1103
rect 1940 1097 1996 1103
rect 2036 1097 2172 1103
rect 2196 1097 2268 1103
rect 3028 1097 3052 1103
rect 3060 1097 3084 1103
rect 3700 1097 3724 1103
rect 4004 1097 4060 1103
rect 4068 1097 4268 1103
rect 4548 1097 4588 1103
rect 5124 1097 5164 1103
rect 5380 1097 5836 1103
rect 5876 1097 5916 1103
rect 6484 1097 6604 1103
rect 6788 1097 6812 1103
rect 6820 1097 6876 1103
rect 260 1077 428 1083
rect 484 1077 508 1083
rect 685 1077 700 1083
rect 685 1063 691 1077
rect 884 1077 1532 1083
rect 1732 1077 1884 1083
rect 1940 1077 2012 1083
rect 2020 1077 2380 1083
rect 2676 1077 2876 1083
rect 3124 1077 3164 1083
rect 3284 1077 3484 1083
rect 3844 1077 3980 1083
rect 4036 1077 4076 1083
rect 4180 1077 4300 1083
rect 4516 1077 4668 1083
rect 4708 1077 4764 1083
rect 4820 1077 5020 1083
rect 5332 1077 5420 1083
rect 5460 1077 5532 1083
rect 5556 1077 5596 1083
rect 5604 1077 5740 1083
rect 5748 1077 5852 1083
rect 5860 1077 5948 1083
rect 6004 1077 6300 1083
rect 6356 1077 6732 1083
rect 356 1057 691 1063
rect 20 1037 60 1043
rect 685 1043 691 1057
rect 708 1057 796 1063
rect 804 1057 1004 1063
rect 1028 1057 1036 1063
rect 1348 1057 1804 1063
rect 1876 1057 1948 1063
rect 2180 1057 2204 1063
rect 2212 1057 2252 1063
rect 2260 1057 2556 1063
rect 2852 1057 3244 1063
rect 3252 1057 3452 1063
rect 3460 1057 3612 1063
rect 3620 1057 3804 1063
rect 3812 1057 3836 1063
rect 4260 1057 4412 1063
rect 4420 1057 4572 1063
rect 4580 1057 4844 1063
rect 4852 1057 4988 1063
rect 4996 1057 5292 1063
rect 5892 1057 6124 1063
rect 6244 1057 6380 1063
rect 6388 1057 6476 1063
rect 685 1037 1260 1043
rect 1268 1037 1372 1043
rect 1444 1037 1580 1043
rect 2253 1037 2316 1043
rect 2253 1024 2259 1037
rect 2324 1037 2428 1043
rect 2660 1037 3036 1043
rect 5252 1037 5468 1043
rect 5476 1037 5628 1043
rect 5636 1037 5772 1043
rect 5780 1037 5836 1043
rect 5908 1037 6012 1043
rect 6308 1037 6812 1043
rect 436 1017 940 1023
rect 948 1017 988 1023
rect 1012 1017 1212 1023
rect 1220 1017 1452 1023
rect 1460 1017 2252 1023
rect 2308 1017 2332 1023
rect 2932 1017 2956 1023
rect 2964 1017 3164 1023
rect 5076 1017 5484 1023
rect 5492 1017 5564 1023
rect 6116 1017 6156 1023
rect 2632 1014 2680 1016
rect 2632 1006 2636 1014
rect 2646 1006 2652 1014
rect 2660 1006 2666 1014
rect 2676 1006 2680 1014
rect 2632 1004 2680 1006
rect 5720 1014 5768 1016
rect 5720 1006 5724 1014
rect 5734 1006 5740 1014
rect 5748 1006 5754 1014
rect 5764 1006 5768 1014
rect 5720 1004 5768 1006
rect 324 997 428 1003
rect 804 997 1276 1003
rect 2244 997 2396 1003
rect 3588 997 3644 1003
rect 4308 997 4524 1003
rect 4532 997 4604 1003
rect 4612 997 4652 1003
rect 4916 997 4956 1003
rect 6100 997 6220 1003
rect 6420 997 6428 1003
rect 276 977 380 983
rect 436 977 460 983
rect 532 977 588 983
rect 1108 977 1308 983
rect 1316 977 1788 983
rect 4292 977 4508 983
rect 4660 977 4716 983
rect 4740 977 5180 983
rect 5844 977 6044 983
rect 6052 977 6252 983
rect 6429 983 6435 996
rect 6429 977 6860 983
rect 228 957 364 963
rect 484 957 652 963
rect 660 957 716 963
rect 724 957 908 963
rect 1012 957 1180 963
rect 1380 957 1756 963
rect 2116 957 2172 963
rect 2180 957 2316 963
rect 2324 957 2380 963
rect 2964 957 3116 963
rect 3124 957 3420 963
rect 3908 957 4284 963
rect 4580 957 4588 963
rect 4756 957 4876 963
rect 5652 957 5756 963
rect 5812 957 5836 963
rect 6004 957 6124 963
rect 6132 957 6515 963
rect 6509 944 6515 957
rect 6580 957 6588 963
rect 100 937 236 943
rect 548 937 636 943
rect 980 937 1340 943
rect 1364 937 1436 943
rect 1476 937 1724 943
rect 1972 937 2044 943
rect 2500 937 2748 943
rect 3060 937 3276 943
rect 3812 937 3916 943
rect 4132 937 4428 943
rect 4596 937 5020 943
rect 5028 937 5084 943
rect 5092 937 5100 943
rect 5108 937 5180 943
rect 5620 937 5676 943
rect 6196 937 6236 943
rect 6308 937 6364 943
rect 6372 937 6444 943
rect 6516 937 6572 943
rect 20 917 172 923
rect 212 917 380 923
rect 388 917 412 923
rect 548 917 684 923
rect 932 917 1027 923
rect 148 897 172 903
rect 180 897 1004 903
rect 1021 903 1027 917
rect 1044 917 1356 923
rect 1364 917 1452 923
rect 1636 917 1932 923
rect 3828 917 3932 923
rect 3956 917 4012 923
rect 4020 917 4115 923
rect 1021 897 1116 903
rect 1236 897 1340 903
rect 1444 897 1564 903
rect 3028 897 3084 903
rect 3876 897 4044 903
rect 4052 897 4092 903
rect 4109 903 4115 917
rect 4516 917 4604 923
rect 5524 917 5644 923
rect 5652 917 5724 923
rect 5748 917 6028 923
rect 6116 917 6204 923
rect 6308 917 6348 923
rect 6372 917 6460 923
rect 4109 897 5356 903
rect 5380 897 5532 903
rect 5604 897 5628 903
rect 5972 897 6204 903
rect 244 877 396 883
rect 532 877 828 883
rect 932 877 972 883
rect 1316 877 1388 883
rect 1492 877 1740 883
rect 1748 877 1836 883
rect 4388 877 4396 883
rect 4404 877 4764 883
rect 5284 877 5532 883
rect 6180 877 6700 883
rect 276 857 508 863
rect 516 857 572 863
rect 596 857 1292 863
rect 1300 857 1324 863
rect 1332 857 1772 863
rect 1780 857 1820 863
rect 5236 857 5676 863
rect 420 837 556 843
rect 564 837 860 843
rect 868 837 908 843
rect 1108 837 1276 843
rect 1300 837 1356 843
rect 1396 837 1692 843
rect 2388 837 2492 843
rect 4580 837 6412 843
rect 6772 837 6828 843
rect 884 817 972 823
rect 1444 817 1500 823
rect 1764 817 1868 823
rect 2573 817 3052 823
rect 1112 814 1160 816
rect 1112 806 1116 814
rect 1126 806 1132 814
rect 1140 806 1146 814
rect 1156 806 1160 814
rect 1112 804 1160 806
rect 1284 797 1548 803
rect 2573 803 2579 817
rect 3060 817 3212 823
rect 4468 817 5564 823
rect 5684 817 5692 823
rect 5732 817 5900 823
rect 4152 814 4200 816
rect 4152 806 4156 814
rect 4166 806 4172 814
rect 4180 806 4186 814
rect 4196 806 4200 814
rect 4152 804 4200 806
rect 1636 797 2579 803
rect 2596 797 2604 803
rect 2724 797 2780 803
rect 5588 797 6172 803
rect 2388 777 2684 783
rect 5572 777 5820 783
rect 6228 777 6332 783
rect 6644 777 6668 783
rect 868 757 1404 763
rect 1732 757 1756 763
rect 2612 757 2636 763
rect 5428 757 5804 763
rect 5828 757 5868 763
rect 5876 757 6124 763
rect 6132 757 6252 763
rect 6708 757 6844 763
rect 349 737 1420 743
rect 349 724 355 737
rect 1453 737 1564 743
rect 196 717 252 723
rect 260 717 348 723
rect 388 717 428 723
rect 468 717 732 723
rect 916 717 940 723
rect 948 717 1260 723
rect 1453 723 1459 737
rect 1700 737 2316 743
rect 2324 737 2908 743
rect 3012 737 3148 743
rect 3156 737 3340 743
rect 3540 737 3612 743
rect 3780 737 3900 743
rect 3972 737 4652 743
rect 5028 737 5132 743
rect 5780 737 5836 743
rect 5860 737 6108 743
rect 6116 737 6236 743
rect 6301 737 6428 743
rect 6301 724 6307 737
rect 6436 737 6444 743
rect 6804 737 6844 743
rect 1332 717 1459 723
rect 1476 717 1532 723
rect 1604 717 1660 723
rect 1668 717 1724 723
rect 1764 717 1852 723
rect 3444 717 3500 723
rect 3988 717 4044 723
rect 4788 717 5084 723
rect 5188 717 5388 723
rect 5444 717 5635 723
rect 308 697 380 703
rect 516 697 604 703
rect 1028 697 1148 703
rect 1284 697 1372 703
rect 1412 697 1628 703
rect 1716 697 1740 703
rect 1844 697 1932 703
rect 2244 697 2300 703
rect 2308 697 2732 703
rect 2740 697 2892 703
rect 2948 697 2988 703
rect 4004 697 4316 703
rect 4500 697 4540 703
rect 5364 697 5388 703
rect 5412 697 5420 703
rect 5540 697 5612 703
rect 5629 703 5635 717
rect 5700 717 6012 723
rect 6276 717 6300 723
rect 6468 717 6636 723
rect 5629 697 5852 703
rect 6356 697 6396 703
rect 6436 697 6524 703
rect 6548 697 6668 703
rect 68 677 316 683
rect 324 677 476 683
rect 484 677 636 683
rect 1076 677 1228 683
rect 1444 677 1715 683
rect 1709 664 1715 677
rect 1732 677 2028 683
rect 2052 677 2124 683
rect 2132 677 2892 683
rect 2964 677 3068 683
rect 3892 677 4636 683
rect 5332 677 6716 683
rect 6724 677 6732 683
rect 100 657 268 663
rect 1140 657 1324 663
rect 1540 657 1612 663
rect 1716 657 1804 663
rect 1812 657 1900 663
rect 1908 657 1916 663
rect 2068 657 2268 663
rect 2276 657 2396 663
rect 2500 657 2524 663
rect 2932 657 3148 663
rect 4628 657 4684 663
rect 4980 657 5036 663
rect 5044 657 5116 663
rect 5684 657 6028 663
rect 6548 657 6684 663
rect 6724 657 6732 663
rect 212 637 524 643
rect 676 637 1116 643
rect 1204 637 1228 643
rect 1604 637 2764 643
rect 2772 637 2867 643
rect 580 617 652 623
rect 660 617 828 623
rect 836 617 876 623
rect 900 617 1260 623
rect 2356 617 2524 623
rect 2861 623 2867 637
rect 2884 637 3052 643
rect 3364 637 3692 643
rect 5364 637 5420 643
rect 5428 637 5516 643
rect 6100 637 6364 643
rect 6372 637 6396 643
rect 2861 617 2988 623
rect 3492 617 3724 623
rect 4516 617 5596 623
rect 5844 617 5996 623
rect 6148 617 6364 623
rect 2632 614 2680 616
rect 2632 606 2636 614
rect 2646 606 2652 614
rect 2660 606 2666 614
rect 2676 606 2680 614
rect 2632 604 2680 606
rect 5720 614 5768 616
rect 5720 606 5724 614
rect 5734 606 5740 614
rect 5748 606 5754 614
rect 5764 606 5768 614
rect 5720 604 5768 606
rect 516 597 588 603
rect 1108 597 1132 603
rect 3796 597 3948 603
rect 4196 597 4460 603
rect 4756 597 4812 603
rect 5684 597 5692 603
rect 5812 597 5932 603
rect 500 577 844 583
rect 948 577 1308 583
rect 1508 577 1644 583
rect 2564 577 2972 583
rect 2980 577 3068 583
rect 3604 577 3868 583
rect 4004 577 4476 583
rect 4916 577 5020 583
rect 5293 577 5516 583
rect 5293 564 5299 577
rect 5524 577 5580 583
rect 5892 577 5996 583
rect 6788 577 6796 583
rect 212 557 220 563
rect 308 557 412 563
rect 548 557 940 563
rect 1140 557 1228 563
rect 1268 557 1404 563
rect 1940 557 2140 563
rect 2148 557 2156 563
rect 2484 557 2572 563
rect 2580 557 2956 563
rect 3028 557 3100 563
rect 3332 557 3756 563
rect 3764 557 4156 563
rect 4164 557 4284 563
rect 5060 557 5180 563
rect 5204 557 5292 563
rect 5412 557 5676 563
rect 5821 563 5827 576
rect 5821 557 5948 563
rect 6276 557 6540 563
rect 6740 557 6860 563
rect 100 537 268 543
rect 308 537 364 543
rect 452 537 915 543
rect 228 517 540 523
rect 612 517 700 523
rect 909 523 915 537
rect 932 537 1180 543
rect 1188 537 1308 543
rect 2772 537 2972 543
rect 3044 537 3276 543
rect 3284 537 3564 543
rect 3572 537 3884 543
rect 3908 537 3932 543
rect 3940 537 4012 543
rect 4420 537 4428 543
rect 4500 537 4540 543
rect 4548 537 4572 543
rect 4724 537 4924 543
rect 5108 537 5244 543
rect 5396 537 5436 543
rect 5620 537 5804 543
rect 5812 537 5852 543
rect 5988 537 6188 543
rect 6196 537 6284 543
rect 6292 537 6348 543
rect 6372 537 6428 543
rect 6468 537 6508 543
rect 6612 537 6668 543
rect 6692 537 6876 543
rect 909 517 956 523
rect 964 517 1052 523
rect 1204 517 1324 523
rect 1396 517 1484 523
rect 1492 517 1516 523
rect 1588 517 1628 523
rect 1652 517 1820 523
rect 2100 517 2156 523
rect 2612 517 2668 523
rect 3588 517 3676 523
rect 4292 517 4396 523
rect 4564 517 4620 523
rect 4948 517 5004 523
rect 5044 517 5148 523
rect 5236 517 5292 523
rect 5316 517 5532 523
rect 5588 517 5964 523
rect 6036 517 6252 523
rect 6420 517 6499 523
rect 196 497 252 503
rect 260 497 492 503
rect 516 497 524 503
rect 884 497 908 503
rect 948 497 1372 503
rect 1380 497 1420 503
rect 1428 497 1452 503
rect 1572 497 1692 503
rect 2068 497 2188 503
rect 2884 497 2956 503
rect 2964 497 3020 503
rect 4996 497 5084 503
rect 5348 497 5404 503
rect 5556 497 5628 503
rect 6004 497 6204 503
rect 6212 497 6444 503
rect 6493 503 6499 517
rect 6516 517 6604 523
rect 6612 517 6780 523
rect 6493 497 6684 503
rect 6724 497 6764 503
rect 6772 497 6812 503
rect 1300 477 1324 483
rect 1364 477 1404 483
rect 1412 477 1436 483
rect 1444 477 1596 483
rect 1684 477 1708 483
rect 1732 477 1756 483
rect 4980 477 5068 483
rect 5076 477 5116 483
rect 5700 477 5836 483
rect 5892 477 5939 483
rect 804 457 2124 463
rect 5156 457 5468 463
rect 5492 457 5916 463
rect 5933 463 5939 477
rect 6132 477 6460 483
rect 6484 477 6508 483
rect 6724 477 6860 483
rect 5933 457 6572 463
rect 6580 457 6636 463
rect 6820 457 6844 463
rect 132 437 172 443
rect 916 437 940 443
rect 6164 437 6332 443
rect 6372 437 6588 443
rect 6740 437 6796 443
rect 916 417 972 423
rect 1188 417 1580 423
rect 1588 417 1756 423
rect 4548 417 4684 423
rect 4692 417 4796 423
rect 6292 417 6380 423
rect 1112 414 1160 416
rect 1112 406 1116 414
rect 1126 406 1132 414
rect 1140 406 1146 414
rect 1156 406 1160 414
rect 1112 404 1160 406
rect 4152 414 4200 416
rect 4152 406 4156 414
rect 4166 406 4172 414
rect 4180 406 4186 414
rect 4196 406 4200 414
rect 4152 404 4200 406
rect 2532 397 2780 403
rect 3716 397 3948 403
rect 4436 397 4780 403
rect 5140 397 5212 403
rect 1012 377 1356 383
rect 1364 377 1468 383
rect 1700 377 1724 383
rect 2340 377 2492 383
rect 2500 377 2796 383
rect 2804 377 2908 383
rect 4276 377 4332 383
rect 4580 377 4636 383
rect 4644 377 4732 383
rect 5156 377 5308 383
rect 5604 377 6092 383
rect 6260 377 6364 383
rect 6388 377 6668 383
rect 1044 357 1068 363
rect 4084 357 4220 363
rect 5508 357 6380 363
rect 6644 357 6668 363
rect 420 337 492 343
rect 500 337 572 343
rect 1044 337 1196 343
rect 3028 337 3484 343
rect 3860 337 4140 343
rect 4788 337 4844 343
rect 4852 337 5052 343
rect 5284 337 5388 343
rect 5396 337 5436 343
rect 5572 337 5676 343
rect 5684 337 5724 343
rect 5940 337 6092 343
rect 6116 337 6268 343
rect 6356 337 6476 343
rect 6484 337 6540 343
rect 6644 337 6844 343
rect 340 317 460 323
rect 596 317 636 323
rect 1108 317 1228 323
rect 1428 317 1564 323
rect 3092 317 3116 323
rect 4116 317 4348 323
rect 4484 317 4620 323
rect 4628 317 4668 323
rect 4836 317 4860 323
rect 5252 317 5516 323
rect 5540 317 6188 323
rect 6228 317 6316 323
rect 6516 317 6604 323
rect 6628 317 6716 323
rect 36 297 412 303
rect 420 297 604 303
rect 996 297 1100 303
rect 1348 297 1372 303
rect 1444 297 1484 303
rect 1508 297 1596 303
rect 1780 297 1868 303
rect 2468 297 2764 303
rect 2900 297 3020 303
rect 3060 297 3084 303
rect 3604 297 3708 303
rect 4116 297 4140 303
rect 4292 297 4348 303
rect 4452 297 4764 303
rect 4772 297 4828 303
rect 4836 297 5036 303
rect 5172 297 5308 303
rect 5476 297 5564 303
rect 5668 297 5836 303
rect 6221 303 6227 316
rect 5988 297 6227 303
rect 6308 297 6492 303
rect 6500 297 6620 303
rect 6628 297 6748 303
rect 148 277 428 283
rect 468 277 588 283
rect 932 277 988 283
rect 996 277 1052 283
rect 1060 277 1372 283
rect 1428 277 1532 283
rect 1773 283 1779 296
rect 1540 277 1779 283
rect 1812 277 1852 283
rect 1860 277 1964 283
rect 1988 277 2188 283
rect 2740 277 2764 283
rect 2772 277 2844 283
rect 2852 277 3036 283
rect 3044 277 3132 283
rect 3668 277 4012 283
rect 4020 277 4156 283
rect 4164 277 4268 283
rect 4452 277 4700 283
rect 5044 277 5372 283
rect 5396 277 5404 283
rect 5508 277 5596 283
rect 5924 277 6044 283
rect 6180 277 6188 283
rect 6196 277 6300 283
rect 6484 277 6588 283
rect 6612 277 6732 283
rect 6756 277 6764 283
rect 388 257 972 263
rect 1124 257 1260 263
rect 1268 257 1420 263
rect 1748 257 1820 263
rect 2580 257 2924 263
rect 3092 257 3340 263
rect 4676 257 4892 263
rect 4900 257 4988 263
rect 4996 257 5340 263
rect 5364 257 5404 263
rect 6372 257 6604 263
rect 6740 257 6876 263
rect 2612 237 2652 243
rect 3156 237 3212 243
rect 3764 237 4044 243
rect 6740 237 6812 243
rect 3380 217 3628 223
rect 6148 217 6492 223
rect 2632 214 2680 216
rect 2632 206 2636 214
rect 2646 206 2652 214
rect 2660 206 2666 214
rect 2676 206 2680 214
rect 2632 204 2680 206
rect 5720 214 5768 216
rect 5720 206 5724 214
rect 5734 206 5740 214
rect 5748 206 5754 214
rect 5764 206 5768 214
rect 5720 204 5768 206
rect 644 197 684 203
rect 948 197 1036 203
rect 1460 197 1644 203
rect 1652 197 1788 203
rect 3540 197 3596 203
rect 3604 197 3772 203
rect 3780 197 3884 203
rect 3892 197 3964 203
rect 4420 197 4476 203
rect 4484 197 4748 203
rect 4756 197 4844 203
rect 4852 197 5132 203
rect 5140 197 5212 203
rect 6260 197 6428 203
rect 1668 177 1836 183
rect 1844 177 2172 183
rect 2676 177 2716 183
rect 2916 177 3004 183
rect 3012 177 3180 183
rect 3188 177 3308 183
rect 5476 177 5756 183
rect 5892 177 5964 183
rect 5972 177 6140 183
rect 6292 177 6412 183
rect 6548 177 6620 183
rect 180 157 204 163
rect 212 157 652 163
rect 916 157 1004 163
rect 1012 157 1244 163
rect 1476 157 1596 163
rect 1604 157 1676 163
rect 1684 157 1740 163
rect 1972 157 2076 163
rect 2148 157 2444 163
rect 2516 157 2764 163
rect 2836 157 3036 163
rect 3940 157 4172 163
rect 5604 157 5820 163
rect 6084 157 6284 163
rect 6308 157 6396 163
rect 36 137 172 143
rect 452 137 508 143
rect 516 137 844 143
rect 852 137 892 143
rect 1572 137 1868 143
rect 2372 137 2396 143
rect 2740 137 2828 143
rect 3236 137 3276 143
rect 3284 137 3292 143
rect 3572 137 3692 143
rect 4132 137 4188 143
rect 4196 137 4300 143
rect 4388 137 4588 143
rect 5188 137 5388 143
rect 6292 137 6316 143
rect 6596 137 6700 143
rect 292 117 572 123
rect 788 117 924 123
rect 2260 117 2348 123
rect 2388 117 2476 123
rect 3140 117 3244 123
rect 3668 117 3788 123
rect 3796 117 3836 123
rect 4052 117 4284 123
rect 4500 117 4764 123
rect 4996 117 5052 123
rect 5060 117 5084 123
rect 5300 117 5468 123
rect 6036 117 6396 123
rect 6564 117 6732 123
rect 6836 117 6844 123
rect 1124 97 2028 103
rect 2452 97 2508 103
rect 2548 97 2604 103
rect 2820 97 2860 103
rect 6020 97 6092 103
rect 6308 97 6540 103
rect 6804 97 6812 103
rect 6244 77 6364 83
rect 4132 37 4156 43
rect 4932 17 4940 23
rect 1112 14 1160 16
rect 1112 6 1116 14
rect 1126 6 1132 14
rect 1140 6 1146 14
rect 1156 6 1160 14
rect 1112 4 1160 6
rect 4152 14 4200 16
rect 4152 6 4156 14
rect 4166 6 4172 14
rect 4180 6 4186 14
rect 4196 6 4200 14
rect 4152 4 4200 6
<< m4contact >>
rect 2636 5006 2638 5014
rect 2638 5006 2644 5014
rect 2652 5006 2660 5014
rect 2668 5006 2674 5014
rect 2674 5006 2676 5014
rect 5724 5006 5726 5014
rect 5726 5006 5732 5014
rect 5740 5006 5748 5014
rect 5756 5006 5762 5014
rect 5762 5006 5764 5014
rect 2252 4996 2260 5004
rect 4844 4996 4852 5004
rect 5516 4996 5524 5004
rect 460 4896 468 4904
rect 5484 4836 5492 4844
rect 1116 4806 1118 4814
rect 1118 4806 1124 4814
rect 1132 4806 1140 4814
rect 1148 4806 1154 4814
rect 1154 4806 1156 4814
rect 4156 4806 4158 4814
rect 4158 4806 4164 4814
rect 4172 4806 4180 4814
rect 4188 4806 4194 4814
rect 4194 4806 4196 4814
rect 2764 4716 2772 4724
rect 3980 4716 3988 4724
rect 6540 4716 6548 4724
rect 6444 4696 6452 4704
rect 6700 4696 6708 4704
rect 940 4676 948 4684
rect 6508 4676 6516 4684
rect 3436 4656 3444 4664
rect 3820 4656 3828 4664
rect 1612 4636 1620 4644
rect 6732 4636 6740 4644
rect 4844 4616 4852 4624
rect 5516 4616 5524 4624
rect 2636 4606 2638 4614
rect 2638 4606 2644 4614
rect 2652 4606 2660 4614
rect 2668 4606 2674 4614
rect 2674 4606 2676 4614
rect 5724 4606 5726 4614
rect 5726 4606 5732 4614
rect 5740 4606 5748 4614
rect 5756 4606 5762 4614
rect 5762 4606 5764 4614
rect 2956 4596 2964 4604
rect 6572 4576 6580 4584
rect 428 4556 436 4564
rect 3052 4556 3060 4564
rect 1644 4536 1652 4544
rect 1708 4536 1716 4544
rect 3692 4516 3700 4524
rect 3884 4516 3892 4524
rect 652 4496 660 4504
rect 4780 4496 4788 4504
rect 5964 4496 5972 4504
rect 6284 4496 6292 4504
rect 6636 4496 6644 4504
rect 6316 4476 6324 4484
rect 2764 4436 2772 4444
rect 6508 4416 6516 4424
rect 1116 4406 1118 4414
rect 1118 4406 1124 4414
rect 1132 4406 1140 4414
rect 1148 4406 1154 4414
rect 1154 4406 1156 4414
rect 4156 4406 4158 4414
rect 4158 4406 4164 4414
rect 4172 4406 4180 4414
rect 4188 4406 4194 4414
rect 4194 4406 4196 4414
rect 3468 4376 3476 4384
rect 3660 4376 3668 4384
rect 428 4356 436 4364
rect 3692 4356 3700 4364
rect 3820 4356 3828 4364
rect 3724 4336 3732 4344
rect 332 4316 340 4324
rect 364 4296 372 4304
rect 3340 4296 3348 4304
rect 5324 4316 5332 4324
rect 5580 4316 5588 4324
rect 1612 4276 1620 4284
rect 2732 4276 2740 4284
rect 2956 4276 2964 4284
rect 3052 4276 3060 4284
rect 6316 4296 6324 4304
rect 3852 4276 3860 4284
rect 5068 4276 5076 4284
rect 5356 4276 5364 4284
rect 5612 4276 5620 4284
rect 3980 4256 3988 4264
rect 5420 4256 5428 4264
rect 876 4236 884 4244
rect 1644 4236 1652 4244
rect 3468 4236 3476 4244
rect 3884 4236 3892 4244
rect 6156 4236 6164 4244
rect 780 4216 788 4224
rect 1708 4216 1716 4224
rect 3436 4216 3444 4224
rect 2636 4206 2638 4214
rect 2638 4206 2644 4214
rect 2652 4206 2660 4214
rect 2668 4206 2674 4214
rect 2674 4206 2676 4214
rect 5724 4206 5726 4214
rect 5726 4206 5732 4214
rect 5740 4206 5748 4214
rect 5756 4206 5762 4214
rect 5762 4206 5764 4214
rect 652 4196 660 4204
rect 908 4196 916 4204
rect 1036 4196 1044 4204
rect 2700 4196 2708 4204
rect 3340 4196 3348 4204
rect 588 4176 596 4184
rect 2924 4176 2932 4184
rect 300 4156 308 4164
rect 1708 4156 1716 4164
rect 3244 4156 3252 4164
rect 3916 4156 3924 4164
rect 5964 4156 5972 4164
rect 6700 4156 6708 4164
rect 6764 4156 6772 4164
rect 3980 4136 3988 4144
rect 5612 4136 5620 4144
rect 5676 4136 5684 4144
rect 6828 4136 6836 4144
rect 1772 4116 1780 4124
rect 3276 4116 3284 4124
rect 3596 4116 3604 4124
rect 3884 4116 3892 4124
rect 620 4096 628 4104
rect 5420 4096 5428 4104
rect 652 4076 660 4084
rect 3724 4076 3732 4084
rect 3852 4076 3860 4084
rect 5484 4076 5492 4084
rect 5516 4076 5524 4084
rect 5676 4076 5684 4084
rect 1260 4056 1268 4064
rect 3148 4056 3156 4064
rect 2860 4036 2868 4044
rect 3404 4036 3412 4044
rect 3660 4036 3668 4044
rect 5324 4036 5332 4044
rect 6380 4016 6388 4024
rect 1116 4006 1118 4014
rect 1118 4006 1124 4014
rect 1132 4006 1140 4014
rect 1148 4006 1154 4014
rect 1154 4006 1156 4014
rect 4156 4006 4158 4014
rect 4158 4006 4164 4014
rect 4172 4006 4180 4014
rect 4188 4006 4194 4014
rect 4194 4006 4196 4014
rect 300 3996 308 4004
rect 6508 3996 6516 4004
rect 684 3976 692 3984
rect 716 3956 724 3964
rect 4780 3956 4788 3964
rect 4812 3956 4820 3964
rect 5900 3956 5908 3964
rect 1420 3936 1428 3944
rect 3628 3936 3636 3944
rect 5196 3936 5204 3944
rect 1036 3916 1044 3924
rect 1772 3916 1780 3924
rect 588 3896 596 3904
rect 2028 3896 2036 3904
rect 5068 3896 5076 3904
rect 6412 3896 6420 3904
rect 652 3876 660 3884
rect 1388 3876 1396 3884
rect 3020 3876 3028 3884
rect 3596 3876 3604 3884
rect 4300 3876 4308 3884
rect 332 3856 340 3864
rect 1420 3856 1428 3864
rect 1516 3856 1524 3864
rect 2412 3856 2420 3864
rect 3468 3856 3476 3864
rect 5196 3856 5204 3864
rect 5356 3856 5364 3864
rect 6348 3856 6356 3864
rect 4940 3836 4948 3844
rect 5612 3836 5620 3844
rect 5868 3836 5876 3844
rect 2252 3816 2260 3824
rect 2572 3816 2580 3824
rect 2956 3816 2964 3824
rect 3180 3816 3188 3824
rect 3980 3816 3988 3824
rect 5676 3816 5684 3824
rect 2636 3806 2638 3814
rect 2638 3806 2644 3814
rect 2652 3806 2660 3814
rect 2668 3806 2674 3814
rect 2674 3806 2676 3814
rect 5724 3806 5726 3814
rect 5726 3806 5732 3814
rect 5740 3806 5748 3814
rect 5756 3806 5762 3814
rect 5762 3806 5764 3814
rect 2124 3796 2132 3804
rect 3660 3796 3668 3804
rect 4908 3796 4916 3804
rect 364 3776 372 3784
rect 3212 3776 3220 3784
rect 5676 3776 5684 3784
rect 6188 3776 6196 3784
rect 716 3756 724 3764
rect 2924 3756 2932 3764
rect 5900 3756 5908 3764
rect 6380 3756 6388 3764
rect 3436 3736 3444 3744
rect 6284 3736 6292 3744
rect 6316 3736 6324 3744
rect 6572 3736 6580 3744
rect 6796 3736 6804 3744
rect 940 3716 948 3724
rect 2860 3716 2868 3724
rect 3404 3716 3412 3724
rect 3628 3716 3636 3724
rect 3852 3696 3860 3704
rect 4108 3676 4116 3684
rect 6476 3676 6484 3684
rect 6572 3676 6580 3684
rect 3244 3656 3252 3664
rect 3756 3616 3764 3624
rect 5548 3616 5556 3624
rect 1116 3606 1118 3614
rect 1118 3606 1124 3614
rect 1132 3606 1140 3614
rect 1148 3606 1154 3614
rect 1154 3606 1156 3614
rect 4156 3606 4158 3614
rect 4158 3606 4164 3614
rect 4172 3606 4180 3614
rect 4188 3606 4194 3614
rect 4194 3606 4196 3614
rect 5388 3596 5396 3604
rect 5644 3596 5652 3604
rect 1516 3576 1524 3584
rect 3340 3576 3348 3584
rect 3500 3576 3508 3584
rect 3660 3576 3668 3584
rect 6700 3576 6708 3584
rect 3148 3556 3156 3564
rect 3468 3556 3476 3564
rect 6060 3556 6068 3564
rect 780 3536 788 3544
rect 1260 3536 1268 3544
rect 2732 3536 2740 3544
rect 3116 3536 3124 3544
rect 3276 3536 3284 3544
rect 3308 3536 3316 3544
rect 5228 3536 5236 3544
rect 6380 3536 6388 3544
rect 908 3516 916 3524
rect 3020 3516 3028 3524
rect 3180 3516 3188 3524
rect 1676 3496 1684 3504
rect 3564 3496 3572 3504
rect 5580 3516 5588 3524
rect 6604 3516 6612 3524
rect 5868 3496 5876 3504
rect 4300 3476 4308 3484
rect 4780 3476 4788 3484
rect 1388 3456 1396 3464
rect 2700 3456 2708 3464
rect 3660 3456 3668 3464
rect 6316 3456 6324 3464
rect 6636 3476 6644 3484
rect 6668 3476 6676 3484
rect 6604 3456 6612 3464
rect 3340 3436 3348 3444
rect 3468 3436 3476 3444
rect 5580 3436 5588 3444
rect 6540 3436 6548 3444
rect 5452 3416 5460 3424
rect 2636 3406 2638 3414
rect 2638 3406 2644 3414
rect 2652 3406 2660 3414
rect 2668 3406 2674 3414
rect 2674 3406 2676 3414
rect 5724 3406 5726 3414
rect 5726 3406 5732 3414
rect 5740 3406 5748 3414
rect 5756 3406 5762 3414
rect 5762 3406 5764 3414
rect 3212 3396 3220 3404
rect 940 3376 948 3384
rect 1548 3376 1556 3384
rect 2412 3376 2420 3384
rect 5388 3396 5396 3404
rect 684 3356 692 3364
rect 3916 3356 3924 3364
rect 4812 3356 4820 3364
rect 5580 3356 5588 3364
rect 6380 3356 6388 3364
rect 6636 3356 6644 3364
rect 1548 3336 1556 3344
rect 3308 3336 3316 3344
rect 2124 3316 2132 3324
rect 172 3296 180 3304
rect 1676 3296 1684 3304
rect 3564 3296 3572 3304
rect 4268 3296 4276 3304
rect 4716 3296 4724 3304
rect 4940 3296 4948 3304
rect 5420 3296 5428 3304
rect 4780 3276 4788 3284
rect 5068 3276 5076 3284
rect 3852 3236 3860 3244
rect 5644 3236 5652 3244
rect 940 3216 948 3224
rect 3500 3216 3508 3224
rect 1116 3206 1118 3214
rect 1118 3206 1124 3214
rect 1132 3206 1140 3214
rect 1148 3206 1154 3214
rect 1154 3206 1156 3214
rect 4156 3206 4158 3214
rect 4158 3206 4164 3214
rect 4172 3206 4180 3214
rect 4188 3206 4194 3214
rect 4194 3206 4196 3214
rect 1900 3176 1908 3184
rect 3372 3176 3380 3184
rect 3756 3176 3764 3184
rect 460 3156 468 3164
rect 4940 3176 4948 3184
rect 5612 3136 5620 3144
rect 2796 3116 2804 3124
rect 3116 3116 3124 3124
rect 5580 3096 5588 3104
rect 5996 3096 6004 3104
rect 2572 3076 2580 3084
rect 2764 3076 2772 3084
rect 3436 3076 3444 3084
rect 3596 3076 3604 3084
rect 6156 3076 6164 3084
rect 172 3056 180 3064
rect 620 3056 628 3064
rect 1868 3056 1876 3064
rect 3532 3056 3540 3064
rect 6412 3056 6420 3064
rect 6540 3056 6548 3064
rect 6668 3056 6676 3064
rect 2156 3036 2164 3044
rect 2636 3006 2638 3014
rect 2638 3006 2644 3014
rect 2652 3006 2660 3014
rect 2668 3006 2674 3014
rect 2674 3006 2676 3014
rect 5724 3006 5726 3014
rect 5726 3006 5732 3014
rect 5740 3006 5748 3014
rect 5756 3006 5762 3014
rect 5762 3006 5764 3014
rect 1900 2976 1908 2984
rect 5580 2976 5588 2984
rect 4364 2956 4372 2964
rect 4556 2956 4564 2964
rect 2796 2936 2804 2944
rect 6700 2936 6708 2944
rect 3788 2916 3796 2924
rect 4044 2916 4052 2924
rect 5228 2916 5236 2924
rect 5452 2916 5460 2924
rect 6028 2916 6036 2924
rect 4716 2896 4724 2904
rect 6700 2896 6708 2904
rect 6764 2896 6772 2904
rect 3724 2856 3732 2864
rect 876 2836 884 2844
rect 2156 2836 2164 2844
rect 5996 2836 6004 2844
rect 1116 2806 1118 2814
rect 1118 2806 1124 2814
rect 1132 2806 1140 2814
rect 1148 2806 1154 2814
rect 1154 2806 1156 2814
rect 4156 2806 4158 2814
rect 4158 2806 4164 2814
rect 4172 2806 4180 2814
rect 4188 2806 4194 2814
rect 4194 2806 4196 2814
rect 3500 2796 3508 2804
rect 5068 2796 5076 2804
rect 1580 2776 1588 2784
rect 2380 2776 2388 2784
rect 3148 2756 3156 2764
rect 3660 2756 3668 2764
rect 3820 2756 3828 2764
rect 4108 2736 4116 2744
rect 2924 2716 2932 2724
rect 3404 2716 3412 2724
rect 3596 2716 3604 2724
rect 6412 2716 6420 2724
rect 3756 2696 3764 2704
rect 3852 2696 3860 2704
rect 6604 2696 6612 2704
rect 2732 2676 2740 2684
rect 2860 2676 2868 2684
rect 3436 2676 3444 2684
rect 6348 2676 6356 2684
rect 172 2656 180 2664
rect 1868 2656 1876 2664
rect 3532 2656 3540 2664
rect 3564 2656 3572 2664
rect 3756 2656 3764 2664
rect 4556 2656 4564 2664
rect 5484 2616 5492 2624
rect 5548 2616 5556 2624
rect 2636 2606 2638 2614
rect 2638 2606 2644 2614
rect 2652 2606 2660 2614
rect 2668 2606 2674 2614
rect 2674 2606 2676 2614
rect 5724 2606 5726 2614
rect 5726 2606 5732 2614
rect 5740 2606 5748 2614
rect 5756 2606 5762 2614
rect 5762 2606 5764 2614
rect 1228 2596 1236 2604
rect 2956 2596 2964 2604
rect 3692 2596 3700 2604
rect 6668 2596 6676 2604
rect 3404 2576 3412 2584
rect 3500 2576 3508 2584
rect 4460 2576 4468 2584
rect 4556 2576 4564 2584
rect 5516 2576 5524 2584
rect 1068 2556 1076 2564
rect 1580 2556 1588 2564
rect 4364 2556 4372 2564
rect 3308 2536 3316 2544
rect 3372 2536 3380 2544
rect 6540 2536 6548 2544
rect 3148 2516 3156 2524
rect 3916 2516 3924 2524
rect 5484 2516 5492 2524
rect 6412 2516 6420 2524
rect 2892 2496 2900 2504
rect 3212 2476 3220 2484
rect 3244 2476 3252 2484
rect 4268 2496 4276 2504
rect 6572 2496 6580 2504
rect 6668 2496 6676 2504
rect 2924 2456 2932 2464
rect 3276 2456 3284 2464
rect 2604 2436 2612 2444
rect 3372 2436 3380 2444
rect 6796 2436 6804 2444
rect 2860 2416 2868 2424
rect 2956 2416 2964 2424
rect 3404 2416 3412 2424
rect 1116 2406 1118 2414
rect 1118 2406 1124 2414
rect 1132 2406 1140 2414
rect 1148 2406 1154 2414
rect 1154 2406 1156 2414
rect 4156 2406 4158 2414
rect 4158 2406 4164 2414
rect 4172 2406 4180 2414
rect 4188 2406 4194 2414
rect 4194 2406 4196 2414
rect 1228 2376 1236 2384
rect 6540 2396 6548 2404
rect 3308 2356 3316 2364
rect 3692 2356 3700 2364
rect 6604 2356 6612 2364
rect 6828 2356 6836 2364
rect 3276 2336 3284 2344
rect 2380 2316 2388 2324
rect 6860 2296 6868 2304
rect 3852 2276 3860 2284
rect 1580 2256 1588 2264
rect 1932 2256 1940 2264
rect 2860 2256 2868 2264
rect 3244 2256 3252 2264
rect 3436 2236 3444 2244
rect 3756 2236 3764 2244
rect 1388 2216 1396 2224
rect 2732 2216 2740 2224
rect 3724 2216 3732 2224
rect 2636 2206 2638 2214
rect 2638 2206 2644 2214
rect 2652 2206 2660 2214
rect 2668 2206 2674 2214
rect 2674 2206 2676 2214
rect 5724 2206 5726 2214
rect 5726 2206 5732 2214
rect 5740 2206 5748 2214
rect 5756 2206 5762 2214
rect 5762 2206 5764 2214
rect 4044 2196 4052 2204
rect 4108 2196 4116 2204
rect 1580 2176 1588 2184
rect 1068 2156 1076 2164
rect 2604 2156 2612 2164
rect 2892 2156 2900 2164
rect 3212 2136 3220 2144
rect 3884 2136 3892 2144
rect 1388 2116 1396 2124
rect 2732 2116 2740 2124
rect 3276 2116 3284 2124
rect 3916 2116 3924 2124
rect 4332 2116 4340 2124
rect 5996 2116 6004 2124
rect 4268 2076 4276 2084
rect 4364 2076 4372 2084
rect 6796 2056 6804 2064
rect 1116 2006 1118 2014
rect 1118 2006 1124 2014
rect 1132 2006 1140 2014
rect 1148 2006 1154 2014
rect 1154 2006 1156 2014
rect 4156 2006 4158 2014
rect 4158 2006 4164 2014
rect 4172 2006 4180 2014
rect 4188 2006 4194 2014
rect 4194 2006 4196 2014
rect 6828 1996 6836 2004
rect 3756 1976 3764 1984
rect 3820 1976 3828 1984
rect 4268 1976 4276 1984
rect 4940 1976 4948 1984
rect 6188 1976 6196 1984
rect 6348 1976 6356 1984
rect 6540 1956 6548 1964
rect 6636 1956 6644 1964
rect 3756 1936 3764 1944
rect 4364 1936 4372 1944
rect 6572 1936 6580 1944
rect 6764 1936 6772 1944
rect 6444 1916 6452 1924
rect 908 1896 916 1904
rect 4044 1896 4052 1904
rect 172 1876 180 1884
rect 4364 1876 4372 1884
rect 4460 1876 4468 1884
rect 6476 1876 6484 1884
rect 3084 1856 3092 1864
rect 4012 1856 4020 1864
rect 6124 1856 6132 1864
rect 6636 1856 6644 1864
rect 140 1836 148 1844
rect 1740 1836 1748 1844
rect 172 1816 180 1824
rect 4108 1836 4116 1844
rect 5676 1836 5684 1844
rect 2636 1806 2638 1814
rect 2638 1806 2644 1814
rect 2652 1806 2660 1814
rect 2668 1806 2674 1814
rect 2674 1806 2676 1814
rect 5724 1806 5726 1814
rect 5726 1806 5732 1814
rect 5740 1806 5748 1814
rect 5756 1806 5762 1814
rect 5762 1806 5764 1814
rect 5324 1796 5332 1804
rect 6636 1776 6644 1784
rect 6668 1776 6676 1784
rect 4844 1756 4852 1764
rect 4908 1756 4916 1764
rect 6796 1756 6804 1764
rect 300 1736 308 1744
rect 2028 1736 2036 1744
rect 2796 1736 2804 1744
rect 3468 1736 3476 1744
rect 1580 1716 1588 1724
rect 524 1696 532 1704
rect 3436 1696 3444 1704
rect 5260 1696 5268 1704
rect 5836 1696 5844 1704
rect 5196 1676 5204 1684
rect 6796 1676 6804 1684
rect 428 1656 436 1664
rect 1932 1656 1940 1664
rect 5676 1656 5684 1664
rect 908 1636 916 1644
rect 1484 1636 1492 1644
rect 5036 1636 5044 1644
rect 5292 1636 5300 1644
rect 5804 1636 5812 1644
rect 6060 1636 6068 1644
rect 6092 1636 6100 1644
rect 6700 1636 6708 1644
rect 5068 1616 5076 1624
rect 1116 1606 1118 1614
rect 1118 1606 1124 1614
rect 1132 1606 1140 1614
rect 1148 1606 1154 1614
rect 1154 1606 1156 1614
rect 4156 1606 4158 1614
rect 4158 1606 4164 1614
rect 4172 1606 4180 1614
rect 4188 1606 4194 1614
rect 4194 1606 4196 1614
rect 4588 1596 4596 1604
rect 5932 1596 5940 1604
rect 364 1576 372 1584
rect 4844 1556 4852 1564
rect 3564 1536 3572 1544
rect 5452 1536 5460 1544
rect 6828 1536 6836 1544
rect 5804 1516 5812 1524
rect 140 1496 148 1504
rect 524 1496 532 1504
rect 5452 1496 5460 1504
rect 5676 1496 5684 1504
rect 5836 1496 5844 1504
rect 6636 1516 6644 1524
rect 6220 1496 6228 1504
rect 172 1476 180 1484
rect 3052 1476 3060 1484
rect 1004 1456 1012 1464
rect 5932 1456 5940 1464
rect 5964 1456 5972 1464
rect 6572 1456 6580 1464
rect 1740 1436 1748 1444
rect 1772 1416 1780 1424
rect 2796 1416 2804 1424
rect 3756 1416 3764 1424
rect 2636 1406 2638 1414
rect 2638 1406 2644 1414
rect 2652 1406 2660 1414
rect 2668 1406 2674 1414
rect 2674 1406 2676 1414
rect 5724 1406 5726 1414
rect 5726 1406 5732 1414
rect 5740 1406 5748 1414
rect 5756 1406 5762 1414
rect 5762 1406 5764 1414
rect 1932 1396 1940 1404
rect 2860 1396 2868 1404
rect 3788 1376 3796 1384
rect 2956 1356 2964 1364
rect 5676 1356 5684 1364
rect 1228 1336 1236 1344
rect 2764 1336 2772 1344
rect 3052 1336 3060 1344
rect 5420 1336 5428 1344
rect 1004 1316 1012 1324
rect 1932 1316 1940 1324
rect 2732 1316 2740 1324
rect 4332 1316 4340 1324
rect 5068 1316 5076 1324
rect 5932 1316 5940 1324
rect 5964 1316 5972 1324
rect 6124 1316 6132 1324
rect 6668 1296 6676 1304
rect 1228 1276 1236 1284
rect 2764 1276 2772 1284
rect 5932 1276 5940 1284
rect 1036 1236 1044 1244
rect 4012 1236 4020 1244
rect 1116 1206 1118 1214
rect 1118 1206 1124 1214
rect 1132 1206 1140 1214
rect 1148 1206 1154 1214
rect 1154 1206 1156 1214
rect 4156 1206 4158 1214
rect 4158 1206 4164 1214
rect 4172 1206 4180 1214
rect 4188 1206 4194 1214
rect 4194 1206 4196 1214
rect 4492 1176 4500 1184
rect 3852 1156 3860 1164
rect 4428 1156 4436 1164
rect 5260 1156 5268 1164
rect 5804 1156 5812 1164
rect 6540 1156 6548 1164
rect 2380 1136 2388 1144
rect 3084 1136 3092 1144
rect 5836 1136 5844 1144
rect 6284 1136 6292 1144
rect 6348 1136 6356 1144
rect 364 1116 372 1124
rect 1260 1116 1268 1124
rect 1900 1116 1908 1124
rect 3212 1116 3220 1124
rect 5196 1116 5204 1124
rect 1932 1096 1940 1104
rect 3052 1096 3060 1104
rect 6348 1096 6356 1104
rect 5324 1076 5332 1084
rect 1004 1056 1012 1064
rect 1036 1056 1044 1064
rect 1580 1036 1588 1044
rect 5836 1036 5844 1044
rect 2636 1006 2638 1014
rect 2638 1006 2644 1014
rect 2652 1006 2660 1014
rect 2668 1006 2674 1014
rect 2674 1006 2676 1014
rect 5724 1006 5726 1014
rect 5726 1006 5732 1014
rect 5740 1006 5748 1014
rect 5756 1006 5762 1014
rect 5762 1006 5764 1014
rect 428 996 436 1004
rect 6092 996 6100 1004
rect 6412 996 6420 1004
rect 6828 996 6836 1004
rect 1004 956 1012 964
rect 2380 956 2388 964
rect 2956 956 2964 964
rect 4588 956 4596 964
rect 5036 956 5044 964
rect 5356 956 5364 964
rect 5836 956 5844 964
rect 6124 956 6132 964
rect 6572 956 6580 964
rect 300 936 308 944
rect 1356 936 1364 944
rect 2476 936 2484 944
rect 6508 936 6516 944
rect 4044 896 4052 904
rect 6348 916 6356 924
rect 1772 856 1780 864
rect 1356 836 1364 844
rect 6412 836 6420 844
rect 1116 806 1118 814
rect 1118 806 1124 814
rect 1132 806 1140 814
rect 1148 806 1154 814
rect 1154 806 1156 814
rect 3212 816 3220 824
rect 5676 816 5684 824
rect 4156 806 4158 814
rect 4158 806 4164 814
rect 4172 806 4180 814
rect 4188 806 4194 814
rect 4194 806 4196 814
rect 2604 796 2612 804
rect 1420 776 1428 784
rect 2380 776 2388 784
rect 6220 776 6228 784
rect 908 716 916 724
rect 1260 716 1268 724
rect 6796 736 6804 744
rect 1932 716 1940 724
rect 204 696 212 704
rect 2732 696 2740 704
rect 4492 696 4500 704
rect 5420 696 5428 704
rect 6540 696 6548 704
rect 1900 656 1908 664
rect 5580 656 5588 664
rect 6732 656 6740 664
rect 2764 636 2772 644
rect 5356 636 5364 644
rect 5996 616 6004 624
rect 2636 606 2638 614
rect 2638 606 2644 614
rect 2652 606 2660 614
rect 2668 606 2674 614
rect 2674 606 2676 614
rect 5724 606 5726 614
rect 5726 606 5732 614
rect 5740 606 5748 614
rect 5756 606 5762 614
rect 5762 606 5764 614
rect 5676 596 5684 604
rect 6124 596 6132 604
rect 6796 576 6804 584
rect 204 556 212 564
rect 1932 556 1940 564
rect 2476 556 2484 564
rect 300 536 308 544
rect 3276 536 3284 544
rect 4428 536 4436 544
rect 5804 536 5812 544
rect 1484 516 1492 524
rect 2156 516 2164 524
rect 5292 516 5300 524
rect 5580 516 5588 524
rect 6412 516 6420 524
rect 524 496 532 504
rect 908 496 916 504
rect 1420 496 1428 504
rect 5836 476 5844 484
rect 6860 476 6868 484
rect 6572 456 6580 464
rect 6732 436 6740 444
rect 1580 416 1588 424
rect 1116 406 1118 414
rect 1118 406 1124 414
rect 1132 406 1140 414
rect 1148 406 1154 414
rect 1154 406 1156 414
rect 4156 406 4158 414
rect 4158 406 4164 414
rect 4172 406 4180 414
rect 4188 406 4194 414
rect 4194 406 4196 414
rect 6636 336 6644 344
rect 5388 276 5396 284
rect 6764 276 6772 284
rect 6604 256 6612 264
rect 6732 236 6740 244
rect 2636 206 2638 214
rect 2638 206 2644 214
rect 2652 206 2660 214
rect 2668 206 2674 214
rect 2674 206 2676 214
rect 5724 206 5726 214
rect 5726 206 5732 214
rect 5740 206 5748 214
rect 5756 206 5762 214
rect 5762 206 5764 214
rect 6284 176 6292 184
rect 3276 136 3284 144
rect 4940 136 4948 144
rect 5388 136 5396 144
rect 6028 116 6036 124
rect 6828 116 6836 124
rect 2604 96 2612 104
rect 6796 96 6804 104
rect 2156 16 2164 24
rect 4940 16 4948 24
rect 1116 6 1118 14
rect 1118 6 1124 14
rect 1132 6 1140 14
rect 1148 6 1154 14
rect 1154 6 1156 14
rect 4156 6 4158 14
rect 4158 6 4164 14
rect 4172 6 4180 14
rect 4188 6 4194 14
rect 4194 6 4196 14
<< metal4 >>
rect 458 4904 470 4906
rect 458 4896 460 4904
rect 468 4896 470 4904
rect 426 4564 438 4566
rect 426 4556 428 4564
rect 436 4556 438 4564
rect 426 4364 438 4556
rect 426 4356 428 4364
rect 436 4356 438 4364
rect 426 4354 438 4356
rect 330 4324 342 4326
rect 330 4316 332 4324
rect 340 4316 342 4324
rect 298 4164 310 4166
rect 298 4156 300 4164
rect 308 4156 310 4164
rect 298 4004 310 4156
rect 298 3996 300 4004
rect 308 3996 310 4004
rect 298 3994 310 3996
rect 330 3864 342 4316
rect 330 3856 332 3864
rect 340 3856 342 3864
rect 330 3854 342 3856
rect 362 4304 374 4306
rect 362 4296 364 4304
rect 372 4296 374 4304
rect 362 3784 374 4296
rect 362 3776 364 3784
rect 372 3776 374 3784
rect 362 3774 374 3776
rect 170 3304 182 3306
rect 170 3296 172 3304
rect 180 3296 182 3304
rect 170 3064 182 3296
rect 458 3164 470 4896
rect 1112 4814 1160 5040
rect 2632 5014 2680 5040
rect 2632 5006 2636 5014
rect 2644 5006 2652 5014
rect 2660 5006 2668 5014
rect 2676 5006 2680 5014
rect 1112 4806 1116 4814
rect 1124 4806 1132 4814
rect 1140 4806 1148 4814
rect 1156 4806 1160 4814
rect 938 4684 950 4686
rect 938 4676 940 4684
rect 948 4676 950 4684
rect 650 4504 662 4506
rect 650 4496 652 4504
rect 660 4496 662 4504
rect 650 4204 662 4496
rect 874 4244 886 4246
rect 874 4236 876 4244
rect 884 4236 886 4244
rect 650 4196 652 4204
rect 660 4196 662 4204
rect 650 4194 662 4196
rect 778 4224 790 4226
rect 778 4216 780 4224
rect 788 4216 790 4224
rect 586 4184 598 4186
rect 586 4176 588 4184
rect 596 4176 598 4184
rect 586 3904 598 4176
rect 586 3896 588 3904
rect 596 3896 598 3904
rect 586 3894 598 3896
rect 618 4104 630 4106
rect 618 4096 620 4104
rect 628 4096 630 4104
rect 458 3156 460 3164
rect 468 3156 470 3164
rect 458 3154 470 3156
rect 170 3056 172 3064
rect 180 3056 182 3064
rect 170 2664 182 3056
rect 618 3064 630 4096
rect 650 4084 662 4086
rect 650 4076 652 4084
rect 660 4076 662 4084
rect 650 3884 662 4076
rect 650 3876 652 3884
rect 660 3876 662 3884
rect 650 3874 662 3876
rect 682 3984 694 3986
rect 682 3976 684 3984
rect 692 3976 694 3984
rect 682 3364 694 3976
rect 714 3964 726 3966
rect 714 3956 716 3964
rect 724 3956 726 3964
rect 714 3764 726 3956
rect 714 3756 716 3764
rect 724 3756 726 3764
rect 714 3754 726 3756
rect 778 3544 790 4216
rect 778 3536 780 3544
rect 788 3536 790 3544
rect 778 3534 790 3536
rect 682 3356 684 3364
rect 692 3356 694 3364
rect 682 3354 694 3356
rect 618 3056 620 3064
rect 628 3056 630 3064
rect 618 3054 630 3056
rect 874 2844 886 4236
rect 906 4204 918 4206
rect 906 4196 908 4204
rect 916 4196 918 4204
rect 906 3524 918 4196
rect 938 3724 950 4676
rect 1112 4414 1160 4806
rect 2250 5004 2262 5006
rect 2250 4996 2252 5004
rect 2260 4996 2262 5004
rect 1112 4406 1116 4414
rect 1124 4406 1132 4414
rect 1140 4406 1148 4414
rect 1156 4406 1160 4414
rect 1034 4204 1046 4206
rect 1034 4196 1036 4204
rect 1044 4196 1046 4204
rect 1034 3924 1046 4196
rect 1034 3916 1036 3924
rect 1044 3916 1046 3924
rect 1034 3914 1046 3916
rect 1112 4014 1160 4406
rect 1610 4644 1622 4646
rect 1610 4636 1612 4644
rect 1620 4636 1622 4644
rect 1610 4284 1622 4636
rect 1610 4276 1612 4284
rect 1620 4276 1622 4284
rect 1610 4274 1622 4276
rect 1642 4544 1654 4546
rect 1642 4536 1644 4544
rect 1652 4536 1654 4544
rect 1642 4244 1654 4536
rect 1642 4236 1644 4244
rect 1652 4236 1654 4244
rect 1642 4234 1654 4236
rect 1706 4544 1718 4546
rect 1706 4536 1708 4544
rect 1716 4536 1718 4544
rect 1706 4224 1718 4536
rect 1706 4216 1708 4224
rect 1716 4216 1718 4224
rect 1706 4164 1718 4216
rect 1706 4156 1708 4164
rect 1716 4156 1718 4164
rect 1706 4154 1718 4156
rect 1770 4124 1782 4126
rect 1770 4116 1772 4124
rect 1780 4116 1782 4124
rect 1112 4006 1116 4014
rect 1124 4006 1132 4014
rect 1140 4006 1148 4014
rect 1156 4006 1160 4014
rect 938 3716 940 3724
rect 948 3716 950 3724
rect 938 3714 950 3716
rect 906 3516 908 3524
rect 916 3516 918 3524
rect 906 3514 918 3516
rect 1112 3614 1160 4006
rect 1112 3606 1116 3614
rect 1124 3606 1132 3614
rect 1140 3606 1148 3614
rect 1156 3606 1160 3614
rect 938 3384 950 3386
rect 938 3376 940 3384
rect 948 3376 950 3384
rect 938 3224 950 3376
rect 938 3216 940 3224
rect 948 3216 950 3224
rect 938 3214 950 3216
rect 1112 3214 1160 3606
rect 1258 4064 1270 4066
rect 1258 4056 1260 4064
rect 1268 4056 1270 4064
rect 1258 3544 1270 4056
rect 1418 3944 1430 3946
rect 1418 3936 1420 3944
rect 1428 3936 1430 3944
rect 1258 3536 1260 3544
rect 1268 3536 1270 3544
rect 1258 3534 1270 3536
rect 1386 3884 1398 3886
rect 1386 3876 1388 3884
rect 1396 3876 1398 3884
rect 1386 3464 1398 3876
rect 1418 3864 1430 3936
rect 1770 3924 1782 4116
rect 1770 3916 1772 3924
rect 1780 3916 1782 3924
rect 1770 3914 1782 3916
rect 2026 3904 2038 3906
rect 2026 3896 2028 3904
rect 2036 3896 2038 3904
rect 1418 3856 1420 3864
rect 1428 3856 1430 3864
rect 1418 3854 1430 3856
rect 1514 3864 1526 3866
rect 1514 3856 1516 3864
rect 1524 3856 1526 3864
rect 1514 3584 1526 3856
rect 1514 3576 1516 3584
rect 1524 3576 1526 3584
rect 1514 3574 1526 3576
rect 1386 3456 1388 3464
rect 1396 3456 1398 3464
rect 1386 3454 1398 3456
rect 1674 3504 1686 3506
rect 1674 3496 1676 3504
rect 1684 3496 1686 3504
rect 1546 3384 1558 3386
rect 1546 3376 1548 3384
rect 1556 3376 1558 3384
rect 1546 3344 1558 3376
rect 1546 3336 1548 3344
rect 1556 3336 1558 3344
rect 1546 3334 1558 3336
rect 1674 3304 1686 3496
rect 1674 3296 1676 3304
rect 1684 3296 1686 3304
rect 1674 3294 1686 3296
rect 874 2836 876 2844
rect 884 2836 886 2844
rect 874 2834 886 2836
rect 1112 3206 1116 3214
rect 1124 3206 1132 3214
rect 1140 3206 1148 3214
rect 1156 3206 1160 3214
rect 170 2656 172 2664
rect 180 2656 182 2664
rect 170 2654 182 2656
rect 1112 2814 1160 3206
rect 1898 3184 1910 3186
rect 1898 3176 1900 3184
rect 1908 3176 1910 3184
rect 1112 2806 1116 2814
rect 1124 2806 1132 2814
rect 1140 2806 1148 2814
rect 1156 2806 1160 2814
rect 1066 2564 1078 2566
rect 1066 2556 1068 2564
rect 1076 2556 1078 2564
rect 1066 2164 1078 2556
rect 1066 2156 1068 2164
rect 1076 2156 1078 2164
rect 1066 2154 1078 2156
rect 1112 2414 1160 2806
rect 1866 3064 1878 3066
rect 1866 3056 1868 3064
rect 1876 3056 1878 3064
rect 1578 2784 1590 2786
rect 1578 2776 1580 2784
rect 1588 2776 1590 2784
rect 1112 2406 1116 2414
rect 1124 2406 1132 2414
rect 1140 2406 1148 2414
rect 1156 2406 1160 2414
rect 1112 2014 1160 2406
rect 1226 2604 1238 2606
rect 1226 2596 1228 2604
rect 1236 2596 1238 2604
rect 1226 2384 1238 2596
rect 1578 2564 1590 2776
rect 1866 2664 1878 3056
rect 1898 2984 1910 3176
rect 1898 2976 1900 2984
rect 1908 2976 1910 2984
rect 1898 2974 1910 2976
rect 1866 2656 1868 2664
rect 1876 2656 1878 2664
rect 1866 2654 1878 2656
rect 1578 2556 1580 2564
rect 1588 2556 1590 2564
rect 1578 2554 1590 2556
rect 1226 2376 1228 2384
rect 1236 2376 1238 2384
rect 1226 2374 1238 2376
rect 1578 2264 1590 2266
rect 1578 2256 1580 2264
rect 1588 2256 1590 2264
rect 1386 2224 1398 2226
rect 1386 2216 1388 2224
rect 1396 2216 1398 2224
rect 1386 2124 1398 2216
rect 1578 2184 1590 2256
rect 1578 2176 1580 2184
rect 1588 2176 1590 2184
rect 1578 2174 1590 2176
rect 1930 2264 1942 2266
rect 1930 2256 1932 2264
rect 1940 2256 1942 2264
rect 1386 2116 1388 2124
rect 1396 2116 1398 2124
rect 1386 2114 1398 2116
rect 1112 2006 1116 2014
rect 1124 2006 1132 2014
rect 1140 2006 1148 2014
rect 1156 2006 1160 2014
rect 906 1904 918 1906
rect 906 1896 908 1904
rect 916 1896 918 1904
rect 170 1884 182 1886
rect 170 1876 172 1884
rect 180 1876 182 1884
rect 138 1844 150 1846
rect 138 1836 140 1844
rect 148 1836 150 1844
rect 138 1504 150 1836
rect 138 1496 140 1504
rect 148 1496 150 1504
rect 138 1494 150 1496
rect 170 1824 182 1876
rect 170 1816 172 1824
rect 180 1816 182 1824
rect 170 1484 182 1816
rect 170 1476 172 1484
rect 180 1476 182 1484
rect 170 1474 182 1476
rect 298 1744 310 1746
rect 298 1736 300 1744
rect 308 1736 310 1744
rect 298 944 310 1736
rect 522 1704 534 1706
rect 522 1696 524 1704
rect 532 1696 534 1704
rect 426 1664 438 1666
rect 426 1656 428 1664
rect 436 1656 438 1664
rect 362 1584 374 1586
rect 362 1576 364 1584
rect 372 1576 374 1584
rect 362 1124 374 1576
rect 362 1116 364 1124
rect 372 1116 374 1124
rect 362 1114 374 1116
rect 426 1004 438 1656
rect 426 996 428 1004
rect 436 996 438 1004
rect 426 994 438 996
rect 522 1504 534 1696
rect 906 1644 918 1896
rect 906 1636 908 1644
rect 916 1636 918 1644
rect 906 1634 918 1636
rect 522 1496 524 1504
rect 532 1496 534 1504
rect 298 936 300 944
rect 308 936 310 944
rect 202 704 214 706
rect 202 696 204 704
rect 212 696 214 704
rect 202 564 214 696
rect 202 556 204 564
rect 212 556 214 564
rect 202 554 214 556
rect 298 544 310 936
rect 298 536 300 544
rect 308 536 310 544
rect 298 534 310 536
rect 522 504 534 1496
rect 1112 1614 1160 2006
rect 1738 1844 1750 1846
rect 1738 1836 1740 1844
rect 1748 1836 1750 1844
rect 1578 1724 1590 1726
rect 1578 1716 1580 1724
rect 1588 1716 1590 1724
rect 1112 1606 1116 1614
rect 1124 1606 1132 1614
rect 1140 1606 1148 1614
rect 1156 1606 1160 1614
rect 1002 1464 1014 1466
rect 1002 1456 1004 1464
rect 1012 1456 1014 1464
rect 1002 1324 1014 1456
rect 1002 1316 1004 1324
rect 1012 1316 1014 1324
rect 1002 1314 1014 1316
rect 1034 1244 1046 1246
rect 1034 1236 1036 1244
rect 1044 1236 1046 1244
rect 1002 1064 1014 1066
rect 1002 1056 1004 1064
rect 1012 1056 1014 1064
rect 1002 964 1014 1056
rect 1034 1064 1046 1236
rect 1034 1056 1036 1064
rect 1044 1056 1046 1064
rect 1034 1054 1046 1056
rect 1112 1214 1160 1606
rect 1482 1644 1494 1646
rect 1482 1636 1484 1644
rect 1492 1636 1494 1644
rect 1226 1344 1238 1346
rect 1226 1336 1228 1344
rect 1236 1336 1238 1344
rect 1226 1284 1238 1336
rect 1226 1276 1228 1284
rect 1236 1276 1238 1284
rect 1226 1274 1238 1276
rect 1112 1206 1116 1214
rect 1124 1206 1132 1214
rect 1140 1206 1148 1214
rect 1156 1206 1160 1214
rect 1002 956 1004 964
rect 1012 956 1014 964
rect 1002 954 1014 956
rect 1112 814 1160 1206
rect 1112 806 1116 814
rect 1124 806 1132 814
rect 1140 806 1148 814
rect 1156 806 1160 814
rect 522 496 524 504
rect 532 496 534 504
rect 522 494 534 496
rect 906 724 918 726
rect 906 716 908 724
rect 916 716 918 724
rect 906 504 918 716
rect 906 496 908 504
rect 916 496 918 504
rect 906 494 918 496
rect 1112 414 1160 806
rect 1258 1124 1270 1126
rect 1258 1116 1260 1124
rect 1268 1116 1270 1124
rect 1258 724 1270 1116
rect 1354 944 1366 946
rect 1354 936 1356 944
rect 1364 936 1366 944
rect 1354 844 1366 936
rect 1354 836 1356 844
rect 1364 836 1366 844
rect 1354 834 1366 836
rect 1258 716 1260 724
rect 1268 716 1270 724
rect 1258 714 1270 716
rect 1418 784 1430 786
rect 1418 776 1420 784
rect 1428 776 1430 784
rect 1418 504 1430 776
rect 1482 524 1494 1636
rect 1482 516 1484 524
rect 1492 516 1494 524
rect 1482 514 1494 516
rect 1578 1044 1590 1716
rect 1738 1444 1750 1836
rect 1738 1436 1740 1444
rect 1748 1436 1750 1444
rect 1738 1434 1750 1436
rect 1930 1664 1942 2256
rect 2026 1744 2038 3896
rect 2250 3824 2262 4996
rect 2632 4614 2680 5006
rect 4152 4814 4200 5040
rect 5720 5014 5768 5040
rect 5720 5006 5724 5014
rect 5732 5006 5740 5014
rect 5748 5006 5756 5014
rect 5764 5006 5768 5014
rect 4152 4806 4156 4814
rect 4164 4806 4172 4814
rect 4180 4806 4188 4814
rect 4196 4806 4200 4814
rect 2632 4606 2636 4614
rect 2644 4606 2652 4614
rect 2660 4606 2668 4614
rect 2676 4606 2680 4614
rect 2632 4214 2680 4606
rect 2762 4724 2774 4726
rect 2762 4716 2764 4724
rect 2772 4716 2774 4724
rect 2762 4444 2774 4716
rect 3978 4724 3990 4726
rect 3978 4716 3980 4724
rect 3988 4716 3990 4724
rect 3434 4664 3446 4666
rect 3434 4656 3436 4664
rect 3444 4656 3446 4664
rect 2762 4436 2764 4444
rect 2772 4436 2774 4444
rect 2762 4434 2774 4436
rect 2954 4604 2966 4606
rect 2954 4596 2956 4604
rect 2964 4596 2966 4604
rect 2632 4206 2636 4214
rect 2644 4206 2652 4214
rect 2660 4206 2668 4214
rect 2676 4206 2680 4214
rect 2730 4284 2742 4286
rect 2730 4276 2732 4284
rect 2740 4276 2742 4284
rect 2250 3816 2252 3824
rect 2260 3816 2262 3824
rect 2250 3814 2262 3816
rect 2410 3864 2422 3866
rect 2410 3856 2412 3864
rect 2420 3856 2422 3864
rect 2122 3804 2134 3806
rect 2122 3796 2124 3804
rect 2132 3796 2134 3804
rect 2122 3324 2134 3796
rect 2410 3384 2422 3856
rect 2410 3376 2412 3384
rect 2420 3376 2422 3384
rect 2410 3374 2422 3376
rect 2570 3824 2582 3826
rect 2570 3816 2572 3824
rect 2580 3816 2582 3824
rect 2122 3316 2124 3324
rect 2132 3316 2134 3324
rect 2122 3314 2134 3316
rect 2570 3084 2582 3816
rect 2570 3076 2572 3084
rect 2580 3076 2582 3084
rect 2570 3074 2582 3076
rect 2632 3814 2680 4206
rect 2632 3806 2636 3814
rect 2644 3806 2652 3814
rect 2660 3806 2668 3814
rect 2676 3806 2680 3814
rect 2632 3414 2680 3806
rect 2698 4204 2710 4206
rect 2698 4196 2700 4204
rect 2708 4196 2710 4204
rect 2698 3464 2710 4196
rect 2730 3544 2742 4276
rect 2954 4284 2966 4596
rect 2954 4276 2956 4284
rect 2964 4276 2966 4284
rect 2922 4184 2934 4186
rect 2922 4176 2924 4184
rect 2932 4176 2934 4184
rect 2858 4044 2870 4046
rect 2858 4036 2860 4044
rect 2868 4036 2870 4044
rect 2858 3724 2870 4036
rect 2922 3764 2934 4176
rect 2954 3824 2966 4276
rect 3050 4564 3062 4566
rect 3050 4556 3052 4564
rect 3060 4556 3062 4564
rect 3050 4284 3062 4556
rect 3050 4276 3052 4284
rect 3060 4276 3062 4284
rect 3050 4274 3062 4276
rect 3338 4304 3350 4306
rect 3338 4296 3340 4304
rect 3348 4296 3350 4304
rect 3338 4204 3350 4296
rect 3434 4224 3446 4656
rect 3818 4664 3830 4666
rect 3818 4656 3820 4664
rect 3828 4656 3830 4664
rect 3690 4524 3702 4526
rect 3690 4516 3692 4524
rect 3700 4516 3702 4524
rect 3466 4384 3478 4386
rect 3466 4376 3468 4384
rect 3476 4376 3478 4384
rect 3466 4244 3478 4376
rect 3466 4236 3468 4244
rect 3476 4236 3478 4244
rect 3466 4234 3478 4236
rect 3658 4384 3670 4386
rect 3658 4376 3660 4384
rect 3668 4376 3670 4384
rect 3434 4216 3436 4224
rect 3444 4216 3446 4224
rect 3434 4214 3446 4216
rect 3338 4196 3340 4204
rect 3348 4196 3350 4204
rect 3338 4194 3350 4196
rect 3242 4164 3254 4166
rect 3242 4156 3244 4164
rect 3252 4156 3254 4164
rect 3146 4064 3158 4066
rect 3146 4056 3148 4064
rect 3156 4056 3158 4064
rect 2954 3816 2956 3824
rect 2964 3816 2966 3824
rect 2954 3814 2966 3816
rect 3018 3884 3030 3886
rect 3018 3876 3020 3884
rect 3028 3876 3030 3884
rect 2922 3756 2924 3764
rect 2932 3756 2934 3764
rect 2922 3754 2934 3756
rect 2858 3716 2860 3724
rect 2868 3716 2870 3724
rect 2858 3714 2870 3716
rect 2730 3536 2732 3544
rect 2740 3536 2742 3544
rect 2730 3534 2742 3536
rect 3018 3524 3030 3876
rect 3146 3564 3158 4056
rect 3146 3556 3148 3564
rect 3156 3556 3158 3564
rect 3146 3554 3158 3556
rect 3178 3824 3190 3826
rect 3178 3816 3180 3824
rect 3188 3816 3190 3824
rect 3018 3516 3020 3524
rect 3028 3516 3030 3524
rect 3018 3514 3030 3516
rect 3114 3544 3126 3546
rect 3114 3536 3116 3544
rect 3124 3536 3126 3544
rect 2698 3456 2700 3464
rect 2708 3456 2710 3464
rect 2698 3454 2710 3456
rect 2632 3406 2636 3414
rect 2644 3406 2652 3414
rect 2660 3406 2668 3414
rect 2676 3406 2680 3414
rect 2154 3044 2166 3046
rect 2154 3036 2156 3044
rect 2164 3036 2166 3044
rect 2154 2844 2166 3036
rect 2154 2836 2156 2844
rect 2164 2836 2166 2844
rect 2154 2834 2166 2836
rect 2632 3014 2680 3406
rect 2794 3124 2806 3126
rect 2794 3116 2796 3124
rect 2804 3116 2806 3124
rect 2632 3006 2636 3014
rect 2644 3006 2652 3014
rect 2660 3006 2668 3014
rect 2676 3006 2680 3014
rect 2378 2784 2390 2786
rect 2378 2776 2380 2784
rect 2388 2776 2390 2784
rect 2378 2324 2390 2776
rect 2632 2614 2680 3006
rect 2762 3084 2774 3086
rect 2762 3076 2764 3084
rect 2772 3076 2774 3084
rect 2632 2606 2636 2614
rect 2644 2606 2652 2614
rect 2660 2606 2668 2614
rect 2676 2606 2680 2614
rect 2378 2316 2380 2324
rect 2388 2316 2390 2324
rect 2378 2314 2390 2316
rect 2602 2444 2614 2446
rect 2602 2436 2604 2444
rect 2612 2436 2614 2444
rect 2602 2164 2614 2436
rect 2602 2156 2604 2164
rect 2612 2156 2614 2164
rect 2602 2154 2614 2156
rect 2632 2214 2680 2606
rect 2632 2206 2636 2214
rect 2644 2206 2652 2214
rect 2660 2206 2668 2214
rect 2676 2206 2680 2214
rect 2026 1736 2028 1744
rect 2036 1736 2038 1744
rect 2026 1734 2038 1736
rect 2632 1814 2680 2206
rect 2730 2684 2742 2686
rect 2730 2676 2732 2684
rect 2740 2676 2742 2684
rect 2730 2224 2742 2676
rect 2730 2216 2732 2224
rect 2740 2216 2742 2224
rect 2730 2124 2742 2216
rect 2730 2116 2732 2124
rect 2740 2116 2742 2124
rect 2730 2114 2742 2116
rect 2632 1806 2636 1814
rect 2644 1806 2652 1814
rect 2660 1806 2668 1814
rect 2676 1806 2680 1814
rect 1930 1656 1932 1664
rect 1940 1656 1942 1664
rect 1578 1036 1580 1044
rect 1588 1036 1590 1044
rect 1418 496 1420 504
rect 1428 496 1430 504
rect 1418 494 1430 496
rect 1578 424 1590 1036
rect 1770 1424 1782 1426
rect 1770 1416 1772 1424
rect 1780 1416 1782 1424
rect 1770 864 1782 1416
rect 1930 1404 1942 1656
rect 1930 1396 1932 1404
rect 1940 1396 1942 1404
rect 1930 1394 1942 1396
rect 2632 1414 2680 1806
rect 2632 1406 2636 1414
rect 2644 1406 2652 1414
rect 2660 1406 2668 1414
rect 2676 1406 2680 1414
rect 1930 1324 1942 1326
rect 1930 1316 1932 1324
rect 1940 1316 1942 1324
rect 1770 856 1772 864
rect 1780 856 1782 864
rect 1770 854 1782 856
rect 1898 1124 1910 1126
rect 1898 1116 1900 1124
rect 1908 1116 1910 1124
rect 1898 664 1910 1116
rect 1930 1104 1942 1316
rect 1930 1096 1932 1104
rect 1940 1096 1942 1104
rect 1930 1094 1942 1096
rect 2378 1144 2390 1146
rect 2378 1136 2380 1144
rect 2388 1136 2390 1144
rect 2378 964 2390 1136
rect 2378 956 2380 964
rect 2388 956 2390 964
rect 2378 784 2390 956
rect 2632 1014 2680 1406
rect 2762 1344 2774 3076
rect 2794 2944 2806 3116
rect 3114 3124 3126 3536
rect 3178 3524 3190 3816
rect 3178 3516 3180 3524
rect 3188 3516 3190 3524
rect 3178 3514 3190 3516
rect 3210 3784 3222 3786
rect 3210 3776 3212 3784
rect 3220 3776 3222 3784
rect 3210 3404 3222 3776
rect 3242 3664 3254 4156
rect 3242 3656 3244 3664
rect 3252 3656 3254 3664
rect 3242 3654 3254 3656
rect 3274 4124 3286 4126
rect 3274 4116 3276 4124
rect 3284 4116 3286 4124
rect 3274 3544 3286 4116
rect 3594 4124 3606 4126
rect 3594 4116 3596 4124
rect 3604 4116 3606 4124
rect 3402 4044 3414 4046
rect 3402 4036 3404 4044
rect 3412 4036 3414 4044
rect 3402 3724 3414 4036
rect 3594 3884 3606 4116
rect 3658 4044 3670 4376
rect 3690 4364 3702 4516
rect 3690 4356 3692 4364
rect 3700 4356 3702 4364
rect 3690 4354 3702 4356
rect 3818 4364 3830 4656
rect 3818 4356 3820 4364
rect 3828 4356 3830 4364
rect 3818 4354 3830 4356
rect 3882 4524 3894 4526
rect 3882 4516 3884 4524
rect 3892 4516 3894 4524
rect 3722 4344 3734 4346
rect 3722 4336 3724 4344
rect 3732 4336 3734 4344
rect 3722 4084 3734 4336
rect 3722 4076 3724 4084
rect 3732 4076 3734 4084
rect 3722 4074 3734 4076
rect 3850 4284 3862 4286
rect 3850 4276 3852 4284
rect 3860 4276 3862 4284
rect 3850 4084 3862 4276
rect 3850 4076 3852 4084
rect 3860 4076 3862 4084
rect 3850 4074 3862 4076
rect 3882 4244 3894 4516
rect 3978 4264 3990 4716
rect 3978 4256 3980 4264
rect 3988 4256 3990 4264
rect 3978 4254 3990 4256
rect 4152 4414 4200 4806
rect 4842 5004 4854 5006
rect 4842 4996 4844 5004
rect 4852 4996 4854 5004
rect 4842 4624 4854 4996
rect 5514 5004 5526 5006
rect 5514 4996 5516 5004
rect 5524 4996 5526 5004
rect 4842 4616 4844 4624
rect 4852 4616 4854 4624
rect 4842 4614 4854 4616
rect 5482 4844 5494 4846
rect 5482 4836 5484 4844
rect 5492 4836 5494 4844
rect 4152 4406 4156 4414
rect 4164 4406 4172 4414
rect 4180 4406 4188 4414
rect 4196 4406 4200 4414
rect 3882 4236 3884 4244
rect 3892 4236 3894 4244
rect 3882 4124 3894 4236
rect 3882 4116 3884 4124
rect 3892 4116 3894 4124
rect 3658 4036 3660 4044
rect 3668 4036 3670 4044
rect 3658 4034 3670 4036
rect 3594 3876 3596 3884
rect 3604 3876 3606 3884
rect 3594 3874 3606 3876
rect 3626 3944 3638 3946
rect 3626 3936 3628 3944
rect 3636 3936 3638 3944
rect 3466 3864 3478 3866
rect 3466 3856 3468 3864
rect 3476 3856 3478 3864
rect 3402 3716 3404 3724
rect 3412 3716 3414 3724
rect 3402 3714 3414 3716
rect 3434 3744 3446 3746
rect 3434 3736 3436 3744
rect 3444 3736 3446 3744
rect 3338 3584 3350 3586
rect 3338 3576 3340 3584
rect 3348 3576 3350 3584
rect 3274 3536 3276 3544
rect 3284 3536 3286 3544
rect 3274 3534 3286 3536
rect 3306 3544 3318 3546
rect 3306 3536 3308 3544
rect 3316 3536 3318 3544
rect 3210 3396 3212 3404
rect 3220 3396 3222 3404
rect 3210 3394 3222 3396
rect 3306 3344 3318 3536
rect 3338 3444 3350 3576
rect 3338 3436 3340 3444
rect 3348 3436 3350 3444
rect 3338 3434 3350 3436
rect 3306 3336 3308 3344
rect 3316 3336 3318 3344
rect 3306 3334 3318 3336
rect 3114 3116 3116 3124
rect 3124 3116 3126 3124
rect 3114 3114 3126 3116
rect 3370 3184 3382 3186
rect 3370 3176 3372 3184
rect 3380 3176 3382 3184
rect 2794 2936 2796 2944
rect 2804 2936 2806 2944
rect 2794 2934 2806 2936
rect 3146 2764 3158 2766
rect 3146 2756 3148 2764
rect 3156 2756 3158 2764
rect 2922 2724 2934 2726
rect 2922 2716 2924 2724
rect 2932 2716 2934 2724
rect 2858 2684 2870 2686
rect 2858 2676 2860 2684
rect 2868 2676 2870 2684
rect 2858 2424 2870 2676
rect 2858 2416 2860 2424
rect 2868 2416 2870 2424
rect 2858 2414 2870 2416
rect 2890 2504 2902 2506
rect 2890 2496 2892 2504
rect 2900 2496 2902 2504
rect 2858 2264 2870 2266
rect 2858 2256 2860 2264
rect 2868 2256 2870 2264
rect 2794 1744 2806 1746
rect 2794 1736 2796 1744
rect 2804 1736 2806 1744
rect 2794 1424 2806 1736
rect 2794 1416 2796 1424
rect 2804 1416 2806 1424
rect 2794 1414 2806 1416
rect 2858 1404 2870 2256
rect 2890 2164 2902 2496
rect 2922 2464 2934 2716
rect 2922 2456 2924 2464
rect 2932 2456 2934 2464
rect 2922 2454 2934 2456
rect 2954 2604 2966 2606
rect 2954 2596 2956 2604
rect 2964 2596 2966 2604
rect 2954 2424 2966 2596
rect 3146 2524 3158 2756
rect 3146 2516 3148 2524
rect 3156 2516 3158 2524
rect 3146 2514 3158 2516
rect 3306 2544 3318 2546
rect 3306 2536 3308 2544
rect 3316 2536 3318 2544
rect 2954 2416 2956 2424
rect 2964 2416 2966 2424
rect 2954 2414 2966 2416
rect 3210 2484 3222 2486
rect 3210 2476 3212 2484
rect 3220 2476 3222 2484
rect 2890 2156 2892 2164
rect 2900 2156 2902 2164
rect 2890 2154 2902 2156
rect 3210 2144 3222 2476
rect 3242 2484 3254 2486
rect 3242 2476 3244 2484
rect 3252 2476 3254 2484
rect 3242 2264 3254 2476
rect 3242 2256 3244 2264
rect 3252 2256 3254 2264
rect 3242 2254 3254 2256
rect 3274 2464 3286 2466
rect 3274 2456 3276 2464
rect 3284 2456 3286 2464
rect 3274 2344 3286 2456
rect 3306 2364 3318 2536
rect 3370 2544 3382 3176
rect 3434 3084 3446 3736
rect 3466 3564 3478 3856
rect 3626 3724 3638 3936
rect 3626 3716 3628 3724
rect 3636 3716 3638 3724
rect 3626 3714 3638 3716
rect 3658 3804 3670 3806
rect 3658 3796 3660 3804
rect 3668 3796 3670 3804
rect 3466 3556 3468 3564
rect 3476 3556 3478 3564
rect 3466 3554 3478 3556
rect 3498 3584 3510 3586
rect 3498 3576 3500 3584
rect 3508 3576 3510 3584
rect 3434 3076 3436 3084
rect 3444 3076 3446 3084
rect 3370 2536 3372 2544
rect 3380 2536 3382 2544
rect 3370 2444 3382 2536
rect 3370 2436 3372 2444
rect 3380 2436 3382 2444
rect 3370 2434 3382 2436
rect 3402 2724 3414 2726
rect 3402 2716 3404 2724
rect 3412 2716 3414 2724
rect 3402 2584 3414 2716
rect 3434 2684 3446 3076
rect 3434 2676 3436 2684
rect 3444 2676 3446 2684
rect 3434 2674 3446 2676
rect 3466 3444 3478 3446
rect 3466 3436 3468 3444
rect 3476 3436 3478 3444
rect 3402 2576 3404 2584
rect 3412 2576 3414 2584
rect 3402 2424 3414 2576
rect 3402 2416 3404 2424
rect 3412 2416 3414 2424
rect 3402 2414 3414 2416
rect 3306 2356 3308 2364
rect 3316 2356 3318 2364
rect 3306 2354 3318 2356
rect 3274 2336 3276 2344
rect 3284 2336 3286 2344
rect 3210 2136 3212 2144
rect 3220 2136 3222 2144
rect 3210 2134 3222 2136
rect 3274 2124 3286 2336
rect 3274 2116 3276 2124
rect 3284 2116 3286 2124
rect 3274 2114 3286 2116
rect 3434 2244 3446 2246
rect 3434 2236 3436 2244
rect 3444 2236 3446 2244
rect 3082 1864 3094 1866
rect 3082 1856 3084 1864
rect 3092 1856 3094 1864
rect 2858 1396 2860 1404
rect 2868 1396 2870 1404
rect 2858 1394 2870 1396
rect 3050 1484 3062 1486
rect 3050 1476 3052 1484
rect 3060 1476 3062 1484
rect 2762 1336 2764 1344
rect 2772 1336 2774 1344
rect 2762 1334 2774 1336
rect 2954 1364 2966 1366
rect 2954 1356 2956 1364
rect 2964 1356 2966 1364
rect 2632 1006 2636 1014
rect 2644 1006 2652 1014
rect 2660 1006 2668 1014
rect 2676 1006 2680 1014
rect 2378 776 2380 784
rect 2388 776 2390 784
rect 2378 774 2390 776
rect 2474 944 2486 946
rect 2474 936 2476 944
rect 2484 936 2486 944
rect 1898 656 1900 664
rect 1908 656 1910 664
rect 1898 654 1910 656
rect 1930 724 1942 726
rect 1930 716 1932 724
rect 1940 716 1942 724
rect 1930 564 1942 716
rect 1930 556 1932 564
rect 1940 556 1942 564
rect 1930 554 1942 556
rect 2474 564 2486 936
rect 2474 556 2476 564
rect 2484 556 2486 564
rect 2474 554 2486 556
rect 2602 804 2614 806
rect 2602 796 2604 804
rect 2612 796 2614 804
rect 1578 416 1580 424
rect 1588 416 1590 424
rect 1578 414 1590 416
rect 2154 524 2166 526
rect 2154 516 2156 524
rect 2164 516 2166 524
rect 1112 406 1116 414
rect 1124 406 1132 414
rect 1140 406 1148 414
rect 1156 406 1160 414
rect 1112 14 1160 406
rect 2154 24 2166 516
rect 2602 104 2614 796
rect 2602 96 2604 104
rect 2612 96 2614 104
rect 2602 94 2614 96
rect 2632 614 2680 1006
rect 2730 1324 2742 1326
rect 2730 1316 2732 1324
rect 2740 1316 2742 1324
rect 2730 704 2742 1316
rect 2730 696 2732 704
rect 2740 696 2742 704
rect 2730 694 2742 696
rect 2762 1284 2774 1286
rect 2762 1276 2764 1284
rect 2772 1276 2774 1284
rect 2762 644 2774 1276
rect 2954 964 2966 1356
rect 3050 1344 3062 1476
rect 3050 1336 3052 1344
rect 3060 1336 3062 1344
rect 3050 1104 3062 1336
rect 3082 1144 3094 1856
rect 3434 1704 3446 2236
rect 3466 1744 3478 3436
rect 3498 3224 3510 3576
rect 3658 3584 3670 3796
rect 3850 3704 3862 3706
rect 3850 3696 3852 3704
rect 3860 3696 3862 3704
rect 3658 3576 3660 3584
rect 3668 3576 3670 3584
rect 3658 3574 3670 3576
rect 3754 3624 3766 3626
rect 3754 3616 3756 3624
rect 3764 3616 3766 3624
rect 3498 3216 3500 3224
rect 3508 3216 3510 3224
rect 3498 3214 3510 3216
rect 3562 3504 3574 3506
rect 3562 3496 3564 3504
rect 3572 3496 3574 3504
rect 3562 3304 3574 3496
rect 3562 3296 3564 3304
rect 3572 3296 3574 3304
rect 3530 3064 3542 3066
rect 3530 3056 3532 3064
rect 3540 3056 3542 3064
rect 3498 2804 3510 2806
rect 3498 2796 3500 2804
rect 3508 2796 3510 2804
rect 3498 2584 3510 2796
rect 3530 2664 3542 3056
rect 3530 2656 3532 2664
rect 3540 2656 3542 2664
rect 3530 2654 3542 2656
rect 3562 2664 3574 3296
rect 3658 3464 3670 3466
rect 3658 3456 3660 3464
rect 3668 3456 3670 3464
rect 3594 3084 3606 3086
rect 3594 3076 3596 3084
rect 3604 3076 3606 3084
rect 3594 2724 3606 3076
rect 3658 2764 3670 3456
rect 3754 3184 3766 3616
rect 3754 3176 3756 3184
rect 3764 3176 3766 3184
rect 3754 3174 3766 3176
rect 3850 3244 3862 3696
rect 3850 3236 3852 3244
rect 3860 3236 3862 3244
rect 3786 2924 3798 2926
rect 3786 2916 3788 2924
rect 3796 2916 3798 2924
rect 3658 2756 3660 2764
rect 3668 2756 3670 2764
rect 3658 2754 3670 2756
rect 3722 2864 3734 2866
rect 3722 2856 3724 2864
rect 3732 2856 3734 2864
rect 3594 2716 3596 2724
rect 3604 2716 3606 2724
rect 3594 2714 3606 2716
rect 3562 2656 3564 2664
rect 3572 2656 3574 2664
rect 3498 2576 3500 2584
rect 3508 2576 3510 2584
rect 3498 2574 3510 2576
rect 3466 1736 3468 1744
rect 3476 1736 3478 1744
rect 3466 1734 3478 1736
rect 3434 1696 3436 1704
rect 3444 1696 3446 1704
rect 3434 1694 3446 1696
rect 3562 1544 3574 2656
rect 3690 2604 3702 2606
rect 3690 2596 3692 2604
rect 3700 2596 3702 2604
rect 3690 2364 3702 2596
rect 3690 2356 3692 2364
rect 3700 2356 3702 2364
rect 3690 2354 3702 2356
rect 3722 2224 3734 2856
rect 3754 2704 3766 2706
rect 3754 2696 3756 2704
rect 3764 2696 3766 2704
rect 3754 2664 3766 2696
rect 3754 2656 3756 2664
rect 3764 2656 3766 2664
rect 3754 2654 3766 2656
rect 3722 2216 3724 2224
rect 3732 2216 3734 2224
rect 3722 2214 3734 2216
rect 3754 2244 3766 2246
rect 3754 2236 3756 2244
rect 3764 2236 3766 2244
rect 3754 1984 3766 2236
rect 3754 1976 3756 1984
rect 3764 1976 3766 1984
rect 3754 1974 3766 1976
rect 3562 1536 3564 1544
rect 3572 1536 3574 1544
rect 3562 1534 3574 1536
rect 3754 1944 3766 1946
rect 3754 1936 3756 1944
rect 3764 1936 3766 1944
rect 3754 1424 3766 1936
rect 3754 1416 3756 1424
rect 3764 1416 3766 1424
rect 3754 1414 3766 1416
rect 3786 1384 3798 2916
rect 3818 2764 3830 2766
rect 3818 2756 3820 2764
rect 3828 2756 3830 2764
rect 3818 1984 3830 2756
rect 3850 2704 3862 3236
rect 3850 2696 3852 2704
rect 3860 2696 3862 2704
rect 3850 2694 3862 2696
rect 3818 1976 3820 1984
rect 3828 1976 3830 1984
rect 3818 1974 3830 1976
rect 3850 2284 3862 2286
rect 3850 2276 3852 2284
rect 3860 2276 3862 2284
rect 3786 1376 3788 1384
rect 3796 1376 3798 1384
rect 3786 1374 3798 1376
rect 3850 1164 3862 2276
rect 3882 2144 3894 4116
rect 3914 4164 3926 4166
rect 3914 4156 3916 4164
rect 3924 4156 3926 4164
rect 3914 3364 3926 4156
rect 3978 4144 3990 4146
rect 3978 4136 3980 4144
rect 3988 4136 3990 4144
rect 3978 3824 3990 4136
rect 3978 3816 3980 3824
rect 3988 3816 3990 3824
rect 3978 3814 3990 3816
rect 4152 4014 4200 4406
rect 4152 4006 4156 4014
rect 4164 4006 4172 4014
rect 4180 4006 4188 4014
rect 4196 4006 4200 4014
rect 3914 3356 3916 3364
rect 3924 3356 3926 3364
rect 3914 3354 3926 3356
rect 4106 3684 4118 3686
rect 4106 3676 4108 3684
rect 4116 3676 4118 3684
rect 4042 2924 4054 2926
rect 4042 2916 4044 2924
rect 4052 2916 4054 2924
rect 3882 2136 3884 2144
rect 3892 2136 3894 2144
rect 3882 2134 3894 2136
rect 3914 2524 3926 2526
rect 3914 2516 3916 2524
rect 3924 2516 3926 2524
rect 3914 2124 3926 2516
rect 4042 2204 4054 2916
rect 4106 2744 4118 3676
rect 4106 2736 4108 2744
rect 4116 2736 4118 2744
rect 4106 2734 4118 2736
rect 4152 3614 4200 4006
rect 4778 4504 4790 4506
rect 4778 4496 4780 4504
rect 4788 4496 4790 4504
rect 4778 3964 4790 4496
rect 5322 4324 5334 4326
rect 5322 4316 5324 4324
rect 5332 4316 5334 4324
rect 5066 4284 5078 4286
rect 5066 4276 5068 4284
rect 5076 4276 5078 4284
rect 4778 3956 4780 3964
rect 4788 3956 4790 3964
rect 4778 3954 4790 3956
rect 4810 3964 4822 3966
rect 4810 3956 4812 3964
rect 4820 3956 4822 3964
rect 4152 3606 4156 3614
rect 4164 3606 4172 3614
rect 4180 3606 4188 3614
rect 4196 3606 4200 3614
rect 4152 3214 4200 3606
rect 4298 3884 4310 3886
rect 4298 3876 4300 3884
rect 4308 3876 4310 3884
rect 4298 3484 4310 3876
rect 4298 3476 4300 3484
rect 4308 3476 4310 3484
rect 4298 3474 4310 3476
rect 4778 3484 4790 3486
rect 4778 3476 4780 3484
rect 4788 3476 4790 3484
rect 4152 3206 4156 3214
rect 4164 3206 4172 3214
rect 4180 3206 4188 3214
rect 4196 3206 4200 3214
rect 4152 2814 4200 3206
rect 4152 2806 4156 2814
rect 4164 2806 4172 2814
rect 4180 2806 4188 2814
rect 4196 2806 4200 2814
rect 4152 2414 4200 2806
rect 4266 3304 4278 3306
rect 4266 3296 4268 3304
rect 4276 3296 4278 3304
rect 4266 2504 4278 3296
rect 4714 3304 4726 3306
rect 4714 3296 4716 3304
rect 4724 3296 4726 3304
rect 4362 2964 4374 2966
rect 4362 2956 4364 2964
rect 4372 2956 4374 2964
rect 4362 2564 4374 2956
rect 4554 2964 4566 2966
rect 4554 2956 4556 2964
rect 4564 2956 4566 2964
rect 4554 2664 4566 2956
rect 4714 2904 4726 3296
rect 4778 3284 4790 3476
rect 4810 3364 4822 3956
rect 5066 3904 5078 4276
rect 5322 4044 5334 4316
rect 5322 4036 5324 4044
rect 5332 4036 5334 4044
rect 5322 4034 5334 4036
rect 5354 4284 5366 4286
rect 5354 4276 5356 4284
rect 5364 4276 5366 4284
rect 5066 3896 5068 3904
rect 5076 3896 5078 3904
rect 5066 3894 5078 3896
rect 5194 3944 5206 3946
rect 5194 3936 5196 3944
rect 5204 3936 5206 3944
rect 5194 3864 5206 3936
rect 5194 3856 5196 3864
rect 5204 3856 5206 3864
rect 5194 3854 5206 3856
rect 5354 3864 5366 4276
rect 5354 3856 5356 3864
rect 5364 3856 5366 3864
rect 5354 3854 5366 3856
rect 5418 4264 5430 4266
rect 5418 4256 5420 4264
rect 5428 4256 5430 4264
rect 5418 4104 5430 4256
rect 5418 4096 5420 4104
rect 5428 4096 5430 4104
rect 4938 3844 4950 3846
rect 4938 3836 4940 3844
rect 4948 3836 4950 3844
rect 4810 3356 4812 3364
rect 4820 3356 4822 3364
rect 4810 3354 4822 3356
rect 4906 3804 4918 3806
rect 4906 3796 4908 3804
rect 4916 3796 4918 3804
rect 4778 3276 4780 3284
rect 4788 3276 4790 3284
rect 4778 3274 4790 3276
rect 4714 2896 4716 2904
rect 4724 2896 4726 2904
rect 4714 2894 4726 2896
rect 4554 2656 4556 2664
rect 4564 2656 4566 2664
rect 4362 2556 4364 2564
rect 4372 2556 4374 2564
rect 4362 2554 4374 2556
rect 4458 2584 4470 2586
rect 4458 2576 4460 2584
rect 4468 2576 4470 2584
rect 4266 2496 4268 2504
rect 4276 2496 4278 2504
rect 4266 2494 4278 2496
rect 4152 2406 4156 2414
rect 4164 2406 4172 2414
rect 4180 2406 4188 2414
rect 4196 2406 4200 2414
rect 4042 2196 4044 2204
rect 4052 2196 4054 2204
rect 4042 2194 4054 2196
rect 4106 2204 4118 2206
rect 4106 2196 4108 2204
rect 4116 2196 4118 2204
rect 3914 2116 3916 2124
rect 3924 2116 3926 2124
rect 3914 2114 3926 2116
rect 4042 1904 4054 1906
rect 4042 1896 4044 1904
rect 4052 1896 4054 1904
rect 4010 1864 4022 1866
rect 4010 1856 4012 1864
rect 4020 1856 4022 1864
rect 4010 1244 4022 1856
rect 4010 1236 4012 1244
rect 4020 1236 4022 1244
rect 4010 1234 4022 1236
rect 3850 1156 3852 1164
rect 3860 1156 3862 1164
rect 3850 1154 3862 1156
rect 3082 1136 3084 1144
rect 3092 1136 3094 1144
rect 3082 1134 3094 1136
rect 3050 1096 3052 1104
rect 3060 1096 3062 1104
rect 3050 1094 3062 1096
rect 3210 1124 3222 1126
rect 3210 1116 3212 1124
rect 3220 1116 3222 1124
rect 2954 956 2956 964
rect 2964 956 2966 964
rect 2954 954 2966 956
rect 3210 824 3222 1116
rect 4042 904 4054 1896
rect 4106 1844 4118 2196
rect 4106 1836 4108 1844
rect 4116 1836 4118 1844
rect 4106 1834 4118 1836
rect 4152 2014 4200 2406
rect 4330 2124 4342 2126
rect 4330 2116 4332 2124
rect 4340 2116 4342 2124
rect 4152 2006 4156 2014
rect 4164 2006 4172 2014
rect 4180 2006 4188 2014
rect 4196 2006 4200 2014
rect 4042 896 4044 904
rect 4052 896 4054 904
rect 4042 894 4054 896
rect 4152 1614 4200 2006
rect 4266 2084 4278 2086
rect 4266 2076 4268 2084
rect 4276 2076 4278 2084
rect 4266 1984 4278 2076
rect 4266 1976 4268 1984
rect 4276 1976 4278 1984
rect 4266 1974 4278 1976
rect 4152 1606 4156 1614
rect 4164 1606 4172 1614
rect 4180 1606 4188 1614
rect 4196 1606 4200 1614
rect 4152 1214 4200 1606
rect 4330 1324 4342 2116
rect 4362 2084 4374 2086
rect 4362 2076 4364 2084
rect 4372 2076 4374 2084
rect 4362 1944 4374 2076
rect 4362 1936 4364 1944
rect 4372 1936 4374 1944
rect 4362 1884 4374 1936
rect 4362 1876 4364 1884
rect 4372 1876 4374 1884
rect 4362 1874 4374 1876
rect 4458 1884 4470 2576
rect 4554 2584 4566 2656
rect 4554 2576 4556 2584
rect 4564 2576 4566 2584
rect 4554 2574 4566 2576
rect 4458 1876 4460 1884
rect 4468 1876 4470 1884
rect 4458 1874 4470 1876
rect 4842 1764 4854 1766
rect 4842 1756 4844 1764
rect 4852 1756 4854 1764
rect 4330 1316 4332 1324
rect 4340 1316 4342 1324
rect 4330 1314 4342 1316
rect 4586 1604 4598 1606
rect 4586 1596 4588 1604
rect 4596 1596 4598 1604
rect 4152 1206 4156 1214
rect 4164 1206 4172 1214
rect 4180 1206 4188 1214
rect 4196 1206 4200 1214
rect 3210 816 3212 824
rect 3220 816 3222 824
rect 3210 814 3222 816
rect 4152 814 4200 1206
rect 4490 1184 4502 1186
rect 4490 1176 4492 1184
rect 4500 1176 4502 1184
rect 2762 636 2764 644
rect 2772 636 2774 644
rect 2762 634 2774 636
rect 4152 806 4156 814
rect 4164 806 4172 814
rect 4180 806 4188 814
rect 4196 806 4200 814
rect 2632 606 2636 614
rect 2644 606 2652 614
rect 2660 606 2668 614
rect 2676 606 2680 614
rect 2632 214 2680 606
rect 2632 206 2636 214
rect 2644 206 2652 214
rect 2660 206 2668 214
rect 2676 206 2680 214
rect 2154 16 2156 24
rect 2164 16 2166 24
rect 2154 14 2166 16
rect 1112 6 1116 14
rect 1124 6 1132 14
rect 1140 6 1148 14
rect 1156 6 1160 14
rect 1112 -40 1160 6
rect 2632 -40 2680 206
rect 3274 544 3286 546
rect 3274 536 3276 544
rect 3284 536 3286 544
rect 3274 144 3286 536
rect 3274 136 3276 144
rect 3284 136 3286 144
rect 3274 134 3286 136
rect 4152 414 4200 806
rect 4426 1164 4438 1166
rect 4426 1156 4428 1164
rect 4436 1156 4438 1164
rect 4426 544 4438 1156
rect 4490 704 4502 1176
rect 4586 964 4598 1596
rect 4842 1564 4854 1756
rect 4906 1764 4918 3796
rect 4938 3304 4950 3836
rect 5386 3604 5398 3606
rect 5386 3596 5388 3604
rect 5396 3596 5398 3604
rect 4938 3296 4940 3304
rect 4948 3296 4950 3304
rect 4938 3294 4950 3296
rect 5226 3544 5238 3546
rect 5226 3536 5228 3544
rect 5236 3536 5238 3544
rect 5066 3284 5078 3286
rect 5066 3276 5068 3284
rect 5076 3276 5078 3284
rect 4938 3184 4950 3186
rect 4938 3176 4940 3184
rect 4948 3176 4950 3184
rect 4938 1984 4950 3176
rect 5066 2804 5078 3276
rect 5226 2924 5238 3536
rect 5386 3404 5398 3596
rect 5386 3396 5388 3404
rect 5396 3396 5398 3404
rect 5386 3394 5398 3396
rect 5418 3304 5430 4096
rect 5482 4084 5494 4836
rect 5514 4624 5526 4996
rect 5514 4616 5516 4624
rect 5524 4616 5526 4624
rect 5514 4614 5526 4616
rect 5720 4614 5768 5006
rect 6538 4724 6550 4726
rect 6538 4716 6540 4724
rect 6548 4716 6550 4724
rect 5720 4606 5724 4614
rect 5732 4606 5740 4614
rect 5748 4606 5756 4614
rect 5764 4606 5768 4614
rect 5578 4324 5590 4326
rect 5578 4316 5580 4324
rect 5588 4316 5590 4324
rect 5482 4076 5484 4084
rect 5492 4076 5494 4084
rect 5482 4074 5494 4076
rect 5514 4084 5526 4086
rect 5514 4076 5516 4084
rect 5524 4076 5526 4084
rect 5418 3296 5420 3304
rect 5428 3296 5430 3304
rect 5418 3294 5430 3296
rect 5450 3424 5462 3426
rect 5450 3416 5452 3424
rect 5460 3416 5462 3424
rect 5226 2916 5228 2924
rect 5236 2916 5238 2924
rect 5226 2914 5238 2916
rect 5450 2924 5462 3416
rect 5450 2916 5452 2924
rect 5460 2916 5462 2924
rect 5450 2914 5462 2916
rect 5066 2796 5068 2804
rect 5076 2796 5078 2804
rect 5066 2794 5078 2796
rect 5482 2624 5494 2626
rect 5482 2616 5484 2624
rect 5492 2616 5494 2624
rect 5482 2524 5494 2616
rect 5514 2584 5526 4076
rect 5546 3624 5558 3626
rect 5546 3616 5548 3624
rect 5556 3616 5558 3624
rect 5546 2624 5558 3616
rect 5578 3524 5590 4316
rect 5610 4284 5622 4286
rect 5610 4276 5612 4284
rect 5620 4276 5622 4284
rect 5610 4144 5622 4276
rect 5720 4214 5768 4606
rect 6442 4704 6454 4706
rect 6442 4696 6444 4704
rect 6452 4696 6454 4704
rect 5720 4206 5724 4214
rect 5732 4206 5740 4214
rect 5748 4206 5756 4214
rect 5764 4206 5768 4214
rect 5610 4136 5612 4144
rect 5620 4136 5622 4144
rect 5610 4134 5622 4136
rect 5674 4144 5686 4146
rect 5674 4136 5676 4144
rect 5684 4136 5686 4144
rect 5674 4084 5686 4136
rect 5674 4076 5676 4084
rect 5684 4076 5686 4084
rect 5674 4074 5686 4076
rect 5578 3516 5580 3524
rect 5588 3516 5590 3524
rect 5578 3514 5590 3516
rect 5610 3844 5622 3846
rect 5610 3836 5612 3844
rect 5620 3836 5622 3844
rect 5578 3444 5590 3446
rect 5578 3436 5580 3444
rect 5588 3436 5590 3444
rect 5578 3364 5590 3436
rect 5578 3356 5580 3364
rect 5588 3356 5590 3364
rect 5578 3354 5590 3356
rect 5610 3144 5622 3836
rect 5674 3824 5686 3826
rect 5674 3816 5676 3824
rect 5684 3816 5686 3824
rect 5674 3784 5686 3816
rect 5674 3776 5676 3784
rect 5684 3776 5686 3784
rect 5674 3774 5686 3776
rect 5720 3814 5768 4206
rect 5962 4504 5974 4506
rect 5962 4496 5964 4504
rect 5972 4496 5974 4504
rect 5962 4164 5974 4496
rect 6282 4504 6294 4506
rect 6282 4496 6284 4504
rect 6292 4496 6294 4504
rect 5962 4156 5964 4164
rect 5972 4156 5974 4164
rect 5962 4154 5974 4156
rect 6154 4244 6166 4246
rect 6154 4236 6156 4244
rect 6164 4236 6166 4244
rect 5898 3964 5910 3966
rect 5898 3956 5900 3964
rect 5908 3956 5910 3964
rect 5720 3806 5724 3814
rect 5732 3806 5740 3814
rect 5748 3806 5756 3814
rect 5764 3806 5768 3814
rect 5642 3604 5654 3606
rect 5642 3596 5644 3604
rect 5652 3596 5654 3604
rect 5642 3244 5654 3596
rect 5642 3236 5644 3244
rect 5652 3236 5654 3244
rect 5642 3234 5654 3236
rect 5720 3414 5768 3806
rect 5866 3844 5878 3846
rect 5866 3836 5868 3844
rect 5876 3836 5878 3844
rect 5866 3504 5878 3836
rect 5898 3764 5910 3956
rect 5898 3756 5900 3764
rect 5908 3756 5910 3764
rect 5898 3754 5910 3756
rect 5866 3496 5868 3504
rect 5876 3496 5878 3504
rect 5866 3494 5878 3496
rect 6058 3564 6070 3566
rect 6058 3556 6060 3564
rect 6068 3556 6070 3564
rect 5720 3406 5724 3414
rect 5732 3406 5740 3414
rect 5748 3406 5756 3414
rect 5764 3406 5768 3414
rect 5610 3136 5612 3144
rect 5620 3136 5622 3144
rect 5610 3134 5622 3136
rect 5578 3104 5590 3106
rect 5578 3096 5580 3104
rect 5588 3096 5590 3104
rect 5578 2984 5590 3096
rect 5578 2976 5580 2984
rect 5588 2976 5590 2984
rect 5578 2974 5590 2976
rect 5720 3014 5768 3406
rect 5720 3006 5724 3014
rect 5732 3006 5740 3014
rect 5748 3006 5756 3014
rect 5764 3006 5768 3014
rect 5546 2616 5548 2624
rect 5556 2616 5558 2624
rect 5546 2614 5558 2616
rect 5720 2614 5768 3006
rect 5994 3104 6006 3106
rect 5994 3096 5996 3104
rect 6004 3096 6006 3104
rect 5994 2844 6006 3096
rect 5994 2836 5996 2844
rect 6004 2836 6006 2844
rect 5994 2834 6006 2836
rect 6026 2924 6038 2926
rect 6026 2916 6028 2924
rect 6036 2916 6038 2924
rect 5514 2576 5516 2584
rect 5524 2576 5526 2584
rect 5514 2574 5526 2576
rect 5720 2606 5724 2614
rect 5732 2606 5740 2614
rect 5748 2606 5756 2614
rect 5764 2606 5768 2614
rect 5482 2516 5484 2524
rect 5492 2516 5494 2524
rect 5482 2514 5494 2516
rect 4938 1976 4940 1984
rect 4948 1976 4950 1984
rect 4938 1974 4950 1976
rect 5720 2214 5768 2606
rect 5720 2206 5724 2214
rect 5732 2206 5740 2214
rect 5748 2206 5756 2214
rect 5764 2206 5768 2214
rect 5674 1844 5686 1846
rect 5674 1836 5676 1844
rect 5684 1836 5686 1844
rect 4906 1756 4908 1764
rect 4916 1756 4918 1764
rect 4906 1754 4918 1756
rect 5322 1804 5334 1806
rect 5322 1796 5324 1804
rect 5332 1796 5334 1804
rect 5258 1704 5270 1706
rect 5258 1696 5260 1704
rect 5268 1696 5270 1704
rect 5194 1684 5206 1686
rect 5194 1676 5196 1684
rect 5204 1676 5206 1684
rect 4842 1556 4844 1564
rect 4852 1556 4854 1564
rect 4842 1554 4854 1556
rect 5034 1644 5046 1646
rect 5034 1636 5036 1644
rect 5044 1636 5046 1644
rect 4586 956 4588 964
rect 4596 956 4598 964
rect 4586 954 4598 956
rect 5034 964 5046 1636
rect 5066 1624 5078 1626
rect 5066 1616 5068 1624
rect 5076 1616 5078 1624
rect 5066 1324 5078 1616
rect 5066 1316 5068 1324
rect 5076 1316 5078 1324
rect 5066 1314 5078 1316
rect 5194 1124 5206 1676
rect 5258 1164 5270 1696
rect 5258 1156 5260 1164
rect 5268 1156 5270 1164
rect 5258 1154 5270 1156
rect 5290 1644 5302 1646
rect 5290 1636 5292 1644
rect 5300 1636 5302 1644
rect 5194 1116 5196 1124
rect 5204 1116 5206 1124
rect 5194 1114 5206 1116
rect 5034 956 5036 964
rect 5044 956 5046 964
rect 5034 954 5046 956
rect 4490 696 4492 704
rect 4500 696 4502 704
rect 4490 694 4502 696
rect 4426 536 4428 544
rect 4436 536 4438 544
rect 4426 534 4438 536
rect 5290 524 5302 1636
rect 5322 1084 5334 1796
rect 5674 1664 5686 1836
rect 5674 1656 5676 1664
rect 5684 1656 5686 1664
rect 5674 1654 5686 1656
rect 5720 1814 5768 2206
rect 5720 1806 5724 1814
rect 5732 1806 5740 1814
rect 5748 1806 5756 1814
rect 5764 1806 5768 1814
rect 5450 1544 5462 1546
rect 5450 1536 5452 1544
rect 5460 1536 5462 1544
rect 5450 1504 5462 1536
rect 5450 1496 5452 1504
rect 5460 1496 5462 1504
rect 5450 1494 5462 1496
rect 5674 1504 5686 1506
rect 5674 1496 5676 1504
rect 5684 1496 5686 1504
rect 5674 1364 5686 1496
rect 5674 1356 5676 1364
rect 5684 1356 5686 1364
rect 5674 1354 5686 1356
rect 5720 1414 5768 1806
rect 5994 2124 6006 2126
rect 5994 2116 5996 2124
rect 6004 2116 6006 2124
rect 5834 1704 5846 1706
rect 5834 1696 5836 1704
rect 5844 1696 5846 1704
rect 5802 1644 5814 1646
rect 5802 1636 5804 1644
rect 5812 1636 5814 1644
rect 5802 1524 5814 1636
rect 5802 1516 5804 1524
rect 5812 1516 5814 1524
rect 5802 1514 5814 1516
rect 5834 1504 5846 1696
rect 5834 1496 5836 1504
rect 5844 1496 5846 1504
rect 5834 1494 5846 1496
rect 5930 1604 5942 1606
rect 5930 1596 5932 1604
rect 5940 1596 5942 1604
rect 5930 1464 5942 1596
rect 5930 1456 5932 1464
rect 5940 1456 5942 1464
rect 5930 1454 5942 1456
rect 5962 1464 5974 1466
rect 5962 1456 5964 1464
rect 5972 1456 5974 1464
rect 5720 1406 5724 1414
rect 5732 1406 5740 1414
rect 5748 1406 5756 1414
rect 5764 1406 5768 1414
rect 5322 1076 5324 1084
rect 5332 1076 5334 1084
rect 5322 1074 5334 1076
rect 5418 1344 5430 1346
rect 5418 1336 5420 1344
rect 5428 1336 5430 1344
rect 5354 964 5366 966
rect 5354 956 5356 964
rect 5364 956 5366 964
rect 5354 644 5366 956
rect 5418 704 5430 1336
rect 5720 1014 5768 1406
rect 5930 1324 5942 1326
rect 5930 1316 5932 1324
rect 5940 1316 5942 1324
rect 5930 1284 5942 1316
rect 5962 1324 5974 1456
rect 5962 1316 5964 1324
rect 5972 1316 5974 1324
rect 5962 1314 5974 1316
rect 5930 1276 5932 1284
rect 5940 1276 5942 1284
rect 5930 1274 5942 1276
rect 5720 1006 5724 1014
rect 5732 1006 5740 1014
rect 5748 1006 5756 1014
rect 5764 1006 5768 1014
rect 5418 696 5420 704
rect 5428 696 5430 704
rect 5418 694 5430 696
rect 5674 824 5686 826
rect 5674 816 5676 824
rect 5684 816 5686 824
rect 5354 636 5356 644
rect 5364 636 5366 644
rect 5354 634 5366 636
rect 5578 664 5590 666
rect 5578 656 5580 664
rect 5588 656 5590 664
rect 5290 516 5292 524
rect 5300 516 5302 524
rect 5290 514 5302 516
rect 5578 524 5590 656
rect 5674 604 5686 816
rect 5674 596 5676 604
rect 5684 596 5686 604
rect 5674 594 5686 596
rect 5720 614 5768 1006
rect 5720 606 5724 614
rect 5732 606 5740 614
rect 5748 606 5756 614
rect 5764 606 5768 614
rect 5578 516 5580 524
rect 5588 516 5590 524
rect 5578 514 5590 516
rect 4152 406 4156 414
rect 4164 406 4172 414
rect 4180 406 4188 414
rect 4196 406 4200 414
rect 4152 14 4200 406
rect 5386 284 5398 286
rect 5386 276 5388 284
rect 5396 276 5398 284
rect 4938 144 4950 146
rect 4938 136 4940 144
rect 4948 136 4950 144
rect 4938 24 4950 136
rect 5386 144 5398 276
rect 5386 136 5388 144
rect 5396 136 5398 144
rect 5386 134 5398 136
rect 5720 214 5768 606
rect 5802 1164 5814 1166
rect 5802 1156 5804 1164
rect 5812 1156 5814 1164
rect 5802 544 5814 1156
rect 5834 1144 5846 1146
rect 5834 1136 5836 1144
rect 5844 1136 5846 1144
rect 5834 1044 5846 1136
rect 5834 1036 5836 1044
rect 5844 1036 5846 1044
rect 5834 1034 5846 1036
rect 5802 536 5804 544
rect 5812 536 5814 544
rect 5802 534 5814 536
rect 5834 964 5846 966
rect 5834 956 5836 964
rect 5844 956 5846 964
rect 5834 484 5846 956
rect 5994 624 6006 2116
rect 5994 616 5996 624
rect 6004 616 6006 624
rect 5994 614 6006 616
rect 5834 476 5836 484
rect 5844 476 5846 484
rect 5834 474 5846 476
rect 5720 206 5724 214
rect 5732 206 5740 214
rect 5748 206 5756 214
rect 5764 206 5768 214
rect 4938 16 4940 24
rect 4948 16 4950 24
rect 4938 14 4950 16
rect 4152 6 4156 14
rect 4164 6 4172 14
rect 4180 6 4188 14
rect 4196 6 4200 14
rect 4152 -40 4200 6
rect 5720 -40 5768 206
rect 6026 124 6038 2916
rect 6058 1644 6070 3556
rect 6154 3084 6166 4236
rect 6154 3076 6156 3084
rect 6164 3076 6166 3084
rect 6154 3074 6166 3076
rect 6186 3784 6198 3786
rect 6186 3776 6188 3784
rect 6196 3776 6198 3784
rect 6186 1984 6198 3776
rect 6282 3744 6294 4496
rect 6314 4484 6326 4486
rect 6314 4476 6316 4484
rect 6324 4476 6326 4484
rect 6314 4304 6326 4476
rect 6314 4296 6316 4304
rect 6324 4296 6326 4304
rect 6314 4294 6326 4296
rect 6378 4024 6390 4026
rect 6378 4016 6380 4024
rect 6388 4016 6390 4024
rect 6346 3864 6358 3866
rect 6346 3856 6348 3864
rect 6356 3856 6358 3864
rect 6282 3736 6284 3744
rect 6292 3736 6294 3744
rect 6282 3734 6294 3736
rect 6314 3744 6326 3746
rect 6314 3736 6316 3744
rect 6324 3736 6326 3744
rect 6314 3464 6326 3736
rect 6314 3456 6316 3464
rect 6324 3456 6326 3464
rect 6314 3454 6326 3456
rect 6346 2684 6358 3856
rect 6378 3764 6390 4016
rect 6378 3756 6380 3764
rect 6388 3756 6390 3764
rect 6378 3754 6390 3756
rect 6410 3904 6422 3906
rect 6410 3896 6412 3904
rect 6420 3896 6422 3904
rect 6378 3544 6390 3546
rect 6378 3536 6380 3544
rect 6388 3536 6390 3544
rect 6378 3364 6390 3536
rect 6378 3356 6380 3364
rect 6388 3356 6390 3364
rect 6378 3354 6390 3356
rect 6410 3064 6422 3896
rect 6410 3056 6412 3064
rect 6420 3056 6422 3064
rect 6410 3054 6422 3056
rect 6346 2676 6348 2684
rect 6356 2676 6358 2684
rect 6346 2674 6358 2676
rect 6410 2724 6422 2726
rect 6410 2716 6412 2724
rect 6420 2716 6422 2724
rect 6410 2524 6422 2716
rect 6410 2516 6412 2524
rect 6420 2516 6422 2524
rect 6410 2514 6422 2516
rect 6186 1976 6188 1984
rect 6196 1976 6198 1984
rect 6186 1974 6198 1976
rect 6346 1984 6358 1986
rect 6346 1976 6348 1984
rect 6356 1976 6358 1984
rect 6122 1864 6134 1866
rect 6122 1856 6124 1864
rect 6132 1856 6134 1864
rect 6058 1636 6060 1644
rect 6068 1636 6070 1644
rect 6058 1634 6070 1636
rect 6090 1644 6102 1646
rect 6090 1636 6092 1644
rect 6100 1636 6102 1644
rect 6090 1004 6102 1636
rect 6122 1324 6134 1856
rect 6122 1316 6124 1324
rect 6132 1316 6134 1324
rect 6122 1314 6134 1316
rect 6218 1504 6230 1506
rect 6218 1496 6220 1504
rect 6228 1496 6230 1504
rect 6090 996 6092 1004
rect 6100 996 6102 1004
rect 6090 994 6102 996
rect 6122 964 6134 966
rect 6122 956 6124 964
rect 6132 956 6134 964
rect 6122 604 6134 956
rect 6218 784 6230 1496
rect 6218 776 6220 784
rect 6228 776 6230 784
rect 6218 774 6230 776
rect 6282 1144 6294 1146
rect 6282 1136 6284 1144
rect 6292 1136 6294 1144
rect 6122 596 6124 604
rect 6132 596 6134 604
rect 6122 594 6134 596
rect 6282 184 6294 1136
rect 6346 1144 6358 1976
rect 6442 1924 6454 4696
rect 6506 4684 6518 4686
rect 6506 4676 6508 4684
rect 6516 4676 6518 4684
rect 6506 4424 6518 4676
rect 6506 4416 6508 4424
rect 6516 4416 6518 4424
rect 6506 4414 6518 4416
rect 6506 4004 6518 4006
rect 6506 3996 6508 4004
rect 6516 3996 6518 4004
rect 6442 1916 6444 1924
rect 6452 1916 6454 1924
rect 6442 1914 6454 1916
rect 6474 3684 6486 3686
rect 6474 3676 6476 3684
rect 6484 3676 6486 3684
rect 6474 1884 6486 3676
rect 6474 1876 6476 1884
rect 6484 1876 6486 1884
rect 6474 1874 6486 1876
rect 6346 1136 6348 1144
rect 6356 1136 6358 1144
rect 6346 1134 6358 1136
rect 6346 1104 6358 1106
rect 6346 1096 6348 1104
rect 6356 1096 6358 1104
rect 6346 924 6358 1096
rect 6346 916 6348 924
rect 6356 916 6358 924
rect 6346 914 6358 916
rect 6410 1004 6422 1006
rect 6410 996 6412 1004
rect 6420 996 6422 1004
rect 6410 844 6422 996
rect 6506 944 6518 3996
rect 6538 3444 6550 4716
rect 6698 4704 6710 4706
rect 6698 4696 6700 4704
rect 6708 4696 6710 4704
rect 6570 4584 6582 4586
rect 6570 4576 6572 4584
rect 6580 4576 6582 4584
rect 6570 3744 6582 4576
rect 6570 3736 6572 3744
rect 6580 3736 6582 3744
rect 6570 3734 6582 3736
rect 6634 4504 6646 4506
rect 6634 4496 6636 4504
rect 6644 4496 6646 4504
rect 6538 3436 6540 3444
rect 6548 3436 6550 3444
rect 6538 3434 6550 3436
rect 6570 3684 6582 3686
rect 6570 3676 6572 3684
rect 6580 3676 6582 3684
rect 6538 3064 6550 3066
rect 6538 3056 6540 3064
rect 6548 3056 6550 3064
rect 6538 2544 6550 3056
rect 6538 2536 6540 2544
rect 6548 2536 6550 2544
rect 6538 2534 6550 2536
rect 6570 2504 6582 3676
rect 6602 3524 6614 3526
rect 6602 3516 6604 3524
rect 6612 3516 6614 3524
rect 6602 3464 6614 3516
rect 6634 3484 6646 4496
rect 6698 4164 6710 4696
rect 6698 4156 6700 4164
rect 6708 4156 6710 4164
rect 6698 4154 6710 4156
rect 6730 4644 6742 4646
rect 6730 4636 6732 4644
rect 6740 4636 6742 4644
rect 6698 3584 6710 3586
rect 6698 3576 6700 3584
rect 6708 3576 6710 3584
rect 6634 3476 6636 3484
rect 6644 3476 6646 3484
rect 6634 3474 6646 3476
rect 6666 3484 6678 3486
rect 6666 3476 6668 3484
rect 6676 3476 6678 3484
rect 6602 3456 6604 3464
rect 6612 3456 6614 3464
rect 6602 2704 6614 3456
rect 6602 2696 6604 2704
rect 6612 2696 6614 2704
rect 6602 2694 6614 2696
rect 6634 3364 6646 3366
rect 6634 3356 6636 3364
rect 6644 3356 6646 3364
rect 6570 2496 6572 2504
rect 6580 2496 6582 2504
rect 6570 2494 6582 2496
rect 6538 2404 6550 2406
rect 6538 2396 6540 2404
rect 6548 2396 6550 2404
rect 6538 1964 6550 2396
rect 6538 1956 6540 1964
rect 6548 1956 6550 1964
rect 6538 1954 6550 1956
rect 6602 2364 6614 2366
rect 6602 2356 6604 2364
rect 6612 2356 6614 2364
rect 6570 1944 6582 1946
rect 6570 1936 6572 1944
rect 6580 1936 6582 1944
rect 6570 1464 6582 1936
rect 6570 1456 6572 1464
rect 6580 1456 6582 1464
rect 6570 1454 6582 1456
rect 6506 936 6508 944
rect 6516 936 6518 944
rect 6506 934 6518 936
rect 6538 1164 6550 1166
rect 6538 1156 6540 1164
rect 6548 1156 6550 1164
rect 6410 836 6412 844
rect 6420 836 6422 844
rect 6410 524 6422 836
rect 6538 704 6550 1156
rect 6538 696 6540 704
rect 6548 696 6550 704
rect 6538 694 6550 696
rect 6570 964 6582 966
rect 6570 956 6572 964
rect 6580 956 6582 964
rect 6410 516 6412 524
rect 6420 516 6422 524
rect 6410 514 6422 516
rect 6570 464 6582 956
rect 6570 456 6572 464
rect 6580 456 6582 464
rect 6570 454 6582 456
rect 6602 264 6614 2356
rect 6634 1964 6646 3356
rect 6666 3064 6678 3476
rect 6666 3056 6668 3064
rect 6676 3056 6678 3064
rect 6666 3054 6678 3056
rect 6698 2944 6710 3576
rect 6698 2936 6700 2944
rect 6708 2936 6710 2944
rect 6698 2934 6710 2936
rect 6698 2904 6710 2906
rect 6698 2896 6700 2904
rect 6708 2896 6710 2904
rect 6666 2604 6678 2606
rect 6666 2596 6668 2604
rect 6676 2596 6678 2604
rect 6666 2504 6678 2596
rect 6666 2496 6668 2504
rect 6676 2496 6678 2504
rect 6666 2494 6678 2496
rect 6634 1956 6636 1964
rect 6644 1956 6646 1964
rect 6634 1954 6646 1956
rect 6634 1864 6646 1866
rect 6634 1856 6636 1864
rect 6644 1856 6646 1864
rect 6634 1784 6646 1856
rect 6634 1776 6636 1784
rect 6644 1776 6646 1784
rect 6634 1774 6646 1776
rect 6666 1784 6678 1786
rect 6666 1776 6668 1784
rect 6676 1776 6678 1784
rect 6634 1524 6646 1526
rect 6634 1516 6636 1524
rect 6644 1516 6646 1524
rect 6634 344 6646 1516
rect 6666 1304 6678 1776
rect 6698 1644 6710 2896
rect 6698 1636 6700 1644
rect 6708 1636 6710 1644
rect 6698 1634 6710 1636
rect 6666 1296 6668 1304
rect 6676 1296 6678 1304
rect 6666 1294 6678 1296
rect 6730 664 6742 4636
rect 6762 4164 6774 4166
rect 6762 4156 6764 4164
rect 6772 4156 6774 4164
rect 6762 2904 6774 4156
rect 6826 4144 6838 4146
rect 6826 4136 6828 4144
rect 6836 4136 6838 4144
rect 6762 2896 6764 2904
rect 6772 2896 6774 2904
rect 6762 2894 6774 2896
rect 6794 3744 6806 3746
rect 6794 3736 6796 3744
rect 6804 3736 6806 3744
rect 6794 2444 6806 3736
rect 6794 2436 6796 2444
rect 6804 2436 6806 2444
rect 6794 2434 6806 2436
rect 6826 2364 6838 4136
rect 6826 2356 6828 2364
rect 6836 2356 6838 2364
rect 6826 2354 6838 2356
rect 6858 2304 6870 2306
rect 6858 2296 6860 2304
rect 6868 2296 6870 2304
rect 6794 2064 6806 2066
rect 6794 2056 6796 2064
rect 6804 2056 6806 2064
rect 6730 656 6732 664
rect 6740 656 6742 664
rect 6730 654 6742 656
rect 6762 1944 6774 1946
rect 6762 1936 6764 1944
rect 6772 1936 6774 1944
rect 6634 336 6636 344
rect 6644 336 6646 344
rect 6634 334 6646 336
rect 6730 444 6742 446
rect 6730 436 6732 444
rect 6740 436 6742 444
rect 6602 256 6604 264
rect 6612 256 6614 264
rect 6602 254 6614 256
rect 6730 244 6742 436
rect 6762 284 6774 1936
rect 6794 1764 6806 2056
rect 6794 1756 6796 1764
rect 6804 1756 6806 1764
rect 6794 1754 6806 1756
rect 6826 2004 6838 2006
rect 6826 1996 6828 2004
rect 6836 1996 6838 2004
rect 6794 1684 6806 1686
rect 6794 1676 6796 1684
rect 6804 1676 6806 1684
rect 6794 744 6806 1676
rect 6826 1544 6838 1996
rect 6826 1536 6828 1544
rect 6836 1536 6838 1544
rect 6826 1534 6838 1536
rect 6794 736 6796 744
rect 6804 736 6806 744
rect 6794 734 6806 736
rect 6826 1004 6838 1006
rect 6826 996 6828 1004
rect 6836 996 6838 1004
rect 6762 276 6764 284
rect 6772 276 6774 284
rect 6762 274 6774 276
rect 6794 584 6806 586
rect 6794 576 6796 584
rect 6804 576 6806 584
rect 6730 236 6732 244
rect 6740 236 6742 244
rect 6730 234 6742 236
rect 6282 176 6284 184
rect 6292 176 6294 184
rect 6282 174 6294 176
rect 6026 116 6028 124
rect 6036 116 6038 124
rect 6026 114 6038 116
rect 6794 104 6806 576
rect 6826 124 6838 996
rect 6858 484 6870 2296
rect 6858 476 6860 484
rect 6868 476 6870 484
rect 6858 474 6870 476
rect 6826 116 6828 124
rect 6836 116 6838 124
rect 6826 114 6838 116
rect 6794 96 6796 104
rect 6804 96 6806 104
rect 6794 94 6806 96
use INVX1  INVX1_97
timestamp 1743127117
transform 1 0 8 0 -1 210
box -4 -6 36 206
use DFFSR  DFFSR_81
timestamp 1743127117
transform 1 0 40 0 -1 210
box -4 -6 356 206
use DFFSR  DFFSR_84
timestamp 1743127117
transform 1 0 8 0 1 210
box -4 -6 356 206
use INVX1  INVX1_99
timestamp 1743127117
transform 1 0 360 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_22
timestamp 1743127117
transform -1 0 440 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_101
timestamp 1743127117
transform 1 0 440 0 -1 210
box -4 -6 36 206
use DFFSR  DFFSR_86
timestamp 1743127117
transform -1 0 824 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_360
timestamp 1743127117
transform 1 0 392 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_359
timestamp 1743127117
transform -1 0 520 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_363
timestamp 1743127117
transform 1 0 520 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_364
timestamp 1743127117
transform 1 0 584 0 1 210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_4
timestamp 1743127117
transform -1 0 792 0 1 210
box -4 -6 148 206
use DFFSR  DFFSR_89
timestamp 1743127117
transform -1 0 1176 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_10
timestamp 1743127117
transform 1 0 792 0 1 210
box -4 -6 148 206
use OAI21X1  OAI21X1_369
timestamp 1743127117
transform -1 0 1000 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_24
timestamp 1743127117
transform -1 0 1064 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_25
timestamp 1743127117
transform -1 0 1128 0 1 210
box -4 -6 68 206
use FILL  FILL_1_0_2
timestamp 1743127117
transform 1 0 1160 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1743127117
transform 1 0 1144 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_0
timestamp 1743127117
transform 1 0 1128 0 1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1743127117
transform 1 0 1208 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1743127117
transform 1 0 1192 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1743127117
transform 1 0 1176 0 -1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_10
timestamp 1743127117
transform -1 0 1480 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_9
timestamp 1743127117
transform 1 0 1368 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_10
timestamp 1743127117
transform -1 0 1464 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1743127117
transform 1 0 1176 0 1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1743127117
transform 1 0 1224 0 -1 210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_2
timestamp 1743127117
transform 1 0 1464 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_4
timestamp 1743127117
transform -1 0 1608 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_3
timestamp 1743127117
transform 1 0 1608 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_16
timestamp 1743127117
transform -1 0 2008 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_10
timestamp 1743127117
transform -1 0 1544 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_21
timestamp 1743127117
transform 1 0 1544 0 1 210
box -4 -6 196 206
use NOR2X1  NOR2X1_7
timestamp 1743127117
transform 1 0 1736 0 1 210
box -4 -6 52 206
use INVX1  INVX1_5
timestamp 1743127117
transform -1 0 1816 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_78
timestamp 1743127117
transform 1 0 2008 0 -1 210
box -4 -6 356 206
use NOR2X1  NOR2X1_8
timestamp 1743127117
transform 1 0 1816 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_1
timestamp 1743127117
transform 1 0 1864 0 1 210
box -4 -6 116 206
use DFFSR  DFFSR_15
timestamp 1743127117
transform -1 0 2328 0 1 210
box -4 -6 356 206
use INVX1  INVX1_105
timestamp 1743127117
transform 1 0 2360 0 -1 210
box -4 -6 36 206
use BUFX2  BUFX2_7
timestamp 1743127117
transform 1 0 2392 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_371
timestamp 1743127117
transform -1 0 2504 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_115
timestamp 1743127117
transform 1 0 2504 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_79
timestamp 1743127117
transform 1 0 2328 0 1 210
box -4 -6 356 206
use FILL  FILL_1_1_1
timestamp 1743127117
transform 1 0 2696 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1743127117
transform 1 0 2680 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_9
timestamp 1743127117
transform -1 0 2728 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_2
timestamp 1743127117
transform -1 0 2680 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1743127117
transform -1 0 2664 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1743127117
transform -1 0 2648 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_106
timestamp 1743127117
transform 1 0 2600 0 -1 210
box -4 -6 36 206
use BUFX2  BUFX2_8
timestamp 1743127117
transform -1 0 2600 0 -1 210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_1
timestamp 1743127117
transform -1 0 3032 0 1 210
box -4 -6 148 206
use NAND2X1  NAND2X1_117
timestamp 1743127117
transform 1 0 2840 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_116
timestamp 1743127117
transform -1 0 2840 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_372
timestamp 1743127117
transform 1 0 2728 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1743127117
transform 1 0 2712 0 1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_373
timestamp 1743127117
transform 1 0 2760 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_107
timestamp 1743127117
transform 1 0 2728 0 -1 210
box -4 -6 36 206
use DFFSR  DFFSR_80
timestamp 1743127117
transform -1 0 3176 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_6
timestamp 1743127117
transform -1 0 3224 0 -1 210
box -4 -6 52 206
use INVX8  INVX8_5
timestamp 1743127117
transform -1 0 3304 0 -1 210
box -4 -6 84 206
use OAI21X1  OAI21X1_370
timestamp 1743127117
transform 1 0 3032 0 1 210
box -4 -6 68 206
use INVX1  INVX1_104
timestamp 1743127117
transform -1 0 3128 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_77
timestamp 1743127117
transform -1 0 3480 0 1 210
box -4 -6 356 206
use BUFX2  BUFX2_13
timestamp 1743127117
transform -1 0 3352 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_94
timestamp 1743127117
transform -1 0 3704 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_17
timestamp 1743127117
transform 1 0 3480 0 1 210
box -4 -6 148 206
use BUFX2  BUFX2_12
timestamp 1743127117
transform 1 0 3704 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_10
timestamp 1743127117
transform 1 0 3752 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_92
timestamp 1743127117
transform 1 0 3800 0 -1 210
box -4 -6 356 206
use INVX1  INVX1_119
timestamp 1743127117
transform 1 0 3624 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_390
timestamp 1743127117
transform 1 0 3656 0 1 210
box -4 -6 68 206
use DFFSR  DFFSR_91
timestamp 1743127117
transform 1 0 3720 0 1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_387
timestamp 1743127117
transform -1 0 4168 0 1 210
box -4 -6 68 206
use INVX1  INVX1_116
timestamp 1743127117
transform 1 0 4072 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_11
timestamp 1743127117
transform -1 0 4200 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_117
timestamp 1743127117
transform -1 0 4312 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_388
timestamp 1743127117
transform -1 0 4280 0 1 210
box -4 -6 68 206
use FILL  FILL_1_2_2
timestamp 1743127117
transform -1 0 4216 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_1
timestamp 1743127117
transform -1 0 4200 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_0
timestamp 1743127117
transform -1 0 4184 0 1 210
box -4 -6 20 206
use FILL  FILL_0_2_2
timestamp 1743127117
transform 1 0 4232 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_1
timestamp 1743127117
transform 1 0 4216 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_0
timestamp 1743127117
transform 1 0 4200 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_99
timestamp 1743127117
transform 1 0 4312 0 1 210
box -4 -6 356 206
use DFFSR  DFFSR_95
timestamp 1743127117
transform 1 0 4248 0 -1 210
box -4 -6 356 206
use INVX1  INVX1_109
timestamp 1743127117
transform -1 0 4632 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_112
timestamp 1743127117
transform 1 0 4632 0 -1 210
box -4 -6 36 206
use DFFSR  DFFSR_100
timestamp 1743127117
transform -1 0 5016 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_379
timestamp 1743127117
transform 1 0 4664 0 1 210
box -4 -6 68 206
use INVX1  INVX1_111
timestamp 1743127117
transform 1 0 5016 0 -1 210
box -4 -6 36 206
use DFFSR  DFFSR_98
timestamp 1743127117
transform 1 0 5048 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_378
timestamp 1743127117
transform -1 0 4792 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_380
timestamp 1743127117
transform -1 0 4856 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_381
timestamp 1743127117
transform -1 0 4920 0 1 210
box -4 -6 68 206
use INVX1  INVX1_113
timestamp 1743127117
transform -1 0 4952 0 1 210
box -4 -6 36 206
use DFFSR  DFFSR_97
timestamp 1743127117
transform -1 0 5304 0 1 210
box -4 -6 356 206
use INVX1  INVX1_110
timestamp 1743127117
transform -1 0 5432 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_375
timestamp 1743127117
transform -1 0 5368 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_377
timestamp 1743127117
transform 1 0 5368 0 1 210
box -4 -6 68 206
use DFFSR  DFFSR_103
timestamp 1743127117
transform 1 0 5432 0 -1 210
box -4 -6 356 206
use OAI21X1  OAI21X1_376
timestamp 1743127117
transform -1 0 5496 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_386
timestamp 1743127117
transform 1 0 5496 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_118
timestamp 1743127117
transform -1 0 5608 0 1 210
box -4 -6 52 206
use MUX2X1  MUX2X1_50
timestamp 1743127117
transform -1 0 5704 0 1 210
box -4 -6 100 206
use FILL  FILL_1_3_0
timestamp 1743127117
transform -1 0 5720 0 1 210
box -4 -6 20 206
use FILL  FILL_1_3_1
timestamp 1743127117
transform -1 0 5736 0 1 210
box -4 -6 20 206
use FILL  FILL_1_3_2
timestamp 1743127117
transform -1 0 5752 0 1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_28
timestamp 1743127117
transform -1 0 5944 0 1 210
box -4 -6 196 206
use FILL  FILL_0_3_0
timestamp 1743127117
transform 1 0 5784 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_3_1
timestamp 1743127117
transform 1 0 5800 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_3_2
timestamp 1743127117
transform 1 0 5816 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_23
timestamp 1743127117
transform 1 0 5832 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_43
timestamp 1743127117
transform -1 0 6072 0 -1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_93
timestamp 1743127117
transform 1 0 6072 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_92
timestamp 1743127117
transform -1 0 6200 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_39
timestamp 1743127117
transform -1 0 5976 0 1 210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_38
timestamp 1743127117
transform -1 0 6168 0 1 210
box -4 -6 196 206
use MUX2X1  MUX2X1_36
timestamp 1743127117
transform -1 0 6392 0 1 210
box -4 -6 100 206
use OAI21X1  OAI21X1_116
timestamp 1743127117
transform -1 0 6296 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_115
timestamp 1743127117
transform 1 0 6168 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_99
timestamp 1743127117
transform -1 0 6328 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_98
timestamp 1743127117
transform 1 0 6200 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_119
timestamp 1743127117
transform 1 0 6488 0 1 210
box -4 -6 68 206
use MUX2X1  MUX2X1_38
timestamp 1743127117
transform 1 0 6392 0 1 210
box -4 -6 100 206
use OAI21X1  OAI21X1_352
timestamp 1743127117
transform -1 0 6424 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_43
timestamp 1743127117
transform -1 0 6360 0 -1 210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_45
timestamp 1743127117
transform -1 0 6616 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_40
timestamp 1743127117
transform -1 0 6808 0 -1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_142
timestamp 1743127117
transform -1 0 6872 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_120
timestamp 1743127117
transform -1 0 6616 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_139
timestamp 1743127117
transform 1 0 6616 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_140
timestamp 1743127117
transform -1 0 6744 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_11
timestamp 1743127117
transform -1 0 6856 0 1 210
box -4 -6 116 206
use FILL  FILL_2_1
timestamp 1743127117
transform 1 0 6856 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1
timestamp 1743127117
transform -1 0 6888 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1743127117
transform 1 0 6872 0 1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1743127117
transform 1 0 8 0 -1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_48
timestamp 1743127117
transform 1 0 200 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_49
timestamp 1743127117
transform -1 0 328 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1743127117
transform -1 0 376 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_4
timestamp 1743127117
transform 1 0 376 0 -1 610
box -4 -6 52 206
use MUX2X1  MUX2X1_21
timestamp 1743127117
transform -1 0 520 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_42
timestamp 1743127117
transform 1 0 520 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_43
timestamp 1743127117
transform -1 0 648 0 -1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1743127117
transform 1 0 648 0 -1 610
box -4 -6 196 206
use NAND2X1  NAND2X1_12
timestamp 1743127117
transform 1 0 840 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_113
timestamp 1743127117
transform -1 0 936 0 -1 610
box -4 -6 52 206
use MUX2X1  MUX2X1_9
timestamp 1743127117
transform 1 0 936 0 -1 610
box -4 -6 100 206
use MUX2X1  MUX2X1_15
timestamp 1743127117
transform -1 0 1128 0 -1 610
box -4 -6 100 206
use FILL  FILL_2_0_0
timestamp 1743127117
transform 1 0 1128 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1743127117
transform 1 0 1144 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1743127117
transform 1 0 1160 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_36
timestamp 1743127117
transform 1 0 1176 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_29
timestamp 1743127117
transform 1 0 1240 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_28
timestamp 1743127117
transform 1 0 1304 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_11
timestamp 1743127117
transform 1 0 1368 0 -1 610
box -4 -6 100 206
use INVX1  INVX1_12
timestamp 1743127117
transform 1 0 1464 0 -1 610
box -4 -6 36 206
use MUX2X1  MUX2X1_3
timestamp 1743127117
transform -1 0 1592 0 -1 610
box -4 -6 100 206
use INVX1  INVX1_17
timestamp 1743127117
transform 1 0 1592 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_69
timestamp 1743127117
transform 1 0 1624 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_4
timestamp 1743127117
transform 1 0 1688 0 -1 610
box -4 -6 68 206
use DFFSR  DFFSR_13
timestamp 1743127117
transform -1 0 2104 0 -1 610
box -4 -6 356 206
use BUFX4  BUFX4_4
timestamp 1743127117
transform -1 0 2168 0 -1 610
box -4 -6 68 206
use DFFSR  DFFSR_5
timestamp 1743127117
transform 1 0 2168 0 -1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_88
timestamp 1743127117
transform -1 0 2584 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_1_0
timestamp 1743127117
transform 1 0 2584 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1743127117
transform 1 0 2600 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1743127117
transform 1 0 2616 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_6
timestamp 1743127117
transform 1 0 2632 0 -1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_28
timestamp 1743127117
transform -1 0 3032 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_89
timestamp 1743127117
transform -1 0 3096 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_114
timestamp 1743127117
transform 1 0 3096 0 -1 610
box -4 -6 52 206
use DFFSR  DFFSR_90
timestamp 1743127117
transform -1 0 3496 0 -1 610
box -4 -6 356 206
use INVX8  INVX8_6
timestamp 1743127117
transform -1 0 3576 0 -1 610
box -4 -6 84 206
use DFFSR  DFFSR_93
timestamp 1743127117
transform -1 0 3928 0 -1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_122
timestamp 1743127117
transform 1 0 3928 0 -1 610
box -4 -6 52 206
use DFFSR  DFFSR_25
timestamp 1743127117
transform -1 0 4328 0 -1 610
box -4 -6 356 206
use FILL  FILL_2_2_0
timestamp 1743127117
transform -1 0 4344 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_1
timestamp 1743127117
transform -1 0 4360 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_2
timestamp 1743127117
transform -1 0 4376 0 -1 610
box -4 -6 20 206
use NAND2X1  NAND2X1_119
timestamp 1743127117
transform -1 0 4424 0 -1 610
box -4 -6 52 206
use OR2X2  OR2X2_10
timestamp 1743127117
transform 1 0 4424 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_32
timestamp 1743127117
transform 1 0 4488 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_31
timestamp 1743127117
transform 1 0 4536 0 -1 610
box -4 -6 52 206
use DFFSR  DFFSR_101
timestamp 1743127117
transform 1 0 4584 0 -1 610
box -4 -6 356 206
use OAI21X1  OAI21X1_383
timestamp 1743127117
transform -1 0 5000 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_382
timestamp 1743127117
transform -1 0 5064 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_29
timestamp 1743127117
transform -1 0 5112 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_374
timestamp 1743127117
transform -1 0 5176 0 -1 610
box -4 -6 68 206
use BUFX4  BUFX4_35
timestamp 1743127117
transform -1 0 5240 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1743127117
transform 1 0 5240 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_113
timestamp 1743127117
transform 1 0 5288 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_114
timestamp 1743127117
transform -1 0 5416 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_35
timestamp 1743127117
transform -1 0 5512 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_143
timestamp 1743127117
transform 1 0 5512 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_47
timestamp 1743127117
transform 1 0 5576 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_144
timestamp 1743127117
transform -1 0 5688 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_3_0
timestamp 1743127117
transform -1 0 5704 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_3_1
timestamp 1743127117
transform -1 0 5720 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_3_2
timestamp 1743127117
transform -1 0 5736 0 -1 610
box -4 -6 20 206
use XOR2X1  XOR2X1_4
timestamp 1743127117
transform -1 0 5848 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_43
timestamp 1743127117
transform -1 0 5896 0 -1 610
box -4 -6 52 206
use MUX2X1  MUX2X1_27
timestamp 1743127117
transform -1 0 5992 0 -1 610
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_44
timestamp 1743127117
transform -1 0 6184 0 -1 610
box -4 -6 196 206
use MUX2X1  MUX2X1_28
timestamp 1743127117
transform 1 0 6184 0 -1 610
box -4 -6 100 206
use BUFX4  BUFX4_32
timestamp 1743127117
transform -1 0 6344 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_29
timestamp 1743127117
transform 1 0 6344 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_95
timestamp 1743127117
transform -1 0 6504 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_96
timestamp 1743127117
transform -1 0 6568 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_48
timestamp 1743127117
transform -1 0 6664 0 -1 610
box -4 -6 100 206
use MUX2X1  MUX2X1_37
timestamp 1743127117
transform 1 0 6664 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_117
timestamp 1743127117
transform 1 0 6760 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_118
timestamp 1743127117
transform -1 0 6888 0 -1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_19
timestamp 1743127117
transform 1 0 8 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_3
timestamp 1743127117
transform 1 0 200 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_4
timestamp 1743127117
transform -1 0 328 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_1
timestamp 1743127117
transform 1 0 328 0 1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_55
timestamp 1743127117
transform -1 0 488 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_24
timestamp 1743127117
transform -1 0 584 0 1 610
box -4 -6 100 206
use MUX2X1  MUX2X1_18
timestamp 1743127117
transform -1 0 680 0 1 610
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1743127117
transform 1 0 680 0 1 610
box -4 -6 196 206
use INVX1  INVX1_20
timestamp 1743127117
transform 1 0 872 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_19
timestamp 1743127117
transform 1 0 904 0 1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1743127117
transform 1 0 952 0 1 610
box -4 -6 196 206
use FILL  FILL_3_0_0
timestamp 1743127117
transform -1 0 1160 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1743127117
transform -1 0 1176 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1743127117
transform -1 0 1192 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_37
timestamp 1743127117
transform -1 0 1256 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_74
timestamp 1743127117
transform 1 0 1256 0 1 610
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1743127117
transform 1 0 1320 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_62
timestamp 1743127117
transform 1 0 1352 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_2
timestamp 1743127117
transform 1 0 1416 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_61
timestamp 1743127117
transform 1 0 1480 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_75
timestamp 1743127117
transform 1 0 1544 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_63
timestamp 1743127117
transform 1 0 1608 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_71
timestamp 1743127117
transform 1 0 1672 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_11
timestamp 1743127117
transform 1 0 1736 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1743127117
transform 1 0 1800 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_13
timestamp 1743127117
transform 1 0 1848 0 1 610
box -4 -6 52 206
use INVX1  INVX1_14
timestamp 1743127117
transform -1 0 1928 0 1 610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_3
timestamp 1743127117
transform -1 0 2040 0 1 610
box -4 -6 116 206
use CLKBUF1  CLKBUF1_8
timestamp 1743127117
transform 1 0 2040 0 1 610
box -4 -6 148 206
use BUFX4  BUFX4_53
timestamp 1743127117
transform -1 0 2248 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_50
timestamp 1743127117
transform -1 0 2312 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_27
timestamp 1743127117
transform -1 0 2360 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_17
timestamp 1743127117
transform 1 0 2360 0 1 610
box -4 -6 356 206
use FILL  FILL_3_1_0
timestamp 1743127117
transform -1 0 2728 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1743127117
transform -1 0 2744 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1743127117
transform -1 0 2760 0 1 610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_6
timestamp 1743127117
transform -1 0 2904 0 1 610
box -4 -6 148 206
use NAND2X1  NAND2X1_18
timestamp 1743127117
transform -1 0 2952 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_68
timestamp 1743127117
transform 1 0 2952 0 1 610
box -4 -6 68 206
use DFFSR  DFFSR_9
timestamp 1743127117
transform 1 0 3016 0 1 610
box -4 -6 356 206
use DFFSR  DFFSR_82
timestamp 1743127117
transform 1 0 3368 0 1 610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_2
timestamp 1743127117
transform 1 0 3720 0 1 610
box -4 -6 148 206
use INVX1  INVX1_118
timestamp 1743127117
transform 1 0 3864 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_389
timestamp 1743127117
transform 1 0 3896 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_121
timestamp 1743127117
transform -1 0 4008 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_120
timestamp 1743127117
transform 1 0 4008 0 1 610
box -4 -6 52 206
use FILL  FILL_3_2_0
timestamp 1743127117
transform -1 0 4072 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_1
timestamp 1743127117
transform -1 0 4088 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_2
timestamp 1743127117
transform -1 0 4104 0 1 610
box -4 -6 20 206
use DFFSR  DFFSR_23
timestamp 1743127117
transform -1 0 4456 0 1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_56
timestamp 1743127117
transform -1 0 4504 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_100
timestamp 1743127117
transform -1 0 4568 0 1 610
box -4 -6 68 206
use INVX8  INVX8_2
timestamp 1743127117
transform -1 0 4648 0 1 610
box -4 -6 84 206
use DFFSR  DFFSR_102
timestamp 1743127117
transform 1 0 4648 0 1 610
box -4 -6 356 206
use INVX1  INVX1_114
timestamp 1743127117
transform -1 0 5032 0 1 610
box -4 -6 36 206
use INVX1  INVX1_115
timestamp 1743127117
transform 1 0 5032 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_385
timestamp 1743127117
transform 1 0 5064 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_384
timestamp 1743127117
transform -1 0 5192 0 1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_13
timestamp 1743127117
transform -1 0 5336 0 1 610
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_37
timestamp 1743127117
transform 1 0 5336 0 1 610
box -4 -6 196 206
use NAND3X1  NAND3X1_9
timestamp 1743127117
transform -1 0 5592 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_127
timestamp 1743127117
transform 1 0 5592 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_128
timestamp 1743127117
transform -1 0 5720 0 1 610
box -4 -6 68 206
use FILL  FILL_3_3_0
timestamp 1743127117
transform -1 0 5736 0 1 610
box -4 -6 20 206
use FILL  FILL_3_3_1
timestamp 1743127117
transform -1 0 5752 0 1 610
box -4 -6 20 206
use FILL  FILL_3_3_2
timestamp 1743127117
transform -1 0 5768 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_154
timestamp 1743127117
transform -1 0 5832 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1743127117
transform -1 0 5896 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_32
timestamp 1743127117
transform -1 0 6088 0 1 610
box -4 -6 196 206
use NAND3X1  NAND3X1_11
timestamp 1743127117
transform -1 0 6152 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_162
timestamp 1743127117
transform 1 0 6152 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_12
timestamp 1743127117
transform -1 0 6280 0 1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_30
timestamp 1743127117
transform 1 0 6280 0 1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_102
timestamp 1743127117
transform 1 0 6376 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_46
timestamp 1743127117
transform -1 0 6632 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_124
timestamp 1743127117
transform -1 0 6696 0 1 610
box -4 -6 68 206
use INVX1  INVX1_41
timestamp 1743127117
transform -1 0 6728 0 1 610
box -4 -6 36 206
use CLKBUF1  CLKBUF1_20
timestamp 1743127117
transform 1 0 6728 0 1 610
box -4 -6 148 206
use FILL  FILL_4_1
timestamp 1743127117
transform 1 0 6872 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_13
timestamp 1743127117
transform -1 0 72 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_4
timestamp 1743127117
transform -1 0 168 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_12
timestamp 1743127117
transform -1 0 232 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_11
timestamp 1743127117
transform -1 0 296 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_5
timestamp 1743127117
transform 1 0 296 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_54
timestamp 1743127117
transform 1 0 360 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_30
timestamp 1743127117
transform 1 0 424 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_31
timestamp 1743127117
transform -1 0 552 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_12
timestamp 1743127117
transform 1 0 552 0 -1 1010
box -4 -6 100 206
use BUFX4  BUFX4_14
timestamp 1743127117
transform -1 0 712 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1743127117
transform -1 0 904 0 -1 1010
box -4 -6 196 206
use INVX1  INVX1_19
timestamp 1743127117
transform 1 0 904 0 -1 1010
box -4 -6 36 206
use BUFX4  BUFX4_76
timestamp 1743127117
transform 1 0 936 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_5
timestamp 1743127117
transform 1 0 1000 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_73
timestamp 1743127117
transform -1 0 1128 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1743127117
transform 1 0 1128 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1743127117
transform 1 0 1144 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1743127117
transform 1 0 1160 0 -1 1010
box -4 -6 20 206
use BUFX4  BUFX4_12
timestamp 1743127117
transform 1 0 1176 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_22
timestamp 1743127117
transform -1 0 1336 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_50
timestamp 1743127117
transform 1 0 1336 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_51
timestamp 1743127117
transform -1 0 1464 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_9
timestamp 1743127117
transform -1 0 1512 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1743127117
transform 1 0 1512 0 -1 1010
box -4 -6 196 206
use NAND2X1  NAND2X1_15
timestamp 1743127117
transform 1 0 1704 0 -1 1010
box -4 -6 52 206
use DFFSR  DFFSR_1
timestamp 1743127117
transform -1 0 2104 0 -1 1010
box -4 -6 356 206
use NAND2X1  NAND2X1_7
timestamp 1743127117
transform 1 0 2104 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_22
timestamp 1743127117
transform 1 0 2152 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_11
timestamp 1743127117
transform 1 0 2216 0 -1 1010
box -4 -6 36 206
use AND2X2  AND2X2_1
timestamp 1743127117
transform 1 0 2248 0 -1 1010
box -4 -6 68 206
use XOR2X1  XOR2X1_1
timestamp 1743127117
transform -1 0 2424 0 -1 1010
box -4 -6 116 206
use OAI21X1  OAI21X1_20
timestamp 1743127117
transform -1 0 2488 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_1_0
timestamp 1743127117
transform -1 0 2504 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1743127117
transform -1 0 2520 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1743127117
transform -1 0 2536 0 -1 1010
box -4 -6 20 206
use DFFSR  DFFSR_19
timestamp 1743127117
transform -1 0 2888 0 -1 1010
box -4 -6 356 206
use BUFX4  BUFX4_51
timestamp 1743127117
transform 1 0 2888 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_86
timestamp 1743127117
transform 1 0 2952 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_25
timestamp 1743127117
transform 1 0 3016 0 -1 1010
box -4 -6 52 206
use DFFSR  DFFSR_3
timestamp 1743127117
transform -1 0 3416 0 -1 1010
box -4 -6 356 206
use INVX1  INVX1_108
timestamp 1743127117
transform 1 0 3416 0 -1 1010
box -4 -6 36 206
use DFFSR  DFFSR_104
timestamp 1743127117
transform 1 0 3448 0 -1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_153
timestamp 1743127117
transform 1 0 3800 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_44
timestamp 1743127117
transform 1 0 3864 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_176
timestamp 1743127117
transform 1 0 3912 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_54
timestamp 1743127117
transform 1 0 3976 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_2_0
timestamp 1743127117
transform -1 0 4040 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_1
timestamp 1743127117
transform -1 0 4056 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_2
timestamp 1743127117
transform -1 0 4072 0 -1 1010
box -4 -6 20 206
use DFFSR  DFFSR_27
timestamp 1743127117
transform -1 0 4424 0 -1 1010
box -4 -6 356 206
use NAND2X1  NAND2X1_48
timestamp 1743127117
transform 1 0 4424 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_178
timestamp 1743127117
transform -1 0 4536 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_97
timestamp 1743127117
transform -1 0 4600 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_177
timestamp 1743127117
transform 1 0 4600 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_24
timestamp 1743127117
transform -1 0 5016 0 -1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_91
timestamp 1743127117
transform 1 0 5016 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_34
timestamp 1743127117
transform 1 0 5080 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_33
timestamp 1743127117
transform -1 0 5176 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_30
timestamp 1743127117
transform 1 0 5176 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_94
timestamp 1743127117
transform 1 0 5208 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_150
timestamp 1743127117
transform -1 0 5336 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_36
timestamp 1743127117
transform -1 0 5368 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_156
timestamp 1743127117
transform -1 0 5432 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_155
timestamp 1743127117
transform -1 0 5496 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_40
timestamp 1743127117
transform -1 0 5528 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_164
timestamp 1743127117
transform -1 0 5592 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_163
timestamp 1743127117
transform -1 0 5656 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_42
timestamp 1743127117
transform -1 0 5752 0 -1 1010
box -4 -6 100 206
use FILL  FILL_4_3_0
timestamp 1743127117
transform -1 0 5768 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_3_1
timestamp 1743127117
transform -1 0 5784 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_3_2
timestamp 1743127117
transform -1 0 5800 0 -1 1010
box -4 -6 20 206
use INVX1  INVX1_44
timestamp 1743127117
transform -1 0 5832 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_34
timestamp 1743127117
transform -1 0 6024 0 -1 1010
box -4 -6 196 206
use MUX2X1  MUX2X1_44
timestamp 1743127117
transform 1 0 6024 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_158
timestamp 1743127117
transform -1 0 6184 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_132
timestamp 1743127117
transform 1 0 6184 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_131
timestamp 1743127117
transform -1 0 6312 0 -1 1010
box -4 -6 68 206
use BUFX4  BUFX4_55
timestamp 1743127117
transform 1 0 6312 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_101
timestamp 1743127117
transform 1 0 6376 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_123
timestamp 1743127117
transform 1 0 6440 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_42
timestamp 1743127117
transform -1 0 6696 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_27
timestamp 1743127117
transform 1 0 6696 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_22
timestamp 1743127117
transform 1 0 8 0 1 1010
box -4 -6 196 206
use BUFX4  BUFX4_74
timestamp 1743127117
transform -1 0 264 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_2
timestamp 1743127117
transform 1 0 264 0 1 1010
box -4 -6 100 206
use BUFX4  BUFX4_42
timestamp 1743127117
transform 1 0 360 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_73
timestamp 1743127117
transform 1 0 424 0 1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1743127117
transform 1 0 488 0 1 1010
box -4 -6 196 206
use MUX2X1  MUX2X1_10
timestamp 1743127117
transform 1 0 680 0 1 1010
box -4 -6 100 206
use INVX1  INVX1_15
timestamp 1743127117
transform 1 0 776 0 1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1743127117
transform 1 0 808 0 1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_59
timestamp 1743127117
transform 1 0 1000 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_58
timestamp 1743127117
transform -1 0 1128 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1743127117
transform 1 0 1128 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1743127117
transform 1 0 1144 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1743127117
transform 1 0 1160 0 1 1010
box -4 -6 20 206
use BUFX4  BUFX4_43
timestamp 1743127117
transform 1 0 1176 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_23
timestamp 1743127117
transform 1 0 1240 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_65
timestamp 1743127117
transform 1 0 1288 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_16
timestamp 1743127117
transform -1 0 1448 0 1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_39
timestamp 1743127117
transform 1 0 1448 0 1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1743127117
transform 1 0 1512 0 1 1010
box -4 -6 196 206
use INVX1  INVX1_16
timestamp 1743127117
transform 1 0 1704 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_66
timestamp 1743127117
transform 1 0 1736 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_67
timestamp 1743127117
transform 1 0 1800 0 1 1010
box -4 -6 68 206
use INVX2  INVX2_1
timestamp 1743127117
transform -1 0 1896 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_84
timestamp 1743127117
transform -1 0 1960 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_85
timestamp 1743127117
transform -1 0 2024 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_2
timestamp 1743127117
transform 1 0 2024 0 1 1010
box -4 -6 52 206
use OR2X2  OR2X2_1
timestamp 1743127117
transform -1 0 2136 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1743127117
transform -1 0 2184 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1743127117
transform -1 0 2216 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_1
timestamp 1743127117
transform -1 0 2264 0 1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_1
timestamp 1743127117
transform 1 0 2264 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_21
timestamp 1743127117
transform 1 0 2328 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_23
timestamp 1743127117
transform 1 0 2392 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1743127117
transform 1 0 2456 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_87
timestamp 1743127117
transform 1 0 2504 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1743127117
transform 1 0 2568 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_1_0
timestamp 1743127117
transform -1 0 2632 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1743127117
transform -1 0 2648 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1743127117
transform -1 0 2664 0 1 1010
box -4 -6 20 206
use DFFSR  DFFSR_4
timestamp 1743127117
transform -1 0 3016 0 1 1010
box -4 -6 356 206
use BUFX4  BUFX4_97
timestamp 1743127117
transform 1 0 3016 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_5
timestamp 1743127117
transform 1 0 3080 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_182
timestamp 1743127117
transform -1 0 3160 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_60
timestamp 1743127117
transform 1 0 3160 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1743127117
transform 1 0 3224 0 1 1010
box -4 -6 52 206
use DFFSR  DFFSR_7
timestamp 1743127117
transform -1 0 3624 0 1 1010
box -4 -6 356 206
use DFFSR  DFFSR_96
timestamp 1743127117
transform -1 0 3976 0 1 1010
box -4 -6 356 206
use INVX1  INVX1_120
timestamp 1743127117
transform -1 0 4008 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_149
timestamp 1743127117
transform -1 0 4072 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_42
timestamp 1743127117
transform 1 0 4072 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_161
timestamp 1743127117
transform -1 0 4184 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_2_0
timestamp 1743127117
transform -1 0 4200 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_1
timestamp 1743127117
transform -1 0 4216 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_2
timestamp 1743127117
transform -1 0 4232 0 1 1010
box -4 -6 20 206
use DFFSR  DFFSR_29
timestamp 1743127117
transform -1 0 4584 0 1 1010
box -4 -6 356 206
use BUFX4  BUFX4_79
timestamp 1743127117
transform -1 0 4648 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_175
timestamp 1743127117
transform 1 0 4648 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_55
timestamp 1743127117
transform 1 0 4712 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_53
timestamp 1743127117
transform 1 0 4760 0 1 1010
box -4 -6 52 206
use DFFSR  DFFSR_22
timestamp 1743127117
transform -1 0 5160 0 1 1010
box -4 -6 356 206
use BUFX4  BUFX4_78
timestamp 1743127117
transform -1 0 5224 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_152
timestamp 1743127117
transform -1 0 5288 0 1 1010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_16
timestamp 1743127117
transform -1 0 5432 0 1 1010
box -4 -6 148 206
use OAI21X1  OAI21X1_151
timestamp 1743127117
transform -1 0 5496 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_40
timestamp 1743127117
transform 1 0 5496 0 1 1010
box -4 -6 52 206
use MUX2X1  MUX2X1_47
timestamp 1743127117
transform -1 0 5640 0 1 1010
box -4 -6 100 206
use BUFX4  BUFX4_56
timestamp 1743127117
transform 1 0 5640 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_3_0
timestamp 1743127117
transform 1 0 5704 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_3_1
timestamp 1743127117
transform 1 0 5720 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_3_2
timestamp 1743127117
transform 1 0 5736 0 1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_41
timestamp 1743127117
transform 1 0 5752 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_38
timestamp 1743127117
transform -1 0 5832 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_160
timestamp 1743127117
transform -1 0 5896 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_159
timestamp 1743127117
transform 1 0 5896 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_45
timestamp 1743127117
transform -1 0 6008 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_42
timestamp 1743127117
transform -1 0 6040 0 1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_33
timestamp 1743127117
transform -1 0 6232 0 1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_130
timestamp 1743127117
transform 1 0 6232 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_129
timestamp 1743127117
transform -1 0 6360 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_43
timestamp 1743127117
transform 1 0 6360 0 1 1010
box -4 -6 100 206
use BUFX4  BUFX4_37
timestamp 1743127117
transform -1 0 6520 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_40
timestamp 1743127117
transform -1 0 6584 0 1 1010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_27
timestamp 1743127117
transform -1 0 6728 0 1 1010
box -4 -6 148 206
use OAI21X1  OAI21X1_141
timestamp 1743127117
transform 1 0 6728 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_49
timestamp 1743127117
transform 1 0 6792 0 1 1010
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_20
timestamp 1743127117
transform 1 0 8 0 -1 1410
box -4 -6 196 206
use OAI21X1  OAI21X1_6
timestamp 1743127117
transform -1 0 264 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_7
timestamp 1743127117
transform -1 0 328 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1743127117
transform 1 0 328 0 -1 1410
box -4 -6 196 206
use OAI21X1  OAI21X1_46
timestamp 1743127117
transform 1 0 520 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_47
timestamp 1743127117
transform -1 0 648 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_20
timestamp 1743127117
transform -1 0 744 0 -1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_27
timestamp 1743127117
transform 1 0 744 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_26
timestamp 1743127117
transform -1 0 872 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1743127117
transform 1 0 872 0 -1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_26
timestamp 1743127117
transform -1 0 1000 0 -1 1410
box -4 -6 100 206
use NAND3X1  NAND3X1_7
timestamp 1743127117
transform 1 0 1000 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_81
timestamp 1743127117
transform -1 0 1128 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_0_0
timestamp 1743127117
transform 1 0 1128 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1743127117
transform 1 0 1144 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1743127117
transform 1 0 1160 0 -1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_17
timestamp 1743127117
transform 1 0 1176 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_70
timestamp 1743127117
transform -1 0 1288 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_18
timestamp 1743127117
transform -1 0 1320 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_3
timestamp 1743127117
transform 1 0 1320 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_24
timestamp 1743127117
transform 1 0 1384 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_82
timestamp 1743127117
transform 1 0 1416 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_38
timestamp 1743127117
transform -1 0 1544 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_83
timestamp 1743127117
transform 1 0 1544 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1743127117
transform -1 0 1640 0 -1 1410
box -4 -6 36 206
use BUFX4  BUFX4_75
timestamp 1743127117
transform 1 0 1640 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_6
timestamp 1743127117
transform -1 0 1768 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_77
timestamp 1743127117
transform -1 0 1832 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1743127117
transform -1 0 1880 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_78
timestamp 1743127117
transform -1 0 1944 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_79
timestamp 1743127117
transform 1 0 1944 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_14
timestamp 1743127117
transform -1 0 2360 0 -1 1410
box -4 -6 356 206
use NAND3X1  NAND3X1_1
timestamp 1743127117
transform -1 0 2424 0 -1 1410
box -4 -6 68 206
use OR2X2  OR2X2_2
timestamp 1743127117
transform -1 0 2488 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_6
timestamp 1743127117
transform -1 0 2536 0 -1 1410
box -4 -6 52 206
use INVX8  INVX8_1
timestamp 1743127117
transform -1 0 2616 0 -1 1410
box -4 -6 84 206
use FILL  FILL_6_1_0
timestamp 1743127117
transform -1 0 2632 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1743127117
transform -1 0 2648 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1743127117
transform -1 0 2664 0 -1 1410
box -4 -6 20 206
use BUFX4  BUFX4_52
timestamp 1743127117
transform -1 0 2728 0 -1 1410
box -4 -6 68 206
use BUFX4  BUFX4_99
timestamp 1743127117
transform -1 0 2792 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_20
timestamp 1743127117
transform -1 0 2840 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_72
timestamp 1743127117
transform -1 0 2904 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1743127117
transform -1 0 2952 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_64
timestamp 1743127117
transform 1 0 2952 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_22
timestamp 1743127117
transform -1 0 3064 0 -1 1410
box -4 -6 52 206
use DFFSR  DFFSR_8
timestamp 1743127117
transform -1 0 3416 0 -1 1410
box -4 -6 356 206
use NOR2X1  NOR2X1_5
timestamp 1743127117
transform -1 0 3464 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_15
timestamp 1743127117
transform 1 0 3464 0 -1 1410
box -4 -6 52 206
use DFFSR  DFFSR_26
timestamp 1743127117
transform 1 0 3512 0 -1 1410
box -4 -6 356 206
use BUFX4  BUFX4_59
timestamp 1743127117
transform -1 0 3928 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_30
timestamp 1743127117
transform -1 0 4280 0 -1 1410
box -4 -6 356 206
use FILL  FILL_6_2_0
timestamp 1743127117
transform -1 0 4296 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_1
timestamp 1743127117
transform -1 0 4312 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_2
timestamp 1743127117
transform -1 0 4328 0 -1 1410
box -4 -6 20 206
use BUFX2  BUFX2_3
timestamp 1743127117
transform -1 0 4376 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_32
timestamp 1743127117
transform 1 0 4376 0 -1 1410
box -4 -6 36 206
use DFFSR  DFFSR_154
timestamp 1743127117
transform 1 0 4408 0 -1 1410
box -4 -6 356 206
use DFFSR  DFFSR_33
timestamp 1743127117
transform 1 0 4760 0 -1 1410
box -4 -6 356 206
use OAI21X1  OAI21X1_106
timestamp 1743127117
transform -1 0 5176 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_25
timestamp 1743127117
transform -1 0 5368 0 -1 1410
box -4 -6 196 206
use BUFX4  BUFX4_54
timestamp 1743127117
transform 1 0 5368 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_138
timestamp 1743127117
transform 1 0 5432 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_137
timestamp 1743127117
transform -1 0 5560 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_19
timestamp 1743127117
transform 1 0 5560 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_48
timestamp 1743127117
transform 1 0 5608 0 -1 1410
box -4 -6 196 206
use FILL  FILL_6_3_0
timestamp 1743127117
transform -1 0 5816 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_3_1
timestamp 1743127117
transform -1 0 5832 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_3_2
timestamp 1743127117
transform -1 0 5848 0 -1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_51
timestamp 1743127117
transform -1 0 5896 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1743127117
transform -1 0 5960 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_170
timestamp 1743127117
transform -1 0 6024 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_52
timestamp 1743127117
transform 1 0 6024 0 -1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_148
timestamp 1743127117
transform 1 0 6120 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_147
timestamp 1743127117
transform 1 0 6184 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_30
timestamp 1743127117
transform -1 0 6440 0 -1 1410
box -4 -6 196 206
use INVX1  INVX1_47
timestamp 1743127117
transform -1 0 6472 0 -1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_40
timestamp 1743127117
transform 1 0 6472 0 -1 1410
box -4 -6 100 206
use BUFX4  BUFX4_38
timestamp 1743127117
transform 1 0 6568 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_134
timestamp 1743127117
transform 1 0 6632 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_35
timestamp 1743127117
transform -1 0 6888 0 -1 1410
box -4 -6 196 206
use INVX1  INVX1_103
timestamp 1743127117
transform -1 0 40 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_368
timestamp 1743127117
transform 1 0 40 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_367
timestamp 1743127117
transform -1 0 168 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_72
timestamp 1743127117
transform -1 0 232 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_44
timestamp 1743127117
transform -1 0 296 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_34
timestamp 1743127117
transform 1 0 296 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_35
timestamp 1743127117
transform -1 0 424 0 1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_14
timestamp 1743127117
transform -1 0 520 0 1 1410
box -4 -6 100 206
use MUX2X1  MUX2X1_6
timestamp 1743127117
transform -1 0 616 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_19
timestamp 1743127117
transform 1 0 616 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_18
timestamp 1743127117
transform -1 0 744 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_10
timestamp 1743127117
transform -1 0 808 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_52
timestamp 1743127117
transform 1 0 808 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_53
timestamp 1743127117
transform -1 0 936 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_24
timestamp 1743127117
transform -1 0 1128 0 1 1410
box -4 -6 196 206
use FILL  FILL_7_0_0
timestamp 1743127117
transform 1 0 1128 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1743127117
transform 1 0 1144 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1743127117
transform 1 0 1160 0 1 1410
box -4 -6 20 206
use MUX2X1  MUX2X1_23
timestamp 1743127117
transform 1 0 1176 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_40
timestamp 1743127117
transform 1 0 1272 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_13
timestamp 1743127117
transform 1 0 1336 0 1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_13
timestamp 1743127117
transform 1 0 1400 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_33
timestamp 1743127117
transform 1 0 1496 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_32
timestamp 1743127117
transform -1 0 1624 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_17
timestamp 1743127117
transform 1 0 1624 0 1 1410
box -4 -6 196 206
use INVX1  INVX1_21
timestamp 1743127117
transform 1 0 1816 0 1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_5
timestamp 1743127117
transform 1 0 1848 0 1 1410
box -4 -6 100 206
use MUX2X1  MUX2X1_25
timestamp 1743127117
transform 1 0 1944 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_56
timestamp 1743127117
transform 1 0 2040 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_57
timestamp 1743127117
transform -1 0 2168 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1743127117
transform -1 0 2360 0 1 1410
box -4 -6 196 206
use MUX2X1  MUX2X1_8
timestamp 1743127117
transform 1 0 2360 0 1 1410
box -4 -6 100 206
use MUX2X1  MUX2X1_7
timestamp 1743127117
transform 1 0 2456 0 1 1410
box -4 -6 100 206
use XOR2X1  XOR2X1_2
timestamp 1743127117
transform 1 0 2552 0 1 1410
box -4 -6 116 206
use FILL  FILL_7_1_0
timestamp 1743127117
transform 1 0 2664 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1743127117
transform 1 0 2680 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1743127117
transform 1 0 2696 0 1 1410
box -4 -6 20 206
use DFFSR  DFFSR_2
timestamp 1743127117
transform 1 0 2712 0 1 1410
box -4 -6 356 206
use OAI21X1  OAI21X1_76
timestamp 1743127117
transform 1 0 3064 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_11
timestamp 1743127117
transform 1 0 3128 0 1 1410
box -4 -6 356 206
use DFFSR  DFFSR_140
timestamp 1743127117
transform -1 0 3832 0 1 1410
box -4 -6 356 206
use DFFSR  DFFSR_156
timestamp 1743127117
transform 1 0 3832 0 1 1410
box -4 -6 356 206
use FILL  FILL_7_2_0
timestamp 1743127117
transform -1 0 4200 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_1
timestamp 1743127117
transform -1 0 4216 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_2
timestamp 1743127117
transform -1 0 4232 0 1 1410
box -4 -6 20 206
use INVX1  INVX1_177
timestamp 1743127117
transform -1 0 4264 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_165
timestamp 1743127117
transform 1 0 4264 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_50
timestamp 1743127117
transform 1 0 4328 0 1 1410
box -4 -6 52 206
use DFFSR  DFFSR_157
timestamp 1743127117
transform 1 0 4376 0 1 1410
box -4 -6 356 206
use INVX1  INVX1_178
timestamp 1743127117
transform -1 0 4760 0 1 1410
box -4 -6 36 206
use DFFSR  DFFSR_144
timestamp 1743127117
transform 1 0 4760 0 1 1410
box -4 -6 356 206
use INVX1  INVX1_33
timestamp 1743127117
transform 1 0 5112 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_103
timestamp 1743127117
transform -1 0 5208 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_174
timestamp 1743127117
transform 1 0 5208 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_173
timestamp 1743127117
transform -1 0 5336 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_14
timestamp 1743127117
transform 1 0 5336 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_26
timestamp 1743127117
transform 1 0 5384 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_90
timestamp 1743127117
transform 1 0 5416 0 1 1410
box -4 -6 68 206
use INVX2  INVX2_2
timestamp 1743127117
transform -1 0 5512 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_39
timestamp 1743127117
transform -1 0 5560 0 1 1410
box -4 -6 52 206
use BUFX4  BUFX4_39
timestamp 1743127117
transform -1 0 5624 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_168
timestamp 1743127117
transform -1 0 5688 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_3_0
timestamp 1743127117
transform -1 0 5704 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_3_1
timestamp 1743127117
transform -1 0 5720 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_3_2
timestamp 1743127117
transform -1 0 5736 0 1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_167
timestamp 1743127117
transform -1 0 5800 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_107
timestamp 1743127117
transform 1 0 5800 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_108
timestamp 1743127117
transform -1 0 5928 0 1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_32
timestamp 1743127117
transform 1 0 5928 0 1 1410
box -4 -6 100 206
use BUFX4  BUFX4_36
timestamp 1743127117
transform 1 0 6024 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_166
timestamp 1743127117
transform 1 0 6088 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_33
timestamp 1743127117
transform -1 0 6216 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_13
timestamp 1743127117
transform -1 0 6280 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_34
timestamp 1743127117
transform 1 0 6280 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_57
timestamp 1743127117
transform 1 0 6344 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_46
timestamp 1743127117
transform -1 0 6440 0 1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_45
timestamp 1743127117
transform 1 0 6440 0 1 1410
box -4 -6 100 206
use MUX2X1  MUX2X1_31
timestamp 1743127117
transform 1 0 6536 0 1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_105
timestamp 1743127117
transform 1 0 6632 0 1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_47
timestamp 1743127117
transform -1 0 6888 0 1 1410
box -4 -6 196 206
use DFFSR  DFFSR_88
timestamp 1743127117
transform 1 0 8 0 -1 1810
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_18
timestamp 1743127117
transform 1 0 360 0 -1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_6
timestamp 1743127117
transform -1 0 600 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_365
timestamp 1743127117
transform 1 0 600 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_366
timestamp 1743127117
transform -1 0 728 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_102
timestamp 1743127117
transform -1 0 760 0 -1 1810
box -4 -6 36 206
use DFFSR  DFFSR_87
timestamp 1743127117
transform 1 0 760 0 -1 1810
box -4 -6 356 206
use FILL  FILL_8_0_0
timestamp 1743127117
transform -1 0 1128 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1743127117
transform -1 0 1144 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1743127117
transform -1 0 1160 0 -1 1810
box -4 -6 20 206
use INVX1  INVX1_6
timestamp 1743127117
transform -1 0 1192 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_5
timestamp 1743127117
transform -1 0 1240 0 -1 1810
box -4 -6 52 206
use BUFX4  BUFX4_41
timestamp 1743127117
transform 1 0 1240 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_41
timestamp 1743127117
transform -1 0 1368 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_17
timestamp 1743127117
transform 1 0 1368 0 -1 1810
box -4 -6 100 206
use NOR2X1  NOR2X1_4
timestamp 1743127117
transform -1 0 1512 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_14
timestamp 1743127117
transform -1 0 1576 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_1
timestamp 1743127117
transform 1 0 1576 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_2
timestamp 1743127117
transform -1 0 1672 0 -1 1810
box -4 -6 36 206
use MUX2X1  MUX2X1_19
timestamp 1743127117
transform 1 0 1672 0 -1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_45
timestamp 1743127117
transform 1 0 1768 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_16
timestamp 1743127117
transform 1 0 1832 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_15
timestamp 1743127117
transform -1 0 1960 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_22
timestamp 1743127117
transform -1 0 1992 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_44
timestamp 1743127117
transform -1 0 2056 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_59
timestamp 1743127117
transform 1 0 2056 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_15
timestamp 1743127117
transform -1 0 2168 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_9
timestamp 1743127117
transform -1 0 2200 0 -1 1810
box -4 -6 36 206
use DFFSR  DFFSR_18
timestamp 1743127117
transform -1 0 2552 0 -1 1810
box -4 -6 356 206
use NOR2X1  NOR2X1_57
timestamp 1743127117
transform -1 0 2600 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_13
timestamp 1743127117
transform -1 0 2664 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_1_0
timestamp 1743127117
transform 1 0 2664 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1743127117
transform 1 0 2680 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1743127117
transform 1 0 2696 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_10
timestamp 1743127117
transform 1 0 2712 0 -1 1810
box -4 -6 356 206
use BUFX4  BUFX4_98
timestamp 1743127117
transform 1 0 3064 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_24
timestamp 1743127117
transform -1 0 3176 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_80
timestamp 1743127117
transform 1 0 3176 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_12
timestamp 1743127117
transform 1 0 3240 0 -1 1810
box -4 -6 356 206
use DFFSR  DFFSR_177
timestamp 1743127117
transform -1 0 3944 0 -1 1810
box -4 -6 356 206
use MUX2X1  MUX2X1_122
timestamp 1743127117
transform 1 0 3944 0 -1 1810
box -4 -6 100 206
use BUFX4  BUFX4_6
timestamp 1743127117
transform 1 0 4040 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_2_0
timestamp 1743127117
transform -1 0 4120 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_1
timestamp 1743127117
transform -1 0 4136 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_2
timestamp 1743127117
transform -1 0 4152 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_31
timestamp 1743127117
transform -1 0 4504 0 -1 1810
box -4 -6 356 206
use NAND2X1  NAND2X1_46
timestamp 1743127117
transform 1 0 4504 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_31
timestamp 1743127117
transform 1 0 4552 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_52
timestamp 1743127117
transform -1 0 4632 0 -1 1810
box -4 -6 52 206
use MUX2X1  MUX2X1_123
timestamp 1743127117
transform 1 0 4632 0 -1 1810
box -4 -6 100 206
use MUX2X1  MUX2X1_120
timestamp 1743127117
transform 1 0 4728 0 -1 1810
box -4 -6 100 206
use INVX1  INVX1_175
timestamp 1743127117
transform -1 0 4856 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_445
timestamp 1743127117
transform -1 0 4920 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_159
timestamp 1743127117
transform -1 0 4952 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_34
timestamp 1743127117
transform 1 0 4952 0 -1 1810
box -4 -6 36 206
use BUFX4  BUFX4_77
timestamp 1743127117
transform -1 0 5048 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_32
timestamp 1743127117
transform 1 0 5048 0 -1 1810
box -4 -6 356 206
use BUFX4  BUFX4_31
timestamp 1743127117
transform -1 0 5464 0 -1 1810
box -4 -6 68 206
use BUFX4  BUFX4_80
timestamp 1743127117
transform 1 0 5464 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_37
timestamp 1743127117
transform -1 0 5560 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_172
timestamp 1743127117
transform -1 0 5624 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_49
timestamp 1743127117
transform 1 0 5624 0 -1 1810
box -4 -6 52 206
use FILL  FILL_8_3_0
timestamp 1743127117
transform -1 0 5688 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_3_1
timestamp 1743127117
transform -1 0 5704 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_3_2
timestamp 1743127117
transform -1 0 5720 0 -1 1810
box -4 -6 20 206
use MUX2X1  MUX2X1_41
timestamp 1743127117
transform -1 0 5816 0 -1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_171
timestamp 1743127117
transform -1 0 5880 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_48
timestamp 1743127117
transform -1 0 5912 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_36
timestamp 1743127117
transform -1 0 6104 0 -1 1810
box -4 -6 196 206
use INVX1  INVX1_45
timestamp 1743127117
transform -1 0 6136 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_135
timestamp 1743127117
transform 1 0 6136 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_136
timestamp 1743127117
transform -1 0 6264 0 -1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_46
timestamp 1743127117
transform 1 0 6264 0 -1 1810
box -4 -6 100 206
use NAND2X1  NAND2X1_38
timestamp 1743127117
transform -1 0 6408 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1743127117
transform 1 0 6408 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_13
timestamp 1743127117
transform -1 0 6504 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_28
timestamp 1743127117
transform -1 0 6536 0 -1 1810
box -4 -6 36 206
use DFFSR  DFFSR_35
timestamp 1743127117
transform -1 0 6888 0 -1 1810
box -4 -6 356 206
use INVX1  INVX1_100
timestamp 1743127117
transform 1 0 8 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_362
timestamp 1743127117
transform 1 0 40 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_357
timestamp 1743127117
transform -1 0 168 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_85
timestamp 1743127117
transform 1 0 168 0 1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_361
timestamp 1743127117
transform -1 0 584 0 1 1810
box -4 -6 68 206
use OR2X2  OR2X2_9
timestamp 1743127117
transform 1 0 584 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1743127117
transform 1 0 648 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_3
timestamp 1743127117
transform 1 0 696 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_2
timestamp 1743127117
transform -1 0 792 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_17
timestamp 1743127117
transform -1 0 856 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1743127117
transform 1 0 856 0 1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_3
timestamp 1743127117
transform -1 0 1096 0 1 1810
box -4 -6 52 206
use FILL  FILL_9_0_0
timestamp 1743127117
transform -1 0 1112 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1743127117
transform -1 0 1128 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1743127117
transform -1 0 1144 0 1 1810
box -4 -6 20 206
use OAI21X1  OAI21X1_8
timestamp 1743127117
transform -1 0 1208 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1743127117
transform 1 0 1208 0 1 1810
box -4 -6 196 206
use INVX1  INVX1_10
timestamp 1743127117
transform -1 0 1432 0 1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1743127117
transform 1 0 1432 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_23
timestamp 1743127117
transform 1 0 1624 0 1 1810
box -4 -6 196 206
use DFFSR  DFFSR_150
timestamp 1743127117
transform -1 0 2168 0 1 1810
box -4 -6 356 206
use NOR2X1  NOR2X1_61
timestamp 1743127117
transform -1 0 2216 0 1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_17
timestamp 1743127117
transform -1 0 2280 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_152
timestamp 1743127117
transform -1 0 2632 0 1 1810
box -4 -6 356 206
use FILL  FILL_9_1_0
timestamp 1743127117
transform -1 0 2648 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1743127117
transform -1 0 2664 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1743127117
transform -1 0 2680 0 1 1810
box -4 -6 20 206
use DFFSR  DFFSR_148
timestamp 1743127117
transform -1 0 3032 0 1 1810
box -4 -6 356 206
use INVX1  INVX1_180
timestamp 1743127117
transform -1 0 3064 0 1 1810
box -4 -6 36 206
use DFFSR  DFFSR_173
timestamp 1743127117
transform 1 0 3064 0 1 1810
box -4 -6 356 206
use NAND2X1  NAND2X1_171
timestamp 1743127117
transform -1 0 3464 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_170
timestamp 1743127117
transform -1 0 3512 0 1 1810
box -4 -6 52 206
use INVX2  INVX2_9
timestamp 1743127117
transform 1 0 3512 0 1 1810
box -4 -6 36 206
use CLKBUF1  CLKBUF1_12
timestamp 1743127117
transform -1 0 3688 0 1 1810
box -4 -6 148 206
use INVX2  INVX2_13
timestamp 1743127117
transform 1 0 3688 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_182
timestamp 1743127117
transform 1 0 3720 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_183
timestamp 1743127117
transform 1 0 3768 0 1 1810
box -4 -6 52 206
use OAI22X1  OAI22X1_7
timestamp 1743127117
transform -1 0 3896 0 1 1810
box -4 -6 84 206
use NAND2X1  NAND2X1_163
timestamp 1743127117
transform -1 0 3944 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_55
timestamp 1743127117
transform 1 0 3944 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_58
timestamp 1743127117
transform 1 0 4008 0 1 1810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_35
timestamp 1743127117
transform -1 0 4216 0 1 1810
box -4 -6 148 206
use FILL  FILL_9_2_0
timestamp 1743127117
transform -1 0 4232 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_1
timestamp 1743127117
transform -1 0 4248 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_2
timestamp 1743127117
transform -1 0 4264 0 1 1810
box -4 -6 20 206
use DFFSR  DFFSR_28
timestamp 1743127117
transform -1 0 4616 0 1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_169
timestamp 1743127117
transform -1 0 4680 0 1 1810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_34
timestamp 1743127117
transform -1 0 4824 0 1 1810
box -4 -6 148 206
use MUX2X1  MUX2X1_124
timestamp 1743127117
transform 1 0 4824 0 1 1810
box -4 -6 100 206
use INVX1  INVX1_179
timestamp 1743127117
transform -1 0 4952 0 1 1810
box -4 -6 36 206
use CLKBUF1  CLKBUF1_28
timestamp 1743127117
transform 1 0 4952 0 1 1810
box -4 -6 148 206
use BUFX4  BUFX4_3
timestamp 1743127117
transform 1 0 5096 0 1 1810
box -4 -6 68 206
use OR2X2  OR2X2_4
timestamp 1743127117
transform 1 0 5160 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1743127117
transform 1 0 5224 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_6
timestamp 1743127117
transform 1 0 5272 0 1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_29
timestamp 1743127117
transform 1 0 5384 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_146
timestamp 1743127117
transform 1 0 5576 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_145
timestamp 1743127117
transform -1 0 5704 0 1 1810
box -4 -6 68 206
use FILL  FILL_9_3_0
timestamp 1743127117
transform 1 0 5704 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_3_1
timestamp 1743127117
transform 1 0 5720 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_3_2
timestamp 1743127117
transform 1 0 5736 0 1 1810
box -4 -6 20 206
use MUX2X1  MUX2X1_51
timestamp 1743127117
transform 1 0 5752 0 1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_126
timestamp 1743127117
transform 1 0 5848 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_125
timestamp 1743127117
transform -1 0 5976 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_31
timestamp 1743127117
transform -1 0 6168 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_121
timestamp 1743127117
transform 1 0 6168 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_122
timestamp 1743127117
transform 1 0 6232 0 1 1810
box -4 -6 68 206
use MUX2X1  MUX2X1_39
timestamp 1743127117
transform -1 0 6392 0 1 1810
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_41
timestamp 1743127117
transform -1 0 6584 0 1 1810
box -4 -6 196 206
use NOR2X1  NOR2X1_18
timestamp 1743127117
transform 1 0 6584 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_29
timestamp 1743127117
transform 1 0 6632 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_20
timestamp 1743127117
transform -1 0 6712 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_133
timestamp 1743127117
transform -1 0 6776 0 1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_5
timestamp 1743127117
transform -1 0 6888 0 1 1810
box -4 -6 116 206
use INVX1  INVX1_98
timestamp 1743127117
transform 1 0 8 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_358
timestamp 1743127117
transform 1 0 40 0 -1 2210
box -4 -6 68 206
use DFFSR  DFFSR_83
timestamp 1743127117
transform 1 0 104 0 -1 2210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_40
timestamp 1743127117
transform -1 0 600 0 -1 2210
box -4 -6 148 206
use DFFSR  DFFSR_147
timestamp 1743127117
transform -1 0 952 0 -1 2210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_31
timestamp 1743127117
transform 1 0 952 0 -1 2210
box -4 -6 148 206
use FILL  FILL_10_0_0
timestamp 1743127117
transform -1 0 1112 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_1
timestamp 1743127117
transform -1 0 1128 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_2
timestamp 1743127117
transform -1 0 1144 0 -1 2210
box -4 -6 20 206
use INVX1  INVX1_7
timestamp 1743127117
transform -1 0 1176 0 -1 2210
box -4 -6 36 206
use DFFSR  DFFSR_149
timestamp 1743127117
transform -1 0 1528 0 -1 2210
box -4 -6 356 206
use DFFSR  DFFSR_162
timestamp 1743127117
transform -1 0 1880 0 -1 2210
box -4 -6 356 206
use DFFSR  DFFSR_151
timestamp 1743127117
transform 1 0 1880 0 -1 2210
box -4 -6 356 206
use NOR2X1  NOR2X1_60
timestamp 1743127117
transform 1 0 2232 0 -1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_16
timestamp 1743127117
transform -1 0 2344 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_161
timestamp 1743127117
transform 1 0 2344 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_55
timestamp 1743127117
transform 1 0 2392 0 -1 2210
box -4 -6 52 206
use BUFX4  BUFX4_68
timestamp 1743127117
transform -1 0 2504 0 -1 2210
box -4 -6 68 206
use BUFX4  BUFX4_66
timestamp 1743127117
transform -1 0 2568 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_157
timestamp 1743127117
transform -1 0 2600 0 -1 2210
box -4 -6 36 206
use FILL  FILL_10_1_0
timestamp 1743127117
transform 1 0 2600 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_1
timestamp 1743127117
transform 1 0 2616 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_2
timestamp 1743127117
transform 1 0 2632 0 -1 2210
box -4 -6 20 206
use DFFSR  DFFSR_171
timestamp 1743127117
transform 1 0 2648 0 -1 2210
box -4 -6 356 206
use NAND2X1  NAND2X1_168
timestamp 1743127117
transform 1 0 3000 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_453
timestamp 1743127117
transform 1 0 3048 0 -1 2210
box -4 -6 68 206
use INVX4  INVX4_3
timestamp 1743127117
transform 1 0 3112 0 -1 2210
box -4 -6 52 206
use INVX4  INVX4_5
timestamp 1743127117
transform -1 0 3208 0 -1 2210
box -4 -6 52 206
use BUFX4  BUFX4_67
timestamp 1743127117
transform 1 0 3208 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_455
timestamp 1743127117
transform -1 0 3336 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_166
timestamp 1743127117
transform -1 0 3384 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_169
timestamp 1743127117
transform -1 0 3432 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_448
timestamp 1743127117
transform 1 0 3432 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_173
timestamp 1743127117
transform -1 0 3544 0 -1 2210
box -4 -6 52 206
use DFFSR  DFFSR_174
timestamp 1743127117
transform -1 0 3896 0 -1 2210
box -4 -6 356 206
use BUFX4  BUFX4_58
timestamp 1743127117
transform -1 0 3960 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_157
timestamp 1743127117
transform 1 0 3960 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_2_0
timestamp 1743127117
transform 1 0 4024 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_1
timestamp 1743127117
transform 1 0 4040 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_2
timestamp 1743127117
transform 1 0 4056 0 -1 2210
box -4 -6 20 206
use DFFSR  DFFSR_158
timestamp 1743127117
transform 1 0 4072 0 -1 2210
box -4 -6 356 206
use BUFX4  BUFX4_60
timestamp 1743127117
transform 1 0 4424 0 -1 2210
box -4 -6 68 206
use DFFSR  DFFSR_21
timestamp 1743127117
transform -1 0 4840 0 -1 2210
box -4 -6 356 206
use INVX1  INVX1_27
timestamp 1743127117
transform 1 0 4840 0 -1 2210
box -4 -6 36 206
use DFFSR  DFFSR_20
timestamp 1743127117
transform 1 0 4872 0 -1 2210
box -4 -6 356 206
use OAI21X1  OAI21X1_109
timestamp 1743127117
transform 1 0 5224 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_37
timestamp 1743127117
transform -1 0 5336 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_112
timestamp 1743127117
transform -1 0 5400 0 -1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_11
timestamp 1743127117
transform 1 0 5400 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_12
timestamp 1743127117
transform -1 0 5496 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_110
timestamp 1743127117
transform 1 0 5496 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_2
timestamp 1743127117
transform -1 0 5624 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_8
timestamp 1743127117
transform -1 0 5688 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_3_0
timestamp 1743127117
transform -1 0 5704 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_3_1
timestamp 1743127117
transform -1 0 5720 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_3_2
timestamp 1743127117
transform -1 0 5736 0 -1 2210
box -4 -6 20 206
use OR2X2  OR2X2_3
timestamp 1743127117
transform -1 0 5800 0 -1 2210
box -4 -6 68 206
use XOR2X1  XOR2X1_3
timestamp 1743127117
transform 1 0 5800 0 -1 2210
box -4 -6 116 206
use MUX2X1  MUX2X1_33
timestamp 1743127117
transform 1 0 5912 0 -1 2210
box -4 -6 100 206
use MUX2X1  MUX2X1_34
timestamp 1743127117
transform 1 0 6008 0 -1 2210
box -4 -6 100 206
use DFFSR  DFFSR_37
timestamp 1743127117
transform -1 0 6456 0 -1 2210
box -4 -6 356 206
use XNOR2X1  XNOR2X1_4
timestamp 1743127117
transform 1 0 6456 0 -1 2210
box -4 -6 116 206
use CLKBUF1  CLKBUF1_15
timestamp 1743127117
transform 1 0 6568 0 -1 2210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_42
timestamp 1743127117
transform 1 0 6712 0 -1 2210
box -4 -6 148 206
use FILL  FILL_11_1
timestamp 1743127117
transform -1 0 6872 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_2
timestamp 1743127117
transform -1 0 6888 0 -1 2210
box -4 -6 20 206
use CLKBUF1  CLKBUF1_11
timestamp 1743127117
transform -1 0 152 0 1 2210
box -4 -6 148 206
use INVX1  INVX1_169
timestamp 1743127117
transform -1 0 184 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_54
timestamp 1743127117
transform 1 0 184 0 1 2210
box -4 -6 36 206
use DFFSR  DFFSR_160
timestamp 1743127117
transform -1 0 568 0 1 2210
box -4 -6 356 206
use MUX2X1  MUX2X1_114
timestamp 1743127117
transform -1 0 664 0 1 2210
box -4 -6 100 206
use NOR2X1  NOR2X1_56
timestamp 1743127117
transform 1 0 664 0 1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_12
timestamp 1743127117
transform -1 0 776 0 1 2210
box -4 -6 68 206
use MUX2X1  MUX2X1_113
timestamp 1743127117
transform 1 0 776 0 1 2210
box -4 -6 100 206
use DFFSR  DFFSR_161
timestamp 1743127117
transform 1 0 872 0 1 2210
box -4 -6 356 206
use FILL  FILL_11_0_0
timestamp 1743127117
transform -1 0 1240 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_1
timestamp 1743127117
transform -1 0 1256 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_2
timestamp 1743127117
transform -1 0 1272 0 1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_58
timestamp 1743127117
transform -1 0 1320 0 1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_14
timestamp 1743127117
transform -1 0 1384 0 1 2210
box -4 -6 68 206
use DFFSR  DFFSR_164
timestamp 1743127117
transform -1 0 1736 0 1 2210
box -4 -6 356 206
use INVX1  INVX1_171
timestamp 1743127117
transform 1 0 1736 0 1 2210
box -4 -6 36 206
use MUX2X1  MUX2X1_116
timestamp 1743127117
transform -1 0 1864 0 1 2210
box -4 -6 100 206
use DFFSR  DFFSR_143
timestamp 1743127117
transform -1 0 2216 0 1 2210
box -4 -6 356 206
use MUX2X1  MUX2X1_117
timestamp 1743127117
transform -1 0 2312 0 1 2210
box -4 -6 100 206
use OAI21X1  OAI21X1_446
timestamp 1743127117
transform -1 0 2376 0 1 2210
box -4 -6 68 206
use DFFSR  DFFSR_172
timestamp 1743127117
transform 1 0 2376 0 1 2210
box -4 -6 356 206
use FILL  FILL_11_1_0
timestamp 1743127117
transform -1 0 2744 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_1
timestamp 1743127117
transform -1 0 2760 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_2
timestamp 1743127117
transform -1 0 2776 0 1 2210
box -4 -6 20 206
use OR2X2  OR2X2_13
timestamp 1743127117
transform -1 0 2840 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_183
timestamp 1743127117
transform -1 0 2872 0 1 2210
box -4 -6 36 206
use INVX2  INVX2_8
timestamp 1743127117
transform 1 0 2872 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_167
timestamp 1743127117
transform 1 0 2904 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_452
timestamp 1743127117
transform -1 0 3016 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_181
timestamp 1743127117
transform 1 0 3016 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_454
timestamp 1743127117
transform 1 0 3048 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_456
timestamp 1743127117
transform 1 0 3112 0 1 2210
box -4 -6 68 206
use DFFSR  DFFSR_178
timestamp 1743127117
transform 1 0 3176 0 1 2210
box -4 -6 356 206
use INVX2  INVX2_10
timestamp 1743127117
transform 1 0 3528 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_174
timestamp 1743127117
transform 1 0 3560 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_457
timestamp 1743127117
transform -1 0 3672 0 1 2210
box -4 -6 68 206
use BUFX4  BUFX4_71
timestamp 1743127117
transform 1 0 3672 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_61
timestamp 1743127117
transform -1 0 3800 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_64
timestamp 1743127117
transform -1 0 3864 0 1 2210
box -4 -6 68 206
use DFFSR  DFFSR_155
timestamp 1743127117
transform 1 0 3864 0 1 2210
box -4 -6 356 206
use FILL  FILL_11_2_0
timestamp 1743127117
transform 1 0 4216 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_1
timestamp 1743127117
transform 1 0 4232 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_2
timestamp 1743127117
transform 1 0 4248 0 1 2210
box -4 -6 20 206
use MUX2X1  MUX2X1_121
timestamp 1743127117
transform 1 0 4264 0 1 2210
box -4 -6 100 206
use INVX1  INVX1_176
timestamp 1743127117
transform 1 0 4360 0 1 2210
box -4 -6 36 206
use CLKBUF1  CLKBUF1_29
timestamp 1743127117
transform 1 0 4392 0 1 2210
box -4 -6 148 206
use DFFSR  DFFSR_153
timestamp 1743127117
transform 1 0 4536 0 1 2210
box -4 -6 356 206
use MUX2X1  MUX2X1_119
timestamp 1743127117
transform 1 0 4888 0 1 2210
box -4 -6 100 206
use INVX1  INVX1_174
timestamp 1743127117
transform -1 0 5016 0 1 2210
box -4 -6 36 206
use DFFSR  DFFSR_38
timestamp 1743127117
transform 1 0 5016 0 1 2210
box -4 -6 356 206
use INVX1  INVX1_35
timestamp 1743127117
transform -1 0 5400 0 1 2210
box -4 -6 36 206
use AND2X2  AND2X2_2
timestamp 1743127117
transform 1 0 5400 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_25
timestamp 1743127117
transform 1 0 5464 0 1 2210
box -4 -6 36 206
use BUFX2  BUFX2_20
timestamp 1743127117
transform -1 0 5544 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_111
timestamp 1743127117
transform -1 0 5608 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_36
timestamp 1743127117
transform 1 0 5608 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_35
timestamp 1743127117
transform -1 0 5704 0 1 2210
box -4 -6 52 206
use FILL  FILL_11_3_0
timestamp 1743127117
transform -1 0 5720 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_3_1
timestamp 1743127117
transform -1 0 5736 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_3_2
timestamp 1743127117
transform -1 0 5752 0 1 2210
box -4 -6 20 206
use DFFSR  DFFSR_36
timestamp 1743127117
transform -1 0 6104 0 1 2210
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_84
timestamp 1743127117
transform -1 0 6296 0 1 2210
box -4 -6 196 206
use DFFSR  DFFSR_34
timestamp 1743127117
transform 1 0 6296 0 1 2210
box -4 -6 356 206
use INVX1  INVX1_77
timestamp 1743127117
transform 1 0 6648 0 1 2210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_26
timestamp 1743127117
transform 1 0 6680 0 1 2210
box -4 -6 196 206
use FILL  FILL_12_1
timestamp 1743127117
transform 1 0 6872 0 1 2210
box -4 -6 20 206
use BUFX2  BUFX2_17
timestamp 1743127117
transform -1 0 56 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_16
timestamp 1743127117
transform -1 0 104 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_130
timestamp 1743127117
transform 1 0 104 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_107
timestamp 1743127117
transform -1 0 488 0 -1 2610
box -4 -6 356 206
use DFFSR  DFFSR_108
timestamp 1743127117
transform -1 0 840 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_168
timestamp 1743127117
transform -1 0 872 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_159
timestamp 1743127117
transform -1 0 1224 0 -1 2610
box -4 -6 356 206
use FILL  FILL_12_0_0
timestamp 1743127117
transform -1 0 1240 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_1
timestamp 1743127117
transform -1 0 1256 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_2
timestamp 1743127117
transform -1 0 1272 0 -1 2610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_24
timestamp 1743127117
transform -1 0 1416 0 -1 2610
box -4 -6 148 206
use CLKBUF1  CLKBUF1_38
timestamp 1743127117
transform 1 0 1416 0 -1 2610
box -4 -6 148 206
use INVX1  INVX1_170
timestamp 1743127117
transform 1 0 1560 0 -1 2610
box -4 -6 36 206
use MUX2X1  MUX2X1_115
timestamp 1743127117
transform -1 0 1688 0 -1 2610
box -4 -6 100 206
use INVX1  INVX1_173
timestamp 1743127117
transform 1 0 1688 0 -1 2610
box -4 -6 36 206
use MUX2X1  MUX2X1_118
timestamp 1743127117
transform -1 0 1816 0 -1 2610
box -4 -6 100 206
use INVX1  INVX1_132
timestamp 1743127117
transform 1 0 1816 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_110
timestamp 1743127117
transform 1 0 1848 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_172
timestamp 1743127117
transform 1 0 2200 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_163
timestamp 1743127117
transform -1 0 2584 0 -1 2610
box -4 -6 356 206
use INVX1  INVX1_161
timestamp 1743127117
transform 1 0 2584 0 -1 2610
box -4 -6 36 206
use FILL  FILL_12_1_0
timestamp 1743127117
transform 1 0 2616 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_1
timestamp 1743127117
transform 1 0 2632 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_2
timestamp 1743127117
transform 1 0 2648 0 -1 2610
box -4 -6 20 206
use OAI21X1  OAI21X1_450
timestamp 1743127117
transform 1 0 2664 0 -1 2610
box -4 -6 68 206
use DFFSR  DFFSR_141
timestamp 1743127117
transform -1 0 3080 0 -1 2610
box -4 -6 356 206
use NAND3X1  NAND3X1_57
timestamp 1743127117
transform 1 0 3080 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_60
timestamp 1743127117
transform 1 0 3144 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_451
timestamp 1743127117
transform -1 0 3272 0 -1 2610
box -4 -6 68 206
use OAI22X1  OAI22X1_9
timestamp 1743127117
transform -1 0 3352 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_164
timestamp 1743127117
transform 1 0 3352 0 -1 2610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_19
timestamp 1743127117
transform -1 0 3544 0 -1 2610
box -4 -6 148 206
use OAI21X1  OAI21X1_449
timestamp 1743127117
transform -1 0 3608 0 -1 2610
box -4 -6 68 206
use OAI22X1  OAI22X1_8
timestamp 1743127117
transform 1 0 3608 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_172
timestamp 1743127117
transform 1 0 3688 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_463
timestamp 1743127117
transform 1 0 3736 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_54
timestamp 1743127117
transform 1 0 3800 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_53
timestamp 1743127117
transform 1 0 3848 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_160
timestamp 1743127117
transform -1 0 3944 0 -1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_175
timestamp 1743127117
transform -1 0 3992 0 -1 2610
box -4 -6 52 206
use BUFX4  BUFX4_9
timestamp 1743127117
transform 1 0 3992 0 -1 2610
box -4 -6 68 206
use OR2X2  OR2X2_14
timestamp 1743127117
transform -1 0 4120 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_59
timestamp 1743127117
transform 1 0 4120 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_2_0
timestamp 1743127117
transform 1 0 4184 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_1
timestamp 1743127117
transform 1 0 4200 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_2
timestamp 1743127117
transform 1 0 4216 0 -1 2610
box -4 -6 20 206
use DFFSR  DFFSR_169
timestamp 1743127117
transform 1 0 4232 0 -1 2610
box -4 -6 356 206
use MUX2X1  MUX2X1_109
timestamp 1743127117
transform 1 0 4584 0 -1 2610
box -4 -6 100 206
use INVX1  INVX1_164
timestamp 1743127117
transform -1 0 4712 0 -1 2610
box -4 -6 36 206
use CLKBUF1  CLKBUF1_30
timestamp 1743127117
transform -1 0 4856 0 -1 2610
box -4 -6 148 206
use MUX2X1  MUX2X1_112
timestamp 1743127117
transform 1 0 4856 0 -1 2610
box -4 -6 100 206
use INVX1  INVX1_167
timestamp 1743127117
transform -1 0 4984 0 -1 2610
box -4 -6 36 206
use MUX2X1  MUX2X1_107
timestamp 1743127117
transform 1 0 4984 0 -1 2610
box -4 -6 100 206
use INVX1  INVX1_162
timestamp 1743127117
transform -1 0 5112 0 -1 2610
box -4 -6 36 206
use DFFSR  DFFSR_165
timestamp 1743127117
transform 1 0 5112 0 -1 2610
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_93
timestamp 1743127117
transform -1 0 5656 0 -1 2610
box -4 -6 196 206
use OAI21X1  OAI21X1_308
timestamp 1743127117
transform 1 0 5656 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_3_0
timestamp 1743127117
transform -1 0 5736 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_3_1
timestamp 1743127117
transform -1 0 5752 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_3_2
timestamp 1743127117
transform -1 0 5768 0 -1 2610
box -4 -6 20 206
use OAI21X1  OAI21X1_307
timestamp 1743127117
transform -1 0 5832 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_81
timestamp 1743127117
transform 1 0 5832 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_88
timestamp 1743127117
transform -1 0 6216 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_75
timestamp 1743127117
transform -1 0 6408 0 -1 2610
box -4 -6 196 206
use OAI21X1  OAI21X1_313
timestamp 1743127117
transform -1 0 6472 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_314
timestamp 1743127117
transform -1 0 6536 0 -1 2610
box -4 -6 68 206
use MUX2X1  MUX2X1_104
timestamp 1743127117
transform -1 0 6632 0 -1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_326
timestamp 1743127117
transform 1 0 6632 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_78
timestamp 1743127117
transform 1 0 6696 0 -1 2610
box -4 -6 196 206
use DFFSR  DFFSR_112
timestamp 1743127117
transform 1 0 8 0 1 2610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_9
timestamp 1743127117
transform -1 0 504 0 1 2610
box -4 -6 148 206
use OAI21X1  OAI21X1_406
timestamp 1743127117
transform -1 0 568 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_131
timestamp 1743127117
transform 1 0 568 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_407
timestamp 1743127117
transform 1 0 600 0 1 2610
box -4 -6 68 206
use DFFSR  DFFSR_115
timestamp 1743127117
transform -1 0 1016 0 1 2610
box -4 -6 356 206
use INVX1  INVX1_58
timestamp 1743127117
transform -1 0 1048 0 1 2610
box -4 -6 36 206
use INVX1  INVX1_57
timestamp 1743127117
transform -1 0 1080 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_126
timestamp 1743127117
transform -1 0 1128 0 1 2610
box -4 -6 52 206
use FILL  FILL_13_0_0
timestamp 1743127117
transform -1 0 1144 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_1
timestamp 1743127117
transform -1 0 1160 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_2
timestamp 1743127117
transform -1 0 1176 0 1 2610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_3
timestamp 1743127117
transform -1 0 1320 0 1 2610
box -4 -6 148 206
use INVX1  INVX1_56
timestamp 1743127117
transform -1 0 1352 0 1 2610
box -4 -6 36 206
use DFFSR  DFFSR_43
timestamp 1743127117
transform -1 0 1704 0 1 2610
box -4 -6 356 206
use NAND2X1  NAND2X1_83
timestamp 1743127117
transform -1 0 1752 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_266
timestamp 1743127117
transform -1 0 1816 0 1 2610
box -4 -6 68 206
use BUFX4  BUFX4_1
timestamp 1743127117
transform -1 0 1880 0 1 2610
box -4 -6 68 206
use DFFSR  DFFSR_118
timestamp 1743127117
transform -1 0 2232 0 1 2610
box -4 -6 356 206
use NOR2X1  NOR2X1_25
timestamp 1743127117
transform -1 0 2280 0 1 2610
box -4 -6 52 206
use DFFSR  DFFSR_145
timestamp 1743127117
transform -1 0 2632 0 1 2610
box -4 -6 356 206
use FILL  FILL_13_1_0
timestamp 1743127117
transform 1 0 2632 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_1
timestamp 1743127117
transform 1 0 2648 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_2
timestamp 1743127117
transform 1 0 2664 0 1 2610
box -4 -6 20 206
use BUFX4  BUFX4_69
timestamp 1743127117
transform 1 0 2680 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_63
timestamp 1743127117
transform -1 0 2808 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_458
timestamp 1743127117
transform -1 0 2872 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_459
timestamp 1743127117
transform 1 0 2872 0 1 2610
box -4 -6 68 206
use DFFSR  DFFSR_176
timestamp 1743127117
transform 1 0 2936 0 1 2610
box -4 -6 356 206
use NAND2X1  NAND2X1_165
timestamp 1743127117
transform 1 0 3288 0 1 2610
box -4 -6 52 206
use INVX2  INVX2_12
timestamp 1743127117
transform -1 0 3368 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_179
timestamp 1743127117
transform 1 0 3368 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_180
timestamp 1743127117
transform 1 0 3416 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_462
timestamp 1743127117
transform -1 0 3528 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_185
timestamp 1743127117
transform -1 0 3560 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_461
timestamp 1743127117
transform 1 0 3560 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_460
timestamp 1743127117
transform -1 0 3688 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_184
timestamp 1743127117
transform -1 0 3720 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_181
timestamp 1743127117
transform 1 0 3720 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_52
timestamp 1743127117
transform 1 0 3768 0 1 2610
box -4 -6 68 206
use INVX8  INVX8_9
timestamp 1743127117
transform 1 0 3832 0 1 2610
box -4 -6 84 206
use BUFX4  BUFX4_70
timestamp 1743127117
transform 1 0 3912 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_1
timestamp 1743127117
transform 1 0 3976 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_65
timestamp 1743127117
transform 1 0 4024 0 1 2610
box -4 -6 68 206
use MUX2X1  MUX2X1_111
timestamp 1743127117
transform 1 0 4088 0 1 2610
box -4 -6 100 206
use FILL  FILL_13_2_0
timestamp 1743127117
transform -1 0 4200 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_1
timestamp 1743127117
transform -1 0 4216 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_2
timestamp 1743127117
transform -1 0 4232 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_166
timestamp 1743127117
transform -1 0 4264 0 1 2610
box -4 -6 36 206
use DFFSR  DFFSR_167
timestamp 1743127117
transform 1 0 4264 0 1 2610
box -4 -6 356 206
use INVX1  INVX1_79
timestamp 1743127117
transform 1 0 4616 0 1 2610
box -4 -6 36 206
use DFFSR  DFFSR_170
timestamp 1743127117
transform 1 0 4648 0 1 2610
box -4 -6 356 206
use INVX1  INVX1_82
timestamp 1743127117
transform 1 0 5000 0 1 2610
box -4 -6 36 206
use INVX1  INVX1_75
timestamp 1743127117
transform -1 0 5064 0 1 2610
box -4 -6 36 206
use CLKBUF1  CLKBUF1_25
timestamp 1743127117
transform 1 0 5064 0 1 2610
box -4 -6 148 206
use OAI21X1  OAI21X1_277
timestamp 1743127117
transform -1 0 5272 0 1 2610
box -4 -6 68 206
use BUFX4  BUFX4_46
timestamp 1743127117
transform -1 0 5336 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_274
timestamp 1743127117
transform 1 0 5336 0 1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_92
timestamp 1743127117
transform 1 0 5400 0 1 2610
box -4 -6 196 206
use NAND2X1  NAND2X1_101
timestamp 1743127117
transform -1 0 5640 0 1 2610
box -4 -6 52 206
use MUX2X1  MUX2X1_95
timestamp 1743127117
transform -1 0 5736 0 1 2610
box -4 -6 100 206
use FILL  FILL_13_3_0
timestamp 1743127117
transform -1 0 5752 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_3_1
timestamp 1743127117
transform -1 0 5768 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_3_2
timestamp 1743127117
transform -1 0 5784 0 1 2610
box -4 -6 20 206
use MUX2X1  MUX2X1_101
timestamp 1743127117
transform -1 0 5880 0 1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_297
timestamp 1743127117
transform -1 0 5944 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_298
timestamp 1743127117
transform -1 0 6008 0 1 2610
box -4 -6 68 206
use BUFX4  BUFX4_47
timestamp 1743127117
transform 1 0 6008 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_319
timestamp 1743127117
transform 1 0 6072 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_320
timestamp 1743127117
transform -1 0 6200 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_96
timestamp 1743127117
transform -1 0 6232 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_107
timestamp 1743127117
transform -1 0 6280 0 1 2610
box -4 -6 52 206
use MUX2X1  MUX2X1_98
timestamp 1743127117
transform 1 0 6280 0 1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_325
timestamp 1743127117
transform 1 0 6376 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_321
timestamp 1743127117
transform 1 0 6440 0 1 2610
box -4 -6 68 206
use MUX2X1  MUX2X1_102
timestamp 1743127117
transform -1 0 6600 0 1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_322
timestamp 1743127117
transform -1 0 6664 0 1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_76
timestamp 1743127117
transform -1 0 6856 0 1 2610
box -4 -6 196 206
use FILL  FILL_14_1
timestamp 1743127117
transform 1 0 6856 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_2
timestamp 1743127117
transform 1 0 6872 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_123
timestamp 1743127117
transform 1 0 8 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_394
timestamp 1743127117
transform 1 0 40 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_393
timestamp 1743127117
transform -1 0 168 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_58
timestamp 1743127117
transform -1 0 216 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_183
timestamp 1743127117
transform -1 0 280 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_399
timestamp 1743127117
transform 1 0 280 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_400
timestamp 1743127117
transform -1 0 408 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_126
timestamp 1743127117
transform -1 0 440 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_61
timestamp 1743127117
transform 1 0 440 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_192
timestamp 1743127117
transform -1 0 552 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_195
timestamp 1743127117
transform -1 0 616 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_46
timestamp 1743127117
transform 1 0 616 0 -1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_72
timestamp 1743127117
transform -1 0 1016 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_242
timestamp 1743127117
transform -1 0 1080 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_82
timestamp 1743127117
transform -1 0 1128 0 -1 3010
box -4 -6 52 206
use FILL  FILL_14_0_0
timestamp 1743127117
transform 1 0 1128 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_1
timestamp 1743127117
transform 1 0 1144 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_2
timestamp 1743127117
transform 1 0 1160 0 -1 3010
box -4 -6 20 206
use DFFSR  DFFSR_47
timestamp 1743127117
transform 1 0 1176 0 -1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_74
timestamp 1743127117
transform -1 0 1576 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_246
timestamp 1743127117
transform -1 0 1640 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_48
timestamp 1743127117
transform 1 0 1640 0 -1 3010
box -4 -6 356 206
use OAI21X1  OAI21X1_250
timestamp 1743127117
transform 1 0 1992 0 -1 3010
box -4 -6 68 206
use DFFSR  DFFSR_175
timestamp 1743127117
transform 1 0 2056 0 -1 3010
box -4 -6 356 206
use INVX2  INVX2_11
timestamp 1743127117
transform 1 0 2408 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_176
timestamp 1743127117
transform 1 0 2440 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_177
timestamp 1743127117
transform 1 0 2488 0 -1 3010
box -4 -6 52 206
use FILL  FILL_14_1_0
timestamp 1743127117
transform 1 0 2536 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_1
timestamp 1743127117
transform 1 0 2552 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_2
timestamp 1743127117
transform 1 0 2568 0 -1 3010
box -4 -6 20 206
use DFFSR  DFFSR_133
timestamp 1743127117
transform 1 0 2584 0 -1 3010
box -4 -6 356 206
use NAND3X1  NAND3X1_54
timestamp 1743127117
transform 1 0 2936 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_26
timestamp 1743127117
transform 1 0 3000 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_66
timestamp 1743127117
transform -1 0 3112 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_69
timestamp 1743127117
transform -1 0 3176 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_67
timestamp 1743127117
transform -1 0 3240 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_178
timestamp 1743127117
transform -1 0 3288 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_71
timestamp 1743127117
transform -1 0 3352 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_56
timestamp 1743127117
transform 1 0 3352 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_70
timestamp 1743127117
transform -1 0 3480 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_62
timestamp 1743127117
transform 1 0 3480 0 -1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_110
timestamp 1743127117
transform -1 0 3640 0 -1 3010
box -4 -6 100 206
use INVX1  INVX1_165
timestamp 1743127117
transform -1 0 3672 0 -1 3010
box -4 -6 36 206
use DFFSR  DFFSR_168
timestamp 1743127117
transform -1 0 4024 0 -1 3010
box -4 -6 356 206
use MUX2X1  MUX2X1_108
timestamp 1743127117
transform 1 0 4024 0 -1 3010
box -4 -6 100 206
use INVX1  INVX1_163
timestamp 1743127117
transform -1 0 4152 0 -1 3010
box -4 -6 36 206
use FILL  FILL_14_2_0
timestamp 1743127117
transform 1 0 4152 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_1
timestamp 1743127117
transform 1 0 4168 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_2
timestamp 1743127117
transform 1 0 4184 0 -1 3010
box -4 -6 20 206
use DFFSR  DFFSR_146
timestamp 1743127117
transform 1 0 4200 0 -1 3010
box -4 -6 356 206
use OAI21X1  OAI21X1_444
timestamp 1743127117
transform -1 0 4616 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_158
timestamp 1743127117
transform -1 0 4648 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_275
timestamp 1743127117
transform 1 0 4648 0 -1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_88
timestamp 1743127117
transform -1 0 4808 0 -1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_294
timestamp 1743127117
transform 1 0 4808 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_86
timestamp 1743127117
transform -1 0 5064 0 -1 3010
box -4 -6 196 206
use INVX1  INVX1_74
timestamp 1743127117
transform 1 0 5064 0 -1 3010
box -4 -6 36 206
use MUX2X1  MUX2X1_81
timestamp 1743127117
transform -1 0 5192 0 -1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_276
timestamp 1743127117
transform -1 0 5256 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_273
timestamp 1743127117
transform 1 0 5256 0 -1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_80
timestamp 1743127117
transform 1 0 5320 0 -1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_337
timestamp 1743127117
transform -1 0 5480 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_90
timestamp 1743127117
transform -1 0 5512 0 -1 3010
box -4 -6 36 206
use BUFX4  BUFX4_22
timestamp 1743127117
transform 1 0 5512 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_74
timestamp 1743127117
transform 1 0 5576 0 -1 3010
box -4 -6 196 206
use FILL  FILL_14_3_0
timestamp 1743127117
transform 1 0 5768 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_3_1
timestamp 1743127117
transform 1 0 5784 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_3_2
timestamp 1743127117
transform 1 0 5800 0 -1 3010
box -4 -6 20 206
use MUX2X1  MUX2X1_90
timestamp 1743127117
transform 1 0 5816 0 -1 3010
box -4 -6 100 206
use MUX2X1  MUX2X1_100
timestamp 1743127117
transform 1 0 5912 0 -1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_318
timestamp 1743127117
transform 1 0 6008 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_317
timestamp 1743127117
transform -1 0 6136 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_349
timestamp 1743127117
transform -1 0 6200 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_341
timestamp 1743127117
transform -1 0 6264 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_103
timestamp 1743127117
transform -1 0 6312 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_92
timestamp 1743127117
transform -1 0 6344 0 -1 3010
box -4 -6 36 206
use MUX2X1  MUX2X1_96
timestamp 1743127117
transform 1 0 6344 0 -1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_309
timestamp 1743127117
transform 1 0 6440 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_82
timestamp 1743127117
transform -1 0 6696 0 -1 3010
box -4 -6 196 206
use CLKBUF1  CLKBUF1_7
timestamp 1743127117
transform 1 0 6696 0 -1 3010
box -4 -6 148 206
use FILL  FILL_15_1
timestamp 1743127117
transform -1 0 6856 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_2
timestamp 1743127117
transform -1 0 6872 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_3
timestamp 1743127117
transform -1 0 6888 0 -1 3010
box -4 -6 20 206
use DFFSR  DFFSR_116
timestamp 1743127117
transform 1 0 8 0 1 3010
box -4 -6 356 206
use OAI21X1  OAI21X1_401
timestamp 1743127117
transform 1 0 360 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_402
timestamp 1743127117
transform -1 0 488 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_127
timestamp 1743127117
transform -1 0 520 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_62
timestamp 1743127117
transform -1 0 568 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_127
timestamp 1743127117
transform 1 0 568 0 1 3010
box -4 -6 52 206
use DFFSR  DFFSR_51
timestamp 1743127117
transform 1 0 616 0 1 3010
box -4 -6 356 206
use INVX1  INVX1_51
timestamp 1743127117
transform -1 0 1000 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_17
timestamp 1743127117
transform 1 0 1000 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_0_0
timestamp 1743127117
transform 1 0 1064 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_1
timestamp 1743127117
transform 1 0 1080 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_2
timestamp 1743127117
transform 1 0 1096 0 1 3010
box -4 -6 20 206
use DFFSR  DFFSR_42
timestamp 1743127117
transform 1 0 1112 0 1 3010
box -4 -6 356 206
use OAI21X1  OAI21X1_265
timestamp 1743127117
transform -1 0 1528 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_125
timestamp 1743127117
transform -1 0 1576 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_55
timestamp 1743127117
transform 1 0 1576 0 1 3010
box -4 -6 36 206
use BUFX4  BUFX4_30
timestamp 1743127117
transform -1 0 1672 0 1 3010
box -4 -6 68 206
use DFFSR  DFFSR_44
timestamp 1743127117
transform -1 0 2024 0 1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_76
timestamp 1743127117
transform 1 0 2024 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_84
timestamp 1743127117
transform -1 0 2120 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_267
timestamp 1743127117
transform -1 0 2184 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_2
timestamp 1743127117
transform -1 0 2232 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_26
timestamp 1743127117
transform 1 0 2232 0 1 3010
box -4 -6 68 206
use INVX8  INVX8_7
timestamp 1743127117
transform -1 0 2376 0 1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_70
timestamp 1743127117
transform -1 0 2424 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_238
timestamp 1743127117
transform 1 0 2424 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_1_0
timestamp 1743127117
transform 1 0 2488 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_1
timestamp 1743127117
transform 1 0 2504 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_2
timestamp 1743127117
transform 1 0 2520 0 1 3010
box -4 -6 20 206
use DFFSR  DFFSR_45
timestamp 1743127117
transform 1 0 2536 0 1 3010
box -4 -6 356 206
use INVX4  INVX4_2
timestamp 1743127117
transform 1 0 2888 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_160
timestamp 1743127117
transform -1 0 2984 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_443
timestamp 1743127117
transform 1 0 2984 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_156
timestamp 1743127117
transform -1 0 3080 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_153
timestamp 1743127117
transform 1 0 3080 0 1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_45
timestamp 1743127117
transform -1 0 3192 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_154
timestamp 1743127117
transform -1 0 3240 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_7
timestamp 1743127117
transform 1 0 3240 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_68
timestamp 1743127117
transform 1 0 3304 0 1 3010
box -4 -6 68 206
use BUFX4  BUFX4_8
timestamp 1743127117
transform -1 0 3432 0 1 3010
box -4 -6 68 206
use INVX4  INVX4_4
timestamp 1743127117
transform 1 0 3432 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_162
timestamp 1743127117
transform 1 0 3480 0 1 3010
box -4 -6 52 206
use OAI22X1  OAI22X1_6
timestamp 1743127117
transform 1 0 3528 0 1 3010
box -4 -6 84 206
use OAI21X1  OAI21X1_447
timestamp 1743127117
transform 1 0 3608 0 1 3010
box -4 -6 68 206
use DFFSR  DFFSR_142
timestamp 1743127117
transform -1 0 4024 0 1 3010
box -4 -6 356 206
use FILL  FILL_15_2_0
timestamp 1743127117
transform 1 0 4024 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_1
timestamp 1743127117
transform 1 0 4040 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_2
timestamp 1743127117
transform 1 0 4056 0 1 3010
box -4 -6 20 206
use DFFSR  DFFSR_166
timestamp 1743127117
transform 1 0 4072 0 1 3010
box -4 -6 356 206
use INVX1  INVX1_80
timestamp 1743127117
transform 1 0 4424 0 1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_87
timestamp 1743127117
transform 1 0 4456 0 1 3010
box -4 -6 196 206
use INVX1  INVX1_81
timestamp 1743127117
transform 1 0 4648 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_278
timestamp 1743127117
transform 1 0 4680 0 1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_89
timestamp 1743127117
transform -1 0 4840 0 1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_296
timestamp 1743127117
transform 1 0 4840 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_295
timestamp 1743127117
transform -1 0 4968 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_293
timestamp 1743127117
transform -1 0 5032 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_89
timestamp 1743127117
transform 1 0 5032 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_268
timestamp 1743127117
transform -1 0 5128 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_34
timestamp 1743127117
transform 1 0 5128 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_81
timestamp 1743127117
transform 1 0 5176 0 1 3010
box -4 -6 68 206
use BUFX4  BUFX4_19
timestamp 1743127117
transform -1 0 5304 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_336
timestamp 1743127117
transform 1 0 5304 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_338
timestamp 1743127117
transform 1 0 5368 0 1 3010
box -4 -6 68 206
use BUFX4  BUFX4_20
timestamp 1743127117
transform 1 0 5432 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_342
timestamp 1743127117
transform -1 0 5560 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_284
timestamp 1743127117
transform 1 0 5560 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_340
timestamp 1743127117
transform -1 0 5688 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_91
timestamp 1743127117
transform -1 0 5720 0 1 3010
box -4 -6 36 206
use FILL  FILL_15_3_0
timestamp 1743127117
transform 1 0 5720 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_3_1
timestamp 1743127117
transform 1 0 5736 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_3_2
timestamp 1743127117
transform 1 0 5752 0 1 3010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_94
timestamp 1743127117
transform 1 0 5768 0 1 3010
box -4 -6 196 206
use OAI21X1  OAI21X1_279
timestamp 1743127117
transform 1 0 5960 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_280
timestamp 1743127117
transform -1 0 6088 0 1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_82
timestamp 1743127117
transform 1 0 6088 0 1 3010
box -4 -6 100 206
use BUFX4  BUFX4_84
timestamp 1743127117
transform 1 0 6184 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_99
timestamp 1743127117
transform 1 0 6248 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_333
timestamp 1743127117
transform -1 0 6360 0 1 3010
box -4 -6 68 206
use OR2X2  OR2X2_7
timestamp 1743127117
transform -1 0 6424 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_88
timestamp 1743127117
transform -1 0 6456 0 1 3010
box -4 -6 36 206
use MUX2X1  MUX2X1_94
timestamp 1743127117
transform -1 0 6552 0 1 3010
box -4 -6 100 206
use OAI21X1  OAI21X1_305
timestamp 1743127117
transform 1 0 6552 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_306
timestamp 1743127117
transform -1 0 6680 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_80
timestamp 1743127117
transform 1 0 6680 0 1 3010
box -4 -6 196 206
use FILL  FILL_16_1
timestamp 1743127117
transform 1 0 6872 0 1 3010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_50
timestamp 1743127117
transform 1 0 8 0 -1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_228
timestamp 1743127117
transform -1 0 264 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_229
timestamp 1743127117
transform -1 0 328 0 -1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_74
timestamp 1743127117
transform -1 0 424 0 -1 3410
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_49
timestamp 1743127117
transform 1 0 424 0 -1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_71
timestamp 1743127117
transform 1 0 616 0 -1 3410
box -4 -6 52 206
use OR2X2  OR2X2_11
timestamp 1743127117
transform -1 0 728 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_68
timestamp 1743127117
transform 1 0 728 0 -1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_243
timestamp 1743127117
transform 1 0 920 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_245
timestamp 1743127117
transform 1 0 984 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_0_0
timestamp 1743127117
transform 1 0 1048 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_1
timestamp 1743127117
transform 1 0 1064 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_2
timestamp 1743127117
transform 1 0 1080 0 -1 3410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_51
timestamp 1743127117
transform 1 0 1096 0 -1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_73
timestamp 1743127117
transform 1 0 1288 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_69
timestamp 1743127117
transform 1 0 1336 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_62
timestamp 1743127117
transform -1 0 1416 0 -1 3410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_9
timestamp 1743127117
transform 1 0 1416 0 -1 3410
box -4 -6 116 206
use INVX2  INVX2_3
timestamp 1743127117
transform 1 0 1528 0 -1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_67
timestamp 1743127117
transform -1 0 1608 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_249
timestamp 1743127117
transform 1 0 1608 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_52
timestamp 1743127117
transform -1 0 2024 0 -1 3410
box -4 -6 356 206
use BUFX4  BUFX4_5
timestamp 1743127117
transform -1 0 2088 0 -1 3410
box -4 -6 68 206
use BUFX4  BUFX4_28
timestamp 1743127117
transform 1 0 2088 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_405
timestamp 1743127117
transform -1 0 2216 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_129
timestamp 1743127117
transform -1 0 2248 0 -1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_26
timestamp 1743127117
transform -1 0 2296 0 -1 3410
box -4 -6 52 206
use DFFSR  DFFSR_106
timestamp 1743127117
transform -1 0 2648 0 -1 3410
box -4 -6 356 206
use FILL  FILL_16_1_0
timestamp 1743127117
transform 1 0 2648 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_1
timestamp 1743127117
transform 1 0 2664 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_2
timestamp 1743127117
transform 1 0 2680 0 -1 3410
box -4 -6 20 206
use DFFSR  DFFSR_134
timestamp 1743127117
transform 1 0 2696 0 -1 3410
box -4 -6 356 206
use OAI21X1  OAI21X1_437
timestamp 1743127117
transform -1 0 3112 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_436
timestamp 1743127117
transform -1 0 3176 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_157
timestamp 1743127117
transform -1 0 3224 0 -1 3410
box -4 -6 52 206
use AOI22X1  AOI22X1_17
timestamp 1743127117
transform -1 0 3304 0 -1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_18
timestamp 1743127117
transform -1 0 3384 0 -1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_11
timestamp 1743127117
transform -1 0 3464 0 -1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_7
timestamp 1743127117
transform -1 0 3544 0 -1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_9
timestamp 1743127117
transform 1 0 3544 0 -1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_151
timestamp 1743127117
transform 1 0 3624 0 -1 3410
box -4 -6 52 206
use AOI22X1  AOI22X1_10
timestamp 1743127117
transform -1 0 3752 0 -1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_149
timestamp 1743127117
transform 1 0 3752 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_150
timestamp 1743127117
transform -1 0 3848 0 -1 3410
box -4 -6 52 206
use AOI22X1  AOI22X1_3
timestamp 1743127117
transform -1 0 3928 0 -1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_148
timestamp 1743127117
transform -1 0 3976 0 -1 3410
box -4 -6 52 206
use AOI22X1  AOI22X1_2
timestamp 1743127117
transform 1 0 3976 0 -1 3410
box -4 -6 84 206
use OAI21X1  OAI21X1_335
timestamp 1743127117
transform -1 0 4120 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_102
timestamp 1743127117
transform 1 0 4120 0 -1 3410
box -4 -6 52 206
use FILL  FILL_16_2_0
timestamp 1743127117
transform 1 0 4168 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_1
timestamp 1743127117
transform 1 0 4184 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_2
timestamp 1743127117
transform 1 0 4200 0 -1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_331
timestamp 1743127117
transform 1 0 4216 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_347
timestamp 1743127117
transform 1 0 4280 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_65
timestamp 1743127117
transform -1 0 4696 0 -1 3410
box -4 -6 356 206
use NAND2X1  NAND2X1_100
timestamp 1743127117
transform 1 0 4696 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_108
timestamp 1743127117
transform 1 0 4744 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_78
timestamp 1743127117
transform 1 0 4792 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_272
timestamp 1743127117
transform 1 0 4824 0 -1 3410
box -4 -6 68 206
use BUFX4  BUFX4_2
timestamp 1743127117
transform -1 0 4952 0 -1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_91
timestamp 1743127117
transform 1 0 4952 0 -1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_300
timestamp 1743127117
transform 1 0 5048 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_299
timestamp 1743127117
transform -1 0 5176 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_87
timestamp 1743127117
transform 1 0 5176 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_282
timestamp 1743127117
transform 1 0 5208 0 -1 3410
box -4 -6 68 206
use BUFX4  BUFX4_83
timestamp 1743127117
transform 1 0 5272 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_25
timestamp 1743127117
transform 1 0 5336 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_332
timestamp 1743127117
transform 1 0 5400 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_24
timestamp 1743127117
transform 1 0 5464 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_334
timestamp 1743127117
transform 1 0 5528 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_77
timestamp 1743127117
transform -1 0 5784 0 -1 3410
box -4 -6 196 206
use FILL  FILL_16_3_0
timestamp 1743127117
transform 1 0 5784 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_3_1
timestamp 1743127117
transform 1 0 5800 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_3_2
timestamp 1743127117
transform 1 0 5816 0 -1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_324
timestamp 1743127117
transform 1 0 5832 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_323
timestamp 1743127117
transform -1 0 5960 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_26
timestamp 1743127117
transform 1 0 5960 0 -1 3410
box -4 -6 68 206
use BUFX4  BUFX4_49
timestamp 1743127117
transform 1 0 6024 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_350
timestamp 1743127117
transform -1 0 6152 0 -1 3410
box -4 -6 68 206
use BUFX4  BUFX4_82
timestamp 1743127117
transform 1 0 6152 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_348
timestamp 1743127117
transform 1 0 6216 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_28
timestamp 1743127117
transform -1 0 6344 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_95
timestamp 1743127117
transform -1 0 6376 0 -1 3410
box -4 -6 36 206
use MUX2X1  MUX2X1_84
timestamp 1743127117
transform 1 0 6376 0 -1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_301
timestamp 1743127117
transform 1 0 6472 0 -1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_92
timestamp 1743127117
transform 1 0 6536 0 -1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_302
timestamp 1743127117
transform -1 0 6696 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_90
timestamp 1743127117
transform 1 0 6696 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_55
timestamp 1743127117
transform 1 0 8 0 1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_214
timestamp 1743127117
transform -1 0 264 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_215
timestamp 1743127117
transform -1 0 328 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_226
timestamp 1743127117
transform 1 0 328 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_52
timestamp 1743127117
transform 1 0 8 0 -1 3810
box -4 -6 196 206
use INVX1  INVX1_60
timestamp 1743127117
transform 1 0 200 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_232
timestamp 1743127117
transform 1 0 232 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_233
timestamp 1743127117
transform -1 0 360 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_67
timestamp 1743127117
transform -1 0 456 0 -1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_76
timestamp 1743127117
transform -1 0 552 0 -1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_73
timestamp 1743127117
transform -1 0 552 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_227
timestamp 1743127117
transform -1 0 456 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_61
timestamp 1743127117
transform 1 0 552 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_68
timestamp 1743127117
transform 1 0 552 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_75
timestamp 1743127117
transform 1 0 648 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_240
timestamp 1743127117
transform -1 0 648 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_54
timestamp 1743127117
transform -1 0 696 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_252
timestamp 1743127117
transform 1 0 728 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_64
timestamp 1743127117
transform 1 0 696 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_244
timestamp 1743127117
transform -1 0 760 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_63
timestamp 1743127117
transform 1 0 792 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_185
timestamp 1743127117
transform 1 0 760 0 1 3410
box -4 -6 68 206
use BUFX4  BUFX4_15
timestamp 1743127117
transform 1 0 824 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_184
timestamp 1743127117
transform -1 0 888 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_253
timestamp 1743127117
transform 1 0 888 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_180
timestamp 1743127117
transform -1 0 952 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_241
timestamp 1743127117
transform 1 0 1016 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_239
timestamp 1743127117
transform 1 0 952 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_231
timestamp 1743127117
transform 1 0 1016 0 1 3410
box -4 -6 68 206
use BUFX4  BUFX4_94
timestamp 1743127117
transform -1 0 1016 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_0_0
timestamp 1743127117
transform 1 0 1080 0 -1 3810
box -4 -6 20 206
use FILL  FILL_17_0_0
timestamp 1743127117
transform 1 0 1080 0 1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_261
timestamp 1743127117
transform -1 0 1256 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_16
timestamp 1743127117
transform 1 0 1128 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_0_2
timestamp 1743127117
transform 1 0 1112 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_1
timestamp 1743127117
transform 1 0 1096 0 -1 3810
box -4 -6 20 206
use MUX2X1  MUX2X1_75
timestamp 1743127117
transform 1 0 1192 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_230
timestamp 1743127117
transform 1 0 1128 0 1 3410
box -4 -6 68 206
use FILL  FILL_17_0_2
timestamp 1743127117
transform 1 0 1112 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_1
timestamp 1743127117
transform 1 0 1096 0 1 3410
box -4 -6 20 206
use BUFX4  BUFX4_95
timestamp 1743127117
transform 1 0 1256 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_50
timestamp 1743127117
transform 1 0 1288 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_257
timestamp 1743127117
transform -1 0 1432 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_24
timestamp 1743127117
transform -1 0 1368 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_248
timestamp 1743127117
transform -1 0 1448 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_179
timestamp 1743127117
transform -1 0 1384 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_66
timestamp 1743127117
transform -1 0 1464 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_247
timestamp 1743127117
transform 1 0 1448 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_262
timestamp 1743127117
transform -1 0 1576 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_263
timestamp 1743127117
transform -1 0 1640 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_186
timestamp 1743127117
transform -1 0 1704 0 1 3410
box -4 -6 68 206
use DFFSR  DFFSR_55
timestamp 1743127117
transform 1 0 1704 0 1 3410
box -4 -6 356 206
use INVX1  INVX1_65
timestamp 1743127117
transform -1 0 1496 0 -1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_57
timestamp 1743127117
transform -1 0 1688 0 -1 3810
box -4 -6 196 206
use BUFX4  BUFX4_29
timestamp 1743127117
transform 1 0 1688 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_78
timestamp 1743127117
transform -1 0 1800 0 -1 3810
box -4 -6 52 206
use DFFSR  DFFSR_49
timestamp 1743127117
transform 1 0 1800 0 -1 3810
box -4 -6 356 206
use XOR2X1  XOR2X1_5
timestamp 1743127117
transform -1 0 2168 0 1 3410
box -4 -6 116 206
use OAI21X1  OAI21X1_198
timestamp 1743127117
transform -1 0 2232 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_254
timestamp 1743127117
transform -1 0 2216 0 -1 3810
box -4 -6 68 206
use OR2X2  OR2X2_6
timestamp 1743127117
transform 1 0 2232 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_264
timestamp 1743127117
transform 1 0 2296 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_81
timestamp 1743127117
transform 1 0 2360 0 1 3410
box -4 -6 52 206
use DFFSR  DFFSR_41
timestamp 1743127117
transform 1 0 2408 0 1 3410
box -4 -6 356 206
use BUFX2  BUFX2_15
timestamp 1743127117
transform 1 0 2216 0 -1 3810
box -4 -6 52 206
use BUFX4  BUFX4_24
timestamp 1743127117
transform 1 0 2264 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_80
timestamp 1743127117
transform -1 0 2376 0 -1 3810
box -4 -6 52 206
use DFFSR  DFFSR_50
timestamp 1743127117
transform 1 0 2376 0 -1 3810
box -4 -6 356 206
use FILL  FILL_17_1_0
timestamp 1743127117
transform 1 0 2760 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_1
timestamp 1743127117
transform 1 0 2776 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_2
timestamp 1743127117
transform 1 0 2792 0 1 3410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_22
timestamp 1743127117
transform 1 0 2808 0 1 3410
box -4 -6 148 206
use FILL  FILL_18_1_0
timestamp 1743127117
transform -1 0 2744 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_1
timestamp 1743127117
transform -1 0 2760 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_2
timestamp 1743127117
transform -1 0 2776 0 -1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_258
timestamp 1743127117
transform -1 0 2840 0 -1 3810
box -4 -6 68 206
use BUFX4  BUFX4_25
timestamp 1743127117
transform 1 0 2840 0 -1 3810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_18
timestamp 1743127117
transform 1 0 2904 0 -1 3810
box -4 -6 148 206
use OAI21X1  OAI21X1_438
timestamp 1743127117
transform -1 0 3096 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_147
timestamp 1743127117
transform 1 0 2984 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_145
timestamp 1743127117
transform -1 0 2984 0 1 3410
box -4 -6 36 206
use AOI22X1  AOI22X1_16
timestamp 1743127117
transform -1 0 3224 0 -1 3810
box -4 -6 84 206
use OAI21X1  OAI21X1_439
timestamp 1743127117
transform 1 0 3080 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_155
timestamp 1743127117
transform 1 0 3048 0 -1 3810
box -4 -6 36 206
use AOI22X1  AOI22X1_15
timestamp 1743127117
transform 1 0 3160 0 1 3410
box -4 -6 84 206
use NAND3X1  NAND3X1_50
timestamp 1743127117
transform -1 0 3160 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_151
timestamp 1743127117
transform -1 0 3256 0 -1 3810
box -4 -6 36 206
use AOI22X1  AOI22X1_14
timestamp 1743127117
transform 1 0 3240 0 1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_8
timestamp 1743127117
transform 1 0 3288 0 -1 3810
box -4 -6 84 206
use INVX1  INVX1_152
timestamp 1743127117
transform 1 0 3256 0 -1 3810
box -4 -6 36 206
use AOI22X1  AOI22X1_6
timestamp 1743127117
transform 1 0 3320 0 1 3410
box -4 -6 84 206
use NAND3X1  NAND3X1_46
timestamp 1743127117
transform 1 0 3368 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_44
timestamp 1743127117
transform 1 0 3400 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_49
timestamp 1743127117
transform -1 0 3560 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_51
timestamp 1743127117
transform 1 0 3432 0 -1 3810
box -4 -6 68 206
use AOI22X1  AOI22X1_12
timestamp 1743127117
transform -1 0 3544 0 1 3410
box -4 -6 84 206
use AOI22X1  AOI22X1_13
timestamp 1743127117
transform -1 0 3672 0 -1 3810
box -4 -6 84 206
use INVX1  INVX1_153
timestamp 1743127117
transform 1 0 3560 0 -1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_48
timestamp 1743127117
transform -1 0 3608 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_155
timestamp 1743127117
transform -1 0 3656 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_156
timestamp 1743127117
transform -1 0 3704 0 1 3410
box -4 -6 52 206
use AOI22X1  AOI22X1_4
timestamp 1743127117
transform 1 0 3704 0 1 3410
box -4 -6 84 206
use NAND3X1  NAND3X1_42
timestamp 1743127117
transform 1 0 3784 0 1 3410
box -4 -6 68 206
use DFFSR  DFFSR_66
timestamp 1743127117
transform -1 0 4200 0 1 3410
box -4 -6 356 206
use INVX1  INVX1_154
timestamp 1743127117
transform 1 0 3672 0 -1 3810
box -4 -6 36 206
use AOI22X1  AOI22X1_5
timestamp 1743127117
transform 1 0 3704 0 -1 3810
box -4 -6 84 206
use NAND3X1  NAND3X1_43
timestamp 1743127117
transform -1 0 3848 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_41
timestamp 1743127117
transform 1 0 3848 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_40
timestamp 1743127117
transform 1 0 3912 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_2_2
timestamp 1743127117
transform -1 0 4152 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_1
timestamp 1743127117
transform -1 0 4136 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_0
timestamp 1743127117
transform -1 0 4120 0 -1 3810
box -4 -6 20 206
use INVX8  INVX8_8
timestamp 1743127117
transform 1 0 4024 0 -1 3810
box -4 -6 84 206
use NOR2X1  NOR2X1_35
timestamp 1743127117
transform 1 0 3976 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_106
timestamp 1743127117
transform 1 0 4312 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_343
timestamp 1743127117
transform -1 0 4312 0 1 3410
box -4 -6 68 206
use FILL  FILL_17_2_2
timestamp 1743127117
transform -1 0 4248 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_1
timestamp 1743127117
transform -1 0 4232 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_0
timestamp 1743127117
transform -1 0 4216 0 1 3410
box -4 -6 20 206
use DFFSR  DFFSR_68
timestamp 1743127117
transform -1 0 4504 0 -1 3810
box -4 -6 356 206
use DFFSR  DFFSR_69
timestamp 1743127117
transform -1 0 4712 0 1 3410
box -4 -6 356 206
use DFFSR  DFFSR_125
timestamp 1743127117
transform 1 0 4504 0 -1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_88
timestamp 1743127117
transform 1 0 4712 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_281
timestamp 1743127117
transform 1 0 4760 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_89
timestamp 1743127117
transform -1 0 5016 0 1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_95
timestamp 1743127117
transform 1 0 5016 0 1 3410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_14
timestamp 1743127117
transform 1 0 4856 0 -1 3810
box -4 -6 148 206
use NAND2X1  NAND2X1_85
timestamp 1743127117
transform 1 0 5000 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_269
timestamp 1743127117
transform -1 0 5112 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_93
timestamp 1743127117
transform 1 0 5208 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_283
timestamp 1743127117
transform -1 0 5304 0 1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_83
timestamp 1743127117
transform 1 0 5304 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_344
timestamp 1743127117
transform 1 0 5400 0 1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_99
timestamp 1743127117
transform -1 0 5208 0 -1 3810
box -4 -6 100 206
use OAI21X1  OAI21X1_291
timestamp 1743127117
transform 1 0 5208 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_292
timestamp 1743127117
transform -1 0 5336 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_27
timestamp 1743127117
transform 1 0 5336 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_87
timestamp 1743127117
transform -1 0 5496 0 -1 3810
box -4 -6 100 206
use INVX1  INVX1_94
timestamp 1743127117
transform -1 0 5624 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_345
timestamp 1743127117
transform -1 0 5592 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_346
timestamp 1743127117
transform 1 0 5464 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_3_2
timestamp 1743127117
transform 1 0 5768 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_3_1
timestamp 1743127117
transform 1 0 5752 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_3_0
timestamp 1743127117
transform 1 0 5736 0 -1 3810
box -4 -6 20 206
use NAND2X1  NAND2X1_96
timestamp 1743127117
transform 1 0 5688 0 -1 3810
box -4 -6 52 206
use MUX2X1  MUX2X1_97
timestamp 1743127117
transform -1 0 5816 0 1 3410
box -4 -6 100 206
use FILL  FILL_17_3_2
timestamp 1743127117
transform -1 0 5720 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_3_1
timestamp 1743127117
transform -1 0 5704 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_3_0
timestamp 1743127117
transform -1 0 5688 0 1 3410
box -4 -6 20 206
use NAND2X1  NAND2X1_105
timestamp 1743127117
transform -1 0 5672 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_83
timestamp 1743127117
transform -1 0 5688 0 -1 3810
box -4 -6 196 206
use BUFX4  BUFX4_45
timestamp 1743127117
transform -1 0 5976 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_311
timestamp 1743127117
transform -1 0 5912 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_312
timestamp 1743127117
transform 1 0 5784 0 -1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_103
timestamp 1743127117
transform -1 0 5912 0 1 3410
box -4 -6 100 206
use INVX1  INVX1_86
timestamp 1743127117
transform 1 0 6120 0 -1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_39
timestamp 1743127117
transform -1 0 6120 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_85
timestamp 1743127117
transform -1 0 6072 0 -1 3810
box -4 -6 36 206
use BUFX4  BUFX4_48
timestamp 1743127117
transform -1 0 6040 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_304
timestamp 1743127117
transform 1 0 6104 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_79
timestamp 1743127117
transform 1 0 5912 0 1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_270
timestamp 1743127117
transform 1 0 6200 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_97
timestamp 1743127117
transform -1 0 6200 0 -1 3810
box -4 -6 52 206
use MUX2X1  MUX2X1_93
timestamp 1743127117
transform 1 0 6232 0 1 3410
box -4 -6 100 206
use OAI21X1  OAI21X1_303
timestamp 1743127117
transform -1 0 6232 0 1 3410
box -4 -6 68 206
use MUX2X1  MUX2X1_79
timestamp 1743127117
transform 1 0 6264 0 -1 3810
box -4 -6 100 206
use OAI21X1  OAI21X1_285
timestamp 1743127117
transform 1 0 6328 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_94
timestamp 1743127117
transform 1 0 6424 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_271
timestamp 1743127117
transform -1 0 6424 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_286
timestamp 1743127117
transform -1 0 6456 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_38
timestamp 1743127117
transform 1 0 6472 0 -1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_37
timestamp 1743127117
transform -1 0 6504 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_96
timestamp 1743127117
transform -1 0 6696 0 1 3410
box -4 -6 196 206
use NOR2X1  NOR2X1_40
timestamp 1743127117
transform -1 0 6744 0 1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_33
timestamp 1743127117
transform -1 0 6792 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_76
timestamp 1743127117
transform 1 0 6792 0 1 3410
box -4 -6 36 206
use FILL  FILL_18_1
timestamp 1743127117
transform 1 0 6824 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2
timestamp 1743127117
transform 1 0 6840 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_3
timestamp 1743127117
transform 1 0 6856 0 1 3410
box -4 -6 20 206
use DFFSR  DFFSR_73
timestamp 1743127117
transform -1 0 6872 0 -1 3810
box -4 -6 356 206
use FILL  FILL_18_4
timestamp 1743127117
transform 1 0 6872 0 1 3410
box -4 -6 20 206
use FILL  FILL_19_1
timestamp 1743127117
transform -1 0 6888 0 -1 3810
box -4 -6 20 206
use BUFX2  BUFX2_24
timestamp 1743127117
transform -1 0 56 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_62
timestamp 1743127117
transform 1 0 56 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_202
timestamp 1743127117
transform -1 0 312 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_17
timestamp 1743127117
transform -1 0 376 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_204
timestamp 1743127117
transform 1 0 376 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_205
timestamp 1743127117
transform -1 0 504 0 1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_62
timestamp 1743127117
transform -1 0 600 0 1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_68
timestamp 1743127117
transform -1 0 696 0 1 3810
box -4 -6 100 206
use INVX1  INVX1_68
timestamp 1743127117
transform 1 0 696 0 1 3810
box -4 -6 36 206
use BUFX4  BUFX4_63
timestamp 1743127117
transform -1 0 792 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_79
timestamp 1743127117
transform 1 0 792 0 1 3810
box -4 -6 52 206
use BUFX4  BUFX4_61
timestamp 1743127117
transform 1 0 840 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_251
timestamp 1743127117
transform -1 0 968 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_96
timestamp 1743127117
transform -1 0 1032 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_260
timestamp 1743127117
transform 1 0 1032 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_0_0
timestamp 1743127117
transform 1 0 1096 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_1
timestamp 1743127117
transform 1 0 1112 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_2
timestamp 1743127117
transform 1 0 1128 0 1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_29
timestamp 1743127117
transform 1 0 1144 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_193
timestamp 1743127117
transform 1 0 1192 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_259
timestamp 1743127117
transform -1 0 1320 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_20
timestamp 1743127117
transform -1 0 1384 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_255
timestamp 1743127117
transform -1 0 1448 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_77
timestamp 1743127117
transform -1 0 1496 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_256
timestamp 1743127117
transform -1 0 1560 0 1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_69
timestamp 1743127117
transform 1 0 1560 0 1 3810
box -4 -6 100 206
use OAI21X1  OAI21X1_219
timestamp 1743127117
transform 1 0 1656 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_218
timestamp 1743127117
transform -1 0 1784 0 1 3810
box -4 -6 68 206
use MUX2X1  MUX2X1_63
timestamp 1743127117
transform 1 0 1784 0 1 3810
box -4 -6 100 206
use OAI21X1  OAI21X1_206
timestamp 1743127117
transform 1 0 1880 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_207
timestamp 1743127117
transform 1 0 1944 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_63
timestamp 1743127117
transform -1 0 2200 0 1 3810
box -4 -6 196 206
use XOR2X1  XOR2X1_6
timestamp 1743127117
transform 1 0 2200 0 1 3810
box -4 -6 116 206
use MUX2X1  MUX2X1_59
timestamp 1743127117
transform 1 0 2312 0 1 3810
box -4 -6 100 206
use MUX2X1  MUX2X1_60
timestamp 1743127117
transform 1 0 2408 0 1 3810
box -4 -6 100 206
use BUFX4  BUFX4_27
timestamp 1743127117
transform 1 0 2504 0 1 3810
box -4 -6 68 206
use INVX8  INVX8_3
timestamp 1743127117
transform 1 0 2568 0 1 3810
box -4 -6 84 206
use FILL  FILL_19_1_0
timestamp 1743127117
transform -1 0 2664 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_1
timestamp 1743127117
transform -1 0 2680 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_2
timestamp 1743127117
transform -1 0 2696 0 1 3810
box -4 -6 20 206
use MUX2X1  MUX2X1_106
timestamp 1743127117
transform -1 0 2792 0 1 3810
box -4 -6 100 206
use DFFSR  DFFSR_137
timestamp 1743127117
transform 1 0 2792 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_152
timestamp 1743127117
transform -1 0 3192 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_440
timestamp 1743127117
transform 1 0 3192 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_159
timestamp 1743127117
transform -1 0 3304 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_441
timestamp 1743127117
transform -1 0 3368 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_442
timestamp 1743127117
transform -1 0 3432 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_11
timestamp 1743127117
transform -1 0 3496 0 1 3810
box -4 -6 68 206
use OAI22X1  OAI22X1_5
timestamp 1743127117
transform -1 0 3576 0 1 3810
box -4 -6 84 206
use NOR2X1  NOR2X1_42
timestamp 1743127117
transform 1 0 3576 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_10
timestamp 1743127117
transform -1 0 3688 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_158
timestamp 1743127117
transform -1 0 3736 0 1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_47
timestamp 1743127117
transform 1 0 3736 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_140
timestamp 1743127117
transform 1 0 3800 0 1 3810
box -4 -6 52 206
use DFFSR  DFFSR_135
timestamp 1743127117
transform 1 0 3848 0 1 3810
box -4 -6 356 206
use FILL  FILL_19_2_0
timestamp 1743127117
transform 1 0 4200 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_1
timestamp 1743127117
transform 1 0 4216 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_2
timestamp 1743127117
transform 1 0 4232 0 1 3810
box -4 -6 20 206
use MUX2X1  MUX2X1_105
timestamp 1743127117
transform 1 0 4248 0 1 3810
box -4 -6 100 206
use BUFX4  BUFX4_91
timestamp 1743127117
transform -1 0 4408 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_339
timestamp 1743127117
transform 1 0 4408 0 1 3810
box -4 -6 68 206
use DFFSR  DFFSR_67
timestamp 1743127117
transform -1 0 4824 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_104
timestamp 1743127117
transform 1 0 4824 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_89
timestamp 1743127117
transform -1 0 4920 0 1 3810
box -4 -6 52 206
use INVX8  INVX8_4
timestamp 1743127117
transform 1 0 4920 0 1 3810
box -4 -6 84 206
use NAND2X1  NAND2X1_86
timestamp 1743127117
transform -1 0 5048 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_416
timestamp 1743127117
transform -1 0 5112 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_408
timestamp 1743127117
transform -1 0 5176 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_414
timestamp 1743127117
transform -1 0 5240 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_86
timestamp 1743127117
transform -1 0 5304 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_87
timestamp 1743127117
transform -1 0 5352 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_315
timestamp 1743127117
transform 1 0 5352 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_316
timestamp 1743127117
transform -1 0 5480 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_73
timestamp 1743127117
transform 1 0 5480 0 1 3810
box -4 -6 196 206
use INVX1  INVX1_84
timestamp 1743127117
transform -1 0 5704 0 1 3810
box -4 -6 36 206
use FILL  FILL_19_3_0
timestamp 1743127117
transform -1 0 5720 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_3_1
timestamp 1743127117
transform -1 0 5736 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_3_2
timestamp 1743127117
transform -1 0 5752 0 1 3810
box -4 -6 20 206
use NAND2X1  NAND2X1_90
timestamp 1743127117
transform -1 0 5800 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_329
timestamp 1743127117
transform -1 0 5864 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_85
timestamp 1743127117
transform 1 0 5864 0 1 3810
box -4 -6 196 206
use NAND3X1  NAND3X1_23
timestamp 1743127117
transform -1 0 6120 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_420
timestamp 1743127117
transform 1 0 6120 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_128
timestamp 1743127117
transform -1 0 6232 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_91
timestamp 1743127117
transform -1 0 6424 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_310
timestamp 1743127117
transform -1 0 6488 0 1 3810
box -4 -6 68 206
use DFFSR  DFFSR_131
timestamp 1743127117
transform 1 0 6488 0 1 3810
box -4 -6 356 206
use FILL  FILL_20_1
timestamp 1743127117
transform 1 0 6840 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_2
timestamp 1743127117
transform 1 0 6856 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_3
timestamp 1743127117
transform 1 0 6872 0 1 3810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_61
timestamp 1743127117
transform 1 0 8 0 -1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_203
timestamp 1743127117
transform 1 0 200 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_61
timestamp 1743127117
transform -1 0 360 0 -1 4210
box -4 -6 100 206
use BUFX4  BUFX4_16
timestamp 1743127117
transform 1 0 360 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_236
timestamp 1743127117
transform 1 0 424 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_237
timestamp 1743127117
transform -1 0 552 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_78
timestamp 1743127117
transform -1 0 648 0 -1 4210
box -4 -6 100 206
use INVX1  INVX1_72
timestamp 1743127117
transform 1 0 648 0 -1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_54
timestamp 1743127117
transform -1 0 872 0 -1 4210
box -4 -6 196 206
use INVX1  INVX1_67
timestamp 1743127117
transform 1 0 872 0 -1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_19
timestamp 1743127117
transform 1 0 904 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_71
timestamp 1743127117
transform 1 0 968 0 -1 4210
box -4 -6 196 206
use FILL  FILL_20_0_0
timestamp 1743127117
transform -1 0 1176 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_1
timestamp 1743127117
transform -1 0 1192 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_2
timestamp 1743127117
transform -1 0 1208 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_194
timestamp 1743127117
transform -1 0 1272 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1743127117
transform 1 0 1272 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_57
timestamp 1743127117
transform 1 0 1336 0 -1 4210
box -4 -6 100 206
use INVX1  INVX1_69
timestamp 1743127117
transform -1 0 1464 0 -1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_18
timestamp 1743127117
transform -1 0 1528 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_70
timestamp 1743127117
transform -1 0 1560 0 -1 4210
box -4 -6 36 206
use BUFX4  BUFX4_18
timestamp 1743127117
transform 1 0 1560 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_234
timestamp 1743127117
transform 1 0 1624 0 -1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_55
timestamp 1743127117
transform 1 0 1688 0 -1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_187
timestamp 1743127117
transform 1 0 1784 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_188
timestamp 1743127117
transform -1 0 1912 0 -1 4210
box -4 -6 68 206
use DFFSR  DFFSR_39
timestamp 1743127117
transform -1 0 2264 0 -1 4210
box -4 -6 356 206
use NAND2X1  NAND2X1_64
timestamp 1743127117
transform 1 0 2264 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_63
timestamp 1743127117
transform -1 0 2360 0 -1 4210
box -4 -6 52 206
use AND2X2  AND2X2_3
timestamp 1743127117
transform 1 0 2360 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_199
timestamp 1743127117
transform 1 0 2424 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_65
timestamp 1743127117
transform -1 0 2536 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_201
timestamp 1743127117
transform -1 0 2600 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_1_0
timestamp 1743127117
transform 1 0 2600 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_1
timestamp 1743127117
transform 1 0 2616 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_2
timestamp 1743127117
transform 1 0 2632 0 -1 4210
box -4 -6 20 206
use DFFSR  DFFSR_40
timestamp 1743127117
transform 1 0 2648 0 -1 4210
box -4 -6 356 206
use NAND2X1  NAND2X1_141
timestamp 1743127117
transform -1 0 3048 0 -1 4210
box -4 -6 52 206
use INVX1  INVX1_148
timestamp 1743127117
transform -1 0 3080 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_143
timestamp 1743127117
transform 1 0 3080 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_50
timestamp 1743127117
transform -1 0 3176 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_51
timestamp 1743127117
transform -1 0 3224 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_431
timestamp 1743127117
transform -1 0 3288 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_6
timestamp 1743127117
transform -1 0 3352 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_142
timestamp 1743127117
transform -1 0 3400 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_432
timestamp 1743127117
transform -1 0 3464 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_5
timestamp 1743127117
transform -1 0 3528 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_48
timestamp 1743127117
transform 1 0 3528 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_135
timestamp 1743127117
transform 1 0 3576 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_30
timestamp 1743127117
transform -1 0 3688 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_29
timestamp 1743127117
transform 1 0 3688 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_31
timestamp 1743127117
transform -1 0 3816 0 -1 4210
box -4 -6 68 206
use INVX2  INVX2_7
timestamp 1743127117
transform -1 0 3848 0 -1 4210
box -4 -6 36 206
use AOI22X1  AOI22X1_1
timestamp 1743127117
transform -1 0 3928 0 -1 4210
box -4 -6 84 206
use NAND3X1  NAND3X1_39
timestamp 1743127117
transform 1 0 3928 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_9
timestamp 1743127117
transform -1 0 4056 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_41
timestamp 1743127117
transform -1 0 4104 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_2_0
timestamp 1743127117
transform -1 0 4120 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_1
timestamp 1743127117
transform -1 0 4136 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_2
timestamp 1743127117
transform -1 0 4152 0 -1 4210
box -4 -6 20 206
use DFFSR  DFFSR_124
timestamp 1743127117
transform -1 0 4504 0 -1 4210
box -4 -6 356 206
use DFFSR  DFFSR_129
timestamp 1743127117
transform 1 0 4504 0 -1 4210
box -4 -6 356 206
use OAI21X1  OAI21X1_409
timestamp 1743127117
transform 1 0 4856 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_417
timestamp 1743127117
transform -1 0 4984 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_138
timestamp 1743127117
transform -1 0 5016 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_415
timestamp 1743127117
transform 1 0 5016 0 -1 4210
box -4 -6 68 206
use DFFSR  DFFSR_128
timestamp 1743127117
transform -1 0 5432 0 -1 4210
box -4 -6 356 206
use BUFX4  BUFX4_21
timestamp 1743127117
transform -1 0 5496 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_419
timestamp 1743127117
transform 1 0 5496 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_139
timestamp 1743127117
transform -1 0 5592 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_418
timestamp 1743127117
transform -1 0 5656 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_328
timestamp 1743127117
transform 1 0 5656 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_3_0
timestamp 1743127117
transform -1 0 5736 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_3_1
timestamp 1743127117
transform -1 0 5752 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_3_2
timestamp 1743127117
transform -1 0 5768 0 -1 4210
box -4 -6 20 206
use DFFSR  DFFSR_130
timestamp 1743127117
transform -1 0 6120 0 -1 4210
box -4 -6 356 206
use XNOR2X1  XNOR2X1_12
timestamp 1743127117
transform 1 0 6120 0 -1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_95
timestamp 1743127117
transform -1 0 6280 0 -1 4210
box -4 -6 52 206
use INVX2  INVX2_4
timestamp 1743127117
transform 1 0 6280 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_351
timestamp 1743127117
transform 1 0 6312 0 -1 4210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_10
timestamp 1743127117
transform 1 0 6376 0 -1 4210
box -4 -6 116 206
use DFFSR  DFFSR_71
timestamp 1743127117
transform -1 0 6840 0 -1 4210
box -4 -6 356 206
use FILL  FILL_21_1
timestamp 1743127117
transform -1 0 6856 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_2
timestamp 1743127117
transform -1 0 6872 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_3
timestamp 1743127117
transform -1 0 6888 0 -1 4210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_56
timestamp 1743127117
transform -1 0 200 0 1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_217
timestamp 1743127117
transform 1 0 200 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_216
timestamp 1743127117
transform -1 0 328 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_70
timestamp 1743127117
transform -1 0 424 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_189
timestamp 1743127117
transform -1 0 488 0 1 4210
box -4 -6 68 206
use BUFX4  BUFX4_65
timestamp 1743127117
transform -1 0 552 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_64
timestamp 1743127117
transform 1 0 552 0 1 4210
box -4 -6 100 206
use MUX2X1  MUX2X1_56
timestamp 1743127117
transform -1 0 744 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_208
timestamp 1743127117
transform 1 0 744 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_209
timestamp 1743127117
transform -1 0 872 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_64
timestamp 1743127117
transform -1 0 1064 0 1 4210
box -4 -6 196 206
use FILL  FILL_21_0_0
timestamp 1743127117
transform -1 0 1080 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_1
timestamp 1743127117
transform -1 0 1096 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_2
timestamp 1743127117
transform -1 0 1112 0 1 4210
box -4 -6 20 206
use MUX2X1  MUX2X1_53
timestamp 1743127117
transform -1 0 1208 0 1 4210
box -4 -6 100 206
use BUFX4  BUFX4_92
timestamp 1743127117
transform 1 0 1208 0 1 4210
box -4 -6 68 206
use BUFX4  BUFX4_62
timestamp 1743127117
transform -1 0 1336 0 1 4210
box -4 -6 68 206
use BUFX4  BUFX4_93
timestamp 1743127117
transform 1 0 1336 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_53
timestamp 1743127117
transform -1 0 1592 0 1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_210
timestamp 1743127117
transform -1 0 1656 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_235
timestamp 1743127117
transform -1 0 1720 0 1 4210
box -4 -6 68 206
use MUX2X1  MUX2X1_77
timestamp 1743127117
transform 1 0 1720 0 1 4210
box -4 -6 100 206
use OAI21X1  OAI21X1_222
timestamp 1743127117
transform -1 0 1880 0 1 4210
box -4 -6 68 206
use BUFX4  BUFX4_64
timestamp 1743127117
transform 1 0 1880 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_69
timestamp 1743127117
transform -1 0 2136 0 1 4210
box -4 -6 196 206
use NOR2X1  NOR2X1_22
timestamp 1743127117
transform 1 0 2136 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_49
timestamp 1743127117
transform -1 0 2216 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_3
timestamp 1743127117
transform -1 0 2280 0 1 4210
box -4 -6 68 206
use OR2X2  OR2X2_5
timestamp 1743127117
transform -1 0 2344 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_21
timestamp 1743127117
transform -1 0 2392 0 1 4210
box -4 -6 52 206
use DFFSR  DFFSR_56
timestamp 1743127117
transform -1 0 2744 0 1 4210
box -4 -6 356 206
use FILL  FILL_21_1_0
timestamp 1743127117
transform -1 0 2760 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_1
timestamp 1743127117
transform -1 0 2776 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_2
timestamp 1743127117
transform -1 0 2792 0 1 4210
box -4 -6 20 206
use NAND2X1  NAND2X1_124
timestamp 1743127117
transform -1 0 2840 0 1 4210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_39
timestamp 1743127117
transform -1 0 2984 0 1 4210
box -4 -6 148 206
use OAI21X1  OAI21X1_434
timestamp 1743127117
transform 1 0 2984 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_433
timestamp 1743127117
transform -1 0 3112 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_150
timestamp 1743127117
transform -1 0 3144 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_45
timestamp 1743127117
transform 1 0 3144 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_49
timestamp 1743127117
transform -1 0 3240 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_144
timestamp 1743127117
transform 1 0 3240 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_145
timestamp 1743127117
transform 1 0 3288 0 1 4210
box -4 -6 52 206
use INVX2  INVX2_5
timestamp 1743127117
transform 1 0 3336 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_427
timestamp 1743127117
transform 1 0 3368 0 1 4210
box -4 -6 68 206
use OAI22X1  OAI22X1_1
timestamp 1743127117
transform -1 0 3512 0 1 4210
box -4 -6 84 206
use INVX1  INVX1_147
timestamp 1743127117
transform -1 0 3544 0 1 4210
box -4 -6 36 206
use OAI22X1  OAI22X1_3
timestamp 1743127117
transform -1 0 3624 0 1 4210
box -4 -6 84 206
use NAND3X1  NAND3X1_37
timestamp 1743127117
transform -1 0 3688 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_146
timestamp 1743127117
transform -1 0 3720 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_33
timestamp 1743127117
transform -1 0 3784 0 1 4210
box -4 -6 68 206
use AND2X2  AND2X2_5
timestamp 1743127117
transform -1 0 3848 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_4
timestamp 1743127117
transform -1 0 3896 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_327
timestamp 1743127117
transform -1 0 3960 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_98
timestamp 1743127117
transform 1 0 3960 0 1 4210
box -4 -6 52 206
use FILL  FILL_21_2_0
timestamp 1743127117
transform 1 0 4008 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_1
timestamp 1743127117
transform 1 0 4024 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_2
timestamp 1743127117
transform 1 0 4040 0 1 4210
box -4 -6 20 206
use DFFSR  DFFSR_132
timestamp 1743127117
transform 1 0 4056 0 1 4210
box -4 -6 356 206
use INVX1  INVX1_144
timestamp 1743127117
transform -1 0 4440 0 1 4210
box -4 -6 36 206
use BUFX4  BUFX4_89
timestamp 1743127117
transform -1 0 4504 0 1 4210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_23
timestamp 1743127117
transform -1 0 4648 0 1 4210
box -4 -6 148 206
use DFFSR  DFFSR_126
timestamp 1743127117
transform 1 0 4648 0 1 4210
box -4 -6 356 206
use OAI21X1  OAI21X1_410
timestamp 1743127117
transform -1 0 5064 0 1 4210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_33
timestamp 1743127117
transform 1 0 5064 0 1 4210
box -4 -6 148 206
use BUFX4  BUFX4_23
timestamp 1743127117
transform -1 0 5272 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_412
timestamp 1743127117
transform 1 0 5272 0 1 4210
box -4 -6 68 206
use OR2X2  OR2X2_12
timestamp 1743127117
transform 1 0 5336 0 1 4210
box -4 -6 68 206
use BUFX4  BUFX4_90
timestamp 1743127117
transform 1 0 5400 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_330
timestamp 1743127117
transform -1 0 5528 0 1 4210
box -4 -6 68 206
use DFFSR  DFFSR_59
timestamp 1743127117
transform -1 0 5880 0 1 4210
box -4 -6 356 206
use FILL  FILL_21_3_0
timestamp 1743127117
transform 1 0 5880 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_3_1
timestamp 1743127117
transform 1 0 5896 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_3_2
timestamp 1743127117
transform 1 0 5912 0 1 4210
box -4 -6 20 206
use BUFX4  BUFX4_85
timestamp 1743127117
transform 1 0 5928 0 1 4210
box -4 -6 68 206
use DFFSR  DFFSR_70
timestamp 1743127117
transform -1 0 6344 0 1 4210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_37
timestamp 1743127117
transform -1 0 6488 0 1 4210
box -4 -6 148 206
use DFFSR  DFFSR_72
timestamp 1743127117
transform -1 0 6840 0 1 4210
box -4 -6 356 206
use FILL  FILL_22_1
timestamp 1743127117
transform 1 0 6840 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_2
timestamp 1743127117
transform 1 0 6856 0 1 4210
box -4 -6 20 206
use FILL  FILL_22_3
timestamp 1743127117
transform 1 0 6872 0 1 4210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_58
timestamp 1743127117
transform -1 0 200 0 -1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_221
timestamp 1743127117
transform 1 0 200 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_220
timestamp 1743127117
transform -1 0 328 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_403
timestamp 1743127117
transform 1 0 328 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_123
timestamp 1743127117
transform -1 0 440 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_224
timestamp 1743127117
transform 1 0 440 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_225
timestamp 1743127117
transform -1 0 568 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_72
timestamp 1743127117
transform -1 0 664 0 -1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_191
timestamp 1743127117
transform -1 0 728 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_190
timestamp 1743127117
transform -1 0 792 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_70
timestamp 1743127117
transform 1 0 792 0 -1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_181
timestamp 1743127117
transform 1 0 984 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_182
timestamp 1743127117
transform -1 0 1112 0 -1 4610
box -4 -6 68 206
use FILL  FILL_22_0_0
timestamp 1743127117
transform -1 0 1128 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_1
timestamp 1743127117
transform -1 0 1144 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_2
timestamp 1743127117
transform -1 0 1160 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_67
timestamp 1743127117
transform -1 0 1352 0 -1 4610
box -4 -6 196 206
use INVX1  INVX1_71
timestamp 1743127117
transform -1 0 1384 0 -1 4610
box -4 -6 36 206
use MUX2X1  MUX2X1_65
timestamp 1743127117
transform 1 0 1384 0 -1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_211
timestamp 1743127117
transform 1 0 1480 0 -1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_71
timestamp 1743127117
transform 1 0 1544 0 -1 4610
box -4 -6 100 206
use NOR2X1  NOR2X1_27
timestamp 1743127117
transform 1 0 1640 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_223
timestamp 1743127117
transform 1 0 1688 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_59
timestamp 1743127117
transform 1 0 1752 0 -1 4610
box -4 -6 196 206
use NOR2X1  NOR2X1_30
timestamp 1743127117
transform 1 0 1944 0 -1 4610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_8
timestamp 1743127117
transform -1 0 2104 0 -1 4610
box -4 -6 116 206
use NAND3X1  NAND3X1_15
timestamp 1743127117
transform -1 0 2168 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_200
timestamp 1743127117
transform 1 0 2168 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_59
timestamp 1743127117
transform 1 0 2232 0 -1 4610
box -4 -6 36 206
use DFFSR  DFFSR_57
timestamp 1743127117
transform -1 0 2616 0 -1 4610
box -4 -6 356 206
use FILL  FILL_22_1_0
timestamp 1743127117
transform 1 0 2616 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_1
timestamp 1743127117
transform 1 0 2632 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_2
timestamp 1743127117
transform 1 0 2648 0 -1 4610
box -4 -6 20 206
use DFFSR  DFFSR_139
timestamp 1743127117
transform 1 0 2664 0 -1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_435
timestamp 1743127117
transform -1 0 3080 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_8
timestamp 1743127117
transform -1 0 3144 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_52
timestamp 1743127117
transform -1 0 3192 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_35
timestamp 1743127117
transform -1 0 3256 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_430
timestamp 1743127117
transform -1 0 3320 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_429
timestamp 1743127117
transform -1 0 3384 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_43
timestamp 1743127117
transform 1 0 3384 0 -1 4610
box -4 -6 52 206
use OAI22X1  OAI22X1_2
timestamp 1743127117
transform 1 0 3432 0 -1 4610
box -4 -6 84 206
use OAI22X1  OAI22X1_4
timestamp 1743127117
transform 1 0 3512 0 -1 4610
box -4 -6 84 206
use INVX1  INVX1_149
timestamp 1743127117
transform -1 0 3624 0 -1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_34
timestamp 1743127117
transform -1 0 3688 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_32
timestamp 1743127117
transform -1 0 3752 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_47
timestamp 1743127117
transform 1 0 3752 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_38
timestamp 1743127117
transform 1 0 3800 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_36
timestamp 1743127117
transform 1 0 3864 0 -1 4610
box -4 -6 68 206
use DFFSR  DFFSR_64
timestamp 1743127117
transform -1 0 4280 0 -1 4610
box -4 -6 356 206
use FILL  FILL_22_2_0
timestamp 1743127117
transform 1 0 4280 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_1
timestamp 1743127117
transform 1 0 4296 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_2
timestamp 1743127117
transform 1 0 4312 0 -1 4610
box -4 -6 20 206
use NAND2X1  NAND2X1_109
timestamp 1743127117
transform 1 0 4328 0 -1 4610
box -4 -6 52 206
use DFFSR  DFFSR_123
timestamp 1743127117
transform 1 0 4376 0 -1 4610
box -4 -6 356 206
use NAND2X1  NAND2X1_110
timestamp 1743127117
transform 1 0 4728 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_133
timestamp 1743127117
transform -1 0 4808 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_411
timestamp 1743127117
transform 1 0 4808 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_134
timestamp 1743127117
transform -1 0 4904 0 -1 4610
box -4 -6 36 206
use BUFX4  BUFX4_88
timestamp 1743127117
transform -1 0 4968 0 -1 4610
box -4 -6 68 206
use DFFSR  DFFSR_127
timestamp 1743127117
transform 1 0 4968 0 -1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_413
timestamp 1743127117
transform -1 0 5384 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_136
timestamp 1743127117
transform -1 0 5416 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_112
timestamp 1743127117
transform 1 0 5416 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_111
timestamp 1743127117
transform 1 0 5464 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_36
timestamp 1743127117
transform 1 0 5512 0 -1 4610
box -4 -6 52 206
use FILL  FILL_22_3_0
timestamp 1743127117
transform -1 0 5576 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_3_1
timestamp 1743127117
transform -1 0 5592 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_3_2
timestamp 1743127117
transform -1 0 5608 0 -1 4610
box -4 -6 20 206
use DFFSR  DFFSR_58
timestamp 1743127117
transform -1 0 5960 0 -1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_290
timestamp 1743127117
transform -1 0 6024 0 -1 4610
box -4 -6 68 206
use BUFX4  BUFX4_87
timestamp 1743127117
transform 1 0 6024 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_4
timestamp 1743127117
transform -1 0 6152 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_31
timestamp 1743127117
transform 1 0 6152 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_32
timestamp 1743127117
transform -1 0 6248 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_73
timestamp 1743127117
transform 1 0 6248 0 -1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_22
timestamp 1743127117
transform -1 0 6344 0 -1 4610
box -4 -6 68 206
use DFFSR  DFFSR_75
timestamp 1743127117
transform -1 0 6696 0 -1 4610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_36
timestamp 1743127117
transform 1 0 6696 0 -1 4610
box -4 -6 148 206
use FILL  FILL_23_1
timestamp 1743127117
transform -1 0 6856 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_2
timestamp 1743127117
transform -1 0 6872 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_3
timestamp 1743127117
transform -1 0 6888 0 -1 4610
box -4 -6 20 206
use DFFSR  DFFSR_117
timestamp 1743127117
transform -1 0 360 0 1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_397
timestamp 1743127117
transform -1 0 424 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_60
timestamp 1743127117
transform -1 0 472 0 1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_60
timestamp 1743127117
transform 1 0 472 0 1 4610
box -4 -6 196 206
use MUX2X1  MUX2X1_58
timestamp 1743127117
transform -1 0 760 0 1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_197
timestamp 1743127117
transform 1 0 760 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_196
timestamp 1743127117
transform -1 0 888 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_57
timestamp 1743127117
transform -1 0 936 0 1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_72
timestamp 1743127117
transform 1 0 936 0 1 4610
box -4 -6 196 206
use FILL  FILL_23_0_0
timestamp 1743127117
transform 1 0 1128 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_1
timestamp 1743127117
transform 1 0 1144 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_2
timestamp 1743127117
transform 1 0 1160 0 1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_212
timestamp 1743127117
transform 1 0 1176 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_213
timestamp 1743127117
transform -1 0 1304 0 1 4610
box -4 -6 68 206
use MUX2X1  MUX2X1_66
timestamp 1743127117
transform 1 0 1304 0 1 4610
box -4 -6 100 206
use DFFPOSX1  DFFPOSX1_65
timestamp 1743127117
transform -1 0 1592 0 1 4610
box -4 -6 196 206
use NAND2X1  NAND2X1_59
timestamp 1743127117
transform 1 0 1592 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_66
timestamp 1743127117
transform 1 0 1640 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_23
timestamp 1743127117
transform -1 0 1736 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_28
timestamp 1743127117
transform 1 0 1736 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_53
timestamp 1743127117
transform -1 0 1816 0 1 4610
box -4 -6 36 206
use INVX1  INVX1_52
timestamp 1743127117
transform -1 0 1848 0 1 4610
box -4 -6 36 206
use DFFSR  DFFSR_54
timestamp 1743127117
transform -1 0 2200 0 1 4610
box -4 -6 356 206
use XNOR2X1  XNOR2X1_7
timestamp 1743127117
transform 1 0 2200 0 1 4610
box -4 -6 116 206
use DFFSR  DFFSR_53
timestamp 1743127117
transform -1 0 2664 0 1 4610
box -4 -6 356 206
use FILL  FILL_23_1_0
timestamp 1743127117
transform 1 0 2664 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_1
timestamp 1743127117
transform 1 0 2680 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_2
timestamp 1743127117
transform 1 0 2696 0 1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_404
timestamp 1743127117
transform 1 0 2712 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_128
timestamp 1743127117
transform -1 0 2808 0 1 4610
box -4 -6 36 206
use CLKBUF1  CLKBUF1_5
timestamp 1743127117
transform 1 0 2808 0 1 4610
box -4 -6 148 206
use NOR2X1  NOR2X1_46
timestamp 1743127117
transform 1 0 2952 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_428
timestamp 1743127117
transform -1 0 3064 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_44
timestamp 1743127117
transform 1 0 3064 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_53
timestamp 1743127117
transform 1 0 3112 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_146
timestamp 1743127117
transform -1 0 3208 0 1 4610
box -4 -6 52 206
use AOI21X1  AOI21X1_7
timestamp 1743127117
transform -1 0 3272 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_133
timestamp 1743127117
transform 1 0 3272 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_134
timestamp 1743127117
transform 1 0 3320 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_425
timestamp 1743127117
transform 1 0 3368 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_136
timestamp 1743127117
transform 1 0 3432 0 1 4610
box -4 -6 52 206
use INVX4  INVX4_1
timestamp 1743127117
transform 1 0 3480 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_137
timestamp 1743127117
transform -1 0 3576 0 1 4610
box -4 -6 52 206
use INVX2  INVX2_6
timestamp 1743127117
transform -1 0 3608 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_139
timestamp 1743127117
transform 1 0 3608 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_426
timestamp 1743127117
transform -1 0 3720 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_138
timestamp 1743127117
transform 1 0 3720 0 1 4610
box -4 -6 52 206
use DFFSR  DFFSR_119
timestamp 1743127117
transform 1 0 3768 0 1 4610
box -4 -6 356 206
use INVX1  INVX1_140
timestamp 1743127117
transform 1 0 4120 0 1 4610
box -4 -6 36 206
use FILL  FILL_23_2_0
timestamp 1743127117
transform -1 0 4168 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_1
timestamp 1743127117
transform -1 0 4184 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_2
timestamp 1743127117
transform -1 0 4200 0 1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_421
timestamp 1743127117
transform -1 0 4264 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_129
timestamp 1743127117
transform -1 0 4312 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_353
timestamp 1743127117
transform -1 0 4376 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_354
timestamp 1743127117
transform 1 0 4376 0 1 4610
box -4 -6 68 206
use DFFSR  DFFSR_60
timestamp 1743127117
transform -1 0 4792 0 1 4610
box -4 -6 356 206
use DFFSR  DFFSR_63
timestamp 1743127117
transform 1 0 4792 0 1 4610
box -4 -6 356 206
use OAI21X1  OAI21X1_356
timestamp 1743127117
transform -1 0 5208 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_355
timestamp 1743127117
transform 1 0 5208 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_131
timestamp 1743127117
transform 1 0 5272 0 1 4610
box -4 -6 52 206
use DFFSR  DFFSR_62
timestamp 1743127117
transform -1 0 5672 0 1 4610
box -4 -6 356 206
use OR2X2  OR2X2_8
timestamp 1743127117
transform 1 0 5672 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_3_0
timestamp 1743127117
transform 1 0 5736 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_3_1
timestamp 1743127117
transform 1 0 5752 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_3_2
timestamp 1743127117
transform 1 0 5768 0 1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_287
timestamp 1743127117
transform 1 0 5784 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_93
timestamp 1743127117
transform 1 0 5848 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_288
timestamp 1743127117
transform -1 0 5960 0 1 4610
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1743127117
transform -1 0 6024 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_83
timestamp 1743127117
transform -1 0 6056 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_289
timestamp 1743127117
transform -1 0 6120 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_92
timestamp 1743127117
transform 1 0 6120 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_91
timestamp 1743127117
transform -1 0 6216 0 1 4610
box -4 -6 52 206
use XOR2X1  XOR2X1_8
timestamp 1743127117
transform -1 0 6328 0 1 4610
box -4 -6 116 206
use MUX2X1  MUX2X1_85
timestamp 1743127117
transform 1 0 6328 0 1 4610
box -4 -6 100 206
use MUX2X1  MUX2X1_86
timestamp 1743127117
transform 1 0 6424 0 1 4610
box -4 -6 100 206
use OAI21X1  OAI21X1_104
timestamp 1743127117
transform -1 0 6584 0 1 4610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_39
timestamp 1743127117
transform -1 0 6776 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_25
timestamp 1743127117
transform 1 0 6776 0 1 4610
box -4 -6 52 206
use FILL  FILL_24_1
timestamp 1743127117
transform 1 0 6824 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_2
timestamp 1743127117
transform 1 0 6840 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_3
timestamp 1743127117
transform 1 0 6856 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_4
timestamp 1743127117
transform 1 0 6872 0 1 4610
box -4 -6 20 206
use DFFSR  DFFSR_114
timestamp 1743127117
transform 1 0 8 0 -1 5010
box -4 -6 356 206
use OAI21X1  OAI21X1_398
timestamp 1743127117
transform -1 0 424 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_125
timestamp 1743127117
transform -1 0 456 0 -1 5010
box -4 -6 36 206
use DFFSR  DFFSR_111
timestamp 1743127117
transform 1 0 456 0 -1 5010
box -4 -6 356 206
use INVX1  INVX1_122
timestamp 1743127117
transform 1 0 808 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_392
timestamp 1743127117
transform 1 0 840 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_391
timestamp 1743127117
transform -1 0 968 0 -1 5010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_21
timestamp 1743127117
transform -1 0 1112 0 -1 5010
box -4 -6 148 206
use FILL  FILL_24_0_0
timestamp 1743127117
transform 1 0 1112 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_1
timestamp 1743127117
transform 1 0 1128 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_2
timestamp 1743127117
transform 1 0 1144 0 -1 5010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_66
timestamp 1743127117
transform 1 0 1160 0 -1 5010
box -4 -6 196 206
use CLKBUF1  CLKBUF1_41
timestamp 1743127117
transform -1 0 1496 0 -1 5010
box -4 -6 148 206
use OAI21X1  OAI21X1_395
timestamp 1743127117
transform 1 0 1496 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_124
timestamp 1743127117
transform 1 0 1560 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_396
timestamp 1743127117
transform 1 0 1592 0 -1 5010
box -4 -6 68 206
use DFFSR  DFFSR_113
timestamp 1743127117
transform -1 0 2008 0 -1 5010
box -4 -6 356 206
use INVX1  INVX1_121
timestamp 1743127117
transform 1 0 2008 0 -1 5010
box -4 -6 36 206
use DFFSR  DFFSR_109
timestamp 1743127117
transform -1 0 2392 0 -1 5010
box -4 -6 356 206
use CLKBUF1  CLKBUF1_26
timestamp 1743127117
transform -1 0 2536 0 -1 5010
box -4 -6 148 206
use FILL  FILL_24_1_0
timestamp 1743127117
transform 1 0 2536 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_1
timestamp 1743127117
transform 1 0 2552 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_2
timestamp 1743127117
transform 1 0 2568 0 -1 5010
box -4 -6 20 206
use DFFSR  DFFSR_105
timestamp 1743127117
transform 1 0 2584 0 -1 5010
box -4 -6 356 206
use BUFX2  BUFX2_14
timestamp 1743127117
transform 1 0 2936 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_136
timestamp 1743127117
transform 1 0 2984 0 -1 5010
box -4 -6 356 206
use XNOR2X1  XNOR2X1_13
timestamp 1743127117
transform 1 0 3336 0 -1 5010
box -4 -6 116 206
use DFFSR  DFFSR_138
timestamp 1743127117
transform -1 0 3800 0 -1 5010
box -4 -6 356 206
use BUFX2  BUFX2_19
timestamp 1743127117
transform -1 0 3848 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_120
timestamp 1743127117
transform -1 0 4200 0 -1 5010
box -4 -6 356 206
use FILL  FILL_24_2_0
timestamp 1743127117
transform 1 0 4200 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_1
timestamp 1743127117
transform 1 0 4216 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_2
timestamp 1743127117
transform 1 0 4232 0 -1 5010
box -4 -6 20 206
use BUFX2  BUFX2_18
timestamp 1743127117
transform 1 0 4248 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_141
timestamp 1743127117
transform 1 0 4296 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_422
timestamp 1743127117
transform 1 0 4328 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_130
timestamp 1743127117
transform 1 0 4392 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_61
timestamp 1743127117
transform -1 0 4792 0 -1 5010
box -4 -6 356 206
use INVX1  INVX1_137
timestamp 1743127117
transform 1 0 4792 0 -1 5010
box -4 -6 36 206
use INVX1  INVX1_135
timestamp 1743127117
transform -1 0 4856 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_21
timestamp 1743127117
transform 1 0 4856 0 -1 5010
box -4 -6 52 206
use DFFSR  DFFSR_122
timestamp 1743127117
transform -1 0 5256 0 -1 5010
box -4 -6 356 206
use INVX1  INVX1_143
timestamp 1743127117
transform 1 0 5256 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_424
timestamp 1743127117
transform 1 0 5288 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_132
timestamp 1743127117
transform -1 0 5400 0 -1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_423
timestamp 1743127117
transform -1 0 5464 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_142
timestamp 1743127117
transform -1 0 5496 0 -1 5010
box -4 -6 36 206
use DFFSR  DFFSR_121
timestamp 1743127117
transform -1 0 5848 0 -1 5010
box -4 -6 356 206
use FILL  FILL_24_3_0
timestamp 1743127117
transform 1 0 5848 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_3_1
timestamp 1743127117
transform 1 0 5864 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_3_2
timestamp 1743127117
transform 1 0 5880 0 -1 5010
box -4 -6 20 206
use DFFSR  DFFSR_76
timestamp 1743127117
transform 1 0 5896 0 -1 5010
box -4 -6 356 206
use XOR2X1  XOR2X1_7
timestamp 1743127117
transform 1 0 6248 0 -1 5010
box -4 -6 116 206
use CLKBUF1  CLKBUF1_32
timestamp 1743127117
transform 1 0 6360 0 -1 5010
box -4 -6 148 206
use DFFSR  DFFSR_74
timestamp 1743127117
transform -1 0 6856 0 -1 5010
box -4 -6 356 206
use FILL  FILL_25_1
timestamp 1743127117
transform -1 0 6872 0 -1 5010
box -4 -6 20 206
use FILL  FILL_25_2
timestamp 1743127117
transform -1 0 6888 0 -1 5010
box -4 -6 20 206
<< labels >>
flabel metal4 s 1112 -40 1160 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 2632 -40 2680 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 2157 -23 2163 -17 7 FreeSans 24 270 0 0 clk
port 2 nsew
flabel metal2 s 3229 -23 3235 -17 7 FreeSans 24 270 0 0 rst
port 3 nsew
flabel metal3 s -19 2097 -13 2103 7 FreeSans 24 0 0 0 ext_data_in[0]
port 4 nsew
flabel metal2 s 365 -23 371 -17 7 FreeSans 24 270 0 0 ext_data_in[1]
port 5 nsew
flabel metal3 s -19 1897 -13 1903 7 FreeSans 24 0 0 0 ext_data_in[2]
port 6 nsew
flabel metal2 s 445 -23 451 -17 7 FreeSans 24 270 0 0 ext_data_in[3]
port 7 nsew
flabel metal2 s 5405 -23 5411 -17 7 FreeSans 24 270 0 0 ext_data_in[4]
port 8 nsew
flabel metal2 s 5021 -23 5027 -17 7 FreeSans 24 270 0 0 ext_data_in[5]
port 9 nsew
flabel metal2 s 4637 -23 4643 -17 7 FreeSans 24 270 0 0 ext_data_in[6]
port 10 nsew
flabel metal2 s 4925 -23 4931 -17 7 FreeSans 24 270 0 0 ext_data_in[7]
port 11 nsew
flabel metal2 s 813 5037 819 5043 3 FreeSans 24 90 0 0 ext_data_in[8]
port 12 nsew
flabel metal3 s -19 2897 -13 2903 7 FreeSans 24 0 0 0 ext_data_in[9]
port 13 nsew
flabel metal2 s 1565 5037 1571 5043 3 FreeSans 24 90 0 0 ext_data_in[10]
port 14 nsew
flabel metal2 s 429 5037 435 5043 3 FreeSans 24 90 0 0 ext_data_in[11]
port 15 nsew
flabel metal2 s 4845 5037 4851 5043 3 FreeSans 24 90 0 0 ext_data_in[12]
port 16 nsew
flabel metal2 s 4877 5037 4883 5043 3 FreeSans 24 90 0 0 ext_data_in[13]
port 17 nsew
flabel metal2 s 5389 5037 5395 5043 3 FreeSans 24 90 0 0 ext_data_in[14]
port 18 nsew
flabel metal2 s 4797 5037 4803 5043 3 FreeSans 24 90 0 0 ext_data_in[15]
port 19 nsew
flabel metal2 s 3197 -23 3203 -17 7 FreeSans 24 270 0 0 ext_data_out[0]
port 20 nsew
flabel metal2 s 2413 -23 2419 -17 7 FreeSans 24 270 0 0 ext_data_out[1]
port 21 nsew
flabel metal2 s 2573 -23 2579 -17 7 FreeSans 24 270 0 0 ext_data_out[2]
port 22 nsew
flabel metal2 s 2701 -23 2707 -17 7 FreeSans 24 270 0 0 ext_data_out[3]
port 23 nsew
flabel metal2 s 3773 -23 3779 -17 7 FreeSans 24 270 0 0 ext_data_out[4]
port 24 nsew
flabel metal2 s 4205 -23 4211 -17 7 FreeSans 24 270 0 0 ext_data_out[5]
port 25 nsew
flabel metal2 s 3725 -23 3731 -17 7 FreeSans 24 270 0 0 ext_data_out[6]
port 26 nsew
flabel metal2 s 3325 -23 3331 -17 7 FreeSans 24 270 0 0 ext_data_out[7]
port 27 nsew
flabel metal2 s 2957 5037 2963 5043 3 FreeSans 24 90 0 0 ext_data_out[8]
port 28 nsew
flabel metal2 s 2237 5037 2243 5043 3 FreeSans 24 90 0 0 ext_data_out[9]
port 29 nsew
flabel metal3 s -19 2537 -13 2543 7 FreeSans 24 0 0 0 ext_data_out[10]
port 30 nsew
flabel metal3 s -19 2497 -13 2503 7 FreeSans 24 0 0 0 ext_data_out[11]
port 31 nsew
flabel metal2 s 4269 5037 4275 5043 3 FreeSans 24 90 0 0 ext_data_out[12]
port 32 nsew
flabel metal2 s 3821 5037 3827 5043 3 FreeSans 24 90 0 0 ext_data_out[13]
port 33 nsew
flabel metal2 s 5517 5037 5523 5043 3 FreeSans 24 90 0 0 ext_data_out[14]
port 34 nsew
flabel metal2 s 4909 5037 4915 5043 3 FreeSans 24 90 0 0 ext_data_out[15]
port 35 nsew
flabel metal2 s 413 -23 419 -17 7 FreeSans 24 270 0 0 pe_busy[0]
port 36 nsew
flabel metal2 s 5853 -23 5859 -17 7 FreeSans 24 270 0 0 pe_busy[1]
port 37 nsew
flabel metal3 s -19 3897 -13 3903 7 FreeSans 24 0 0 0 pe_busy[2]
port 38 nsew
flabel metal3 s 6909 4697 6915 4703 3 FreeSans 24 0 0 0 pe_busy[3]
port 39 nsew
<< end >>

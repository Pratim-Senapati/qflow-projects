magic
tech scmos
magscale 1 2
timestamp 1739819275
<< checkpaint >>
rect -76 -66 140 270
<< nwell >>
rect -16 96 80 210
<< ntransistor >>
rect 14 12 18 72
rect 24 12 28 72
rect 34 12 38 72
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
rect 46 148 50 188
<< ndiffusion >>
rect 4 71 14 72
rect 12 13 14 71
rect 4 12 14 13
rect 18 12 24 72
rect 28 12 34 72
rect 38 71 48 72
rect 38 13 40 71
rect 38 12 48 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 30 188
rect 18 149 20 187
rect 28 149 30 187
rect 18 148 30 149
rect 34 184 46 188
rect 34 156 36 184
rect 44 156 46 184
rect 34 148 46 156
rect 50 187 60 188
rect 50 149 52 187
rect 50 148 60 149
<< ndcontact >>
rect 4 13 12 71
rect 40 13 48 71
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 36 156 44 184
rect 52 149 60 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 14 106 18 148
rect 30 146 34 148
rect 12 98 18 106
rect 14 72 18 98
rect 24 142 34 146
rect 24 72 28 142
rect 46 126 50 148
rect 44 118 50 126
rect 46 78 50 118
rect 34 74 50 78
rect 34 72 38 74
rect 14 8 18 12
rect 24 8 28 12
rect 34 8 38 12
<< polycontact >>
rect 4 98 12 106
rect 36 118 44 126
rect 28 86 36 94
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 4 187 12 194
rect 4 148 12 149
rect 20 187 28 188
rect 36 184 44 194
rect 36 152 44 156
rect 52 187 60 188
rect 20 148 28 149
rect 22 146 28 148
rect 52 148 60 149
rect 52 146 58 148
rect 22 140 58 146
rect 36 126 44 134
rect 52 114 58 140
rect 4 106 12 114
rect 52 106 60 114
rect 20 86 28 94
rect 52 74 58 106
rect 42 72 58 74
rect 4 71 12 72
rect 4 6 12 13
rect 40 71 58 72
rect 48 68 58 71
rect 40 12 48 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 36 126 44 134
rect 4 106 12 114
rect 52 106 60 114
rect 20 86 28 94
<< labels >>
rlabel metal1 24 90 24 90 4 B
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 110 8 110 4 A
rlabel metal1 40 130 40 130 4 C
rlabel metal1 56 110 56 110 4 Y
<< end >>

* NGSPICE file created from sincos.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt sincos vdd gnd clk rst theta[0] theta[1] theta[2] theta[3] theta[4] theta[5]
+ theta[6] theta[7] sine[0] sine[1] sine[2] sine[3] sine[4] sine[5] sine[6] sine[7]
+ cosine[0] cosine[1] cosine[2] cosine[3] cosine[4] cosine[5] cosine[6] cosine[7]
+ done
XFILL_5_1_2 gnd vdd FILL
XAND2X2_5 OR2X2_8/A OR2X2_8/B gnd AND2X2_5/Y vdd AND2X2
XFILL_13_0_2 gnd vdd FILL
XDFFSR_9 DFFSR_9/Q DFFSR_6/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XOAI21X1_190 NOR2X1_109/Y NOR2X1_108/Y BUFX2_5/Y gnd OAI21X1_190/Y vdd OAI21X1
XNAND2X1_21 NAND2X1_21/A NAND2X1_21/B gnd NAND2X1_21/Y vdd NAND2X1
XNAND2X1_10 INVX1_11/A INVX2_1/A gnd NAND2X1_10/Y vdd NAND2X1
XNAND2X1_32 INVX2_2/A NOR2X1_22/B gnd OAI21X1_42/A vdd NAND2X1
XNAND2X1_43 INVX4_1/Y NOR2X1_30/Y gnd NAND2X1_43/Y vdd NAND2X1
XNAND2X1_87 NAND2X1_85/Y AOI21X1_19/B gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_98 INVX1_82/Y INVX1_85/Y gnd AOI22X1_11/B vdd NAND2X1
XNAND2X1_54 INVX2_4/A INVX1_48/Y gnd NAND2X1_54/Y vdd NAND2X1
XNAND2X1_76 INVX4_5/Y INVX1_68/Y gnd INVX1_69/A vdd NAND2X1
XNAND2X1_65 OR2X2_5/Y NAND2X1_65/B gnd OAI21X1_76/B vdd NAND2X1
XAOI22X1_30 BUFX4_24/Y AOI22X1_28/B INVX1_166/Y AOI22X1_30/D gnd AOI21X1_56/A vdd
+ AOI22X1
XOAI22X1_3 OAI22X1_3/A OAI22X1_3/B BUFX4_1/Y INVX1_24/Y gnd OAI22X1_3/Y vdd OAI22X1
XFILL_20_1_0 gnd vdd FILL
XINVX2_23 INVX2_23/A gnd INVX2_23/Y vdd INVX2
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XOAI21X1_19 INVX1_16/Y OAI21X1_17/Y INVX8_1/A gnd AOI21X1_1/B vdd OAI21X1
XFILL_19_2_0 gnd vdd FILL
XDFFPOSX1_103 DFFPOSX1_40/D CLKBUF1_10/Y XNOR2X1_69/Y gnd vdd DFFPOSX1
XFILL_12_3 gnd vdd FILL
XDFFPOSX1_114 OR2X2_9/A CLKBUF1_9/Y NOR2X1_89/Y gnd vdd DFFPOSX1
XNAND2X1_228 rst theta[2] gnd DFFSR_3/S vdd NAND2X1
XDFFPOSX1_136 BUFX2_6/A CLKBUF1_1/Y NAND2X1_67/Y gnd vdd DFFPOSX1
XNAND2X1_206 NOR2X1_141/Y XOR2X1_30/Y gnd OAI21X1_273/A vdd NAND2X1
XDFFPOSX1_147 INVX1_25/A CLKBUF1_5/Y XNOR2X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_125 INVX2_6/A CLKBUF1_6/Y XNOR2X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_169 INVX1_13/A DFFSR_8/CLK INVX1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 DFFPOSX1_49/D DFFSR_8/CLK NAND2X1_34/Y gnd vdd DFFPOSX1
XNAND2X1_217 OAI21X1_296/A NAND2X1_217/B gnd NOR2X1_155/A vdd NAND2X1
XOR2X2_22 OR2X2_18/A theta[7] gnd DFFSR_8/R vdd OR2X2
XOR2X2_11 OR2X2_11/A OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XXNOR2X1_6 XNOR2X1_6/A XNOR2X1_6/B gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_8_1_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XAND2X2_6 OR2X2_9/A OR2X2_9/B gnd AND2X2_6/Y vdd AND2X2
XOAI21X1_191 INVX1_122/A XNOR2X1_65/Y INVX1_129/Y gnd AOI22X1_20/D vdd OAI21X1
XOAI21X1_180 INVX1_125/A INVX1_124/A BUFX4_16/Y gnd OAI21X1_180/Y vdd OAI21X1
XAOI22X1_1 INVX2_2/Y INVX1_29/A AOI22X1_1/C NOR2X1_25/Y gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_66 OAI21X1_77/Y NAND3X1_5/Y gnd MUX2X1_1/B vdd NAND2X1
XNAND2X1_55 NAND2X1_55/A NAND2X1_54/Y gnd NOR2X1_42/B vdd NAND2X1
XNAND2X1_77 OR2X2_7/B INVX1_68/A gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_22 NAND2X1_21/Y OAI21X1_28/Y gnd NAND2X1_22/Y vdd NAND2X1
XNAND2X1_11 OAI21X1_12/C NAND2X1_11/B gnd NAND2X1_11/Y vdd NAND2X1
XNAND2X1_33 NOR2X1_22/B INVX1_29/A gnd NOR2X1_24/A vdd NAND2X1
XNAND2X1_44 INVX4_1/Y OAI21X1_57/Y gnd NAND2X1_44/Y vdd NAND2X1
XNAND2X1_99 INVX1_83/A INVX4_6/Y gnd NAND2X1_99/Y vdd NAND2X1
XNAND2X1_88 OR2X2_8/A OR2X2_8/B gnd NAND2X1_89/A vdd NAND2X1
XAOI22X1_20 BUFX4_17/Y AOI22X1_19/B NOR2X1_110/Y AOI22X1_20/D gnd AOI22X1_20/Y vdd
+ AOI22X1
XAOI22X1_31 AOI22X1_31/A AOI21X1_63/Y INVX8_2/A AOI22X1_31/D gnd AOI22X1_31/Y vdd
+ AOI22X1
XOAI22X1_4 INVX4_4/A OAI22X1_4/B OAI22X1_5/A INVX1_26/Y gnd XOR2X1_2/B vdd OAI22X1
XFILL_20_1_1 gnd vdd FILL
XINVX2_24 INVX2_24/A gnd INVX2_24/Y vdd INVX2
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_104 DFFPOSX1_41/D CLKBUF1_7/Y XNOR2X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_137 INVX1_62/A CLKBUF1_5/Y NAND2X1_87/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 INVX1_54/A CLKBUF1_6/Y XNOR2X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 INVX1_102/A CLKBUF1_9/Y XNOR2X1_54/Y gnd vdd DFFPOSX1
XNAND2X1_229 rst theta[3] gnd DFFSR_4/S vdd NAND2X1
XNAND2X1_218 AOI21X1_67/B AOI21X1_67/A gnd NAND2X1_218/Y vdd NAND2X1
XDFFPOSX1_148 NOR2X1_21/A CLKBUF1_5/Y XNOR2X1_35/Y gnd vdd DFFPOSX1
XNAND2X1_207 INVX1_44/Y INVX1_57/Y gnd AOI22X1_32/B vdd NAND2X1
XDFFPOSX1_159 DFFPOSX1_50/D CLKBUF1_10/Y XNOR2X1_16/Y gnd vdd DFFPOSX1
XBUFX4_20 INVX8_4/Y gnd DFFSR_9/R vdd BUFX4
XFILL_10_1 gnd vdd FILL
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 XNOR2X1_7/A INVX1_16/A gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A INVX2_14/A gnd AND2X2_7/Y vdd AND2X2
XAOI22X1_2 INVX2_3/A INVX1_34/A AOI22X1_2/C AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XOAI21X1_192 OR2X2_12/A OR2X2_12/B BUFX4_18/Y gnd OAI21X1_192/Y vdd OAI21X1
XOAI21X1_181 OAI21X1_181/A AOI21X1_37/Y OAI21X1_180/Y gnd AOI21X1_40/A vdd OAI21X1
XOAI21X1_170 INVX2_19/A INVX4_7/A NAND3X1_12/C gnd MUX2X1_9/A vdd OAI21X1
XNAND2X1_67 NAND3X1_6/Y OAI21X1_86/Y gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_78 NAND2X1_77/Y INVX1_69/A gnd NOR2X1_56/B vdd NAND2X1
XNAND2X1_56 OAI21X1_66/Y NOR2X1_42/B gnd AOI22X1_4/D vdd NAND2X1
XNAND2X1_89 NAND2X1_89/A OR2X2_8/Y gnd XOR2X1_10/B vdd NAND2X1
XNAND2X1_12 NAND2X1_11/Y OAI21X1_13/Y gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_23 DFFPOSX1_8/Q BUFX4_1/Y gnd NAND2X1_23/Y vdd NAND2X1
XNAND2X1_34 OAI21X1_41/Y AOI22X1_1/Y gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_45 INVX1_42/Y AOI21X1_7/Y gnd INVX1_43/A vdd NAND2X1
XAOI22X1_21 BUFX4_17/Y OR2X2_12/Y INVX1_133/Y AOI21X1_40/A gnd AOI22X1_21/Y vdd AOI22X1
XAOI22X1_32 INVX2_27/A AOI22X1_32/B INVX1_180/A AOI22X1_32/D gnd MUX2X1_12/A vdd AOI22X1
XAOI22X1_10 OR2X2_7/B AOI22X1_8/B NAND2X1_80/B INVX1_72/Y gnd AOI22X1_10/Y vdd AOI22X1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B INVX4_4/A OAI22X1_5/D gnd OAI22X1_5/Y vdd OAI22X1
XFILL_20_1_2 gnd vdd FILL
XINVX2_25 INVX2_25/A gnd INVX2_25/Y vdd INVX2
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XFILL_3_2_2 gnd vdd FILL
XFILL_11_1_2 gnd vdd FILL
XFILL_19_2_2 gnd vdd FILL
XDFFPOSX1_138 OR2X2_7/A CLKBUF1_3/Y XOR2X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 INVX1_52/A CLKBUF1_6/Y XNOR2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 NOR2X1_22/B CLKBUF1_10/Y XNOR2X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 DFFPOSX1_42/D CLKBUF1_7/Y XNOR2X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 INVX2_14/A CLKBUF1_9/Y XNOR2X1_55/Y gnd vdd DFFPOSX1
XNAND2X1_219 BUFX4_9/Y AOI21X1_69/A gnd OAI21X1_290/C vdd NAND2X1
XNAND2X1_208 XNOR2X1_94/Y INVX1_177/Y gnd INVX1_178/A vdd NAND2X1
XINVX8_1 INVX8_1/A gnd BUFX4_8/A vdd INVX8
XBUFX4_21 INVX8_4/Y gnd OR2X2_18/A vdd BUFX4
XBUFX4_10 BUFX4_8/A gnd BUFX4_10/Y vdd BUFX4
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XXNOR2X1_8 XNOR2X1_8/A XNOR2X1_8/B gnd XNOR2X1_8/Y vdd XNOR2X1
XFILL_0_0_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_8_1_2 gnd vdd FILL
XFILL_16_0_2 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XXOR2X1_30 INVX2_27/A XOR2X1_30/B gnd XOR2X1_30/Y vdd XOR2X1
XOAI21X1_182 INVX1_125/A INVX1_124/A INVX4_8/Y gnd OAI21X1_182/Y vdd OAI21X1
XOAI21X1_160 INVX1_108/A AOI21X1_27/Y OAI21X1_160/C gnd OAI21X1_162/B vdd OAI21X1
XAOI22X1_3 INVX1_43/A DFFSR_7/Q INVX4_1/Y AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_171 INVX2_19/A INVX4_7/Y AOI21X1_36/A gnd AOI21X1_35/C vdd OAI21X1
XOAI21X1_193 NOR2X1_99/Y NOR2X1_101/B INVX1_128/Y gnd INVX1_133/A vdd OAI21X1
XNAND2X1_68 INVX1_62/A INVX2_7/Y gnd NAND2X1_68/Y vdd NAND2X1
XNAND2X1_57 BUFX4_6/Y OAI21X1_69/Y gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_79 NOR2X1_56/A NOR2X1_56/B gnd NAND2X1_79/Y vdd NAND2X1
XNAND2X1_46 INVX1_45/A INVX1_44/Y gnd NAND2X1_48/A vdd NAND2X1
XNAND2X1_35 INVX2_2/A NOR2X1_23/B gnd OAI22X1_5/D vdd NAND2X1
XNAND2X1_24 DFFPOSX1_8/Q NOR2X1_16/Y gnd INVX1_24/A vdd NAND2X1
XNAND2X1_13 INVX1_12/Y INVX1_13/Y gnd OR2X2_1/A vdd NAND2X1
XAOI22X1_11 INVX4_6/Y AOI22X1_11/B AOI22X1_11/C NOR2X1_65/Y gnd AOI22X1_11/Y vdd AOI22X1
XAOI22X1_33 INVX2_27/Y AOI22X1_32/B INVX1_178/Y AOI22X1_33/D gnd AOI22X1_33/Y vdd
+ AOI22X1
XAOI22X1_22 INVX4_4/Y INVX1_134/Y AOI22X1_22/C INVX2_22/A gnd XNOR2X1_67/A vdd AOI22X1
XOAI22X1_6 INVX1_35/Y OAI22X1_7/D INVX2_3/Y OR2X2_4/Y gnd XOR2X1_4/A vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XINVX2_26 BUFX4_26/Y gnd INVX2_26/Y vdd INVX2
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XDFFPOSX1_139 INVX1_65/A CLKBUF1_3/Y XNOR2X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 INVX2_27/A CLKBUF1_6/Y NAND2X1_123/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 DFFPOSX1_43/D DFFSR_2/CLK XNOR2X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 INVX2_13/A CLKBUF1_9/Y XNOR2X1_56/Y gnd vdd DFFPOSX1
XNAND2X1_209 NAND3X1_19/Y OAI21X1_282/Y gnd NAND2X1_209/Y vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd BUFX2_1/A vdd INVX8
XBUFX4_22 INVX8_4/Y gnd BUFX4_22/Y vdd BUFX4
XBUFX4_11 BUFX4_8/A gnd BUFX4_11/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XOR2X2_14 OR2X2_14/A OR2X2_14/B gnd OR2X2_14/Y vdd OR2X2
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XXNOR2X1_9 XNOR2X1_9/A INVX1_19/A gnd XNOR2X1_9/Y vdd XNOR2X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_9_2 gnd vdd FILL
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XXOR2X1_20 XOR2X1_20/A XOR2X1_20/B gnd XOR2X1_20/Y vdd XOR2X1
XXOR2X1_31 OR2X2_5/B INVX2_27/A gnd XOR2X1_31/Y vdd XOR2X1
XOAI21X1_194 INVX1_133/A AOI22X1_20/Y OAI21X1_192/Y gnd XNOR2X1_66/A vdd OAI21X1
XOAI21X1_183 AND2X2_8/Y OAI21X1_183/B OAI21X1_182/Y gnd AOI22X1_18/C vdd OAI21X1
XAOI22X1_4 INVX1_49/Y INVX2_5/Y AOI22X1_4/C AOI22X1_4/D gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_161 INVX2_15/A INVX2_12/Y INVX8_3/A gnd INVX1_112/A vdd OAI21X1
XOAI21X1_150 BUFX4_3/Y AOI21X1_26/A NAND2X1_117/Y gnd XNOR2X1_49/A vdd OAI21X1
XOAI21X1_172 INVX4_7/A INVX2_19/Y INVX8_1/A gnd OAI21X1_173/A vdd OAI21X1
XNAND2X1_14 BUFX4_10/Y NOR2X1_8/Y gnd OAI22X1_2/B vdd NAND2X1
XNAND2X1_25 OAI21X1_35/Y OAI21X1_34/Y gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_69 INVX2_7/A INVX1_62/Y gnd OAI21X1_89/C vdd NAND2X1
XNAND2X1_58 INVX2_5/Y INVX2_6/Y gnd NAND2X1_60/B vdd NAND2X1
XNAND2X1_47 INVX1_44/A INVX1_45/Y gnd AOI21X1_8/B vdd NAND2X1
XNAND2X1_36 INVX2_3/Y INVX1_33/A gnd AOI22X1_2/C vdd NAND2X1
XAOI22X1_12 INVX4_6/Y AOI22X1_12/B INVX1_90/A AOI22X1_12/D gnd MUX2X1_7/A vdd AOI22X1
XAOI22X1_23 NOR2X1_116/B NOR2X1_111/Y NOR2X1_115/A INVX2_22/Y gnd XOR2X1_20/A vdd
+ AOI22X1
XOAI22X1_7 INVX2_3/A INVX1_37/Y OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XINVX2_27 INVX2_27/A gnd INVX2_27/Y vdd INVX2
XDFFPOSX1_107 INVX1_94/A DFFSR_8/CLK INVX4_1/Y gnd vdd DFFPOSX1
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_129 INVX1_79/A CLKBUF1_1/Y NAND2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_118 AND2X2_10/A CLKBUF1_13/Y XNOR2X1_57/Y gnd vdd DFFPOSX1
XFILL_3_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd BUFX4_3/A vdd INVX8
XBUFX4_23 INVX8_4/Y gnd DFFSR_11/R vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_12 BUFX4_13/A gnd OR2X2_7/B vdd BUFX4
XOR2X2_15 BUFX4_22/Y theta[0] gnd DFFSR_1/R vdd OR2X2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XFILL_9_3 gnd vdd FILL
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B gnd XOR2X1_10/Y vdd XOR2X1
XXOR2X1_21 INVX2_21/A XOR2X1_21/B gnd XOR2X1_21/Y vdd XOR2X1
XXOR2X1_32 BUFX2_57/A BUFX2_58/A gnd XOR2X1_32/Y vdd XOR2X1
XOAI21X1_140 INVX8_3/A INVX1_99/Y OAI21X1_140/C gnd XOR2X1_14/A vdd OAI21X1
XOAI21X1_195 BUFX2_2/Y XNOR2X1_66/Y OAI21X1_190/Y gnd OAI21X1_195/Y vdd OAI21X1
XAOI22X1_5 INVX2_5/Y AOI22X1_6/B INVX1_55/Y AOI22X1_5/D gnd MUX2X1_1/A vdd AOI22X1
XOAI21X1_184 BUFX2_2/Y AOI21X1_40/A NAND2X1_146/Y gnd XNOR2X1_62/A vdd OAI21X1
XOAI21X1_162 NOR2X1_82/Y OAI21X1_162/B INVX1_112/Y gnd NAND3X1_11/C vdd OAI21X1
XOAI21X1_173 OAI21X1_173/A AOI21X1_35/Y OAI21X1_173/C gnd OAI21X1_173/Y vdd OAI21X1
XOAI21X1_151 BUFX4_2/Y AOI21X1_26/Y NAND3X1_9/Y gnd XNOR2X1_51/A vdd OAI21X1
XNAND2X1_59 INVX2_5/A INVX2_6/A gnd NAND3X1_4/B vdd NAND2X1
XNAND2X1_48 NAND2X1_48/A AOI21X1_8/B gnd NAND2X1_48/Y vdd NAND2X1
XNAND2X1_26 OR2X2_3/A OR2X2_3/B gnd INVX1_26/A vdd NAND2X1
XNAND2X1_15 OR2X2_1/B NOR2X1_8/Y gnd NOR2X1_10/B vdd NAND2X1
XNAND2X1_37 XOR2X1_4/B OR2X2_4/B gnd OAI22X1_7/C vdd NAND2X1
XNAND2X1_190 INVX1_78/Y INVX1_156/Y gnd AOI22X1_28/B vdd NAND2X1
XAOI22X1_13 INVX4_6/A AOI22X1_11/B NAND2X1_92/A NOR2X1_70/Y gnd AOI22X1_13/Y vdd AOI22X1
XAOI22X1_24 INVX2_22/Y AOI22X1_24/B NOR2X1_111/Y AOI22X1_24/D gnd AOI22X1_24/Y vdd
+ AOI22X1
XXNOR2X1_90 XNOR2X1_90/A XOR2X1_29/Y gnd XNOR2X1_90/Y vdd XNOR2X1
XOAI22X1_8 OAI22X1_8/A BUFX2_58/A BUFX2_57/A NOR2X1_90/Y gnd OAI22X1_8/Y vdd OAI22X1
XFILL_6_2_2 gnd vdd FILL
XFILL_14_1_2 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B INVX8_2/A gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_108 BUFX2_55/A CLKBUF1_12/Y BUFX2_40/A gnd vdd DFFPOSX1
XDFFPOSX1_119 INVX2_15/A CLKBUF1_13/Y XOR2X1_16/Y gnd vdd DFFPOSX1
XCLKBUF1_2 clk gnd DFFSR_6/CLK vdd CLKBUF1
XFILL_3_0_2 gnd vdd FILL
XINVX8_4 rst gnd INVX8_4/Y vdd INVX8
XDFFPOSX1_90 BUFX4_13/A CLKBUF1_5/Y NAND2X1_192/Y gnd vdd DFFPOSX1
XFILL_19_0_2 gnd vdd FILL
XBUFX4_24 BUFX2_6/A gnd BUFX4_24/Y vdd BUFX4
XBUFX4_13 BUFX4_13/A gnd BUFX4_13/Y vdd BUFX4
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XOR2X2_16 BUFX4_22/Y theta[1] gnd DFFSR_2/R vdd OR2X2
XFILL_12_2_0 gnd vdd FILL
XXOR2X1_11 INVX4_6/A INVX1_85/A gnd XOR2X1_11/Y vdd XOR2X1
XXOR2X1_22 INVX2_14/A XOR2X1_22/B gnd XOR2X1_22/Y vdd XOR2X1
XXOR2X1_33 INVX1_118/A INVX4_7/A gnd XOR2X1_33/Y vdd XOR2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 INVX4_4/Y INVX1_25/Y NAND3X1_2/C gnd NAND3X1_1/Y vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 INVX4_6/Y INVX2_10/Y BUFX2_7/Y gnd INVX1_89/A vdd OAI21X1
XOAI21X1_141 NOR2X1_75/Y AND2X2_6/Y AOI21X1_23/B gnd OAI21X1_142/C vdd OAI21X1
XOAI21X1_152 INVX1_100/Y INVX1_110/Y INVX1_99/A gnd OAI21X1_152/Y vdd OAI21X1
XOAI21X1_196 INVX4_8/A INVX2_7/Y BUFX2_5/Y gnd INVX1_130/A vdd OAI21X1
XAOI22X1_6 INVX2_5/A AOI22X1_6/B NAND3X1_5/B AOI22X1_4/Y gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_185 NOR2X1_102/Y AND2X2_9/Y BUFX2_2/Y gnd OAI21X1_186/C vdd OAI21X1
XOAI21X1_174 XOR2X1_17/B INVX2_8/Y BUFX2_4/Y gnd OAI21X1_174/Y vdd OAI21X1
XOAI21X1_163 AOI21X1_28/Y AOI21X1_29/Y INVX1_113/Y gnd NAND2X1_123/B vdd OAI21X1
XNAND2X1_180 BUFX2_6/Y INVX1_154/Y gnd AOI22X1_29/C vdd NAND2X1
XNAND2X1_191 INVX1_157/A INVX1_161/Y gnd INVX1_162/A vdd NAND2X1
XNAND2X1_49 OR2X2_5/A OR2X2_5/B gnd OAI21X1_66/C vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_27 INVX4_4/A INVX2_2/A gnd OAI22X1_5/A vdd NAND2X1
XNAND2X1_16 BUFX4_11/Y NOR2X1_11/B gnd NAND2X1_16/Y vdd NAND2X1
XNAND2X1_38 INVX2_3/A NOR2X1_28/Y gnd NAND2X1_38/Y vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_14 INVX4_6/A AOI22X1_12/B NAND2X1_97/B INVX1_88/Y gnd AOI22X1_14/Y vdd AOI22X1
XAOI22X1_25 INVX2_25/A AOI22X1_25/B INVX1_149/A AOI21X1_48/A gnd MUX2X1_10/A vdd AOI22X1
XXNOR2X1_91 INVX1_54/A XOR2X1_29/B gnd XNOR2X1_91/Y vdd XNOR2X1
XXNOR2X1_80 XNOR2X1_80/A INVX2_24/Y gnd XNOR2X1_80/Y vdd XNOR2X1
XOAI22X1_9 XOR2X1_17/B INVX2_8/Y INVX4_8/Y OAI22X1_9/D gnd AND2X2_8/A vdd OAI22X1
XFILL_19_2 gnd vdd FILL
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 OR2X2_3/A INVX2_2/A gnd XOR2X1_1/Y vdd XOR2X1
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B INVX4_2/A gnd MUX2X1_2/Y vdd MUX2X1
XDFFPOSX1_109 BUFX2_57/A DFFSR_8/CLK BUFX2_18/Y gnd vdd DFFPOSX1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XBUFX4_25 BUFX2_6/A gnd BUFX4_25/Y vdd BUFX4
XBUFX4_14 BUFX4_13/A gnd XOR2X1_8/A vdd BUFX4
XDFFPOSX1_91 INVX1_134/A CLKBUF1_7/Y XOR2X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_80 INVX1_78/A CLKBUF1_1/Y XNOR2X1_97/Y gnd vdd DFFPOSX1
XOR2X2_17 OR2X2_18/A theta[2] gnd DFFSR_3/R vdd OR2X2
XFILL_12_2_1 gnd vdd FILL
XXOR2X1_12 INVX1_82/A INVX4_6/A gnd NOR2X1_65/B vdd XOR2X1
XXOR2X1_23 INVX2_13/A XOR2X1_23/B gnd XOR2X1_23/Y vdd XOR2X1
XXOR2X1_34 XOR2X1_34/A XOR2X1_34/B gnd XOR2X1_34/Y vdd XOR2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 INVX1_29/Y NOR2X1_22/Y NAND3X1_2/C gnd NOR2X1_23/B vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_142 INVX1_100/Y OR2X2_9/B OAI21X1_142/C gnd AOI21X1_27/B vdd OAI21X1
XOAI21X1_131 INVX1_87/A AOI22X1_14/Y INVX1_89/Y gnd NAND3X1_8/B vdd OAI21X1
XOAI21X1_120 INVX1_82/Y INVX4_6/Y NAND2X1_92/Y gnd MUX2X1_5/B vdd OAI21X1
XAOI22X1_7 INVX4_5/Y AOI22X1_7/B AOI22X1_7/C AOI22X1_7/D gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_153 XNOR2X1_47/B OAI21X1_153/B AOI21X1_25/Y gnd NAND3X1_10/C vdd OAI21X1
XOAI21X1_164 INVX1_116/A INVX1_117/Y OAI22X1_8/Y gnd AOI21X1_32/A vdd OAI21X1
XOAI21X1_197 INVX1_127/A NOR2X1_108/B INVX1_130/Y gnd NAND3X1_13/B vdd OAI21X1
XOAI21X1_186 BUFX2_2/Y XNOR2X1_64/Y OAI21X1_186/C gnd OAI21X1_186/Y vdd OAI21X1
XOAI21X1_175 BUFX2_4/Y INVX1_122/Y OAI21X1_174/Y gnd XNOR2X1_58/A vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_181 NAND2X1_181/A AOI22X1_29/C gnd XNOR2X1_84/B vdd NAND2X1
XNAND2X1_192 NAND3X1_18/Y OAI21X1_257/Y gnd NAND2X1_192/Y vdd NAND2X1
XNAND2X1_28 INVX2_2/A INVX1_25/Y gnd OAI21X1_38/B vdd NAND2X1
XNAND2X1_17 INVX8_1/A OAI21X1_17/Y gnd NAND2X1_17/Y vdd NAND2X1
XNAND2X1_39 OAI21X1_49/Y OAI21X1_50/Y gnd NAND2X1_40/A vdd NAND2X1
XNAND2X1_170 XOR2X1_23/B INVX2_13/Y gnd AOI21X1_44/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_26 INVX2_25/Y AOI22X1_25/B INVX1_147/Y AOI22X1_26/D gnd AOI22X1_26/Y vdd
+ AOI22X1
XAOI22X1_15 INVX1_103/Y INVX2_14/Y AOI21X1_25/Y AOI22X1_15/D gnd AOI22X1_15/Y vdd
+ AOI22X1
XXNOR2X1_92 XNOR2X1_92/A NOR2X1_141/Y gnd XNOR2X1_92/Y vdd XNOR2X1
XXNOR2X1_70 XNOR2X1_70/A INVX2_23/Y gnd XNOR2X1_70/Y vdd XNOR2X1
XXNOR2X1_81 MUX2X1_10/Y INVX1_144/Y gnd XNOR2X1_81/Y vdd XNOR2X1
XAOI21X1_70 INVX1_118/A INVX4_7/A MUX2X1_13/B gnd AOI21X1_70/Y vdd AOI21X1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B INVX4_2/A gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 clk gnd DFFSR_2/CLK vdd CLKBUF1
XDFFPOSX1_81 OR2X2_8/B CLKBUF1_1/Y XNOR2X1_98/Y gnd vdd DFFPOSX1
XDFFPOSX1_70 XOR2X1_30/B CLKBUF1_13/Y XNOR2X1_76/Y gnd vdd DFFPOSX1
XBUFX4_26 BUFX2_6/A gnd BUFX4_26/Y vdd BUFX4
XBUFX4_15 BUFX4_13/A gnd INVX4_5/A vdd BUFX4
XDFFPOSX1_92 INVX1_135/A CLKBUF1_7/Y XNOR2X1_58/Y gnd vdd DFFPOSX1
XOR2X2_18 OR2X2_18/A theta[3] gnd DFFSR_4/R vdd OR2X2
XFILL_12_2_2 gnd vdd FILL
XXOR2X1_13 MUX2X1_6/Y XOR2X1_13/B gnd XOR2X1_13/Y vdd XOR2X1
XXOR2X1_24 NOR2X1_78/A INVX2_25/A gnd INVX2_24/A vdd XOR2X1
XNAND3X1_3 INVX2_3/Y INVX1_36/A INVX1_33/Y gnd OAI22X1_7/D vdd NAND3X1
XFILL_1_1_2 gnd vdd FILL
XOAI21X1_165 INVX1_116/A BUFX2_58/A BUFX2_57/A gnd OAI21X1_166/B vdd OAI21X1
XOAI21X1_143 INVX1_99/A NOR2X1_75/Y NAND2X1_106/A gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_198 INVX2_7/A BUFX4_16/Y INVX4_2/A gnd INVX1_131/A vdd OAI21X1
XOAI21X1_132 INVX1_83/A INVX2_9/A INVX4_6/Y gnd OAI21X1_132/Y vdd OAI21X1
XOAI21X1_176 INVX4_2/A AND2X2_8/Y NAND2X1_136/Y gnd XNOR2X1_59/A vdd OAI21X1
XOAI21X1_187 OR2X2_12/A OR2X2_12/B INVX4_8/Y gnd OAI21X1_187/Y vdd OAI21X1
XOAI21X1_121 INVX1_82/A INVX1_85/A INVX4_6/Y gnd OAI21X1_121/Y vdd OAI21X1
XAOI22X1_8 INVX4_5/Y AOI22X1_8/B INVX1_74/A AOI22X1_8/D gnd MUX2X1_4/A vdd AOI22X1
XOAI21X1_110 INVX1_77/A OAI21X1_110/B INVX1_75/Y gnd NAND3X1_7/C vdd OAI21X1
XOAI21X1_154 INVX2_13/A AND2X2_10/A INVX2_12/A gnd NAND2X1_122/A vdd OAI21X1
XFILL_9_2_2 gnd vdd FILL
XNAND2X1_193 INVX1_167/A INVX2_6/Y gnd NAND2X1_195/A vdd NAND2X1
XNAND2X1_182 BUFX4_24/Y XOR2X1_27/B gnd OAI21X1_236/C vdd NAND2X1
XNAND2X1_160 OR2X2_13/A OR2X2_13/B gnd NOR2X1_115/B vdd NAND2X1
XNAND2X1_18 INVX1_19/Y NOR2X1_13/Y gnd INVX1_20/A vdd NAND2X1
XNAND2X1_29 OAI21X1_38/Y OAI21X1_39/Y gnd NAND2X1_29/Y vdd NAND2X1
XNAND2X1_171 BUFX4_3/Y OAI21X1_216/Y gnd OAI21X1_218/C vdd NAND2X1
XFILL_17_1_2 gnd vdd FILL
XAOI22X1_27 BUFX4_26/Y AOI22X1_29/B AOI22X1_27/C AOI22X1_27/D gnd AOI22X1_27/Y vdd
+ AOI22X1
XAOI22X1_16 INVX2_12/Y AOI22X1_17/B INVX1_108/Y AOI21X1_26/A gnd MUX2X1_8/A vdd AOI22X1
XXNOR2X1_60 XNOR2X1_60/A XNOR2X1_60/B gnd XNOR2X1_60/Y vdd XNOR2X1
XXNOR2X1_93 XNOR2X1_93/A XOR2X1_30/Y gnd XNOR2X1_93/Y vdd XNOR2X1
XXNOR2X1_82 XNOR2X1_82/A XOR2X1_26/Y gnd XNOR2X1_82/Y vdd XNOR2X1
XXNOR2X1_71 AOI22X1_24/Y XOR2X1_21/Y gnd XNOR2X1_71/Y vdd XNOR2X1
XAOI21X1_60 AOI21X1_60/A AOI21X1_59/Y AOI21X1_60/C gnd AOI21X1_60/Y vdd AOI21X1
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B INVX4_2/A gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_17_1 gnd vdd FILL
XDFFPOSX1_82 INVX4_6/A CLKBUF1_1/Y NAND2X1_209/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 OR2X2_13/A CLKBUF1_7/Y XNOR2X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 INVX1_44/A CLKBUF1_6/Y XNOR2X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_60 XOR2X1_23/B CLKBUF1_9/Y XNOR2X1_99/Y gnd vdd DFFPOSX1
XBUFX4_16 BUFX4_16/A gnd BUFX4_16/Y vdd BUFX4
XBUFX4_27 INVX4_3/Y gnd BUFX4_27/Y vdd BUFX4
XFILL_15_2_0 gnd vdd FILL
XOR2X2_19 DFFSR_11/R theta[4] gnd DFFSR_5/R vdd OR2X2
XXOR2X1_14 XOR2X1_14/A XOR2X1_14/B gnd XOR2X1_14/Y vdd XOR2X1
XXOR2X1_25 INVX2_9/A XOR2X1_25/B gnd XOR2X1_25/Y vdd XOR2X1
XBUFX4_1 BUFX4_3/A gnd BUFX4_1/Y vdd BUFX4
XFILL_4_1_0 gnd vdd FILL
XINVX4_1 DFFSR_8/Q gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_4 BUFX2_1/Y NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_166 NOR2X1_90/Y OAI21X1_166/B NAND2X1_125/Y gnd AOI21X1_33/B vdd OAI21X1
XOAI21X1_144 BUFX4_4/Y AOI21X1_27/B OAI21X1_144/C gnd XNOR2X1_47/A vdd OAI21X1
XOAI21X1_199 INVX1_132/A XNOR2X1_66/A INVX1_131/Y gnd NAND3X1_13/C vdd OAI21X1
XOAI21X1_188 INVX4_8/Y OR2X2_12/B INVX2_20/A gnd OAI21X1_189/A vdd OAI21X1
XOAI21X1_177 NOR2X1_110/B AOI21X1_37/Y OAI21X1_177/C gnd OAI21X1_177/Y vdd OAI21X1
XOAI21X1_133 AOI22X1_11/Y INVX1_90/Y OAI21X1_132/Y gnd OAI21X1_135/B vdd OAI21X1
XOAI21X1_122 NAND2X1_96/Y AOI21X1_19/Y OAI21X1_121/Y gnd AOI22X1_12/D vdd OAI21X1
XAOI22X1_9 OR2X2_7/B AOI22X1_7/B AOI22X1_9/C NOR2X1_56/Y gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_111 AOI21X1_17/Y AOI21X1_18/Y INVX1_76/Y gnd NAND2X1_84/B vdd OAI21X1
XOAI21X1_100 BUFX2_3/Y AOI22X1_8/D NAND2X1_80/Y gnd XNOR2X1_36/A vdd OAI21X1
XOAI21X1_155 INVX2_12/Y INVX2_15/Y BUFX4_1/Y gnd INVX1_111/A vdd OAI21X1
XNAND2X1_161 NAND3X1_15/Y NAND3X1_14/Y gnd XNOR2X1_70/A vdd NAND2X1
XNAND2X1_19 INVX1_19/A NOR2X1_14/Y gnd NAND2X1_19/Y vdd NAND2X1
XNAND2X1_150 INVX2_21/A INVX1_134/Y gnd AOI22X1_22/C vdd NAND2X1
XNAND2X1_194 INVX2_6/A INVX1_167/Y gnd AOI21X1_58/B vdd NAND2X1
XNAND2X1_183 INVX2_26/Y INVX1_155/Y gnd NAND2X1_183/Y vdd NAND2X1
XNAND2X1_172 AOI21X1_44/C AOI21X1_47/A gnd NAND2X1_172/Y vdd NAND2X1
XAOI22X1_28 INVX2_26/Y AOI22X1_28/B AOI22X1_28/C INVX1_162/Y gnd NOR2X1_138/B vdd
+ AOI22X1
XAOI22X1_17 INVX2_12/A AOI22X1_17/B NOR2X1_84/Y AOI22X1_15/Y gnd AOI22X1_17/Y vdd
+ AOI22X1
XXNOR2X1_61 BUFX4_17/Y INVX1_124/A gnd XNOR2X1_61/Y vdd XNOR2X1
XXNOR2X1_83 XNOR2X1_83/A XOR2X1_27/Y gnd XNOR2X1_83/Y vdd XNOR2X1
XFILL_5_1 gnd vdd FILL
XXNOR2X1_94 INVX1_44/A INVX2_27/A gnd XNOR2X1_94/Y vdd XNOR2X1
XXNOR2X1_72 XNOR2X1_72/A XOR2X1_3/B gnd XNOR2X1_72/Y vdd XNOR2X1
XXNOR2X1_50 INVX2_12/A AND2X2_10/A gnd INVX1_104/A vdd XNOR2X1
XAOI21X1_61 AOI21X1_61/A AOI21X1_61/B AOI21X1_61/C gnd AOI21X1_61/Y vdd AOI21X1
XOAI21X1_1 INVX1_5/Y OAI21X1_1/B INVX4_2/A gnd OAI21X1_1/Y vdd OAI21X1
XAOI21X1_50 MUX2X1_10/B INVX1_144/Y INVX1_148/A gnd AOI21X1_50/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B INVX4_3/A gnd MUX2X1_5/Y vdd MUX2X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XFILL_17_2 gnd vdd FILL
XDFFPOSX1_83 XOR2X1_17/B CLKBUF1_5/Y XOR2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 OR2X2_13/B CLKBUF1_7/Y XNOR2X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 OR2X2_5/B CLKBUF1_6/Y XNOR2X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 BUFX2_34/A CLKBUF1_10/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_61 AND2X2_10/B CLKBUF1_13/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XBUFX4_17 BUFX4_16/A gnd BUFX4_17/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XXOR2X1_26 INVX2_10/A XOR2X1_26/B gnd XOR2X1_26/Y vdd XOR2X1
XBUFX4_2 BUFX4_3/A gnd BUFX4_2/Y vdd BUFX4
XXOR2X1_15 INVX2_19/A INVX4_7/A gnd XOR2X1_34/B vdd XOR2X1
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 INVX1_56/Y NAND3X1_5/B NAND3X1_5/C gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_112 INVX1_79/A INVX1_78/Y INVX4_3/A gnd OAI21X1_112/Y vdd OAI21X1
XOAI21X1_101 INVX1_67/A AOI22X1_7/Y NAND2X1_82/Y gnd MUX2X1_3/A vdd OAI21X1
XOAI21X1_134 INVX2_10/A INVX4_6/Y INVX4_3/A gnd INVX1_91/A vdd OAI21X1
XOAI21X1_189 OAI21X1_189/A AOI22X1_19/Y OAI21X1_187/Y gnd NOR2X1_109/B vdd OAI21X1
XOAI21X1_178 NOR2X1_98/Y AOI21X1_38/Y BUFX2_5/Y gnd OAI21X1_178/Y vdd OAI21X1
XOAI21X1_123 INVX1_82/A INVX1_85/A INVX4_6/A gnd OAI21X1_124/C vdd OAI21X1
XOAI21X1_156 NOR2X1_83/Y AOI22X1_17/Y INVX1_111/Y gnd NAND3X1_11/B vdd OAI21X1
XOAI21X1_145 NOR2X1_86/B AOI21X1_23/Y NAND2X1_111/A gnd OAI21X1_147/B vdd OAI21X1
XOAI21X1_167 BUFX4_11/Y AOI21X1_32/A OAI21X1_167/C gnd XNOR2X1_56/A vdd OAI21X1
XNAND2X1_195 NAND2X1_195/A AOI21X1_58/B gnd DFFPOSX1_75/D vdd NAND2X1
XNAND2X1_140 NAND2X1_140/A AOI22X1_19/C gnd XNOR2X1_60/B vdd NAND2X1
XNAND2X1_184 OAI21X1_236/C NAND2X1_183/Y gnd NOR2X1_134/B vdd NAND2X1
XNAND2X1_162 NOR2X1_117/Y NOR2X1_115/Y gnd AOI22X1_24/B vdd NAND2X1
XNAND2X1_151 NAND2X1_149/Y AOI22X1_22/C gnd NAND2X1_151/Y vdd NAND2X1
XNAND2X1_173 INVX1_110/Y INVX1_101/Y gnd AOI22X1_25/B vdd NAND2X1
XAOI22X1_18 INVX4_8/Y OR2X2_12/Y AOI22X1_18/C AOI22X1_18/D gnd NOR2X1_108/B vdd AOI22X1
XAOI22X1_29 INVX2_26/Y AOI22X1_29/B AOI22X1_29/C AOI22X1_29/D gnd AOI22X1_29/Y vdd
+ AOI22X1
XXNOR2X1_62 XNOR2X1_62/A INVX2_20/Y gnd XNOR2X1_62/Y vdd XNOR2X1
XXNOR2X1_84 XNOR2X1_84/A XNOR2X1_84/B gnd XNOR2X1_84/Y vdd XNOR2X1
XFILL_5_2 gnd vdd FILL
XXNOR2X1_95 INVX2_27/A XOR2X1_30/B gnd XNOR2X1_95/Y vdd XNOR2X1
XXNOR2X1_40 XNOR2X1_40/A NOR2X1_70/A gnd XNOR2X1_40/Y vdd XNOR2X1
XXNOR2X1_51 XNOR2X1_51/A INVX1_104/Y gnd XNOR2X1_51/Y vdd XNOR2X1
XXNOR2X1_73 XNOR2X1_73/A XOR2X1_23/Y gnd XNOR2X1_73/Y vdd XNOR2X1
XBUFX2_50 vdd gnd BUFX2_50/Y vdd BUFX2
XAOI21X1_40 AOI21X1_40/A INVX2_20/Y NOR2X1_103/Y gnd XNOR2X1_64/A vdd AOI21X1
XAOI21X1_62 XNOR2X1_95/Y INVX1_175/Y INVX1_173/A gnd AOI21X1_62/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 INVX1_5/A OAI21X1_2/B BUFX2_3/Y gnd INVX1_7/A vdd OAI21X1
XAOI21X1_51 MUX2X1_10/A INVX1_151/Y INVX1_150/A gnd AOI21X1_51/Y vdd AOI21X1
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B INVX4_3/A gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XDFFPOSX1_62 INVX1_97/A CLKBUF1_9/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XDFFPOSX1_95 INVX1_137/A CLKBUF1_7/Y XNOR2X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 OAI22X1_9/D CLKBUF1_5/Y XNOR2X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 BUFX2_23/A CLKBUF1_10/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_73 INVX2_4/A CLKBUF1_6/Y XNOR2X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 BUFX2_35/A DFFSR_2/CLK DFFPOSX1_51/D gnd vdd DFFPOSX1
XBUFX4_18 BUFX4_16/A gnd BUFX4_18/Y vdd BUFX4
XFILL_15_2_2 gnd vdd FILL
XBUFX4_3 BUFX4_3/A gnd BUFX4_3/Y vdd BUFX4
XXOR2X1_27 BUFX4_25/Y XOR2X1_27/B gnd XOR2X1_27/Y vdd XOR2X1
XXOR2X1_16 MUX2X1_9/Y XOR2X1_16/B gnd XOR2X1_16/Y vdd XOR2X1
XFILL_4_1_2 gnd vdd FILL
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XFILL_12_0_2 gnd vdd FILL
XNAND3X1_6 INVX1_60/A NAND3X1_6/B NAND3X1_6/C gnd NAND3X1_6/Y vdd NAND3X1
XOAI21X1_135 INVX1_93/A OAI21X1_135/B INVX1_91/Y gnd NAND3X1_8/C vdd OAI21X1
XOAI21X1_124 INVX1_86/Y NAND2X1_92/Y OAI21X1_124/C gnd NAND2X1_97/B vdd OAI21X1
XOAI21X1_113 INVX4_3/A INVX1_80/Y OAI21X1_112/Y gnd XOR2X1_10/A vdd OAI21X1
XOAI21X1_102 INVX1_66/A INVX1_70/A BUFX4_13/Y gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_146 INVX1_102/Y INVX1_101/Y AOI22X1_15/D gnd OAI21X1_146/Y vdd OAI21X1
XOAI21X1_179 BUFX2_5/Y OAI21X1_177/Y OAI21X1_178/Y gnd XNOR2X1_60/A vdd OAI21X1
XOAI21X1_168 BUFX4_11/Y AOI21X1_32/Y OAI21X1_168/C gnd XNOR2X1_57/A vdd OAI21X1
XOAI21X1_157 OR2X2_10/B AND2X2_7/Y NOR2X1_78/Y gnd OAI21X1_158/C vdd OAI21X1
XNAND2X1_196 INVX2_6/A INVX1_167/A gnd INVX1_168/A vdd NAND2X1
XNAND2X1_141 BUFX4_17/Y INVX1_125/A gnd OAI21X1_177/C vdd NAND2X1
XNAND2X1_185 XOR2X1_27/Y XNOR2X1_84/B gnd NAND2X1_185/Y vdd NAND2X1
XNAND2X1_163 OAI21X1_206/Y AOI22X1_24/Y gnd XNOR2X1_72/A vdd NAND2X1
XNAND2X1_152 INVX2_21/A INVX4_4/Y gnd INVX2_22/A vdd NAND2X1
XNAND2X1_174 INVX1_143/A INVX2_24/Y gnd INVX1_147/A vdd NAND2X1
XNAND2X1_130 BUFX4_11/Y AOI21X1_33/Y gnd OAI21X1_168/C vdd NAND2X1
XAOI22X1_19 INVX4_8/Y AOI22X1_19/B AOI22X1_19/C AOI21X1_38/Y gnd AOI22X1_19/Y vdd
+ AOI22X1
XXNOR2X1_30 OAI21X1_74/Y INVX1_50/Y gnd XNOR2X1_30/Y vdd XNOR2X1
XFILL_5_3 gnd vdd FILL
XXNOR2X1_41 MUX2X1_5/Y XOR2X1_11/Y gnd XNOR2X1_41/Y vdd XNOR2X1
XBUFX2_40 BUFX2_40/A gnd BUFX2_40/Y vdd BUFX2
XBUFX2_51 BUFX2_55/A gnd BUFX2_51/Y vdd BUFX2
XXNOR2X1_63 BUFX4_18/Y OR2X2_12/B gnd AND2X2_9/B vdd XNOR2X1
XXNOR2X1_85 BUFX4_24/Y INVX1_154/A gnd XNOR2X1_85/Y vdd XNOR2X1
XXNOR2X1_96 XNOR2X1_96/A XNOR2X1_94/Y gnd XNOR2X1_96/Y vdd XNOR2X1
XXNOR2X1_52 MUX2X1_8/Y INVX1_106/Y gnd XNOR2X1_52/Y vdd XNOR2X1
XXNOR2X1_74 INVX2_13/A XOR2X1_23/B gnd XNOR2X1_74/Y vdd XNOR2X1
XAOI21X1_30 BUFX4_8/Y INVX2_16/A NOR2X1_87/Y gnd XNOR2X1_54/A vdd AOI21X1
XAOI21X1_41 NOR2X1_109/B INVX1_127/Y INVX1_130/A gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_52 XOR2X1_26/Y INVX1_152/Y INVX1_158/A gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_63 INVX2_27/Y INVX1_44/A INVX8_2/A gnd AOI21X1_63/Y vdd AOI21X1
XFILL_9_0_2 gnd vdd FILL
XOAI21X1_3 OAI21X1_3/A INVX1_7/Y OAI21X1_1/Y gnd OAI21X1_3/Y vdd OAI21X1
XXNOR2X1_100 XNOR2X1_100/A NOR2X1_91/B gnd DFFPOSX1_61/D vdd XNOR2X1
XFILL_2_2_0 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_6/B gnd XOR2X1_6/Y vdd XOR2X1
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B INVX4_3/A gnd MUX2X1_7/Y vdd MUX2X1
XCLKBUF1_8 clk gnd DFFSR_8/CLK vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_63 OR2X2_9/B CLKBUF1_9/Y DFFPOSX1_63/D gnd vdd DFFPOSX1
XDFFPOSX1_52 BUFX2_58/A CLKBUF1_12/Y INVX2_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 BUFX2_24/A CLKBUF1_7/Y DFFPOSX1_41/D gnd vdd DFFPOSX1
XDFFPOSX1_30 INVX1_4/A CLKBUF1_3/Y XNOR2X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_96 INVX2_23/A CLKBUF1_7/Y OAI21X1_186/Y gnd vdd DFFPOSX1
XBUFX4_19 BUFX4_16/A gnd INVX4_8/A vdd BUFX4
XDFFPOSX1_85 INVX1_125/A CLKBUF1_5/Y XNOR2X1_83/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX2_5/A CLKBUF1_6/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XFILL_15_1 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XBUFX4_4 BUFX4_3/A gnd BUFX4_4/Y vdd BUFX4
XXOR2X1_28 INVX1_78/A BUFX4_25/Y gnd XOR2X1_28/Y vdd XOR2X1
XXOR2X1_17 INVX2_8/A XOR2X1_17/B gnd XOR2X1_17/Y vdd XOR2X1
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 INVX1_76/A NAND3X1_7/B NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_136 AOI21X1_21/Y AOI21X1_22/Y INVX1_92/Y gnd OAI21X1_136/Y vdd OAI21X1
XOAI21X1_125 BUFX4_27/Y AOI22X1_12/D NAND2X1_97/Y gnd XNOR2X1_42/A vdd OAI21X1
XOAI21X1_114 NOR2X1_57/Y AND2X2_5/Y AOI21X1_19/B gnd OAI21X1_115/C vdd OAI21X1
XOAI21X1_103 XOR2X1_8/A INVX1_70/A INVX1_67/A gnd INVX1_72/A vdd OAI21X1
XOAI21X1_169 INVX2_19/Y INVX4_7/Y AOI21X1_33/Y gnd NAND3X1_12/C vdd OAI21X1
XOAI21X1_147 BUFX4_4/Y OAI21X1_147/B OAI21X1_147/C gnd XNOR2X1_48/A vdd OAI21X1
XOAI21X1_158 AND2X2_7/A INVX2_14/Y OAI21X1_158/C gnd AOI21X1_27/C vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd BUFX2_1/Y vdd BUFX2
XNAND2X1_197 BUFX4_7/Y AOI21X1_60/A gnd OAI21X1_263/C vdd NAND2X1
XNAND2X1_142 INVX4_8/Y NOR2X1_98/B gnd NAND2X1_142/Y vdd NAND2X1
XNAND2X1_186 XNOR2X1_85/Y NOR2X1_134/B gnd NAND2X1_186/Y vdd NAND2X1
XNAND2X1_153 INVX2_21/Y INVX1_136/Y gnd NAND2X1_155/B vdd NAND2X1
XNAND2X1_175 NAND3X1_17/Y OAI21X1_232/Y gnd DFFPOSX1_74/D vdd NAND2X1
XNAND2X1_120 INVX1_104/A INVX1_105/A gnd INVX1_108/A vdd NAND2X1
XNAND2X1_164 INVX2_14/A XOR2X1_22/B gnd INVX1_138/A vdd NAND2X1
XNAND2X1_131 INVX2_19/A INVX2_18/Y gnd AOI21X1_36/A vdd NAND2X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 XNOR2X1_8/B AOI21X1_1/B AOI21X1_1/C gnd AOI21X1_1/Y vdd AOI21X1
XXNOR2X1_64 XNOR2X1_64/A AND2X2_9/B gnd XNOR2X1_64/Y vdd XNOR2X1
XXNOR2X1_31 MUX2X1_1/Y INVX1_53/Y gnd XNOR2X1_31/Y vdd XNOR2X1
XXNOR2X1_42 XNOR2X1_42/A INVX1_84/Y gnd XNOR2X1_42/Y vdd XNOR2X1
XXNOR2X1_75 XNOR2X1_75/A AOI21X1_44/C gnd XNOR2X1_75/Y vdd XNOR2X1
XXNOR2X1_53 INVX2_12/A INVX2_25/A gnd INVX1_113/A vdd XNOR2X1
XXNOR2X1_20 XNOR2X1_20/A INVX1_37/A gnd XNOR2X1_20/Y vdd XNOR2X1
XBUFX2_52 BUFX2_55/A gnd BUFX2_52/Y vdd BUFX2
XBUFX2_41 BUFX2_40/A gnd BUFX2_41/Y vdd BUFX2
XXNOR2X1_86 XNOR2X1_86/A INVX1_157/Y gnd XNOR2X1_86/Y vdd XNOR2X1
XXNOR2X1_97 AOI22X1_31/Y XOR2X1_31/Y gnd XNOR2X1_97/Y vdd XNOR2X1
XBUFX2_30 BUFX2_30/A gnd sine[2] vdd BUFX2
XAOI21X1_42 AOI22X1_21/Y INVX1_132/Y INVX1_131/A gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_53 AND2X2_11/B AND2X2_11/A XOR2X1_27/Y gnd AOI22X1_29/D vdd AOI21X1
XAOI21X1_64 XOR2X1_30/Y AND2X2_12/Y INVX1_174/A gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_20 NAND2X1_97/B INVX1_84/A NOR2X1_60/Y gnd MUX2X1_6/B vdd AOI21X1
XAOI21X1_31 AOI21X1_31/A AOI21X1_31/B NOR2X1_90/Y gnd AOI21X1_31/Y vdd AOI21X1
XXNOR2X1_101 XNOR2X1_101/A AOI21X1_67/A gnd DFFPOSX1_62/D vdd XNOR2X1
XOAI21X1_4 NOR2X1_5/Y NOR2X1_6/Y BUFX2_9/Y gnd OAI21X1_6/C vdd OAI21X1
XFILL_3_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_8/A INVX1_68/A gnd XOR2X1_7/Y vdd XOR2X1
XFILL_10_1_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B INVX8_3/A gnd MUX2X1_8/Y vdd MUX2X1
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_18_2_1 gnd vdd FILL
XDFFPOSX1_53 INVX1_183/A CLKBUF1_12/Y NOR2X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 NOR2X1_78/A CLKBUF1_9/Y DFFPOSX1_64/D gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_124/A CLKBUF1_5/Y XNOR2X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 XOR2X1_25/B CLKBUF1_1/Y DFFPOSX1_75/D gnd vdd DFFPOSX1
XDFFPOSX1_42 BUFX2_25/A CLKBUF1_10/Y DFFPOSX1_42/D gnd vdd DFFPOSX1
XDFFPOSX1_20 INVX1_8/A CLKBUF1_11/Y BUFX2_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_6/A CLKBUF1_3/Y XNOR2X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_97 XOR2X1_21/B CLKBUF1_7/Y OAI21X1_195/Y gnd vdd DFFPOSX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XXOR2X1_18 BUFX4_17/Y OAI22X1_9/D gnd XOR2X1_18/Y vdd XOR2X1
XBUFX4_5 BUFX2_1/A gnd BUFX4_5/Y vdd BUFX4
XXOR2X1_29 INVX1_54/A XOR2X1_29/B gnd XOR2X1_29/Y vdd XOR2X1
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XNAND3X1_8 INVX1_92/A NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_137 BUFX2_55/A INVX1_94/Y INVX2_3/A gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_126 INVX1_84/A AOI22X1_11/Y NAND2X1_99/Y gnd MUX2X1_6/A vdd OAI21X1
XOAI21X1_115 INVX1_81/Y OR2X2_8/B OAI21X1_115/C gnd AOI22X1_11/C vdd OAI21X1
XOAI21X1_104 INVX1_72/A AOI22X1_9/Y OAI21X1_102/Y gnd MUX2X1_4/B vdd OAI21X1
XOAI21X1_159 INVX2_13/A AND2X2_10/A INVX2_12/Y gnd OAI21X1_160/C vdd OAI21X1
XOAI21X1_148 OR2X2_10/B AND2X2_7/Y XNOR2X1_47/B gnd OAI21X1_148/Y vdd OAI21X1
XNAND2X1_121 OR2X2_9/Y OAI21X1_152/Y gnd OAI21X1_153/B vdd NAND2X1
XNAND2X1_110 NOR2X1_78/A INVX1_102/Y gnd NAND2X1_110/Y vdd NAND2X1
XBUFX2_2 INVX4_2/Y gnd BUFX2_2/Y vdd BUFX2
XNAND2X1_143 OAI21X1_177/C NAND2X1_142/Y gnd NOR2X1_110/B vdd NAND2X1
XNAND2X1_132 INVX2_18/A INVX2_19/Y gnd AOI21X1_35/B vdd NAND2X1
XNAND2X1_187 BUFX2_8/Y AOI22X1_28/C gnd OAI21X1_243/C vdd NAND2X1
XNAND2X1_176 INVX2_9/A XOR2X1_25/B gnd INVX1_152/A vdd NAND2X1
XNAND2X1_198 INVX1_52/A AND2X2_12/B gnd AOI21X1_59/B vdd NAND2X1
XNAND2X1_154 INVX2_21/A OR2X2_13/A gnd OAI21X1_201/A vdd NAND2X1
XNAND2X1_165 BUFX4_2/Y INVX1_145/A gnd OAI21X1_211/C vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 INVX1_20/Y INVX1_21/Y INVX8_2/A gnd AOI21X1_2/Y vdd AOI21X1
XXNOR2X1_54 XNOR2X1_54/A INVX2_17/Y gnd XNOR2X1_54/Y vdd XNOR2X1
XXNOR2X1_65 BUFX4_16/Y OAI22X1_9/D gnd XNOR2X1_65/Y vdd XNOR2X1
XXNOR2X1_87 INVX2_10/A XOR2X1_26/B gnd XNOR2X1_87/Y vdd XNOR2X1
XXNOR2X1_43 MUX2X1_7/Y INVX1_87/Y gnd XNOR2X1_43/Y vdd XNOR2X1
XXNOR2X1_32 INVX2_5/A INVX2_27/A gnd INVX1_60/A vdd XNOR2X1
XXNOR2X1_98 MUX2X1_12/Y INVX1_176/Y gnd XNOR2X1_98/Y vdd XNOR2X1
XXNOR2X1_10 XNOR2X1_10/A INVX1_21/A gnd XNOR2X1_10/Y vdd XNOR2X1
XXNOR2X1_76 XNOR2X1_76/A AOI21X1_47/A gnd XNOR2X1_76/Y vdd XNOR2X1
XXNOR2X1_21 XNOR2X1_21/A DFFSR_4/Q gnd XNOR2X1_21/Y vdd XNOR2X1
XBUFX2_53 BUFX2_55/A gnd BUFX2_53/Y vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd sine[3] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd cosine[1] vdd BUFX2
XBUFX2_42 INVX4_1/Y gnd BUFX2_42/Y vdd BUFX2
XAOI21X1_21 MUX2X1_7/B INVX1_87/Y INVX1_89/A gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_54 AOI22X1_28/C INVX1_157/A AOI21X1_54/C gnd MUX2X1_11/B vdd AOI21X1
XAOI21X1_65 MUX2X1_12/B INVX1_176/Y INVX1_179/A gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_10 INVX1_48/A INVX2_4/A OR2X2_6/A gnd AOI22X1_4/C vdd AOI21X1
XOAI21X1_5 INVX1_9/Y INVX1_8/Y INVX4_3/A gnd OAI21X1_6/B vdd OAI21X1
XAOI21X1_43 XOR2X1_23/Y INVX1_138/Y INVX1_140/A gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_32 AOI21X1_32/A OR2X2_11/Y NOR2X1_93/Y gnd AOI21X1_32/Y vdd AOI21X1
XXNOR2X1_102 XNOR2X1_102/A NOR2X1_155/A gnd DFFPOSX1_63/D vdd XNOR2X1
XFILL_3_2 gnd vdd FILL
XFILL_2_2_2 gnd vdd FILL
XXOR2X1_8 XOR2X1_8/A INVX1_65/A gnd XOR2X1_8/Y vdd XOR2X1
XFILL_10_1_2 gnd vdd FILL
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B BUFX4_11/Y gnd MUX2X1_9/Y vdd MUX2X1
XFILL_18_2_2 gnd vdd FILL
XDFFPOSX1_54 INVX2_16/A CLKBUF1_9/Y INVX1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 OR2X2_12/A CLKBUF1_5/Y XNOR2X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 XOR2X1_26/B CLKBUF1_1/Y XNOR2X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX2_2/A CLKBUF1_7/Y NAND2X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 INVX1_9/A CLKBUF1_13/Y INVX1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_5/A CLKBUF1_3/Y XNOR2X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 INVX8_3/A CLKBUF1_11/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 BUFX2_26/A DFFSR_2/CLK DFFPOSX1_43/D gnd vdd DFFPOSX1
XDFFPOSX1_65 AND2X2_7/A CLKBUF1_9/Y DFFPOSX1_65/D gnd vdd DFFPOSX1
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XFILL_7_1_2 gnd vdd FILL
XFILL_15_0_2 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XBUFX4_6 BUFX2_1/A gnd BUFX4_6/Y vdd BUFX4
XXOR2X1_19 BUFX4_18/Y INVX1_125/A gnd XOR2X1_19/Y vdd XOR2X1
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XNAND3X1_9 BUFX4_3/Y NAND3X1_9/B NAND3X1_9/C gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_138 INVX2_11/Y INVX1_94/A OAI21X1_137/Y gnd BUFX2_47/A vdd OAI21X1
XOAI21X1_127 INVX1_83/A INVX2_9/A INVX4_6/A gnd OAI21X1_127/Y vdd OAI21X1
XBUFX2_3 INVX4_2/Y gnd BUFX2_3/Y vdd BUFX2
XOAI21X1_105 INVX4_5/Y INVX2_8/Y BUFX2_3/Y gnd INVX1_73/A vdd OAI21X1
XOAI21X1_116 INVX1_80/A NOR2X1_57/Y NAND2X1_89/A gnd NAND2X1_92/A vdd OAI21X1
XOAI21X1_149 OAI21X1_148/Y AOI21X1_23/Y AOI21X1_24/Y gnd AOI21X1_26/A vdd OAI21X1
XNAND2X1_111 NAND2X1_111/A NAND2X1_110/Y gnd NOR2X1_86/B vdd NAND2X1
XNAND2X1_100 INVX1_83/Y INVX2_9/Y gnd AOI22X1_12/B vdd NAND2X1
XNAND2X1_144 XOR2X1_19/Y XNOR2X1_60/B gnd OAI21X1_181/A vdd NAND2X1
XNAND2X1_177 INVX4_3/A AOI21X1_52/Y gnd NAND2X1_177/Y vdd NAND2X1
XNAND2X1_155 OAI21X1_201/A NAND2X1_155/B gnd XOR2X1_20/B vdd NAND2X1
XNAND2X1_166 INVX2_15/A INVX1_97/Y gnd AOI21X1_49/B vdd NAND2X1
XNAND2X1_122 NAND2X1_122/A NAND3X1_10/Y gnd MUX2X1_8/B vdd NAND2X1
XNAND2X1_133 AOI21X1_36/A AOI21X1_35/B gnd XOR2X1_16/B vdd NAND2X1
XNAND2X1_188 INVX1_155/Y INVX1_154/Y gnd AOI22X1_29/B vdd NAND2X1
XNAND2X1_199 INVX1_52/Y INVX1_171/Y gnd AOI21X1_59/A vdd NAND2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XAOI21X1_3 INVX4_4/Y OR2X2_3/A INVX2_2/Y gnd AOI21X1_3/Y vdd AOI21X1
XXNOR2X1_99 XNOR2X1_99/A INVX1_183/Y gnd XNOR2X1_99/Y vdd XNOR2X1
XXNOR2X1_55 AOI21X1_31/Y XNOR2X1_55/B gnd XNOR2X1_55/Y vdd XNOR2X1
XXNOR2X1_22 OAI21X1_56/Y DFFSR_5/Q gnd XNOR2X1_22/Y vdd XNOR2X1
XXNOR2X1_66 XNOR2X1_66/A INVX1_127/A gnd XNOR2X1_66/Y vdd XNOR2X1
XXNOR2X1_44 INVX4_6/A BUFX4_24/Y gnd INVX1_92/A vdd XNOR2X1
XXNOR2X1_88 MUX2X1_11/Y XOR2X1_28/Y gnd XNOR2X1_88/Y vdd XNOR2X1
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XXNOR2X1_33 XOR2X1_8/A INVX1_65/A gnd NOR2X1_56/A vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd BUFX2_10/Y vdd BUFX2
XXNOR2X1_11 XNOR2X1_11/A DFFPOSX1_8/Q gnd XNOR2X1_11/Y vdd XNOR2X1
XXNOR2X1_77 OR2X2_9/B INVX2_25/A gnd INVX1_143/A vdd XNOR2X1
XBUFX2_32 BUFX2_32/A gnd sine[4] vdd BUFX2
XBUFX2_43 BUFX2_40/A gnd BUFX2_43/Y vdd BUFX2
XBUFX2_54 INVX1_94/A gnd BUFX2_54/Y vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd cosine[2] vdd BUFX2
XNOR2X1_1 INVX1_1/Y INVX1_2/Y gnd NOR2X1_1/Y vdd NOR2X1
XAOI21X1_55 AOI21X1_55/A INVX1_160/Y INVX1_163/A gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_22 MUX2X1_7/A INVX1_93/Y INVX1_91/A gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_11 AOI22X1_5/D INVX1_51/A NOR2X1_36/Y gnd OAI21X1_74/B vdd AOI21X1
XAOI21X1_66 MUX2X1_12/A INVX1_182/Y INVX1_181/A gnd AOI21X1_66/Y vdd AOI21X1
XOAI21X1_6 NOR2X1_5/Y OAI21X1_6/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_44 AOI21X1_44/A OAI22X1_10/Y AOI21X1_44/C gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_33 NOR2X1_94/Y AOI21X1_33/B OR2X2_11/A gnd AOI21X1_33/Y vdd AOI21X1
XXNOR2X1_103 XNOR2X1_103/A AOI21X1_68/A gnd DFFPOSX1_64/D vdd XNOR2X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XFILL_3_3 gnd vdd FILL
XXOR2X1_9 MUX2X1_3/Y XOR2X1_9/B gnd XOR2X1_9/Y vdd XOR2X1
XDFFPOSX1_11 BUFX2_11/A CLKBUF1_10/Y BUFX2_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX2_17/A CLKBUF1_9/Y INVX1_186/A gnd vdd DFFPOSX1
XDFFPOSX1_77 XOR2X1_27/B CLKBUF1_1/Y XNOR2X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 OR2X2_12/B CLKBUF1_5/Y XNOR2X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 NOR2X1_7/A CLKBUF1_13/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 OAI21X1_3/A CLKBUF1_10/Y NAND2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 DFFPOSX1_99/Q DFFSR_2/CLK NAND2X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 BUFX2_28/A DFFSR_6/CLK DFFPOSX1_44/D gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX2_12/A CLKBUF1_9/Y XOR2X1_34/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XINVX1_171 AND2X2_12/B gnd INVX1_171/Y vdd INVX1
XFILL_20_2 gnd vdd FILL
XBUFX4_7 BUFX2_1/A gnd BUFX4_7/Y vdd BUFX4
XFILL_13_1 gnd vdd FILL
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XOAI21X1_128 INVX4_6/A INVX2_9/A INVX1_84/A gnd INVX1_88/A vdd OAI21X1
XOAI21X1_117 BUFX4_27/Y AOI22X1_11/C NAND2X1_91/Y gnd XNOR2X1_40/A vdd OAI21X1
XOAI21X1_106 INVX1_71/A AOI22X1_10/Y INVX1_73/Y gnd NAND3X1_7/B vdd OAI21X1
XOAI21X1_139 INVX1_98/A INVX1_97/Y INVX8_3/A gnd OAI21X1_140/C vdd OAI21X1
XBUFX2_4 INVX4_2/Y gnd BUFX2_4/Y vdd BUFX2
XNAND2X1_112 OAI21X1_143/Y NOR2X1_86/B gnd AOI22X1_15/D vdd NAND2X1
XNAND2X1_101 NAND3X1_8/Y OAI21X1_136/Y gnd NAND2X1_101/Y vdd NAND2X1
XNAND2X1_145 XNOR2X1_61/Y NOR2X1_110/B gnd OAI21X1_183/B vdd NAND2X1
XNAND2X1_178 XOR2X1_26/B INVX2_10/Y gnd AND2X2_11/B vdd NAND2X1
XNAND2X1_189 BUFX2_6/Y INVX1_156/A gnd NAND2X1_189/Y vdd NAND2X1
XNAND2X1_156 INVX1_134/A INVX1_135/A gnd NOR2X1_115/A vdd NAND2X1
XNAND2X1_123 NAND3X1_11/Y NAND2X1_123/B gnd NAND2X1_123/Y vdd NAND2X1
XNAND2X1_167 INVX1_97/A INVX2_15/Y gnd INVX1_146/A vdd NAND2X1
XNAND2X1_134 AOI21X1_36/Y NAND3X1_12/Y gnd OAI21X1_173/C vdd NAND2X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XAOI21X1_4 NAND3X1_2/C NOR2X1_22/Y INVX1_29/Y gnd AOI21X1_4/Y vdd AOI21X1
XXNOR2X1_12 OAI21X1_36/Y OR2X2_3/B gnd XNOR2X1_12/Y vdd XNOR2X1
XXNOR2X1_23 OAI21X1_58/Y DFFSR_6/Q gnd XNOR2X1_23/Y vdd XNOR2X1
XBUFX2_44 vdd gnd BUFX2_44/Y vdd BUFX2
XXNOR2X1_45 INVX1_95/A INVX2_3/Y gnd INVX1_96/A vdd XNOR2X1
XXNOR2X1_89 XNOR2X1_89/A INVX1_160/A gnd XNOR2X1_89/Y vdd XNOR2X1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XBUFX2_22 BUFX2_22/A gnd cosine[3] vdd BUFX2
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XXNOR2X1_34 OAI21X1_92/Y NOR2X1_56/A gnd XNOR2X1_34/Y vdd XNOR2X1
XBUFX2_11 BUFX2_11/A gnd BUFX2_11/Y vdd BUFX2
XXNOR2X1_67 XNOR2X1_67/A INVX1_135/Y gnd XNOR2X1_67/Y vdd XNOR2X1
XXNOR2X1_78 INVX1_97/A INVX2_15/A gnd NOR2X1_122/A vdd XNOR2X1
XBUFX2_33 BUFX2_33/A gnd sine[5] vdd BUFX2
XXNOR2X1_56 XNOR2X1_56/A OR2X2_11/Y gnd XNOR2X1_56/Y vdd XNOR2X1
XBUFX2_55 BUFX2_55/A gnd BUFX2_55/Y vdd BUFX2
XNOR2X1_2 INVX1_1/A INVX1_2/A gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_23 XOR2X1_14/B AOI21X1_23/B NOR2X1_77/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_12 NOR2X1_42/Y OAI21X1_65/Y OAI21X1_81/Y gnd OAI21X1_83/B vdd AOI21X1
XAOI21X1_34 AOI21X1_32/Y INVX1_120/Y NOR2X1_95/Y gnd MUX2X1_9/B vdd AOI21X1
XAOI21X1_67 AOI21X1_67/A AOI21X1_67/B NOR2X1_152/Y gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_56 AOI21X1_56/A INVX1_165/Y INVX1_164/A gnd AOI21X1_56/Y vdd AOI21X1
XOAI21X1_7 INVX4_3/A NOR2X1_5/Y OAI21X1_6/B gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B AOI21X1_45/C gnd AOI21X1_45/Y vdd AOI21X1
XFILL_5_2_1 gnd vdd FILL
XXNOR2X1_104 MUX2X1_13/Y XOR2X1_33/Y gnd DFFPOSX1_65/D vdd XNOR2X1
XFILL_13_1_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_23 INVX2_1/A CLKBUF1_3/Y XNOR2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX4_2/A CLKBUF1_3/Y NAND2X1_11/B gnd vdd DFFPOSX1
XDFFPOSX1_12 BUFX2_12/A CLKBUF1_11/Y BUFX2_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_45 BUFX2_29/A DFFSR_2/CLK DFFPOSX1_45/D gnd vdd DFFPOSX1
XDFFPOSX1_56 INVX1_116/A CLKBUF1_9/Y INVX1_95/A gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX2_7/A CLKBUF1_5/Y OAI21X1_252/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 INVX1_154/A CLKBUF1_1/Y XNOR2X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_167/A CLKBUF1_6/Y XOR2X1_22/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_161 XOR2X1_28/Y gnd INVX1_161/Y vdd INVX1
XINVX1_172 XOR2X1_30/B gnd INVX1_172/Y vdd INVX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XFILL_20_3 gnd vdd FILL
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XOAI21X1_129 INVX1_88/A AOI22X1_13/Y OAI21X1_127/Y gnd MUX2X1_7/B vdd OAI21X1
XOAI21X1_118 INVX1_82/Y INVX4_6/A AOI21X1_19/Y gnd OAI21X1_118/Y vdd OAI21X1
XOAI21X1_107 INVX1_66/A INVX1_70/A INVX4_5/Y gnd OAI21X1_107/Y vdd OAI21X1
XBUFX2_5 INVX4_2/Y gnd BUFX2_5/Y vdd BUFX2
XNAND2X1_102 INVX1_98/A INVX1_97/Y gnd NAND2X1_104/A vdd NAND2X1
XNAND2X1_135 INVX2_8/A XOR2X1_17/B gnd INVX1_122/A vdd NAND2X1
XNAND2X1_146 BUFX2_2/Y AOI22X1_18/C gnd NAND2X1_146/Y vdd NAND2X1
XNAND2X1_179 INVX1_154/A INVX2_26/Y gnd NAND2X1_181/A vdd NAND2X1
XNAND2X1_157 INVX1_134/Y INVX1_135/Y gnd NOR2X1_116/B vdd NAND2X1
XNAND2X1_168 AOI21X1_49/B INVX1_146/A gnd AOI21X1_47/A vdd NAND2X1
XNAND2X1_113 BUFX4_4/Y OAI21X1_146/Y gnd OAI21X1_147/C vdd NAND2X1
XNAND2X1_124 OAI22X1_8/A INVX1_117/Y gnd NAND2X1_124/Y vdd NAND2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XAOI21X1_5 AOI21X1_5/A AOI21X1_5/B OAI22X1_5/Y gnd XOR2X1_3/A vdd AOI21X1
XXNOR2X1_35 MUX2X1_2/Y XOR2X1_7/Y gnd XNOR2X1_35/Y vdd XNOR2X1
XXNOR2X1_13 NAND2X1_29/Y NOR2X1_21/A gnd XNOR2X1_13/Y vdd XNOR2X1
XXNOR2X1_24 XNOR2X1_24/A INVX1_41/Y gnd XNOR2X1_24/Y vdd XNOR2X1
XXNOR2X1_57 XNOR2X1_57/A XOR2X1_34/B gnd XNOR2X1_57/Y vdd XNOR2X1
XXNOR2X1_46 INVX1_102/A NOR2X1_78/A gnd XNOR2X1_47/B vdd XNOR2X1
XBUFX2_56 vdd gnd BUFX2_56/Y vdd BUFX2
XBUFX2_45 BUFX2_18/Y gnd BUFX2_45/Y vdd BUFX2
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XXNOR2X1_68 XNOR2X1_68/A OR2X2_13/B gnd XNOR2X1_68/Y vdd XNOR2X1
XINVX1_81 OR2X2_8/A gnd INVX1_81/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XBUFX2_23 BUFX2_23/A gnd cosine[4] vdd BUFX2
XBUFX2_34 BUFX2_34/A gnd sine[6] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd BUFX2_12/Y vdd BUFX2
XXNOR2X1_79 XNOR2X1_79/A INVX1_143/A gnd XNOR2X1_79/Y vdd XNOR2X1
XNOR2X1_3 INVX1_4/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_68 AOI21X1_68/A NOR2X1_153/Y AOI21X1_68/C gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_57 XOR2X1_29/Y INVX1_168/Y INVX1_170/A gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_13 MUX2X1_1/B INVX1_53/Y INVX1_58/A gnd OAI21X1_86/A vdd AOI21X1
XAOI21X1_46 INVX2_25/Y OR2X2_9/B INVX8_3/A gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_35 INVX1_121/Y AOI21X1_35/B AOI21X1_35/C gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_24 OR2X2_10/Y NOR2X1_78/Y NOR2X1_79/Y gnd AOI21X1_24/Y vdd AOI21X1
XOAI21X1_8 BUFX2_9/Y OAI21X1_9/B NAND2X1_6/Y gnd OAI21X1_8/Y vdd OAI21X1
XFILL_5_2_2 gnd vdd FILL
XFILL_13_1_2 gnd vdd FILL
XOAI22X1_10 XOR2X1_22/B INVX2_14/Y INVX2_13/Y XOR2X1_23/B gnd OAI22X1_10/Y vdd OAI22X1
XOAI21X1_290 BUFX4_9/Y OAI21X1_288/Y OAI21X1_290/C gnd XNOR2X1_102/A vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XDFFPOSX1_57 INVX1_118/A CLKBUF1_12/Y INVX1_186/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 INVX1_11/A CLKBUF1_3/Y XNOR2X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 XOR2X1_29/B CLKBUF1_6/Y XNOR2X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 INVX4_4/A CLKBUF1_10/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 INVX1_17/A CLKBUF1_11/Y BUFX2_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_46 BUFX2_30/A DFFSR_2/CLK DFFPOSX1_46/D gnd vdd DFFPOSX1
XDFFPOSX1_79 INVX1_156/A CLKBUF1_1/Y XNOR2X1_96/Y gnd vdd DFFPOSX1
XFILL_2_0_2 gnd vdd FILL
XFILL_18_0_2 gnd vdd FILL
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XFILL_20_2_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XBUFX4_9 BUFX4_8/A gnd BUFX4_9/Y vdd BUFX4
XNOR2X1_90 INVX2_16/A INVX2_17/A gnd NOR2X1_90/Y vdd NOR2X1
XOAI21X1_119 INVX1_82/A INVX4_6/Y OAI21X1_118/Y gnd MUX2X1_5/A vdd OAI21X1
XOAI21X1_108 AOI22X1_7/Y INVX1_74/Y OAI21X1_107/Y gnd OAI21X1_110/B vdd OAI21X1
XNAND2X1_125 INVX1_116/A BUFX2_58/A gnd NAND2X1_125/Y vdd NAND2X1
XNAND2X1_103 INVX1_97/A INVX1_98/Y gnd AOI21X1_23/B vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd BUFX2_6/Y vdd BUFX2
XNAND2X1_114 INVX2_12/Y INVX2_13/Y gnd NAND2X1_116/B vdd NAND2X1
XNAND2X1_136 INVX4_2/A AOI21X1_37/Y gnd NAND2X1_136/Y vdd NAND2X1
XNAND2X1_147 NOR2X1_98/B INVX1_124/Y gnd AOI22X1_19/B vdd NAND2X1
XNAND2X1_158 INVX2_21/A INVX1_136/Y gnd NAND2X1_158/Y vdd NAND2X1
XNAND2X1_1 INVX1_3/A NOR2X1_1/Y gnd NOR2X1_4/B vdd NAND2X1
XNAND2X1_169 AND2X2_10/A AND2X2_10/B gnd OAI21X1_217/A vdd NAND2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 INVX1_33/Y INVX2_3/A INVX1_34/A gnd AOI22X1_2/D vdd AOI21X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XXNOR2X1_58 XNOR2X1_58/A XOR2X1_18/Y gnd XNOR2X1_58/Y vdd XNOR2X1
XXNOR2X1_25 INVX1_48/A INVX2_4/A gnd OAI21X1_71/C vdd XNOR2X1
XFILL_8_2_0 gnd vdd FILL
XXNOR2X1_69 XNOR2X1_69/A NOR2X1_114/Y gnd XNOR2X1_69/Y vdd XNOR2X1
XXNOR2X1_36 XNOR2X1_36/A INVX1_67/Y gnd XNOR2X1_36/Y vdd XNOR2X1
XXNOR2X1_14 NAND2X1_31/Y NOR2X1_22/B gnd XNOR2X1_14/Y vdd XNOR2X1
XXNOR2X1_47 XNOR2X1_47/A XNOR2X1_47/B gnd XNOR2X1_47/Y vdd XNOR2X1
XBUFX2_57 BUFX2_57/A gnd BUFX2_57/Y vdd BUFX2
XBUFX2_46 INVX2_11/Y gnd BUFX2_46/Y vdd BUFX2
XBUFX2_24 BUFX2_24/A gnd cosine[5] vdd BUFX2
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XBUFX2_13 BUFX2_13/A gnd BUFX2_13/Y vdd BUFX2
XBUFX2_35 BUFX2_35/A gnd sine[7] vdd BUFX2
XDFFPOSX1_1 XNOR2X1_8/B CLKBUF1_11/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_16_1_0 gnd vdd FILL
XNOR2X1_4 INVX1_4/Y NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_58 XNOR2X1_91/Y AOI21X1_58/B NOR2X1_143/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_14 MUX2X1_1/A INVX1_61/Y INVX1_59/A gnd OAI21X1_86/B vdd AOI21X1
XAOI21X1_47 AOI21X1_47/A OR2X2_14/A INVX1_142/A gnd AOI21X1_47/Y vdd AOI21X1
XAOI21X1_36 AOI21X1_36/A INVX4_7/Y INVX8_1/A gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_25 INVX1_102/A NOR2X1_78/A AND2X2_7/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_69 AOI21X1_69/A NOR2X1_155/Y AOI21X1_69/C gnd MUX2X1_13/A vdd AOI21X1
XOAI21X1_9 INVX2_1/Y OAI21X1_9/B INVX4_3/A gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_11 XOR2X1_25/B INVX2_9/Y INVX2_10/Y XOR2X1_26/B gnd AND2X2_11/A vdd OAI22X1
XFILL_5_0_0 gnd vdd FILL
XOAI21X1_291 INVX2_17/Y INVX2_18/Y OAI21X1_291/C gnd OAI21X1_294/B vdd OAI21X1
XOAI21X1_280 INVX2_4/A INVX2_27/A INVX8_2/A gnd INVX1_181/A vdd OAI21X1
XDFFPOSX1_25 OAI21X1_13/C CLKBUF1_3/Y NAND2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 AND2X2_12/B CLKBUF1_6/Y XNOR2X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_18/A CLKBUF1_13/Y INVX1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 BUFX2_31/A CLKBUF1_10/Y DFFPOSX1_47/D gnd vdd DFFPOSX1
XDFFPOSX1_36 BUFX2_19/A DFFSR_2/CLK DFFPOSX1_99/Q gnd vdd DFFPOSX1
XDFFPOSX1_58 INVX2_19/A CLKBUF1_11/Y gnd gnd vdd DFFPOSX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_141 AND2X2_10/B gnd INVX1_141/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XFILL_20_2_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XNOR2X1_91 INVX1_118/A NOR2X1_91/B gnd OR2X2_11/B vdd NOR2X1
XNOR2X1_80 INVX2_12/A INVX2_13/Y gnd NOR2X1_80/Y vdd NOR2X1
XBUFX2_7 INVX4_3/Y gnd BUFX2_7/Y vdd BUFX2
XOAI21X1_109 INVX2_8/A INVX4_5/Y INVX4_2/A gnd INVX1_75/A vdd OAI21X1
XNAND2X1_126 NAND2X1_125/Y NAND2X1_124/Y gnd XNOR2X1_55/B vdd NAND2X1
XNAND2X1_104 NAND2X1_104/A AOI21X1_23/B gnd NAND2X1_104/Y vdd NAND2X1
XNAND2X1_137 OAI22X1_9/D INVX4_8/Y gnd AND2X2_8/B vdd NAND2X1
XNAND2X1_148 NAND3X1_13/Y OAI21X1_200/Y gnd NAND2X1_148/Y vdd NAND2X1
XNAND2X1_159 OAI21X1_201/Y NAND2X1_159/B gnd XNOR2X1_68/A vdd NAND2X1
XNAND2X1_115 INVX2_12/A INVX2_13/A gnd NAND3X1_9/B vdd NAND2X1
XNAND2X1_2 INVX1_3/Y NOR2X1_2/Y gnd NOR2X1_3/B vdd NAND2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_7 AOI21X1_7/A DFFSR_4/Q DFFSR_5/Q gnd AOI21X1_7/Y vdd AOI21X1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XXNOR2X1_59 XNOR2X1_59/A XOR2X1_19/Y gnd XNOR2X1_59/Y vdd XNOR2X1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XXNOR2X1_26 OAI21X1_67/Y OAI21X1_71/C gnd XNOR2X1_26/Y vdd XNOR2X1
XFILL_8_2_1 gnd vdd FILL
XXNOR2X1_37 MUX2X1_4/Y INVX1_71/Y gnd XNOR2X1_37/Y vdd XNOR2X1
XXNOR2X1_15 INVX2_2/A INVX1_30/A gnd XNOR2X1_15/Y vdd XNOR2X1
XXNOR2X1_48 XNOR2X1_48/A OR2X2_10/Y gnd XNOR2X1_48/Y vdd XNOR2X1
XBUFX2_58 BUFX2_58/A gnd BUFX2_58/Y vdd BUFX2
XBUFX2_47 BUFX2_47/A gnd BUFX2_47/Y vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd cosine[6] vdd BUFX2
XBUFX2_14 BUFX2_14/A gnd BUFX2_14/Y vdd BUFX2
XBUFX2_36 gnd gnd BUFX2_36/Y vdd BUFX2
XDFFPOSX1_2 INVX8_1/A CLKBUF1_11/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 INVX1_9/A INVX1_8/A gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_37 XOR2X1_18/Y INVX1_122/Y INVX1_129/A gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_59 AOI21X1_59/A AOI21X1_59/B XOR2X1_30/Y gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_15 XOR2X1_6/B OAI21X1_89/C NOR2X1_44/Y gnd OAI21X1_97/B vdd AOI21X1
XAOI21X1_48 AOI21X1_48/A INVX1_143/Y AOI21X1_48/C gnd AOI21X1_48/Y vdd AOI21X1
XAOI21X1_26 AOI21X1_26/A INVX1_105/A NOR2X1_80/Y gnd AOI21X1_26/Y vdd AOI21X1
XOAI22X1_12 OAI22X1_12/A AOI21X1_70/Y OAI22X1_12/C NOR2X1_156/Y gnd XOR2X1_34/A vdd
+ OAI22X1
XFILL_5_0_1 gnd vdd FILL
XOAI21X1_292 INVX2_17/A INVX2_18/Y AOI21X1_69/A gnd OAI21X1_293/C vdd OAI21X1
XOAI21X1_281 INVX1_182/A OAI21X1_281/B INVX1_181/Y gnd NAND3X1_19/C vdd OAI21X1
XOAI21X1_270 NOR2X1_140/Y AND2X2_12/Y XNOR2X1_95/Y gnd OAI21X1_271/A vdd OAI21X1
XDFFPOSX1_48 BUFX2_32/A DFFSR_6/CLK DFFPOSX1_48/D gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX4_3/A CLKBUF1_13/Y NAND2X1_21/B gnd vdd DFFPOSX1
XDFFPOSX1_15 INVX1_19/A CLKBUF1_13/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 BUFX2_20/A CLKBUF1_10/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XDFFPOSX1_59 XOR2X1_22/B CLKBUF1_9/Y XOR2X1_32/Y gnd vdd DFFPOSX1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_153 XOR2X1_26/B gnd INVX1_153/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_120 NOR2X1_96/Y gnd INVX1_120/Y vdd INVX1
XFILL_20_2_2 gnd vdd FILL
XFILL_11_2_2 gnd vdd FILL
XNOR2X1_92 INVX1_118/Y INVX1_119/Y gnd OR2X2_11/A vdd NOR2X1
XNOR2X1_70 NOR2X1_70/A NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_81 INVX2_15/A INVX2_12/Y gnd NOR2X1_83/A vdd NOR2X1
XBUFX2_8 INVX4_3/Y gnd BUFX2_8/Y vdd BUFX2
XNAND2X1_105 OR2X2_9/A OR2X2_9/B gnd NAND2X1_106/A vdd NAND2X1
XNAND2X1_138 INVX1_124/A INVX4_8/Y gnd NAND2X1_140/A vdd NAND2X1
XNAND2X1_149 INVX1_134/A INVX2_21/Y gnd NAND2X1_149/Y vdd NAND2X1
XNAND2X1_3 INVX1_6/Y NOR2X1_3/Y gnd OAI21X1_2/B vdd NAND2X1
XNAND2X1_116 NAND3X1_9/B NAND2X1_116/B gnd INVX1_105/A vdd NAND2X1
XNAND2X1_127 BUFX2_57/A BUFX4_8/Y gnd AOI21X1_31/A vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XAOI21X1_8 XOR2X1_5/B AOI21X1_8/B AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XBUFX2_26 BUFX2_26/A gnd cosine[7] vdd BUFX2
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XXNOR2X1_38 INVX4_5/A BUFX4_16/Y gnd INVX1_76/A vdd XNOR2X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XXNOR2X1_27 OAI21X1_70/Y OR2X2_6/Y gnd XNOR2X1_27/Y vdd XNOR2X1
XFILL_8_2_2 gnd vdd FILL
XXNOR2X1_16 OAI22X1_5/Y XNOR2X1_15/Y gnd XNOR2X1_16/Y vdd XNOR2X1
XBUFX2_15 BUFX2_15/A gnd BUFX2_15/Y vdd BUFX2
XXNOR2X1_49 XNOR2X1_49/A INVX1_105/A gnd XNOR2X1_49/Y vdd XNOR2X1
XBUFX2_48 vdd gnd BUFX2_48/Y vdd BUFX2
XDFFPOSX1_3 BUFX2_13/A DFFSR_8/CLK INVX1_13/Y gnd vdd DFFPOSX1
XBUFX2_37 gnd gnd BUFX2_37/Y vdd BUFX2
XBUFX2_59 INVX4_7/A gnd BUFX2_59/Y vdd BUFX2
XFILL_16_1_2 gnd vdd FILL
XNOR2X1_6 INVX1_9/Y INVX1_8/Y gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 NAND2X1_80/B INVX1_67/A NOR2X1_47/B gnd MUX2X1_3/B vdd AOI21X1
XAOI21X1_27 NOR2X1_86/Y AOI21X1_27/B AOI21X1_27/C gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_38 AND2X2_8/B AND2X2_8/A XOR2X1_19/Y gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_49 AOI21X1_49/A AOI21X1_49/B INVX1_146/Y gnd AOI21X1_49/Y vdd AOI21X1
XOAI21X1_90 INVX1_64/Y BUFX4_13/Y OAI21X1_89/Y gnd AOI22X1_7/C vdd OAI21X1
XFILL_5_0_2 gnd vdd FILL
XOAI21X1_293 INVX2_17/Y INVX2_18/A OAI21X1_293/C gnd NAND2X1_224/B vdd OAI21X1
XOAI21X1_260 INVX1_168/A XNOR2X1_91/Y INVX1_170/Y gnd AOI21X1_61/A vdd OAI21X1
XOAI21X1_282 AOI21X1_65/Y AOI21X1_66/Y INVX1_60/A gnd OAI21X1_282/Y vdd OAI21X1
XOAI21X1_271 OAI21X1_271/A AOI21X1_58/Y AOI21X1_62/Y gnd AOI22X1_33/D vdd OAI21X1
XDFFPOSX1_16 INVX1_21/A CLKBUF1_13/Y XNOR2X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_27 INVX1_2/A CLKBUF1_3/Y BUFX2_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 BUFX2_21/A CLKBUF1_7/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 BUFX2_33/A DFFSR_2/CLK DFFPOSX1_49/D gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_121 MUX2X1_9/B gnd INVX1_121/Y vdd INVX1
XINVX1_110 OR2X2_9/B gnd INVX1_110/Y vdd INVX1
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_71 INVX2_3/A INVX2_11/Y gnd NOR2X1_71/Y vdd NOR2X1
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_60 INVX4_6/Y INVX1_83/Y gnd NOR2X1_60/Y vdd NOR2X1
XNOR2X1_82 INVX2_12/A INVX2_15/Y gnd NOR2X1_82/Y vdd NOR2X1
XNOR2X1_93 INVX1_118/A INVX1_119/Y gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 INVX4_3/Y gnd BUFX2_9/Y vdd BUFX2
XNAND2X1_128 INVX8_1/A NOR2X1_88/A gnd AOI21X1_31/B vdd NAND2X1
XNAND2X1_106 NAND2X1_106/A OR2X2_9/Y gnd XOR2X1_14/B vdd NAND2X1
XNAND2X1_139 BUFX4_16/Y INVX1_124/Y gnd AOI22X1_19/C vdd NAND2X1
XNAND2X1_4 INVX1_6/A NOR2X1_4/Y gnd OAI21X1_1/B vdd NAND2X1
XNAND2X1_117 BUFX4_3/Y AOI22X1_15/Y gnd NAND2X1_117/Y vdd NAND2X1
XNOR2X1_150 XNOR2X1_94/Y INVX1_177/Y gnd INVX1_180/A vdd NOR2X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XAOI21X1_9 OR2X2_6/Y AOI21X1_9/B NOR2X1_35/Y gnd AOI21X1_9/Y vdd AOI21X1
XXNOR2X1_28 XNOR2X1_28/A INVX1_51/A gnd XNOR2X1_28/Y vdd XNOR2X1
XXNOR2X1_39 INVX1_82/A INVX4_6/A gnd NOR2X1_70/A vdd XNOR2X1
XXNOR2X1_17 INVX2_2/A INVX2_21/A gnd XOR2X1_3/B vdd XNOR2X1
XBUFX2_16 DFFSR_8/Q gnd BUFX2_40/A vdd BUFX2
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XBUFX2_38 vdd gnd BUFX2_38/Y vdd BUFX2
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XBUFX2_49 gnd gnd BUFX2_49/Y vdd BUFX2
XINVX1_41 DFFSR_7/Q gnd INVX1_41/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XBUFX2_27 DFFSR_9/Q gnd done vdd BUFX2
XDFFPOSX1_4 BUFX2_14/A CLKBUF1_11/Y OAI22X1_1/Y gnd vdd DFFPOSX1
XNOR2X1_7 NOR2X1_7/A INVX1_10/Y gnd NOR2X1_7/Y vdd NOR2X1
XAOI21X1_39 AOI22X1_18/C INVX2_20/A NOR2X1_99/Y gnd AND2X2_9/A vdd AOI21X1
XAOI21X1_17 MUX2X1_4/B INVX1_71/Y INVX1_73/A gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 MUX2X1_8/B INVX1_106/Y INVX1_111/A gnd AOI21X1_28/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_91 INVX1_63/A NOR2X1_43/Y NAND2X1_71/Y gnd AOI22X1_9/C vdd OAI21X1
XOAI21X1_80 OR2X2_6/B OR2X2_6/A AOI21X1_9/B gnd OAI21X1_81/C vdd OAI21X1
XOAI21X1_250 AOI21X1_54/C NOR2X1_132/Y XOR2X1_28/Y gnd INVX1_166/A vdd OAI21X1
XOAI21X1_294 BUFX4_9/Y OAI21X1_294/B OAI21X1_294/C gnd XNOR2X1_103/A vdd OAI21X1
XOAI21X1_261 INVX1_54/Y XOR2X1_29/B AOI21X1_58/B gnd OAI21X1_261/Y vdd OAI21X1
XOAI21X1_272 XNOR2X1_94/Y AOI21X1_61/Y NAND2X1_205/Y gnd AOI22X1_31/D vdd OAI21X1
XOAI21X1_283 BUFX2_57/A INVX1_117/Y AOI21X1_31/A gnd XNOR2X1_99/A vdd OAI21X1
XDFFPOSX1_39 BUFX2_22/A CLKBUF1_7/Y DFFPOSX1_39/D gnd vdd DFFPOSX1
XDFFPOSX1_17 OAI21X1_27/A CLKBUF1_13/Y NAND2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 INVX1_1/A CLKBUF1_11/Y INVX1_8/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 OR2X2_9/A gnd INVX1_100/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XINVX1_166 INVX1_166/A gnd INVX1_166/Y vdd INVX1
XINVX1_155 XOR2X1_27/B gnd INVX1_155/Y vdd INVX1
XINVX1_177 XOR2X1_31/Y gnd INVX1_177/Y vdd INVX1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_72 BUFX2_55/A INVX1_94/Y gnd NOR2X1_74/A vdd NOR2X1
XNOR2X1_61 NOR2X1_59/Y NOR2X1_60/Y gnd INVX1_84/A vdd NOR2X1
XNOR2X1_50 NOR2X1_48/Y NOR2X1_50/B gnd XOR2X1_9/B vdd NOR2X1
XNOR2X1_83 NOR2X1_83/A NOR2X1_82/Y gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_94 OR2X2_11/B OR2X2_11/A gnd NOR2X1_94/Y vdd NOR2X1
XNAND2X1_107 INVX1_98/A INVX1_97/A gnd INVX1_99/A vdd NAND2X1
XNAND2X1_5 NOR2X1_7/A NOR2X1_6/Y gnd OAI21X1_9/B vdd NAND2X1
XNAND2X1_118 INVX1_105/Y AOI22X1_15/Y gnd NAND3X1_9/C vdd NAND2X1
XNAND2X1_129 BUFX4_8/Y AOI21X1_33/B gnd OAI21X1_167/C vdd NAND2X1
XNOR2X1_151 INVX1_119/Y INVX1_184/A gnd AOI21X1_67/B vdd NOR2X1
XNOR2X1_140 INVX1_52/A AND2X2_12/B gnd NOR2X1_140/Y vdd NOR2X1
XXNOR2X1_29 INVX2_5/A INVX1_54/A gnd INVX1_50/A vdd XNOR2X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XXNOR2X1_18 XNOR2X1_18/A INVX1_36/A gnd XNOR2X1_18/Y vdd XNOR2X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_42 DFFSR_6/Q gnd INVX1_42/Y vdd INVX1
XBUFX2_28 BUFX2_28/A gnd sine[0] vdd BUFX2
XBUFX2_39 BUFX2_40/A gnd BUFX2_39/Y vdd BUFX2
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XINVX1_64 OR2X2_7/A gnd INVX1_64/Y vdd INVX1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XDFFPOSX1_5 BUFX2_15/A CLKBUF1_11/Y XNOR2X1_4/Y gnd vdd DFFPOSX1
XBUFX2_17 DFFSR_1/Q gnd BUFX2_17/Y vdd BUFX2
XNOR2X1_8 INVX1_12/Y INVX1_13/Y gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 MUX2X1_4/A INVX1_77/Y INVX1_75/A gnd AOI21X1_18/Y vdd AOI21X1
XAOI21X1_29 MUX2X1_8/A INVX1_114/Y INVX1_112/A gnd AOI21X1_29/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 INVX1_49/Y INVX2_5/A OAI21X1_81/C gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_70 BUFX4_6/Y OAI21X1_68/Y NAND2X1_57/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 BUFX2_4/Y AOI22X1_7/C NAND2X1_74/Y gnd OAI21X1_92/Y vdd OAI21X1
XOAI21X1_262 INVX1_54/A INVX1_169/Y OAI21X1_261/Y gnd AOI21X1_60/A vdd OAI21X1
XOAI21X1_240 NAND2X1_185/Y AOI21X1_52/Y OAI21X1_240/C gnd AOI22X1_30/D vdd OAI21X1
XOAI21X1_251 INVX1_166/A AOI22X1_27/Y OAI21X1_249/Y gnd XNOR2X1_89/A vdd OAI21X1
XOAI21X1_273 OAI21X1_273/A AOI21X1_57/Y AOI21X1_64/Y gnd AOI22X1_32/D vdd OAI21X1
XOAI21X1_284 BUFX2_57/A INVX1_183/A BUFX2_58/A gnd INVX1_184/A vdd OAI21X1
XOAI21X1_295 NAND2X1_225/Y AOI21X1_67/Y AOI21X1_68/Y gnd MUX2X1_13/B vdd OAI21X1
XDFFPOSX1_29 INVX1_3/A CLKBUF1_3/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 INVX8_2/A CLKBUF1_13/Y OAI22X1_3/Y gnd vdd DFFPOSX1
XFILL_14_2_2 gnd vdd FILL
XINVX1_123 OAI22X1_9/D gnd INVX1_123/Y vdd INVX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_101 NOR2X1_78/A gnd INVX1_101/Y vdd INVX1
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XFILL_20_0_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XFILL_11_0_2 gnd vdd FILL
XNOR2X1_73 INVX1_94/A INVX2_11/Y gnd NOR2X1_73/Y vdd NOR2X1
XFILL_19_1_2 gnd vdd FILL
XNOR2X1_40 INVX1_50/A INVX1_51/A gnd NAND3X1_5/B vdd NOR2X1
XNOR2X1_62 INVX4_6/A INVX2_9/A gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_51 XOR2X1_7/Y XOR2X1_8/Y gnd AOI22X1_7/D vdd NOR2X1
XNOR2X1_84 INVX1_104/A INVX1_105/A gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_95 INVX4_7/A INVX2_19/Y gnd NOR2X1_95/Y vdd NOR2X1
XNAND2X1_108 BUFX4_4/Y OAI21X1_143/Y gnd OAI21X1_144/C vdd NAND2X1
XNAND2X1_119 INVX2_13/Y INVX1_107/Y gnd AOI22X1_17/B vdd NAND2X1
XNAND2X1_6 BUFX2_9/Y NOR2X1_7/Y gnd NAND2X1_6/Y vdd NAND2X1
XNOR2X1_152 INVX2_16/Y INVX4_7/Y gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_130 BUFX4_25/Y INVX1_155/Y gnd NOR2X1_130/Y vdd NOR2X1
XNOR2X1_141 NOR2X1_140/Y AND2X2_12/Y gnd NOR2X1_141/Y vdd NOR2X1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 NOR2X1_5/Y gnd INVX1_10/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XXNOR2X1_19 XNOR2X1_19/A INVX1_35/Y gnd XNOR2X1_19/Y vdd XNOR2X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XBUFX2_18 BUFX2_55/A gnd BUFX2_18/Y vdd BUFX2
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XDFFPOSX1_6 INVX1_22/A CLKBUF1_11/Y XNOR2X1_5/Y gnd vdd DFFPOSX1
XBUFX2_29 BUFX2_29/A gnd sine[1] vdd BUFX2
XNOR2X1_9 BUFX4_10/Y NOR2X1_8/Y gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 XOR2X1_10/B AOI21X1_19/B NOR2X1_58/Y gnd AOI21X1_19/Y vdd AOI21X1
XFILL_8_0_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XOAI21X1_82 INVX2_6/A INVX1_54/A INVX2_5/Y gnd OAI21X1_83/C vdd OAI21X1
XOAI21X1_93 BUFX4_13/Y INVX1_65/Y OAI21X1_97/B gnd OAI21X1_94/C vdd OAI21X1
XOAI21X1_71 OR2X2_6/B OR2X2_6/A OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_60 INVX4_1/Y INVX1_43/Y OAI21X1_60/C gnd XNOR2X1_24/A vdd OAI21X1
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_285 BUFX2_57/A BUFX2_58/A INVX1_183/Y gnd OAI21X1_285/Y vdd OAI21X1
XOAI21X1_252 BUFX2_8/Y XNOR2X1_89/Y OAI21X1_248/Y gnd OAI21X1_252/Y vdd OAI21X1
XOAI21X1_263 BUFX4_7/Y AOI21X1_61/A OAI21X1_263/C gnd XNOR2X1_92/A vdd OAI21X1
XOAI21X1_241 XOR2X1_27/B INVX1_154/A INVX2_26/Y gnd OAI21X1_241/Y vdd OAI21X1
XOAI21X1_274 INVX1_44/A OR2X2_5/B INVX2_27/Y gnd OAI21X1_274/Y vdd OAI21X1
XOAI21X1_230 AND2X2_7/A INVX2_25/A INVX8_3/A gnd INVX1_150/A vdd OAI21X1
XOAI21X1_296 OAI21X1_296/A AOI21X1_68/A NAND2X1_220/Y gnd AOI21X1_69/C vdd OAI21X1
XFILL_17_2_0 gnd vdd FILL
XDFFPOSX1_19 BUFX2_10/A CLKBUF1_3/Y BUFX2_11/Y gnd vdd DFFPOSX1
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XFILL_6_1_0 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_30 DFFSR_4/Q INVX1_40/A gnd NOR2X1_30/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_74/A NOR2X1_73/Y gnd INVX1_95/A vdd NOR2X1
XNOR2X1_63 INVX4_6/Y INVX2_9/Y gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_41 OR2X2_6/B OR2X2_6/A gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_52 INVX2_8/A INVX4_5/Y gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_96 INVX2_19/A INVX4_7/Y gnd NOR2X1_96/Y vdd NOR2X1
XNOR2X1_85 OR2X2_10/B AND2X2_7/Y gnd NOR2X1_85/Y vdd NOR2X1
XNAND2X1_7 INVX2_1/Y NOR2X1_7/Y gnd NAND2X1_7/Y vdd NAND2X1
XNAND2X1_109 INVX1_102/A INVX1_101/Y gnd NAND2X1_111/A vdd NAND2X1
XNOR2X1_142 INVX1_54/Y INVX1_169/Y gnd INVX1_170/A vdd NOR2X1
XNOR2X1_131 BUFX4_26/Y INVX1_156/Y gnd AOI21X1_54/C vdd NOR2X1
XNOR2X1_120 INVX2_13/Y INVX1_139/Y gnd INVX1_140/A vdd NOR2X1
XNOR2X1_153 INVX2_17/Y INVX2_18/Y gnd NOR2X1_153/Y vdd NOR2X1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd cosine[0] vdd BUFX2
XDFFPOSX1_7 INVX1_23/A CLKBUF1_11/Y XNOR2X1_6/Y gnd vdd DFFPOSX1
XFILL_8_2 gnd vdd FILL
XOAI21X1_83 INVX1_55/A OAI21X1_83/B OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_94 INVX4_5/Y INVX1_65/A OAI21X1_94/C gnd MUX2X1_2/A vdd OAI21X1
XOAI21X1_72 OAI21X1_71/Y AOI21X1_8/Y AOI21X1_9/Y gnd AOI22X1_5/D vdd OAI21X1
XOAI21X1_50 OAI21X1_50/A OAI22X1_7/Y OAI21X1_49/Y gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 INVX1_42/Y OAI21X1_57/Y INVX1_41/Y gnd AOI22X1_3/D vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_297 INVX4_7/A INVX1_118/Y BUFX4_8/Y gnd OAI22X1_12/C vdd OAI21X1
XOAI21X1_286 BUFX4_8/Y INVX1_184/Y OAI21X1_286/C gnd XNOR2X1_100/A vdd OAI21X1
XOAI21X1_253 BUFX4_26/Y INVX1_159/Y BUFX4_27/Y gnd INVX1_163/A vdd OAI21X1
XOAI21X1_242 AND2X2_11/Y NAND2X1_186/Y OAI21X1_241/Y gnd AOI22X1_28/C vdd OAI21X1
XOAI21X1_264 NOR2X1_145/B AOI21X1_57/Y AOI21X1_59/B gnd OAI21X1_266/B vdd OAI21X1
XOAI21X1_275 INVX1_178/A AOI21X1_60/Y OAI21X1_274/Y gnd MUX2X1_12/B vdd OAI21X1
XOAI21X1_220 NAND2X1_172/Y AOI21X1_43/Y AOI21X1_47/Y gnd AOI21X1_48/A vdd OAI21X1
XOAI21X1_231 INVX1_151/A OAI21X1_231/B INVX1_150/Y gnd NAND3X1_17/C vdd OAI21X1
XFILL_17_2_1 gnd vdd FILL
XINVX1_169 XOR2X1_29/B gnd INVX1_169/Y vdd INVX1
XINVX1_125 INVX1_125/A gnd NOR2X1_98/B vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_136 OR2X2_13/A gnd INVX1_136/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XINVX1_114 NOR2X1_82/Y gnd INVX1_114/Y vdd INVX1
XINVX1_103 AND2X2_7/A gnd INVX1_103/Y vdd INVX1
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XNOR2X1_64 NOR2X1_62/Y NOR2X1_63/Y gnd XOR2X1_13/B vdd NOR2X1
XNOR2X1_42 NOR2X1_41/Y NOR2X1_42/B gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_53 INVX4_5/A INVX2_8/Y gnd INVX1_77/A vdd NOR2X1
XNOR2X1_31 OR2X2_5/A OR2X2_5/B gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_20 INVX1_26/A NOR2X1_20/B gnd INVX1_28/A vdd NOR2X1
XNOR2X1_75 OR2X2_9/A OR2X2_9/B gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_86 NOR2X1_85/Y NOR2X1_86/B gnd NOR2X1_86/Y vdd NOR2X1
XNOR2X1_97 INVX4_8/Y INVX1_123/Y gnd INVX1_129/A vdd NOR2X1
XNAND2X1_8 BUFX2_9/Y NAND2X1_7/Y gnd NAND2X1_9/B vdd NAND2X1
XNOR2X1_154 OAI22X1_8/A INVX4_7/Y gnd AOI21X1_68/C vdd NOR2X1
XNOR2X1_143 INVX1_54/A INVX1_169/Y gnd NOR2X1_143/Y vdd NOR2X1
XNOR2X1_110 XNOR2X1_61/Y NOR2X1_110/B gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_132 INVX1_156/A INVX2_26/Y gnd NOR2X1_132/Y vdd NOR2X1
XNOR2X1_121 AND2X2_10/A INVX1_141/Y gnd AOI21X1_49/A vdd NOR2X1
XINVX1_56 OR2X2_6/B gnd INVX1_56/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XDFFPOSX1_8 DFFPOSX1_8/Q CLKBUF1_11/Y XNOR2X1_7/Y gnd vdd DFFPOSX1
XOAI21X1_84 INVX1_52/A INVX2_5/Y INVX8_2/A gnd INVX1_59/A vdd OAI21X1
XOAI21X1_73 BUFX2_1/Y AOI22X1_5/D NAND2X1_61/Y gnd XNOR2X1_28/A vdd OAI21X1
XOAI21X1_95 INVX4_5/Y INVX1_65/Y OAI21X1_95/C gnd MUX2X1_2/B vdd OAI21X1
XOAI21X1_62 INVX1_45/A INVX1_44/Y INVX8_2/A gnd OAI21X1_63/C vdd OAI21X1
XOAI21X1_40 INVX4_4/Y INVX1_28/Y NAND3X1_1/Y gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_51 OAI22X1_7/Y OAI21X1_50/Y OAI21X1_50/A gnd NAND2X1_40/B vdd OAI21X1
XFILL_1_2_2 gnd vdd FILL
XOAI21X1_221 BUFX4_3/Y AOI21X1_48/Y OAI21X1_221/C gnd XNOR2X1_80/A vdd OAI21X1
XOAI21X1_210 INVX2_13/A INVX1_139/Y OAI22X1_10/Y gnd INVX1_145/A vdd OAI21X1
XOAI21X1_287 BUFX4_9/Y AOI21X1_67/B OAI21X1_287/C gnd XNOR2X1_101/A vdd OAI21X1
XOAI21X1_254 INVX1_160/A NOR2X1_138/B INVX1_163/Y gnd NAND3X1_18/B vdd OAI21X1
XOAI21X1_265 NOR2X1_141/Y AOI21X1_58/Y INVX1_175/A gnd OAI21X1_265/Y vdd OAI21X1
XOAI21X1_243 BUFX2_8/Y AOI22X1_30/D OAI21X1_243/C gnd XNOR2X1_86/A vdd OAI21X1
XOAI21X1_276 INVX2_27/A INVX2_4/Y BUFX4_6/Y gnd INVX1_179/A vdd OAI21X1
XOAI21X1_232 AOI21X1_50/Y AOI21X1_51/Y INVX1_113/A gnd OAI21X1_232/Y vdd OAI21X1
XAND2X2_10 AND2X2_10/A AND2X2_10/B gnd OR2X2_14/A vdd AND2X2
XOAI21X1_298 INVX1_118/A INVX4_7/A INVX8_1/A gnd OAI22X1_12/A vdd OAI21X1
XFILL_17_2_2 gnd vdd FILL
XDFFSR_10 DFFSR_10/Q DFFSR_6/CLK DFFSR_11/R vdd vdd gnd vdd DFFSR
XINVX1_115 BUFX2_57/A gnd NOR2X1_88/A vdd INVX1
XINVX1_159 OR2X2_8/B gnd INVX1_159/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_126 OR2X2_12/A gnd INVX1_126/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XFILL_6_1_2 gnd vdd FILL
XFILL_14_0_2 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XNAND3X1_10 INVX1_109/Y NOR2X1_84/Y NAND3X1_10/C gnd NAND3X1_10/Y vdd NAND3X1
XNOR2X1_87 BUFX2_57/A INVX2_16/A gnd NOR2X1_87/Y vdd NOR2X1
XNOR2X1_43 OR2X2_7/A INVX4_5/A gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_32 AND2X2_3/A INVX2_5/A gnd OR2X2_6/B vdd NOR2X1
XNOR2X1_54 NOR2X1_52/Y INVX1_77/A gnd INVX1_71/A vdd NOR2X1
XNOR2X1_65 XOR2X1_11/Y NOR2X1_65/B gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_21 NOR2X1_21/A OR2X2_3/Y gnd NAND3X1_2/C vdd NOR2X1
XNOR2X1_10 INVX1_15/Y NOR2X1_10/B gnd NOR2X1_11/B vdd NOR2X1
XNOR2X1_76 AND2X2_7/A INVX2_14/A gnd OR2X2_10/B vdd NOR2X1
XNOR2X1_98 BUFX4_18/Y NOR2X1_98/B gnd NOR2X1_98/Y vdd NOR2X1
XNAND2X1_9 OAI21X1_9/Y NAND2X1_9/B gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_100 OR2X2_12/A INVX4_8/Y gnd NOR2X1_101/B vdd NOR2X1
XNOR2X1_133 AOI21X1_54/C NOR2X1_132/Y gnd INVX1_157/A vdd NOR2X1
XNOR2X1_144 INVX2_27/A INVX1_172/Y gnd INVX1_173/A vdd NOR2X1
XNOR2X1_111 INVX4_4/Y INVX2_21/Y gnd NOR2X1_111/Y vdd NOR2X1
XNOR2X1_122 NOR2X1_122/A OR2X2_14/Y gnd AOI21X1_45/A vdd NOR2X1
XNOR2X1_155 NOR2X1_155/A AOI21X1_68/A gnd NOR2X1_155/Y vdd NOR2X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_57 OR2X2_5/B gnd INVX1_57/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XDFFPOSX1_9 OAI22X1_3/A CLKBUF1_13/Y XNOR2X1_8/Y gnd vdd DFFPOSX1
XINVX1_35 OR2X2_4/B gnd INVX1_35/Y vdd INVX1
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_52 AOI21X1_7/A INVX1_40/Y INVX4_1/Y gnd OAI21X1_54/C vdd OAI21X1
XOAI21X1_63 INVX8_2/A INVX1_46/Y OAI21X1_63/C gnd XOR2X1_5/A vdd OAI21X1
XOAI21X1_30 INVX1_23/Y INVX1_22/Y INVX8_3/A gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_41 AOI21X1_4/Y NOR2X1_23/Y INVX4_4/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_85 INVX1_61/A OAI21X1_83/Y INVX1_59/Y gnd NAND3X1_6/C vdd OAI21X1
XOAI21X1_74 BUFX2_1/Y OAI21X1_74/B NAND3X1_4/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 INVX1_65/A INVX1_68/A INVX4_5/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_200 AOI21X1_41/Y AOI21X1_42/Y INVX1_76/A gnd OAI21X1_200/Y vdd OAI21X1
XOAI21X1_255 OR2X2_8/B BUFX2_6/Y INVX4_3/A gnd INVX1_164/A vdd OAI21X1
XOAI21X1_244 INVX1_152/A XNOR2X1_87/Y INVX1_158/Y gnd AOI22X1_27/D vdd OAI21X1
XOAI21X1_233 XOR2X1_25/B INVX2_9/Y BUFX2_7/Y gnd OAI21X1_234/C vdd OAI21X1
XOAI21X1_211 BUFX4_1/Y AOI21X1_45/B OAI21X1_211/C gnd XNOR2X1_75/A vdd OAI21X1
XOAI21X1_222 OR2X2_9/B NOR2X1_78/A INVX2_25/Y gnd OAI21X1_223/C vdd OAI21X1
XOAI21X1_288 INVX2_16/Y INVX4_7/Y NAND2X1_218/Y gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_299 INVX2_3/A NOR2X1_73/Y OAI21X1_137/Y gnd INVX1_186/A vdd OAI21X1
XOAI21X1_266 BUFX4_5/Y OAI21X1_266/B NAND2X1_202/Y gnd XNOR2X1_93/A vdd OAI21X1
XAND2X2_11 AND2X2_11/A AND2X2_11/B gnd AND2X2_11/Y vdd AND2X2
XOAI21X1_277 INVX1_176/A AOI22X1_33/Y INVX1_179/Y gnd NAND3X1_19/B vdd OAI21X1
XFILL_6_1 gnd vdd FILL
XDFFSR_11 DFFSR_11/Q DFFSR_6/CLK DFFSR_11/R vdd DFFSR_10/Q gnd vdd DFFSR
XFILL_1_0_0 gnd vdd FILL
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XINVX1_116 INVX1_116/A gnd OAI22X1_8/A vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XFILL_17_0_0 gnd vdd FILL
XNAND3X1_11 INVX1_113/A NAND3X1_11/B NAND3X1_11/C gnd NAND3X1_11/Y vdd NAND3X1
XNOR2X1_88 NOR2X1_88/A INVX2_16/Y gnd NOR2X1_89/B vdd NOR2X1
XNOR2X1_77 OR2X2_9/B INVX1_100/Y gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_66 INVX2_10/A INVX4_6/Y gnd NOR2X1_68/A vdd NOR2X1
XNOR2X1_99 INVX4_8/A INVX1_126/Y gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_44 OR2X2_7/B INVX1_64/Y gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_33 OR2X2_5/B INVX1_47/Y gnd AOI21X1_8/C vdd NOR2X1
XNOR2X1_55 INVX1_67/A XOR2X1_9/B gnd INVX1_74/A vdd NOR2X1
XNOR2X1_11 XNOR2X1_6/B NOR2X1_11/B gnd AND2X2_1/A vdd NOR2X1
XNOR2X1_22 INVX1_25/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_101 NOR2X1_99/Y NOR2X1_101/B gnd INVX2_20/A vdd NOR2X1
XNOR2X1_134 XNOR2X1_85/Y NOR2X1_134/B gnd AOI22X1_27/C vdd NOR2X1
XNOR2X1_145 XNOR2X1_95/Y NOR2X1_145/B gnd AOI21X1_61/B vdd NOR2X1
XNOR2X1_112 INVX2_21/A INVX1_137/Y gnd NOR2X1_112/Y vdd NOR2X1
XNOR2X1_123 INVX1_97/Y INVX2_15/Y gnd INVX1_142/A vdd NOR2X1
XNOR2X1_156 XOR2X1_33/Y MUX2X1_13/A gnd NOR2X1_156/Y vdd NOR2X1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_47 OR2X2_5/A gnd INVX1_47/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_14 OR2X2_1/B gnd INVX1_14/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_53 INVX1_39/Y INVX1_38/Y DFFSR_8/Q gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_86 OAI21X1_86/A OAI21X1_86/B INVX1_60/Y gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_64 NOR2X1_31/Y AND2X2_2/Y AOI21X1_8/B gnd OAI21X1_65/C vdd OAI21X1
XOAI21X1_75 INVX1_47/Y INVX1_57/Y INVX1_46/A gnd NAND2X1_65/B vdd OAI21X1
XOAI21X1_31 NOR2X1_15/Y OAI21X1_30/Y OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_42 OAI21X1_42/A INVX1_28/Y INVX1_29/Y gnd AOI22X1_1/C vdd OAI21X1
XOAI21X1_20 INVX8_1/A AND2X2_1/Y AOI21X1_1/B gnd XNOR2X1_8/A vdd OAI21X1
XOAI21X1_97 NAND2X1_79/Y OAI21X1_97/B OAI21X1_96/Y gnd AOI22X1_8/D vdd OAI21X1
XOAI21X1_289 INVX1_185/Y OAI21X1_287/C NAND2X1_211/Y gnd AOI21X1_69/A vdd OAI21X1
XOAI21X1_256 INVX1_165/A XNOR2X1_89/A INVX1_164/Y gnd NAND3X1_18/C vdd OAI21X1
XOAI21X1_234 BUFX2_7/Y INVX1_152/Y OAI21X1_234/C gnd XNOR2X1_82/A vdd OAI21X1
XOAI21X1_245 INVX1_157/A AOI22X1_27/Y NAND2X1_189/Y gnd MUX2X1_11/A vdd OAI21X1
XOAI21X1_267 INVX1_175/A XOR2X1_30/Y INVX1_173/Y gnd AOI21X1_60/C vdd OAI21X1
XOAI21X1_278 INVX1_44/A OR2X2_5/B INVX2_27/A gnd OAI21X1_278/Y vdd OAI21X1
XOAI21X1_201 OAI21X1_201/A NOR2X1_115/A INVX4_4/Y gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_223 INVX1_147/A OAI21X1_216/Y OAI21X1_223/C gnd MUX2X1_10/B vdd OAI21X1
XOAI21X1_212 OR2X2_14/Y AOI21X1_43/Y OAI21X1_217/A gnd OAI21X1_214/B vdd OAI21X1
XAND2X2_12 INVX1_52/A AND2X2_12/B gnd AND2X2_12/Y vdd AND2X2
XDFFPOSX1_170 INVX1_12/A DFFSR_8/CLK AOI22X1_2/Y gnd vdd DFFPOSX1
XFILL_6_2 gnd vdd FILL
XDFFSR_12 DFFSR_13/D DFFSR_6/CLK DFFSR_9/R vdd DFFSR_11/Q gnd vdd DFFSR
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XINVX1_128 AND2X2_9/B gnd INVX1_128/Y vdd INVX1
XINVX1_106 NOR2X1_83/Y gnd INVX1_106/Y vdd INVX1
XINVX1_139 XOR2X1_23/B gnd INVX1_139/Y vdd INVX1
XINVX1_117 BUFX2_58/A gnd INVX1_117/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XNOR2X1_12 INVX8_1/A AND2X2_1/Y gnd AOI21X1_1/C vdd NOR2X1
XNAND3X1_12 XOR2X1_34/B XOR2X1_16/B NAND3X1_12/C gnd NAND3X1_12/Y vdd NAND3X1
XNOR2X1_89 NOR2X1_87/Y NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_67 INVX4_6/A INVX2_10/Y gnd INVX1_93/A vdd NOR2X1
XNOR2X1_34 INVX2_4/A INVX1_48/Y gnd AOI21X1_9/B vdd NOR2X1
XNOR2X1_56 NOR2X1_56/A NOR2X1_56/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_45 INVX4_5/A INVX1_66/A gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_23 INVX2_2/Y NOR2X1_23/B gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A INVX1_102/Y gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_102 AND2X2_9/B AND2X2_9/A gnd NOR2X1_102/Y vdd NOR2X1
XNOR2X1_113 INVX1_137/A INVX2_21/Y gnd NOR2X1_114/B vdd NOR2X1
XNOR2X1_124 INVX1_110/Y INVX2_25/Y gnd AOI21X1_48/C vdd NOR2X1
XNOR2X1_135 OR2X2_8/B BUFX4_24/Y gnd NOR2X1_135/Y vdd NOR2X1
XNOR2X1_146 INVX2_27/Y INVX1_172/Y gnd INVX1_174/A vdd NOR2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_15 OR2X2_2/B gnd INVX1_15/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XFILL_4_2_2 gnd vdd FILL
XFILL_12_1_2 gnd vdd FILL
XOAI21X1_54 INVX1_40/Y OAI21X1_53/Y OAI21X1_54/C gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_87 INVX1_62/A INVX2_7/Y INVX4_2/A gnd OAI21X1_88/C vdd OAI21X1
XOAI21X1_98 INVX1_65/A INVX1_68/A BUFX4_13/Y gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_76 OAI21X1_71/C OAI21X1_76/B AOI22X1_4/C gnd NAND3X1_5/C vdd OAI21X1
XOAI21X1_65 INVX1_47/Y OR2X2_5/B OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_10 INVX4_3/A INVX1_11/Y NAND2X1_9/B gnd OAI21X1_13/A vdd OAI21X1
XOAI21X1_21 NOR2X1_13/Y NOR2X1_14/Y BUFX4_5/Y gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_43 INVX4_4/Y INVX2_2/Y INVX1_30/Y gnd AOI21X1_5/A vdd OAI21X1
XOAI21X1_32 INVX8_3/A NOR2X1_15/Y OAI21X1_30/Y gnd XNOR2X1_11/A vdd OAI21X1
XOAI21X1_257 AOI21X1_55/Y AOI21X1_56/Y INVX1_92/A gnd OAI21X1_257/Y vdd OAI21X1
XOAI21X1_235 INVX4_3/A AND2X2_11/Y NAND2X1_177/Y gnd XNOR2X1_83/A vdd OAI21X1
XOAI21X1_246 INVX1_78/A INVX1_156/A INVX2_26/Y gnd OAI21X1_246/Y vdd OAI21X1
XOAI21X1_268 AOI21X1_59/B XNOR2X1_95/Y INVX1_174/Y gnd AOI21X1_61/C vdd OAI21X1
XOAI21X1_279 AOI21X1_61/Y INVX1_180/Y OAI21X1_278/Y gnd OAI21X1_281/B vdd OAI21X1
XOAI21X1_202 NAND2X1_158/Y NOR2X1_116/B INVX4_4/A gnd NAND2X1_159/B vdd OAI21X1
XOAI21X1_224 OR2X2_14/B OR2X2_14/A NOR2X1_122/A gnd OAI21X1_225/A vdd OAI21X1
XOAI21X1_213 AOI21X1_49/A AOI21X1_44/Y BUFX4_2/Y gnd OAI21X1_213/Y vdd OAI21X1
XNAND2X1_230 rst theta[4] gnd DFFSR_5/S vdd NAND2X1
XDFFPOSX1_171 OR2X2_1/B DFFSR_8/CLK XNOR2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_160 DFFPOSX1_51/D DFFSR_2/CLK XOR2X1_3/Y gnd vdd DFFPOSX1
XDFFSR_13 DFFSR_14/D DFFSR_6/CLK DFFSR_9/R vdd DFFSR_13/D gnd vdd DFFSR
XCLKBUF1_11 clk gnd CLKBUF1_11/Y vdd CLKBUF1
XFILL_1_0_2 gnd vdd FILL
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XINVX1_107 AND2X2_10/A gnd INVX1_107/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XFILL_17_0_2 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XNAND3X1_13 INVX1_76/Y NAND3X1_13/B NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XNOR2X1_35 INVX2_5/A INVX1_49/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_46 INVX4_5/Y INVX1_66/Y gnd NOR2X1_47/B vdd NOR2X1
XNOR2X1_13 INVX1_18/A INVX1_17/A gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A INVX1_28/Y gnd OAI22X1_5/B vdd NOR2X1
XNOR2X1_68 NOR2X1_68/A INVX1_93/A gnd INVX1_87/A vdd NOR2X1
XNOR2X1_57 OR2X2_8/A OR2X2_8/B gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_79 AND2X2_7/A INVX2_14/Y gnd NOR2X1_79/Y vdd NOR2X1
XNOR2X1_147 INVX2_4/A INVX2_27/A gnd NOR2X1_147/Y vdd NOR2X1
XNOR2X1_136 INVX1_159/Y INVX2_26/Y gnd INVX1_165/A vdd NOR2X1
XNOR2X1_103 INVX4_8/Y INVX1_126/Y gnd NOR2X1_103/Y vdd NOR2X1
XNOR2X1_114 NOR2X1_112/Y NOR2X1_114/B gnd NOR2X1_114/Y vdd NOR2X1
XNOR2X1_125 AND2X2_7/A INVX2_25/A gnd NOR2X1_125/Y vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XDFFSR_1 DFFSR_1/Q DFFSR_2/CLK DFFSR_1/R DFFSR_1/S theta[0] gnd vdd DFFSR
XINVX1_49 AND2X2_3/A gnd INVX1_49/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_38 DFFSR_2/Q gnd INVX1_38/Y vdd INVX1
XNAND2X1_90 INVX1_79/A INVX1_78/A gnd INVX1_80/A vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_11 NAND2X1_10/Y OAI21X1_9/B INVX4_3/A gnd OAI21X1_12/C vdd OAI21X1
XOAI21X1_55 DFFSR_8/Q INVX1_40/Y OAI21X1_53/Y gnd XNOR2X1_21/A vdd OAI21X1
XOAI21X1_88 INVX4_2/A INVX1_63/Y OAI21X1_88/C gnd XOR2X1_6/A vdd OAI21X1
XOAI21X1_77 INVX2_6/A INVX1_54/A INVX2_5/A gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_99 INVX1_69/Y OAI21X1_95/C OAI21X1_98/Y gnd NAND2X1_80/B vdd OAI21X1
XOAI21X1_66 INVX1_46/A NOR2X1_31/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_44 INVX4_4/A INVX2_2/Y INVX1_30/A gnd AOI21X1_5/B vdd OAI21X1
XOAI21X1_22 INVX1_18/Y INVX1_17/Y INVX8_2/A gnd OAI21X1_24/C vdd OAI21X1
XOAI21X1_33 INVX8_3/A NOR2X1_15/Y NAND2X1_23/Y gnd OAI22X1_3/B vdd OAI21X1
XOAI21X1_203 OR2X2_13/Y NOR2X1_116/B NOR2X1_111/Y gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_258 INVX1_167/A INVX2_6/Y BUFX4_7/Y gnd OAI21X1_259/C vdd OAI21X1
XOAI21X1_236 NOR2X1_134/B AOI21X1_52/Y OAI21X1_236/C gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_247 INVX1_162/A AOI22X1_29/Y OAI21X1_246/Y gnd AOI21X1_55/A vdd OAI21X1
XOAI21X1_269 BUFX4_5/Y AOI21X1_61/Y NAND2X1_203/Y gnd XNOR2X1_96/A vdd OAI21X1
XOAI21X1_225 OAI21X1_225/A INVX1_145/Y AOI21X1_49/Y gnd AOI22X1_26/D vdd OAI21X1
XOAI21X1_214 BUFX4_2/Y OAI21X1_214/B OAI21X1_213/Y gnd XNOR2X1_76/A vdd OAI21X1
XNAND2X1_231 rst theta[5] gnd DFFSR_6/S vdd NAND2X1
XDFFPOSX1_150 INVX1_29/A CLKBUF1_10/Y XOR2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_161 INVX1_32/A DFFSR_8/CLK BUFX2_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_172 OR2X2_2/B CLKBUF1_12/Y XNOR2X1_19/Y gnd vdd DFFPOSX1
XNAND2X1_220 INVX1_116/A INVX4_7/Y gnd NAND2X1_220/Y vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XDFFSR_14 DFFSR_14/Q DFFSR_6/CLK DFFSR_9/R vdd DFFSR_14/D gnd vdd DFFSR
XCLKBUF1_12 clk gnd CLKBUF1_12/Y vdd CLKBUF1
XINVX1_119 NOR2X1_91/B gnd INVX1_119/Y vdd INVX1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNAND3X1_14 INVX4_4/A NOR2X1_114/B NAND3X1_14/C gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_36 INVX2_5/A INVX2_6/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_69 INVX1_84/A XOR2X1_13/B gnd INVX1_90/A vdd NOR2X1
XNOR2X1_58 OR2X2_8/B INVX1_81/Y gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_47 NOR2X1_45/Y NOR2X1_47/B gnd INVX1_67/A vdd NOR2X1
XNOR2X1_14 INVX1_18/Y INVX1_17/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_25 INVX4_4/Y OAI22X1_5/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_137 NOR2X1_135/Y INVX1_165/A gnd INVX1_160/A vdd NOR2X1
XNOR2X1_104 INVX2_7/A INVX4_8/A gnd NOR2X1_104/Y vdd NOR2X1
XNOR2X1_148 INVX2_4/Y INVX2_27/Y gnd INVX1_182/A vdd NOR2X1
XNOR2X1_115 NOR2X1_115/A NOR2X1_115/B gnd NOR2X1_115/Y vdd NOR2X1
XMUX2X1_10 MUX2X1_10/A MUX2X1_10/B INVX8_3/A gnd MUX2X1_10/Y vdd MUX2X1
XNOR2X1_126 INVX1_103/Y INVX2_25/Y gnd INVX1_151/A vdd NOR2X1
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_2/R DFFSR_2/S theta[1] gnd vdd DFFSR
XFILL_16_2 gnd vdd FILL
XINVX1_39 DFFSR_3/Q gnd INVX1_39/Y vdd INVX1
XNAND2X1_91 BUFX4_27/Y NAND2X1_92/A gnd NAND2X1_91/Y vdd NAND2X1
XNAND2X1_80 BUFX2_3/Y NAND2X1_80/B gnd NAND2X1_80/Y vdd NAND2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_12 OAI21X1_13/C OAI21X1_13/A OAI21X1_12/C gnd NAND2X1_11/B vdd OAI21X1
XOAI21X1_23 NOR2X1_13/Y OAI21X1_24/C OAI21X1_21/Y gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_34 OAI22X1_3/B OAI22X1_3/Y OAI22X1_3/A gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 INVX2_3/Y INVX1_34/Y AOI22X1_2/C gnd XNOR2X1_18/A vdd OAI21X1
XOAI21X1_78 INVX2_5/Y INVX1_52/Y BUFX4_7/Y gnd INVX1_58/A vdd OAI21X1
XOAI21X1_89 NOR2X1_43/Y AND2X2_4/Y OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XOAI21X1_67 BUFX4_6/Y OAI21X1_65/Y OAI21X1_67/C gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_56 INVX4_1/Y OAI21X1_56/B NAND2X1_43/Y gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_237 NOR2X1_130/Y AOI22X1_29/D BUFX2_7/Y gnd OAI21X1_238/C vdd OAI21X1
XOAI21X1_204 INVX2_22/A NOR2X1_115/Y OAI21X1_203/Y gnd XNOR2X1_69/A vdd OAI21X1
XOAI21X1_226 INVX2_25/A INVX1_103/Y BUFX4_4/Y gnd INVX1_148/A vdd OAI21X1
XOAI21X1_215 AND2X2_10/A INVX1_141/Y INVX1_146/A gnd OAI21X1_216/A vdd OAI21X1
XOAI21X1_248 NOR2X1_139/Y NOR2X1_138/Y BUFX2_8/Y gnd OAI21X1_248/Y vdd OAI21X1
XOAI21X1_259 BUFX4_7/Y INVX1_168/Y OAI21X1_259/C gnd XNOR2X1_90/A vdd OAI21X1
XDFFPOSX1_140 INVX1_68/A CLKBUF1_3/Y XNOR2X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_151 INVX1_30/A CLKBUF1_10/Y XNOR2X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 INVX1_31/A DFFSR_8/CLK INVX1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_173 XNOR2X1_6/B CLKBUF1_12/Y XOR2X1_4/Y gnd vdd DFFPOSX1
XNAND2X1_232 rst theta[6] gnd DFFSR_7/S vdd NAND2X1
XNAND2X1_210 BUFX4_8/Y OAI21X1_285/Y gnd OAI21X1_286/C vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_221 INVX4_7/A OAI22X1_8/A gnd NAND2X1_221/Y vdd NAND2X1
XDFFSR_15 DFFSR_16/D DFFSR_6/CLK BUFX4_22/Y vdd DFFSR_14/Q gnd vdd DFFSR
XCLKBUF1_13 clk gnd CLKBUF1_13/Y vdd CLKBUF1
XINVX1_109 OR2X2_10/B gnd INVX1_109/Y vdd INVX1
XFILL_10_2_2 gnd vdd FILL
XNAND3X1_15 INVX1_137/A NOR2X1_115/Y INVX2_22/Y gnd NAND3X1_15/Y vdd NAND3X1
XNOR2X1_37 INVX1_52/A INVX2_5/Y gnd NOR2X1_39/A vdd NOR2X1
XNOR2X1_59 INVX4_6/A INVX1_83/A gnd NOR2X1_59/Y vdd NOR2X1
XNOR2X1_48 XOR2X1_8/A INVX1_70/A gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_15 INVX1_23/A INVX1_22/A gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_26 INVX1_31/Y INVX1_32/Y gnd INVX1_34/A vdd NOR2X1
XMUX2X1_11 MUX2X1_11/A MUX2X1_11/B INVX4_3/A gnd MUX2X1_11/Y vdd MUX2X1
XNOR2X1_105 INVX2_7/Y INVX4_8/Y gnd INVX1_132/A vdd NOR2X1
XNOR2X1_138 INVX1_160/Y NOR2X1_138/B gnd NOR2X1_138/Y vdd NOR2X1
XNOR2X1_149 NOR2X1_147/Y INVX1_182/A gnd INVX1_176/A vdd NOR2X1
XNOR2X1_116 OR2X2_13/Y NOR2X1_116/B gnd NAND3X1_14/C vdd NOR2X1
XNOR2X1_127 NOR2X1_125/Y INVX1_151/A gnd INVX1_144/A vdd NOR2X1
XDFFSR_3 DFFSR_3/Q DFFSR_8/CLK DFFSR_3/R DFFSR_3/S theta[2] gnd vdd DFFSR
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XNAND2X1_70 NAND2X1_68/Y OAI21X1_89/C gnd NAND2X1_70/Y vdd NAND2X1
XNAND2X1_81 INVX1_65/Y INVX1_68/Y gnd AOI22X1_7/B vdd NAND2X1
XNAND2X1_92 NAND2X1_92/A NOR2X1_65/B gnd NAND2X1_92/Y vdd NAND2X1
XFILL_7_2_2 gnd vdd FILL
XFILL_15_1_2 gnd vdd FILL
XFILL_21_1 gnd vdd FILL
XOAI21X1_68 NOR2X1_42/B AOI21X1_8/Y NAND2X1_55/A gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_13 OAI21X1_13/A NAND2X1_11/B OAI21X1_13/C gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_24 INVX8_2/A NOR2X1_13/Y OAI21X1_24/C gnd XNOR2X1_9/A vdd OAI21X1
XOAI21X1_35 BUFX4_1/Y INVX1_24/Y OAI22X1_3/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_46 INVX1_31/Y INVX1_32/Y INVX1_36/Y gnd OR2X2_4/A vdd OAI21X1
XOAI21X1_57 DFFSR_4/Q INVX1_40/A DFFSR_5/Q gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_79 INVX1_53/A AOI22X1_6/Y INVX1_58/Y gnd NAND3X1_6/B vdd OAI21X1
XOAI21X1_238 BUFX2_7/Y OAI21X1_236/Y OAI21X1_238/C gnd XNOR2X1_84/A vdd OAI21X1
XOAI21X1_249 INVX1_78/A INVX1_156/A BUFX4_25/Y gnd OAI21X1_249/Y vdd OAI21X1
XOAI21X1_205 INVX4_4/Y INVX2_21/Y XOR2X1_21/B gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_227 INVX1_144/A AOI22X1_26/Y INVX1_148/Y gnd NAND3X1_17/B vdd OAI21X1
XOAI21X1_216 OAI21X1_216/A AOI21X1_44/Y AOI21X1_49/B gnd OAI21X1_216/Y vdd OAI21X1
XNAND2X1_211 INVX2_16/A INVX4_7/Y gnd NAND2X1_211/Y vdd NAND2X1
XDFFPOSX1_163 INVX1_36/A CLKBUF1_12/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XNAND2X1_200 AOI21X1_59/B AOI21X1_59/A gnd NOR2X1_145/B vdd NAND2X1
XDFFPOSX1_141 INVX1_66/A CLKBUF1_3/Y XNOR2X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 INVX2_21/A CLKBUF1_10/Y NAND2X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_130 OR2X2_8/A CLKBUF1_6/Y XOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_174 INVX1_16/A CLKBUF1_11/Y XNOR2X1_20/Y gnd vdd DFFPOSX1
XNAND2X1_233 rst theta[7] gnd DFFSR_8/S vdd NAND2X1
XFILL_4_0_2 gnd vdd FILL
XNAND2X1_222 NAND2X1_220/Y NAND2X1_221/Y gnd AOI21X1_68/A vdd NAND2X1
XDFFSR_16 DFFSR_16/Q DFFSR_6/CLK BUFX4_22/Y vdd DFFSR_16/D gnd vdd DFFSR
XFILL_13_2_0 gnd vdd FILL
XNAND3X1_16 INVX1_137/Y INVX2_23/Y NAND3X1_14/C gnd AOI22X1_24/D vdd NAND3X1
XNOR2X1_38 INVX2_5/A INVX1_52/Y gnd INVX1_61/A vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_49 INVX4_5/Y INVX1_70/Y gnd NOR2X1_50/B vdd NOR2X1
XNOR2X1_16 INVX1_23/Y INVX1_22/Y gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_27 INVX1_31/A INVX1_32/A gnd INVX1_33/A vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XNOR2X1_106 NOR2X1_104/Y INVX1_132/A gnd INVX1_127/A vdd NOR2X1
XMUX2X1_12 MUX2X1_12/A MUX2X1_12/B INVX8_2/A gnd MUX2X1_12/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_139 INVX1_160/A AOI21X1_55/A gnd NOR2X1_139/Y vdd NOR2X1
XNOR2X1_117 INVX1_137/Y INVX2_23/Y gnd NOR2X1_117/Y vdd NOR2X1
XNOR2X1_128 INVX1_143/A INVX2_24/Y gnd INVX1_149/A vdd NOR2X1
XDFFSR_4 DFFSR_4/Q DFFSR_6/CLK DFFSR_4/R DFFSR_4/S theta[3] gnd vdd DFFSR
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 NAND3X1_4/B NAND2X1_60/B gnd INVX1_51/A vdd NAND2X1
XNAND2X1_93 INVX4_6/Y INVX1_85/Y gnd INVX1_86/A vdd NAND2X1
XNAND2X1_71 OR2X2_7/A BUFX4_13/Y gnd NAND2X1_71/Y vdd NAND2X1
XNAND2X1_82 INVX1_66/A INVX4_5/Y gnd NAND2X1_82/Y vdd NAND2X1
XFILL_21_2 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_69 INVX1_48/Y INVX2_4/Y AOI22X1_4/D gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_25 INVX8_2/A INVX1_20/Y OAI21X1_25/C gnd XNOR2X1_10/A vdd OAI21X1
XOAI21X1_36 INVX4_4/Y OR2X2_3/A AOI21X1_3/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_14 INVX1_12/A INVX1_13/A OAI22X1_2/B gnd OAI22X1_1/D vdd OAI21X1
XOAI21X1_47 INVX2_3/Y OR2X2_4/A OAI22X1_7/D gnd XNOR2X1_19/A vdd OAI21X1
XOAI21X1_58 INVX4_1/Y AOI21X1_7/Y NAND2X1_44/Y gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_239 XOR2X1_27/B INVX1_154/A BUFX2_6/Y gnd OAI21X1_240/C vdd OAI21X1
XOAI21X1_206 XOR2X1_21/B INVX2_22/Y OAI21X1_205/Y gnd OAI21X1_206/Y vdd OAI21X1
XOAI21X1_228 OR2X2_9/B NOR2X1_78/A INVX2_25/A gnd OAI21X1_228/Y vdd OAI21X1
XOAI21X1_217 OAI21X1_217/A NOR2X1_122/A INVX1_142/Y gnd AOI21X1_45/C vdd OAI21X1
XNAND2X1_223 NOR2X1_155/A OAI21X1_288/Y gnd OAI21X1_291/C vdd NAND2X1
XNAND2X1_212 INVX4_7/A INVX2_16/Y gnd INVX1_185/A vdd NAND2X1
XNAND2X1_201 AND2X2_12/B INVX1_52/Y gnd INVX1_175/A vdd NAND2X1
XDFFPOSX1_142 INVX1_70/A CLKBUF1_3/Y XOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 INVX1_82/A CLKBUF1_1/Y XNOR2X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 INVX2_25/A CLKBUF1_13/Y OAI21X1_173/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 DFFPOSX1_44/D DFFSR_2/CLK XOR2X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_164 OR2X2_4/B CLKBUF1_12/Y XNOR2X1_21/Y gnd vdd DFFPOSX1
XDFFSR_17 DFFSR_9/D DFFSR_6/CLK DFFSR_11/R vdd DFFSR_16/Q gnd vdd DFFSR
XXNOR2X1_1 OAI21X1_7/Y NOR2X1_7/A gnd XNOR2X1_1/Y vdd XNOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XAND2X2_1 AND2X2_1/A INVX1_16/Y gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_17 INVX2_2/A INVX1_25/A gnd NOR2X1_17/Y vdd NOR2X1
XNAND3X1_17 INVX1_113/Y NAND3X1_17/B NAND3X1_17/C gnd NAND3X1_17/Y vdd NAND3X1
XNOR2X1_28 XOR2X1_4/B OR2X2_4/Y gnd NOR2X1_28/Y vdd NOR2X1
XNOR2X1_39 NOR2X1_39/A INVX1_61/A gnd INVX1_53/A vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_107 INVX1_128/Y INVX2_20/Y gnd AOI22X1_18/D vdd NOR2X1
XNOR2X1_129 INVX2_10/Y INVX1_153/Y gnd INVX1_158/A vdd NOR2X1
XNOR2X1_118 AND2X2_10/A AND2X2_10/B gnd OR2X2_14/B vdd NOR2X1
XMUX2X1_13 MUX2X1_13/A MUX2X1_13/B BUFX4_9/Y gnd MUX2X1_13/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XDFFSR_5 DFFSR_5/Q DFFSR_6/CLK DFFSR_5/R DFFSR_5/S theta[4] gnd vdd DFFSR
XNAND2X1_61 BUFX2_1/Y AOI22X1_4/Y gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_50 OAI21X1_66/C OR2X2_5/Y gnd XOR2X1_5/B vdd NAND2X1
XNAND2X1_72 NAND2X1_71/Y OR2X2_7/Y gnd XOR2X1_6/B vdd NAND2X1
XNAND2X1_94 INVX4_6/A INVX1_85/A gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_83 INVX1_66/Y INVX1_70/Y gnd AOI22X1_8/B vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_26 INVX1_21/Y NAND2X1_19/Y INVX8_2/A gnd NAND2X1_21/A vdd OAI21X1
XOAI21X1_37 OR2X2_3/A OR2X2_3/B INVX2_2/A gnd OAI22X1_4/B vdd OAI21X1
XOAI21X1_15 BUFX4_10/Y OR2X2_1/A OAI22X1_2/B gnd XNOR2X1_4/A vdd OAI21X1
XOAI21X1_59 INVX1_42/Y OAI21X1_57/Y INVX4_1/Y gnd OAI21X1_60/C vdd OAI21X1
XOAI21X1_48 OAI22X1_7/D OAI22X1_7/C NAND2X1_38/Y gnd XNOR2X1_20/A vdd OAI21X1
XOAI21X1_229 INVX1_149/Y AOI21X1_45/Y OAI21X1_228/Y gnd OAI21X1_231/B vdd OAI21X1
XOAI21X1_218 BUFX4_3/Y AOI21X1_45/Y OAI21X1_218/C gnd XNOR2X1_79/A vdd OAI21X1
XOAI21X1_207 XOR2X1_22/B INVX2_14/Y BUFX4_2/Y gnd OAI21X1_207/Y vdd OAI21X1
XDFFPOSX1_110 NOR2X1_91/B CLKBUF1_12/Y INVX1_96/A gnd vdd DFFPOSX1
XDFFPOSX1_121 INVX1_45/A CLKBUF1_9/Y NAND2X1_104/Y gnd vdd DFFPOSX1
XNAND2X1_213 NAND2X1_211/Y INVX1_185/A gnd AOI21X1_67/A vdd NAND2X1
XNAND2X1_224 BUFX4_9/Y NAND2X1_224/B gnd OAI21X1_294/C vdd NAND2X1
XNAND2X1_202 BUFX4_5/Y OAI21X1_265/Y gnd NAND2X1_202/Y vdd NAND2X1
XDFFPOSX1_143 INVX2_8/A CLKBUF1_5/Y XNOR2X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_132 INVX1_85/A CLKBUF1_1/Y XNOR2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 DFFPOSX1_45/D DFFSR_8/CLK XNOR2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_165 XOR2X1_4/B CLKBUF1_12/Y XNOR2X1_22/Y gnd vdd DFFPOSX1
XXNOR2X1_2 OAI21X1_8/Y INVX2_1/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XFILL_13_2_2 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XAND2X2_2 OR2X2_5/A OR2X2_5/B gnd AND2X2_2/Y vdd AND2X2
XFILL_2_2 gnd vdd FILL
XNOR2X1_29 INVX1_39/Y INVX1_38/Y gnd AOI21X1_7/A vdd NOR2X1
XNAND3X1_18 INVX1_92/Y NAND3X1_18/B NAND3X1_18/C gnd NAND3X1_18/Y vdd NAND3X1
XNOR2X1_18 INVX2_2/Y INVX1_25/Y gnd INVX1_27/A vdd NOR2X1
XFILL_2_1_2 gnd vdd FILL
XFILL_10_0_2 gnd vdd FILL
XNOR2X1_108 INVX1_127/Y NOR2X1_108/B gnd NOR2X1_108/Y vdd NOR2X1
XNOR2X1_119 OR2X2_14/B OR2X2_14/A gnd AOI21X1_44/C vdd NOR2X1
XFILL_18_1_2 gnd vdd FILL
XDFFSR_6 DFFSR_6/Q DFFSR_6/CLK DFFSR_6/R DFFSR_6/S theta[5] gnd vdd DFFSR
XNAND2X1_73 INVX1_62/A INVX2_7/A gnd INVX1_63/A vdd NAND2X1
XNAND2X1_62 INVX1_51/Y AOI22X1_4/Y gnd NAND3X1_4/C vdd NAND2X1
XNAND2X1_95 NAND2X1_94/Y INVX1_86/A gnd NOR2X1_70/B vdd NAND2X1
XNAND2X1_84 NAND3X1_7/Y NAND2X1_84/B gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_51 INVX1_45/A INVX1_44/A gnd INVX1_46/A vdd NAND2X1
XNAND2X1_40 NAND2X1_40/A NAND2X1_40/B gnd DFFPOSX1_1/D vdd NAND2X1
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XFILL_7_0_2 gnd vdd FILL
XOAI21X1_16 BUFX4_10/Y OR2X2_2/Y NAND2X1_16/Y gnd XNOR2X1_6/A vdd OAI21X1
XOAI21X1_27 OAI21X1_27/A AOI21X1_2/Y NAND2X1_21/A gnd NAND2X1_21/B vdd OAI21X1
XOAI21X1_38 OR2X2_3/Y OAI21X1_38/B INVX4_4/Y gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_49 INVX1_37/Y NOR2X1_28/Y INVX2_3/A gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_219 INVX1_143/Y OAI21X1_216/Y AOI21X1_46/Y gnd OAI21X1_221/C vdd OAI21X1
XOAI21X1_208 BUFX4_2/Y INVX1_138/Y OAI21X1_207/Y gnd XNOR2X1_73/A vdd OAI21X1
XDFFPOSX1_111 INVX4_7/A CLKBUF1_12/Y BUFX2_47/A gnd vdd DFFPOSX1
XDFFPOSX1_144 BUFX4_16/A CLKBUF1_5/Y NAND2X1_101/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 INVX1_83/A CLKBUF1_1/Y XNOR2X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 OR2X2_5/A CLKBUF1_6/Y XOR2X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 DFFPOSX1_37/D DFFSR_2/CLK XNOR2X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_155 DFFPOSX1_46/D DFFSR_2/CLK XOR2X1_2/Y gnd vdd DFFPOSX1
XNAND2X1_214 INVX1_119/Y OAI21X1_285/Y gnd OAI21X1_287/C vdd NAND2X1
XNAND2X1_203 BUFX4_5/Y AOI21X1_60/Y gnd NAND2X1_203/Y vdd NAND2X1
XDFFPOSX1_166 INVX1_37/A CLKBUF1_12/Y XNOR2X1_23/Y gnd vdd DFFPOSX1
XNAND2X1_225 NOR2X1_155/A AOI21X1_68/A gnd NAND2X1_225/Y vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XXNOR2X1_3 NAND2X1_9/Y INVX1_11/A gnd XNOR2X1_3/Y vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_2/A vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XAND2X2_3 AND2X2_3/A INVX2_5/A gnd OR2X2_6/A vdd AND2X2
XNAND3X1_19 INVX1_60/Y NAND3X1_19/B NAND3X1_19/C gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_19 NOR2X1_17/Y INVX1_27/A gnd XOR2X1_2/A vdd NOR2X1
XNOR2X1_109 INVX1_127/A NOR2X1_109/B gnd NOR2X1_109/Y vdd NOR2X1
XDFFSR_7 DFFSR_7/Q DFFSR_8/CLK DFFSR_7/R DFFSR_7/S theta[6] gnd vdd DFFSR
XNAND2X1_41 INVX1_39/Y INVX1_38/Y gnd INVX1_40/A vdd NAND2X1
XNAND2X1_63 INVX2_6/Y INVX1_54/Y gnd AOI22X1_6/B vdd NAND2X1
XNAND2X1_85 INVX1_79/A INVX1_78/Y gnd NAND2X1_85/Y vdd NAND2X1
XNAND2X1_74 BUFX2_4/Y AOI22X1_9/C gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_96 NOR2X1_70/A NOR2X1_70/B gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_52 BUFX4_6/Y OAI21X1_66/Y gnd OAI21X1_67/C vdd NAND2X1
XNAND2X1_30 INVX1_25/A NOR2X1_21/A gnd NOR2X1_20/B vdd NAND2X1
XOAI22X1_1 BUFX4_10/Y OR2X2_1/A NOR2X1_9/Y OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XOAI21X1_28 AOI21X1_2/Y NAND2X1_21/B OAI21X1_27/A gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_39 INVX1_26/A INVX1_27/Y INVX4_4/A gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_17 OR2X2_2/B OR2X2_2/A XNOR2X1_6/B gnd OAI21X1_17/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XOAI21X1_209 INVX1_138/A XNOR2X1_74/Y INVX1_140/Y gnd AOI21X1_45/B vdd OAI21X1
XDFFPOSX1_134 INVX2_9/A CLKBUF1_1/Y XNOR2X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 OR2X2_3/A CLKBUF1_5/Y NAND2X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 DFFPOSX1_38/D CLKBUF1_7/Y XOR2X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 INVX1_48/A CLKBUF1_6/Y XNOR2X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 DFFPOSX1_47/D DFFSR_2/CLK XNOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_167 OAI21X1_50/A CLKBUF1_12/Y XNOR2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 INVX2_18/A CLKBUF1_12/Y INVX1_96/Y gnd vdd DFFPOSX1
XNAND2X1_204 XNOR2X1_94/Y AOI22X1_33/D gnd AOI22X1_31/A vdd NAND2X1
XNAND2X1_226 rst theta[0] gnd DFFSR_1/S vdd NAND2X1
XNAND2X1_215 INVX2_17/A INVX2_18/Y gnd OAI21X1_296/A vdd NAND2X1
XFILL_0_2_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XOR2X2_20 DFFSR_9/R theta[5] gnd DFFSR_6/R vdd OR2X2
XXNOR2X1_4 XNOR2X1_4/A INVX1_14/Y gnd XNOR2X1_4/Y vdd XNOR2X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XAND2X2_4 OR2X2_7/A OR2X2_7/B gnd AND2X2_4/Y vdd AND2X2
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_8/R DFFSR_8/S theta[7] gnd vdd DFFSR
XNAND2X1_42 DFFSR_4/Q AOI21X1_7/A gnd OAI21X1_56/B vdd NAND2X1
XNAND2X1_64 INVX1_50/A INVX1_51/A gnd INVX1_55/A vdd NAND2X1
XNAND2X1_86 INVX1_78/A INVX1_79/Y gnd AOI21X1_19/B vdd NAND2X1
XNAND2X1_97 BUFX4_27/Y NAND2X1_97/B gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_53 INVX1_48/A INVX2_4/Y gnd NAND2X1_55/A vdd NAND2X1
XNAND2X1_75 AOI22X1_9/C XOR2X1_8/Y gnd OAI21X1_95/C vdd NAND2X1
XNAND2X1_20 INVX8_2/A NAND2X1_19/Y gnd OAI21X1_25/C vdd NAND2X1
XNAND2X1_31 INVX2_2/A OAI21X1_40/Y gnd NAND2X1_31/Y vdd NAND2X1
XOAI22X1_2 INVX1_14/Y OAI22X1_2/B BUFX4_10/Y OR2X2_2/A gnd XNOR2X1_5/A vdd OAI22X1
XINVX2_11 BUFX2_55/A gnd INVX2_11/Y vdd INVX2
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XOAI21X1_29 NOR2X1_15/Y NOR2X1_16/Y BUFX4_1/Y gnd OAI21X1_31/C vdd OAI21X1
XOAI21X1_18 INVX8_1/A AND2X2_1/A NAND2X1_17/Y gnd XNOR2X1_7/A vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_113 INVX1_98/A DFFSR_8/CLK vdd gnd vdd DFFPOSX1
XNAND2X1_216 INVX2_18/A INVX2_17/Y gnd NAND2X1_217/B vdd NAND2X1
XDFFPOSX1_135 INVX2_10/A CLKBUF1_1/Y XNOR2X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_102 DFFPOSX1_39/D CLKBUF1_7/Y XNOR2X1_68/Y gnd vdd DFFPOSX1
XNAND2X1_205 INVX1_44/A INVX2_27/A gnd NAND2X1_205/Y vdd NAND2X1
XDFFPOSX1_124 AND2X2_3/A CLKBUF1_6/Y XNOR2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_146 OR2X2_3/B CLKBUF1_5/Y XOR2X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 INVX2_3/A DFFSR_8/CLK AOI22X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 DFFPOSX1_48/D DFFSR_6/CLK XNOR2X1_14/Y gnd vdd DFFPOSX1
XNAND2X1_227 rst theta[1] gnd DFFSR_2/S vdd NAND2X1
XFILL_0_2_2 gnd vdd FILL
XFILL_16_2_2 gnd vdd FILL
XOR2X2_21 OR2X2_18/A theta[6] gnd DFFSR_7/R vdd OR2X2
XOR2X2_10 AND2X2_7/Y OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XXNOR2X1_5 XNOR2X1_5/A INVX1_15/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends


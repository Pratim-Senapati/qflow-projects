VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO noc_top
  CLASS BLOCK ;
  FOREIGN noc_top ;
  ORIGIN 1.900 4.000 ;
  SIZE 693.400 BY 508.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 30.600 490.800 31.400 491.000 ;
        RECT 75.400 490.800 76.200 491.000 ;
        RECT 4.400 490.200 31.400 490.800 ;
        RECT 49.200 490.200 76.200 490.800 ;
        RECT 170.200 490.800 171.000 491.000 ;
        RECT 208.600 490.800 209.400 491.000 ;
        RECT 288.200 490.800 289.000 491.000 ;
        RECT 328.200 490.800 329.000 491.000 ;
        RECT 170.200 490.200 197.200 490.800 ;
        RECT 208.600 490.200 235.600 490.800 ;
        RECT 262.000 490.200 289.000 490.800 ;
        RECT 302.000 490.200 329.000 490.800 ;
        RECT 349.400 490.800 350.200 491.000 ;
        RECT 389.400 490.800 390.200 491.000 ;
        RECT 448.600 490.800 449.400 491.000 ;
        RECT 495.000 490.800 495.800 491.000 ;
        RECT 554.200 490.800 555.000 491.000 ;
        RECT 619.400 490.800 620.200 491.000 ;
        RECT 349.400 490.200 376.400 490.800 ;
        RECT 389.400 490.200 416.400 490.800 ;
        RECT 448.600 490.200 475.600 490.800 ;
        RECT 495.000 490.200 522.000 490.800 ;
        RECT 554.200 490.200 581.200 490.800 ;
        RECT 4.400 489.600 5.200 490.200 ;
        RECT 7.800 490.000 8.600 490.200 ;
        RECT 1.200 481.600 2.000 486.200 ;
        RECT 4.400 481.600 5.200 486.200 ;
        RECT 7.600 481.600 8.400 486.200 ;
        RECT 14.000 481.600 14.800 486.200 ;
        RECT 17.200 481.600 18.000 486.200 ;
        RECT 25.200 481.600 26.000 486.200 ;
        RECT 28.400 481.600 29.200 486.200 ;
        RECT 31.600 481.600 32.400 486.200 ;
        RECT 34.800 481.600 35.600 486.200 ;
        RECT 37.000 481.600 37.800 486.200 ;
        RECT 41.200 481.600 42.000 490.200 ;
        RECT 49.200 489.600 50.000 490.200 ;
        RECT 52.400 490.000 53.400 490.200 ;
        RECT 44.400 481.600 45.200 486.200 ;
        RECT 46.000 481.600 46.800 486.200 ;
        RECT 49.200 481.600 50.000 486.200 ;
        RECT 52.400 481.600 53.200 486.200 ;
        RECT 58.800 481.600 59.600 486.200 ;
        RECT 62.000 481.600 62.800 486.200 ;
        RECT 70.000 481.600 70.800 486.200 ;
        RECT 73.200 481.600 74.000 486.200 ;
        RECT 76.400 481.600 77.200 486.200 ;
        RECT 79.600 481.600 80.400 486.200 ;
        RECT 81.200 481.600 82.000 486.200 ;
        RECT 84.400 481.600 85.200 490.200 ;
        RECT 88.600 481.600 89.400 486.200 ;
        RECT 91.400 481.600 92.200 486.200 ;
        RECT 95.600 481.600 96.400 490.200 ;
        RECT 97.200 481.600 98.000 490.200 ;
        RECT 100.400 481.600 101.200 490.200 ;
        RECT 103.600 481.600 104.400 490.200 ;
        RECT 106.800 481.600 107.600 490.200 ;
        RECT 110.000 481.600 110.800 490.200 ;
        RECT 118.000 481.600 118.800 490.000 ;
        RECT 123.600 481.600 124.400 486.200 ;
        RECT 126.800 481.600 127.600 486.200 ;
        RECT 132.400 481.600 133.200 490.200 ;
        RECT 135.600 481.600 136.400 490.200 ;
        RECT 138.800 481.600 139.600 490.200 ;
        RECT 142.000 481.600 142.800 490.200 ;
        RECT 145.200 481.600 146.000 490.200 ;
        RECT 148.400 481.600 149.200 490.200 ;
        RECT 150.000 481.600 150.800 490.200 ;
        RECT 154.200 481.600 155.000 486.200 ;
        RECT 156.400 481.600 157.200 486.200 ;
        RECT 159.600 481.600 160.400 490.200 ;
        RECT 193.000 490.000 193.800 490.200 ;
        RECT 196.400 489.600 197.200 490.200 ;
        RECT 231.400 490.000 232.200 490.200 ;
        RECT 234.800 489.600 235.600 490.200 ;
        RECT 163.800 481.600 164.600 486.200 ;
        RECT 166.000 481.600 166.800 486.200 ;
        RECT 169.200 481.600 170.000 486.200 ;
        RECT 172.400 481.600 173.200 486.200 ;
        RECT 175.600 481.600 176.400 486.200 ;
        RECT 183.600 481.600 184.400 486.200 ;
        RECT 186.800 481.600 187.600 486.200 ;
        RECT 193.200 481.600 194.000 486.200 ;
        RECT 196.400 481.600 197.200 486.200 ;
        RECT 199.600 481.600 200.400 486.200 ;
        RECT 201.200 481.600 202.000 486.200 ;
        RECT 204.400 481.600 205.200 486.200 ;
        RECT 207.600 481.600 208.400 486.200 ;
        RECT 210.800 481.600 211.600 486.200 ;
        RECT 214.000 481.600 214.800 486.200 ;
        RECT 222.000 481.600 222.800 486.200 ;
        RECT 225.200 481.600 226.000 486.200 ;
        RECT 231.600 481.600 232.400 486.200 ;
        RECT 234.800 481.600 235.600 486.200 ;
        RECT 238.000 481.600 238.800 486.200 ;
        RECT 239.600 481.600 240.400 490.200 ;
        RECT 242.800 481.600 243.600 490.200 ;
        RECT 246.000 481.600 246.800 490.200 ;
        RECT 249.200 481.600 250.000 490.200 ;
        RECT 252.400 481.600 253.200 490.200 ;
        RECT 262.000 489.600 262.800 490.200 ;
        RECT 265.400 490.000 266.200 490.200 ;
        RECT 302.000 489.600 302.800 490.200 ;
        RECT 305.400 490.000 306.200 490.200 ;
        RECT 372.200 490.000 373.200 490.200 ;
        RECT 375.600 489.600 376.400 490.200 ;
        RECT 412.200 490.000 413.200 490.200 ;
        RECT 415.600 489.600 416.400 490.200 ;
        RECT 258.800 481.600 259.600 486.200 ;
        RECT 262.000 481.600 262.800 486.200 ;
        RECT 265.200 481.600 266.000 486.200 ;
        RECT 271.600 481.600 272.400 486.200 ;
        RECT 274.800 481.600 275.600 486.200 ;
        RECT 282.800 481.600 283.600 486.200 ;
        RECT 286.000 481.600 286.800 486.200 ;
        RECT 289.200 481.600 290.000 486.200 ;
        RECT 292.400 481.600 293.200 486.200 ;
        RECT 295.600 481.600 296.400 489.000 ;
        RECT 298.800 481.600 299.600 486.200 ;
        RECT 302.000 481.600 302.800 486.200 ;
        RECT 305.200 481.600 306.000 486.200 ;
        RECT 311.600 481.600 312.400 486.200 ;
        RECT 314.800 481.600 315.600 486.200 ;
        RECT 322.800 481.600 323.600 486.200 ;
        RECT 326.000 481.600 326.800 486.200 ;
        RECT 329.200 481.600 330.000 486.200 ;
        RECT 332.400 481.600 333.200 486.200 ;
        RECT 335.600 482.200 336.600 488.800 ;
        RECT 335.800 481.600 336.600 482.200 ;
        RECT 341.800 481.600 342.800 488.800 ;
        RECT 345.200 481.600 346.000 486.200 ;
        RECT 348.400 481.600 349.200 486.200 ;
        RECT 351.600 481.600 352.400 486.200 ;
        RECT 354.800 481.600 355.600 486.200 ;
        RECT 362.800 481.600 363.600 486.200 ;
        RECT 366.000 481.600 366.800 486.200 ;
        RECT 372.400 481.600 373.200 486.200 ;
        RECT 375.600 481.600 376.400 486.200 ;
        RECT 378.800 481.600 379.600 486.200 ;
        RECT 382.000 481.600 382.800 489.000 ;
        RECT 385.200 481.600 386.000 486.200 ;
        RECT 388.400 481.600 389.200 486.200 ;
        RECT 391.600 481.600 392.400 486.200 ;
        RECT 394.800 481.600 395.600 486.200 ;
        RECT 402.800 481.600 403.600 486.200 ;
        RECT 406.000 481.600 406.800 486.200 ;
        RECT 412.400 481.600 413.200 486.200 ;
        RECT 415.600 481.600 416.400 486.200 ;
        RECT 418.800 481.600 419.600 486.200 ;
        RECT 426.800 481.600 427.600 489.000 ;
        RECT 430.000 481.600 430.800 486.200 ;
        RECT 433.200 481.600 434.000 490.200 ;
        RECT 471.400 490.000 472.200 490.200 ;
        RECT 474.800 489.600 475.600 490.200 ;
        RECT 517.800 490.000 518.800 490.200 ;
        RECT 521.200 489.600 522.000 490.200 ;
        RECT 437.400 481.600 438.200 486.200 ;
        RECT 439.600 481.600 440.400 486.200 ;
        RECT 442.800 481.600 443.600 486.200 ;
        RECT 444.400 481.600 445.200 486.200 ;
        RECT 447.600 481.600 448.400 486.200 ;
        RECT 450.800 481.600 451.600 486.200 ;
        RECT 454.000 481.600 454.800 486.200 ;
        RECT 462.000 481.600 462.800 486.200 ;
        RECT 465.200 481.600 466.000 486.200 ;
        RECT 471.600 481.600 472.400 486.200 ;
        RECT 474.800 481.600 475.600 486.200 ;
        RECT 478.000 481.600 478.800 486.200 ;
        RECT 479.600 481.600 480.400 486.200 ;
        RECT 484.400 481.600 485.200 486.200 ;
        RECT 487.600 481.600 488.400 489.000 ;
        RECT 490.800 481.600 491.600 486.200 ;
        RECT 494.000 481.600 494.800 486.200 ;
        RECT 497.200 481.600 498.000 486.200 ;
        RECT 500.400 481.600 501.200 486.200 ;
        RECT 508.400 481.600 509.200 486.200 ;
        RECT 511.600 481.600 512.400 486.200 ;
        RECT 518.000 481.600 518.800 486.200 ;
        RECT 521.200 481.600 522.000 486.200 ;
        RECT 524.400 481.600 525.200 486.200 ;
        RECT 526.000 481.600 526.800 486.200 ;
        RECT 529.200 481.600 530.000 490.200 ;
        RECT 533.400 481.600 534.200 486.200 ;
        RECT 535.600 481.600 536.400 486.200 ;
        RECT 538.800 481.600 539.600 486.200 ;
        RECT 541.000 481.600 541.800 486.200 ;
        RECT 545.200 481.600 546.000 490.200 ;
        RECT 577.000 490.000 578.000 490.200 ;
        RECT 580.400 489.600 581.200 490.200 ;
        RECT 593.200 490.200 620.200 490.800 ;
        RECT 655.000 490.800 655.800 491.000 ;
        RECT 655.000 490.200 682.000 490.800 ;
        RECT 593.200 489.600 594.000 490.200 ;
        RECT 596.600 490.000 597.400 490.200 ;
        RECT 548.400 481.600 549.200 486.200 ;
        RECT 550.000 481.600 550.800 486.200 ;
        RECT 553.200 481.600 554.000 486.200 ;
        RECT 556.400 481.600 557.200 486.200 ;
        RECT 559.600 481.600 560.400 486.200 ;
        RECT 567.600 481.600 568.400 486.200 ;
        RECT 570.800 481.600 571.600 486.200 ;
        RECT 577.200 481.600 578.000 486.200 ;
        RECT 580.400 481.600 581.200 486.200 ;
        RECT 583.600 481.600 584.400 486.200 ;
        RECT 590.000 481.600 590.800 486.200 ;
        RECT 593.200 481.600 594.000 486.200 ;
        RECT 596.400 481.600 597.200 486.200 ;
        RECT 602.800 481.600 603.600 486.200 ;
        RECT 606.000 481.600 606.800 486.200 ;
        RECT 614.000 481.600 614.800 486.200 ;
        RECT 617.200 481.600 618.000 486.200 ;
        RECT 620.400 481.600 621.200 486.200 ;
        RECT 623.600 481.600 624.400 486.200 ;
        RECT 626.800 482.200 627.800 488.800 ;
        RECT 627.000 481.600 627.800 482.200 ;
        RECT 633.000 481.600 634.000 488.800 ;
        RECT 636.400 481.600 637.200 490.200 ;
        RECT 639.600 481.600 640.400 490.200 ;
        RECT 642.800 481.600 643.600 490.200 ;
        RECT 646.000 481.600 646.800 490.200 ;
        RECT 649.200 481.600 650.000 490.200 ;
        RECT 677.800 490.000 678.600 490.200 ;
        RECT 681.200 489.600 682.000 490.200 ;
        RECT 650.800 481.600 651.600 486.200 ;
        RECT 654.000 481.600 654.800 486.200 ;
        RECT 657.200 481.600 658.000 486.200 ;
        RECT 660.400 481.600 661.200 486.200 ;
        RECT 668.400 481.600 669.200 486.200 ;
        RECT 671.600 481.600 672.400 486.200 ;
        RECT 678.000 481.600 678.800 486.200 ;
        RECT 681.200 481.600 682.000 486.200 ;
        RECT 684.400 481.600 685.200 486.200 ;
        RECT 0.400 480.400 689.200 481.600 ;
        RECT 1.200 475.800 2.000 480.400 ;
        RECT 4.400 475.800 5.200 480.400 ;
        RECT 7.600 475.800 8.400 480.400 ;
        RECT 10.800 475.800 11.600 480.400 ;
        RECT 18.800 475.800 19.600 480.400 ;
        RECT 22.000 475.800 22.800 480.400 ;
        RECT 28.400 475.800 29.200 480.400 ;
        RECT 31.600 475.800 32.400 480.400 ;
        RECT 34.800 475.800 35.600 480.400 ;
        RECT 37.000 475.800 37.800 480.400 ;
        RECT 28.200 471.800 29.000 472.000 ;
        RECT 31.600 471.800 32.400 472.400 ;
        RECT 41.200 471.800 42.000 480.400 ;
        RECT 42.800 475.800 43.600 480.400 ;
        RECT 46.000 475.800 46.800 480.400 ;
        RECT 49.200 472.000 50.000 480.400 ;
        RECT 54.800 475.800 55.600 480.400 ;
        RECT 58.000 475.800 58.800 480.400 ;
        RECT 63.600 471.800 64.400 480.400 ;
        RECT 68.000 471.800 68.800 480.400 ;
        RECT 73.200 472.200 74.000 480.400 ;
        RECT 76.400 471.800 77.200 480.400 ;
        RECT 80.600 475.800 81.400 480.400 ;
        RECT 83.400 475.800 84.200 480.400 ;
        RECT 87.600 471.800 88.400 480.400 ;
        RECT 89.200 475.800 90.000 480.400 ;
        RECT 92.400 475.800 93.200 480.400 ;
        RECT 95.600 472.000 96.400 480.400 ;
        RECT 101.200 475.800 102.000 480.400 ;
        RECT 104.400 475.800 105.200 480.400 ;
        RECT 110.000 471.800 110.800 480.400 ;
        RECT 118.000 471.800 118.800 480.400 ;
        RECT 122.200 475.800 123.000 480.400 ;
        RECT 125.000 475.800 125.800 480.400 ;
        RECT 129.200 471.800 130.000 480.400 ;
        RECT 132.400 472.200 133.200 480.400 ;
        RECT 137.600 471.800 138.400 480.400 ;
        RECT 142.000 471.800 142.800 480.400 ;
        RECT 147.600 475.800 148.400 480.400 ;
        RECT 150.800 475.800 151.600 480.400 ;
        RECT 156.400 472.000 157.200 480.400 ;
        RECT 159.600 475.800 160.400 480.400 ;
        RECT 162.800 475.800 163.600 480.400 ;
        RECT 164.400 475.800 165.200 480.400 ;
        RECT 167.600 475.800 168.400 480.400 ;
        RECT 172.400 471.800 173.200 480.400 ;
        RECT 174.000 471.800 174.800 480.400 ;
        RECT 180.400 475.800 181.200 480.400 ;
        RECT 183.600 475.800 184.400 480.400 ;
        RECT 185.200 475.800 186.000 480.400 ;
        RECT 188.400 475.800 189.200 480.400 ;
        RECT 191.600 475.800 192.400 480.400 ;
        RECT 194.800 475.800 195.600 480.400 ;
        RECT 202.800 475.800 203.600 480.400 ;
        RECT 206.000 475.800 206.800 480.400 ;
        RECT 212.400 475.800 213.200 480.400 ;
        RECT 215.600 475.800 216.400 480.400 ;
        RECT 218.800 475.800 219.600 480.400 ;
        RECT 222.200 479.800 223.000 480.400 ;
        RECT 222.000 473.200 223.000 479.800 ;
        RECT 228.200 473.200 229.200 480.400 ;
        RECT 231.600 475.800 232.400 480.400 ;
        RECT 234.800 475.800 235.600 480.400 ;
        RECT 238.000 475.800 238.800 480.400 ;
        RECT 241.200 475.800 242.000 480.400 ;
        RECT 249.200 475.800 250.000 480.400 ;
        RECT 252.400 475.800 253.200 480.400 ;
        RECT 258.800 475.800 259.600 480.400 ;
        RECT 262.000 475.800 262.800 480.400 ;
        RECT 265.200 475.800 266.000 480.400 ;
        RECT 212.200 471.800 213.000 472.000 ;
        RECT 215.600 471.800 216.400 472.400 ;
        RECT 258.600 471.800 259.600 472.000 ;
        RECT 262.000 471.800 262.800 472.400 ;
        RECT 271.600 471.800 272.400 480.400 ;
        RECT 275.800 475.800 276.600 480.400 ;
        RECT 279.600 475.800 280.400 480.400 ;
        RECT 281.200 471.800 282.000 480.400 ;
        RECT 284.400 471.800 285.200 480.400 ;
        RECT 287.600 471.800 288.400 480.400 ;
        RECT 290.800 471.800 291.600 480.400 ;
        RECT 294.000 471.800 294.800 480.400 ;
        RECT 295.600 471.800 296.400 480.400 ;
        RECT 301.000 475.800 301.800 480.400 ;
        RECT 305.200 471.800 306.000 480.400 ;
        RECT 306.800 471.800 307.600 480.400 ;
        RECT 311.600 471.800 312.400 480.400 ;
        RECT 316.400 475.800 317.200 480.400 ;
        RECT 319.600 475.800 320.400 480.400 ;
        RECT 324.400 473.000 325.200 480.400 ;
        RECT 327.600 475.800 328.400 480.400 ;
        RECT 330.800 475.800 331.600 480.400 ;
        RECT 332.400 475.800 333.200 480.400 ;
        RECT 335.600 475.800 336.400 480.400 ;
        RECT 337.200 471.800 338.000 480.400 ;
        RECT 341.400 475.800 342.200 480.400 ;
        RECT 343.600 475.800 344.400 480.400 ;
        RECT 346.800 475.800 347.600 480.400 ;
        RECT 348.400 471.800 349.200 480.400 ;
        RECT 351.600 471.800 352.400 480.400 ;
        RECT 353.200 475.800 354.000 480.400 ;
        RECT 356.400 475.800 357.200 480.400 ;
        RECT 359.600 471.800 360.400 480.400 ;
        RECT 361.200 475.800 362.000 480.400 ;
        RECT 364.400 475.800 365.200 480.400 ;
        RECT 366.600 475.800 367.400 480.400 ;
        RECT 370.800 471.800 371.600 480.400 ;
        RECT 372.400 475.800 373.200 480.400 ;
        RECT 375.600 475.800 376.400 480.400 ;
        RECT 377.200 475.800 378.000 480.400 ;
        RECT 380.400 475.800 381.200 480.400 ;
        RECT 383.600 475.800 384.400 480.400 ;
        RECT 390.000 475.800 390.800 480.400 ;
        RECT 393.200 475.800 394.000 480.400 ;
        RECT 401.200 475.800 402.000 480.400 ;
        RECT 404.400 475.800 405.200 480.400 ;
        RECT 407.600 475.800 408.400 480.400 ;
        RECT 410.800 475.800 411.600 480.400 ;
        RECT 412.400 475.800 413.200 480.400 ;
        RECT 421.000 475.800 421.800 480.400 ;
        RECT 380.400 471.800 381.200 472.400 ;
        RECT 383.800 471.800 384.600 472.000 ;
        RECT 425.200 471.800 426.000 480.400 ;
        RECT 426.800 475.800 427.600 480.400 ;
        RECT 430.000 475.800 430.800 480.400 ;
        RECT 432.200 475.800 433.000 480.400 ;
        RECT 436.400 471.800 437.200 480.400 ;
        RECT 438.000 471.800 438.800 480.400 ;
        RECT 442.200 475.800 443.000 480.400 ;
        RECT 444.400 475.800 445.200 480.400 ;
        RECT 447.600 475.800 448.400 480.400 ;
        RECT 450.800 475.800 451.600 480.400 ;
        RECT 454.000 475.800 454.800 480.400 ;
        RECT 462.000 475.800 462.800 480.400 ;
        RECT 465.200 475.800 466.000 480.400 ;
        RECT 471.600 475.800 472.400 480.400 ;
        RECT 474.800 475.800 475.600 480.400 ;
        RECT 478.000 475.800 478.800 480.400 ;
        RECT 479.600 475.800 480.400 480.400 ;
        RECT 482.800 475.800 483.600 480.400 ;
        RECT 486.000 475.800 486.800 480.400 ;
        RECT 492.400 475.800 493.200 480.400 ;
        RECT 495.600 475.800 496.400 480.400 ;
        RECT 503.600 475.800 504.400 480.400 ;
        RECT 506.800 475.800 507.600 480.400 ;
        RECT 510.000 475.800 510.800 480.400 ;
        RECT 513.200 475.800 514.000 480.400 ;
        RECT 515.400 475.800 516.200 480.400 ;
        RECT 471.400 471.800 472.200 472.000 ;
        RECT 474.800 471.800 475.600 472.400 ;
        RECT 5.400 471.200 32.400 471.800 ;
        RECT 189.400 471.200 216.400 471.800 ;
        RECT 235.800 471.200 262.800 471.800 ;
        RECT 380.400 471.200 407.400 471.800 ;
        RECT 5.400 471.000 6.200 471.200 ;
        RECT 189.400 471.000 190.200 471.200 ;
        RECT 235.800 471.000 236.600 471.200 ;
        RECT 406.600 471.000 407.400 471.200 ;
        RECT 448.600 471.200 475.600 471.800 ;
        RECT 482.800 471.800 483.600 472.400 ;
        RECT 486.000 471.800 487.000 472.000 ;
        RECT 519.600 471.800 520.400 480.400 ;
        RECT 521.200 471.800 522.000 480.400 ;
        RECT 525.400 475.800 526.200 480.400 ;
        RECT 527.600 475.800 528.400 480.400 ;
        RECT 530.800 475.800 531.600 480.400 ;
        RECT 532.400 475.800 533.200 480.400 ;
        RECT 535.600 475.800 536.400 480.400 ;
        RECT 538.800 475.800 539.600 480.400 ;
        RECT 542.000 475.800 542.800 480.400 ;
        RECT 550.000 475.800 550.800 480.400 ;
        RECT 553.200 475.800 554.000 480.400 ;
        RECT 559.600 475.800 560.400 480.400 ;
        RECT 562.800 475.800 563.600 480.400 ;
        RECT 566.000 475.800 566.800 480.400 ;
        RECT 559.400 471.800 560.200 472.000 ;
        RECT 562.800 471.800 563.600 472.400 ;
        RECT 570.200 471.800 571.000 480.400 ;
        RECT 578.800 471.800 579.600 480.400 ;
        RECT 583.000 475.800 583.800 480.400 ;
        RECT 585.200 475.800 586.000 480.400 ;
        RECT 588.400 475.800 589.200 480.400 ;
        RECT 590.600 475.800 591.400 480.400 ;
        RECT 594.800 471.800 595.600 480.400 ;
        RECT 598.000 472.200 598.800 480.400 ;
        RECT 601.200 475.800 602.000 480.400 ;
        RECT 604.400 475.800 605.200 480.400 ;
        RECT 606.600 475.800 607.400 480.400 ;
        RECT 610.800 471.800 611.600 480.400 ;
        RECT 612.400 475.800 613.200 480.400 ;
        RECT 615.600 475.800 616.400 480.400 ;
        RECT 617.200 475.800 618.000 480.400 ;
        RECT 620.400 475.800 621.200 480.400 ;
        RECT 623.600 473.200 624.600 480.400 ;
        RECT 629.800 479.800 630.600 480.400 ;
        RECT 629.800 473.200 630.800 479.800 ;
        RECT 634.800 472.200 635.600 480.400 ;
        RECT 640.000 471.800 640.800 480.400 ;
        RECT 644.400 472.200 645.200 480.400 ;
        RECT 649.600 471.800 650.400 480.400 ;
        RECT 653.000 475.800 653.800 480.400 ;
        RECT 657.200 471.800 658.000 480.400 ;
        RECT 660.400 471.800 661.200 480.400 ;
        RECT 666.000 475.800 666.800 480.400 ;
        RECT 669.200 475.800 670.000 480.400 ;
        RECT 674.800 472.000 675.600 480.400 ;
        RECT 679.600 473.000 680.400 480.400 ;
        RECT 482.800 471.200 509.800 471.800 ;
        RECT 448.600 471.000 449.400 471.200 ;
        RECT 509.000 471.000 509.800 471.200 ;
        RECT 536.600 471.200 563.600 471.800 ;
        RECT 536.600 471.000 537.400 471.200 ;
        RECT 231.000 450.800 231.800 451.000 ;
        RECT 296.200 450.800 297.000 451.000 ;
        RECT 231.000 450.200 258.000 450.800 ;
        RECT 2.800 441.600 3.600 450.200 ;
        RECT 8.400 441.600 9.200 446.200 ;
        RECT 11.600 441.600 12.400 446.200 ;
        RECT 17.200 441.600 18.000 450.000 ;
        RECT 20.400 441.600 21.200 450.200 ;
        RECT 24.600 441.600 25.400 446.200 ;
        RECT 27.400 441.600 28.200 446.200 ;
        RECT 31.600 441.600 32.400 450.200 ;
        RECT 33.200 441.600 34.000 450.200 ;
        RECT 37.400 441.600 38.200 446.200 ;
        RECT 39.600 441.600 40.400 446.200 ;
        RECT 42.800 441.600 43.600 446.200 ;
        RECT 44.400 441.600 45.200 450.200 ;
        RECT 48.600 441.600 49.400 446.200 ;
        RECT 51.400 441.600 52.200 446.200 ;
        RECT 55.600 441.600 56.400 450.200 ;
        RECT 58.400 441.600 59.200 450.200 ;
        RECT 63.600 441.600 64.400 449.800 ;
        RECT 67.400 441.600 68.200 446.200 ;
        RECT 71.600 441.600 72.400 450.200 ;
        RECT 73.800 441.600 74.600 446.200 ;
        RECT 78.000 441.600 78.800 450.200 ;
        RECT 81.200 441.600 82.000 450.000 ;
        RECT 86.800 441.600 87.600 446.200 ;
        RECT 90.000 441.600 90.800 446.200 ;
        RECT 95.600 441.600 96.400 450.200 ;
        RECT 98.800 441.600 99.600 450.200 ;
        RECT 103.000 441.600 103.800 446.200 ;
        RECT 105.800 441.600 106.600 446.200 ;
        RECT 110.000 441.600 110.800 450.200 ;
        RECT 118.000 441.600 118.800 450.200 ;
        RECT 123.600 441.600 124.400 446.200 ;
        RECT 126.800 441.600 127.600 446.200 ;
        RECT 132.400 441.600 133.200 450.000 ;
        RECT 137.200 441.600 138.000 446.200 ;
        RECT 140.400 441.600 141.200 449.800 ;
        RECT 145.600 441.600 146.400 450.200 ;
        RECT 148.400 441.600 149.200 450.200 ;
        RECT 152.600 441.600 153.400 446.200 ;
        RECT 156.400 441.600 157.200 449.800 ;
        RECT 161.600 441.600 162.400 450.200 ;
        RECT 164.400 441.600 165.200 450.200 ;
        RECT 169.200 441.600 170.000 450.200 ;
        RECT 173.400 441.600 174.200 446.200 ;
        RECT 177.200 441.600 178.000 450.000 ;
        RECT 182.800 441.600 183.600 446.200 ;
        RECT 186.000 441.600 186.800 446.200 ;
        RECT 191.600 441.600 192.400 450.200 ;
        RECT 194.800 441.600 195.600 450.200 ;
        RECT 201.200 441.600 202.200 448.800 ;
        RECT 207.400 442.200 208.400 448.800 ;
        RECT 207.400 441.600 208.200 442.200 ;
        RECT 212.400 441.600 213.200 445.800 ;
        RECT 215.600 441.600 216.400 446.200 ;
        RECT 217.200 441.600 218.000 450.200 ;
        RECT 253.800 450.000 254.800 450.200 ;
        RECT 257.200 449.600 258.000 450.200 ;
        RECT 270.000 450.200 297.000 450.800 ;
        RECT 397.400 450.800 398.200 451.000 ;
        RECT 467.400 450.800 468.200 451.000 ;
        RECT 526.600 450.800 527.400 451.000 ;
        RECT 397.400 450.200 424.400 450.800 ;
        RECT 270.000 449.600 270.800 450.200 ;
        RECT 273.200 450.000 274.200 450.200 ;
        RECT 221.400 441.600 222.200 446.200 ;
        RECT 223.600 441.600 224.400 446.200 ;
        RECT 226.800 441.600 227.600 446.200 ;
        RECT 230.000 441.600 230.800 446.200 ;
        RECT 233.200 441.600 234.000 446.200 ;
        RECT 236.400 441.600 237.200 446.200 ;
        RECT 244.400 441.600 245.200 446.200 ;
        RECT 247.600 441.600 248.400 446.200 ;
        RECT 254.000 441.600 254.800 446.200 ;
        RECT 257.200 441.600 258.000 446.200 ;
        RECT 260.400 441.600 261.200 446.200 ;
        RECT 266.800 441.600 267.600 446.200 ;
        RECT 270.000 441.600 270.800 446.200 ;
        RECT 273.200 441.600 274.000 446.200 ;
        RECT 279.600 441.600 280.400 446.200 ;
        RECT 282.800 441.600 283.600 446.200 ;
        RECT 290.800 441.600 291.600 446.200 ;
        RECT 294.000 441.600 294.800 446.200 ;
        RECT 297.200 441.600 298.000 446.200 ;
        RECT 300.400 441.600 301.200 446.200 ;
        RECT 302.600 441.600 303.400 446.200 ;
        RECT 306.800 441.600 307.600 450.200 ;
        RECT 311.600 441.600 312.400 449.000 ;
        RECT 318.000 441.600 318.800 450.200 ;
        RECT 321.200 441.600 322.000 445.800 ;
        RECT 324.400 441.600 325.200 446.200 ;
        RECT 326.600 441.600 327.400 446.200 ;
        RECT 330.800 441.600 331.600 450.200 ;
        RECT 333.000 441.600 333.800 446.200 ;
        RECT 337.200 441.600 338.000 450.200 ;
        RECT 338.800 441.600 339.600 450.200 ;
        RECT 343.600 441.600 344.400 450.200 ;
        RECT 350.000 441.600 350.800 450.200 ;
        RECT 351.600 441.600 352.400 450.200 ;
        RECT 358.000 441.600 358.800 450.200 ;
        RECT 361.200 441.600 362.000 446.200 ;
        RECT 364.400 441.600 365.200 445.800 ;
        RECT 367.600 441.600 368.400 446.200 ;
        RECT 370.800 441.600 371.600 445.800 ;
        RECT 374.000 441.600 374.800 446.200 ;
        RECT 375.600 441.600 376.400 450.200 ;
        RECT 420.200 450.000 421.200 450.200 ;
        RECT 423.600 449.600 424.400 450.200 ;
        RECT 441.200 450.200 468.200 450.800 ;
        RECT 500.400 450.200 527.400 450.800 ;
        RECT 565.400 450.800 566.200 451.000 ;
        RECT 639.000 450.800 639.800 451.000 ;
        RECT 565.400 450.200 592.400 450.800 ;
        RECT 639.000 450.200 666.000 450.800 ;
        RECT 441.200 449.600 442.000 450.200 ;
        RECT 444.400 450.000 445.400 450.200 ;
        RECT 380.400 441.600 381.200 446.200 ;
        RECT 383.600 441.600 384.400 445.800 ;
        RECT 386.800 441.600 387.600 446.200 ;
        RECT 390.000 441.600 390.800 445.800 ;
        RECT 393.200 441.600 394.000 446.200 ;
        RECT 396.400 441.600 397.200 446.200 ;
        RECT 399.600 441.600 400.400 446.200 ;
        RECT 402.800 441.600 403.600 446.200 ;
        RECT 410.800 441.600 411.600 446.200 ;
        RECT 414.000 441.600 414.800 446.200 ;
        RECT 420.400 441.600 421.200 446.200 ;
        RECT 423.600 441.600 424.400 446.200 ;
        RECT 426.800 441.600 427.600 446.200 ;
        RECT 433.200 441.600 434.000 446.200 ;
        RECT 436.400 441.600 437.200 446.200 ;
        RECT 438.000 441.600 438.800 446.200 ;
        RECT 441.200 441.600 442.000 446.200 ;
        RECT 444.400 441.600 445.200 446.200 ;
        RECT 450.800 441.600 451.600 446.200 ;
        RECT 454.000 441.600 454.800 446.200 ;
        RECT 462.000 441.600 462.800 446.200 ;
        RECT 465.200 441.600 466.000 446.200 ;
        RECT 468.400 441.600 469.200 446.200 ;
        RECT 471.600 441.600 472.400 446.200 ;
        RECT 473.200 441.600 474.000 446.200 ;
        RECT 476.400 441.600 477.200 446.200 ;
        RECT 479.600 441.600 480.400 446.200 ;
        RECT 481.200 441.600 482.000 450.200 ;
        RECT 485.400 441.600 486.200 446.200 ;
        RECT 489.200 441.600 490.000 446.200 ;
        RECT 490.800 441.600 491.600 450.200 ;
        RECT 500.400 449.600 501.200 450.200 ;
        RECT 503.800 450.000 504.600 450.200 ;
        RECT 494.000 441.600 494.800 449.000 ;
        RECT 497.200 441.600 498.000 446.200 ;
        RECT 500.400 441.600 501.200 446.200 ;
        RECT 503.600 441.600 504.400 446.200 ;
        RECT 510.000 441.600 510.800 446.200 ;
        RECT 513.200 441.600 514.000 446.200 ;
        RECT 521.200 441.600 522.000 446.200 ;
        RECT 524.400 441.600 525.200 446.200 ;
        RECT 527.600 441.600 528.400 446.200 ;
        RECT 530.800 441.600 531.600 446.200 ;
        RECT 533.000 441.600 533.800 446.200 ;
        RECT 537.200 441.600 538.000 450.200 ;
        RECT 540.400 441.600 541.200 446.200 ;
        RECT 542.000 441.600 542.800 446.200 ;
        RECT 545.200 441.600 546.000 446.200 ;
        RECT 546.800 441.600 547.600 446.200 ;
        RECT 550.000 441.600 550.800 446.200 ;
        RECT 551.600 441.600 552.400 450.200 ;
        RECT 588.200 450.000 589.200 450.200 ;
        RECT 591.600 449.600 592.400 450.200 ;
        RECT 561.200 441.600 562.000 446.200 ;
        RECT 564.400 441.600 565.200 446.200 ;
        RECT 567.600 441.600 568.400 446.200 ;
        RECT 570.800 441.600 571.600 446.200 ;
        RECT 578.800 441.600 579.600 446.200 ;
        RECT 582.000 441.600 582.800 446.200 ;
        RECT 588.400 441.600 589.200 446.200 ;
        RECT 591.600 441.600 592.400 446.200 ;
        RECT 594.800 441.600 595.600 446.200 ;
        RECT 597.000 441.600 597.800 446.200 ;
        RECT 601.200 441.600 602.000 450.200 ;
        RECT 604.400 441.600 605.200 449.000 ;
        RECT 607.600 441.600 608.400 450.200 ;
        RECT 612.400 441.600 613.200 449.000 ;
        RECT 615.600 441.600 616.400 450.200 ;
        RECT 623.600 441.600 624.400 450.200 ;
        RECT 661.800 450.000 662.600 450.200 ;
        RECT 665.200 449.600 666.000 450.200 ;
        RECT 625.200 441.600 626.000 446.200 ;
        RECT 630.000 441.600 630.800 445.800 ;
        RECT 633.200 441.600 634.000 446.200 ;
        RECT 634.800 441.600 635.600 446.200 ;
        RECT 638.000 441.600 638.800 446.200 ;
        RECT 641.200 441.600 642.000 446.200 ;
        RECT 644.400 441.600 645.200 446.200 ;
        RECT 652.400 441.600 653.200 446.200 ;
        RECT 655.600 441.600 656.400 446.200 ;
        RECT 662.000 441.600 662.800 446.200 ;
        RECT 665.200 441.600 666.000 446.200 ;
        RECT 668.400 441.600 669.200 446.200 ;
        RECT 670.000 441.600 670.800 450.200 ;
        RECT 673.200 441.600 674.000 450.200 ;
        RECT 676.400 441.600 677.200 450.200 ;
        RECT 679.600 441.600 680.400 450.200 ;
        RECT 682.800 441.600 683.600 450.200 ;
        RECT 0.400 440.400 689.200 441.600 ;
        RECT 2.800 431.800 3.600 440.400 ;
        RECT 8.400 435.800 9.200 440.400 ;
        RECT 11.600 435.800 12.400 440.400 ;
        RECT 17.200 432.000 18.000 440.400 ;
        RECT 20.400 431.800 21.200 440.400 ;
        RECT 24.600 435.800 25.400 440.400 ;
        RECT 27.400 435.800 28.200 440.400 ;
        RECT 31.600 431.800 32.400 440.400 ;
        RECT 34.400 431.800 35.200 440.400 ;
        RECT 39.600 432.200 40.400 440.400 ;
        RECT 43.400 435.800 44.200 440.400 ;
        RECT 47.600 431.800 48.400 440.400 ;
        RECT 49.200 431.800 50.000 440.400 ;
        RECT 52.400 433.000 53.200 440.400 ;
        RECT 57.200 432.200 58.000 440.400 ;
        RECT 62.400 431.800 63.200 440.400 ;
        RECT 66.400 431.800 67.200 440.400 ;
        RECT 71.600 432.200 72.400 440.400 ;
        RECT 74.800 431.800 75.600 440.400 ;
        RECT 79.000 435.800 79.800 440.400 ;
        RECT 81.800 435.800 82.600 440.400 ;
        RECT 86.000 431.800 86.800 440.400 ;
        RECT 89.200 431.800 90.000 440.400 ;
        RECT 94.800 435.800 95.600 440.400 ;
        RECT 98.000 435.800 98.800 440.400 ;
        RECT 103.600 432.000 104.400 440.400 ;
        RECT 112.800 431.800 113.600 440.400 ;
        RECT 118.000 432.200 118.800 440.400 ;
        RECT 122.800 433.000 123.600 440.400 ;
        RECT 126.000 431.800 126.800 440.400 ;
        RECT 127.600 431.800 128.400 440.400 ;
        RECT 130.800 433.000 131.600 440.400 ;
        RECT 135.600 433.000 136.400 440.400 ;
        RECT 138.800 431.800 139.600 440.400 ;
        RECT 142.000 431.800 142.800 440.400 ;
        RECT 147.600 435.800 148.400 440.400 ;
        RECT 150.800 435.800 151.600 440.400 ;
        RECT 156.400 432.000 157.200 440.400 ;
        RECT 160.200 435.800 161.000 440.400 ;
        RECT 164.400 431.800 165.200 440.400 ;
        RECT 166.600 435.800 167.400 440.400 ;
        RECT 170.800 431.800 171.600 440.400 ;
        RECT 174.000 432.200 174.800 440.400 ;
        RECT 179.200 431.800 180.000 440.400 ;
        RECT 182.600 435.800 183.400 440.400 ;
        RECT 186.800 431.800 187.600 440.400 ;
        RECT 190.000 433.000 190.800 440.400 ;
        RECT 193.200 431.800 194.000 440.400 ;
        RECT 196.400 431.800 197.200 440.400 ;
        RECT 202.000 435.800 202.800 440.400 ;
        RECT 205.200 435.800 206.000 440.400 ;
        RECT 210.800 432.000 211.600 440.400 ;
        RECT 214.000 431.800 214.800 440.400 ;
        RECT 220.400 435.800 221.200 440.400 ;
        RECT 225.200 433.000 226.000 440.400 ;
        RECT 230.600 431.800 231.400 440.400 ;
        RECT 238.000 431.800 238.800 440.400 ;
        RECT 239.600 435.800 240.400 440.400 ;
        RECT 242.800 435.800 243.600 440.400 ;
        RECT 246.000 435.800 246.800 440.400 ;
        RECT 249.200 435.800 250.000 440.400 ;
        RECT 257.200 435.800 258.000 440.400 ;
        RECT 260.400 435.800 261.200 440.400 ;
        RECT 266.800 435.800 267.600 440.400 ;
        RECT 270.000 435.800 270.800 440.400 ;
        RECT 273.200 435.800 274.000 440.400 ;
        RECT 279.600 435.800 280.400 440.400 ;
        RECT 282.800 435.800 283.600 440.400 ;
        RECT 266.600 431.800 267.600 432.000 ;
        RECT 270.000 431.800 270.800 432.400 ;
        RECT 284.400 431.800 285.200 440.400 ;
        RECT 287.600 431.800 288.400 440.400 ;
        RECT 290.800 431.800 291.600 440.400 ;
        RECT 294.000 431.800 294.800 440.400 ;
        RECT 297.200 431.800 298.000 440.400 ;
        RECT 298.800 431.800 299.600 440.400 ;
        RECT 303.000 435.800 303.800 440.400 ;
        RECT 305.800 435.800 306.600 440.400 ;
        RECT 310.000 431.800 310.800 440.400 ;
        RECT 313.200 435.800 314.000 440.400 ;
        RECT 314.800 431.800 315.600 440.400 ;
        RECT 322.800 431.800 323.600 440.400 ;
        RECT 324.400 435.800 325.200 440.400 ;
        RECT 327.600 435.800 328.400 440.400 ;
        RECT 329.200 435.800 330.000 440.400 ;
        RECT 332.400 435.800 333.200 440.400 ;
        RECT 334.000 431.800 334.800 440.400 ;
        RECT 337.200 431.800 338.000 440.400 ;
        RECT 341.400 435.800 342.200 440.400 ;
        RECT 343.600 431.800 344.400 440.400 ;
        RECT 350.000 431.800 350.800 440.400 ;
        RECT 353.200 435.800 354.000 440.400 ;
        RECT 354.800 431.800 355.600 440.400 ;
        RECT 361.200 431.800 362.000 440.400 ;
        RECT 364.400 436.200 365.200 440.400 ;
        RECT 367.600 435.800 368.400 440.400 ;
        RECT 370.800 435.800 371.600 440.400 ;
        RECT 374.000 436.200 374.800 440.400 ;
        RECT 377.200 435.800 378.000 440.400 ;
        RECT 380.400 432.200 381.200 440.400 ;
        RECT 383.600 435.800 384.400 440.400 ;
        RECT 386.800 433.000 387.600 440.400 ;
        RECT 390.600 435.800 391.400 440.400 ;
        RECT 394.800 431.800 395.600 440.400 ;
        RECT 396.400 435.800 397.200 440.400 ;
        RECT 399.600 435.800 400.400 440.400 ;
        RECT 406.000 435.800 406.800 440.400 ;
        RECT 409.200 435.800 410.000 440.400 ;
        RECT 412.400 435.800 413.200 440.400 ;
        RECT 418.800 435.800 419.600 440.400 ;
        RECT 422.000 435.800 422.800 440.400 ;
        RECT 430.000 435.800 430.800 440.400 ;
        RECT 433.200 435.800 434.000 440.400 ;
        RECT 436.400 435.800 437.200 440.400 ;
        RECT 439.600 435.800 440.400 440.400 ;
        RECT 442.800 435.800 443.600 440.400 ;
        RECT 409.200 431.800 410.000 432.400 ;
        RECT 412.400 431.800 413.400 432.000 ;
        RECT 444.400 431.800 445.200 440.400 ;
        RECT 447.600 433.000 448.400 440.400 ;
        RECT 450.800 431.800 451.600 440.400 ;
        RECT 454.000 431.800 454.800 440.400 ;
        RECT 457.200 431.800 458.000 440.400 ;
        RECT 460.400 431.800 461.200 440.400 ;
        RECT 463.600 431.800 464.400 440.400 ;
        RECT 465.200 435.800 466.000 440.400 ;
        RECT 468.400 435.800 469.200 440.400 ;
        RECT 471.600 435.800 472.400 440.400 ;
        RECT 478.000 435.800 478.800 440.400 ;
        RECT 481.200 435.800 482.000 440.400 ;
        RECT 489.200 435.800 490.000 440.400 ;
        RECT 492.400 435.800 493.200 440.400 ;
        RECT 495.600 435.800 496.400 440.400 ;
        RECT 498.800 435.800 499.600 440.400 ;
        RECT 501.000 435.800 501.800 440.400 ;
        RECT 468.400 431.800 469.200 432.400 ;
        RECT 471.800 431.800 472.600 432.000 ;
        RECT 505.200 431.800 506.000 440.400 ;
        RECT 506.800 431.800 507.600 440.400 ;
        RECT 510.000 431.800 510.800 440.400 ;
        RECT 513.200 431.800 514.000 440.400 ;
        RECT 516.400 431.800 517.200 440.400 ;
        RECT 519.600 431.800 520.400 440.400 ;
        RECT 521.200 431.800 522.000 440.400 ;
        RECT 524.400 433.000 525.200 440.400 ;
        RECT 527.600 431.800 528.400 440.400 ;
        RECT 531.800 435.800 532.600 440.400 ;
        RECT 536.600 431.800 537.400 440.400 ;
        RECT 542.000 433.000 542.800 440.400 ;
        RECT 545.200 431.800 546.000 440.400 ;
        RECT 547.400 435.800 548.200 440.400 ;
        RECT 551.600 431.800 552.400 440.400 ;
        RECT 553.200 435.800 554.000 440.400 ;
        RECT 556.400 435.800 557.200 440.400 ;
        RECT 559.600 435.800 560.400 440.400 ;
        RECT 562.800 435.800 563.600 440.400 ;
        RECT 570.800 435.800 571.600 440.400 ;
        RECT 574.000 435.800 574.800 440.400 ;
        RECT 580.400 435.800 581.200 440.400 ;
        RECT 583.600 435.800 584.400 440.400 ;
        RECT 586.800 435.800 587.600 440.400 ;
        RECT 594.800 433.000 595.600 440.400 ;
        RECT 598.000 431.800 598.800 440.400 ;
        RECT 599.600 435.800 600.400 440.400 ;
        RECT 602.800 435.800 603.600 440.400 ;
        RECT 606.000 435.800 606.800 440.400 ;
        RECT 609.200 435.800 610.000 440.400 ;
        RECT 617.200 435.800 618.000 440.400 ;
        RECT 620.400 435.800 621.200 440.400 ;
        RECT 626.800 435.800 627.600 440.400 ;
        RECT 630.000 435.800 630.800 440.400 ;
        RECT 633.200 435.800 634.000 440.400 ;
        RECT 626.600 431.800 627.400 432.000 ;
        RECT 630.000 431.800 630.800 432.400 ;
        RECT 634.800 431.800 635.600 440.400 ;
        RECT 638.000 431.800 638.800 440.400 ;
        RECT 641.200 431.800 642.000 440.400 ;
        RECT 644.400 431.800 645.200 440.400 ;
        RECT 647.600 431.800 648.400 440.400 ;
        RECT 649.200 435.800 650.000 440.400 ;
        RECT 652.400 435.800 653.200 440.400 ;
        RECT 655.600 435.800 656.400 440.400 ;
        RECT 658.800 435.800 659.600 440.400 ;
        RECT 666.800 435.800 667.600 440.400 ;
        RECT 670.000 435.800 670.800 440.400 ;
        RECT 676.400 435.800 677.200 440.400 ;
        RECT 679.600 435.800 680.400 440.400 ;
        RECT 682.800 435.800 683.600 440.400 ;
        RECT 676.200 431.800 677.200 432.000 ;
        RECT 679.600 431.800 680.400 432.400 ;
        RECT 243.800 431.200 270.800 431.800 ;
        RECT 409.200 431.200 436.200 431.800 ;
        RECT 468.400 431.200 495.400 431.800 ;
        RECT 243.800 431.000 244.600 431.200 ;
        RECT 435.400 431.000 436.200 431.200 ;
        RECT 494.600 431.000 495.400 431.200 ;
        RECT 603.800 431.200 630.800 431.800 ;
        RECT 653.400 431.200 680.400 431.800 ;
        RECT 603.800 431.000 604.600 431.200 ;
        RECT 653.400 431.000 654.200 431.200 ;
        RECT 562.800 430.000 586.200 430.600 ;
        RECT 562.800 429.400 563.600 430.000 ;
        RECT 580.400 429.600 581.200 430.000 ;
        RECT 585.400 429.800 586.200 430.000 ;
        RECT 266.600 412.000 267.400 412.200 ;
        RECT 271.600 412.000 272.400 412.400 ;
        RECT 278.000 412.000 278.800 412.400 ;
        RECT 289.200 412.000 290.000 412.600 ;
        RECT 266.600 411.400 290.000 412.000 ;
        RECT 195.800 410.800 196.600 411.000 ;
        RECT 419.800 410.800 420.600 411.000 ;
        RECT 480.200 410.800 481.000 411.000 ;
        RECT 195.800 410.200 222.800 410.800 ;
        RECT 419.800 410.200 446.800 410.800 ;
        RECT 2.800 401.600 3.600 410.000 ;
        RECT 8.400 401.600 9.200 406.200 ;
        RECT 11.600 401.600 12.400 406.200 ;
        RECT 17.200 401.600 18.000 410.200 ;
        RECT 20.400 401.600 21.200 410.200 ;
        RECT 24.600 401.600 25.400 406.200 ;
        RECT 28.000 401.600 28.800 410.200 ;
        RECT 33.200 401.600 34.000 409.800 ;
        RECT 38.000 401.600 38.800 409.000 ;
        RECT 41.200 401.600 42.000 410.200 ;
        RECT 42.800 401.600 43.600 410.200 ;
        RECT 47.000 401.600 47.800 406.200 ;
        RECT 49.800 401.600 50.600 406.200 ;
        RECT 54.000 401.600 54.800 410.200 ;
        RECT 56.800 401.600 57.600 410.200 ;
        RECT 62.000 401.600 62.800 409.800 ;
        RECT 65.200 401.600 66.000 406.200 ;
        RECT 70.000 401.600 70.800 410.200 ;
        RECT 75.600 401.600 76.400 406.200 ;
        RECT 78.800 401.600 79.600 406.200 ;
        RECT 84.400 401.600 85.200 410.000 ;
        RECT 87.600 401.600 88.400 406.200 ;
        RECT 90.800 401.600 91.600 406.200 ;
        RECT 94.000 401.600 94.800 405.800 ;
        RECT 98.800 401.600 99.600 410.000 ;
        RECT 104.400 401.600 105.200 406.200 ;
        RECT 107.600 401.600 108.400 406.200 ;
        RECT 113.200 401.600 114.000 410.200 ;
        RECT 121.800 401.600 122.600 406.200 ;
        RECT 126.000 401.600 126.800 410.200 ;
        RECT 127.600 401.600 128.400 406.200 ;
        RECT 130.800 401.600 131.600 405.800 ;
        RECT 135.600 401.600 136.400 409.800 ;
        RECT 140.800 401.600 141.600 410.200 ;
        RECT 145.200 401.600 146.000 406.200 ;
        RECT 148.400 401.600 149.200 405.800 ;
        RECT 151.600 401.600 152.400 406.200 ;
        RECT 154.800 401.600 155.600 406.200 ;
        RECT 158.000 401.600 158.800 409.000 ;
        RECT 161.200 401.600 162.000 410.200 ;
        RECT 162.800 401.600 163.600 410.200 ;
        RECT 167.000 401.600 167.800 406.200 ;
        RECT 170.800 401.600 171.600 409.800 ;
        RECT 176.000 401.600 176.800 410.200 ;
        RECT 178.800 401.600 179.600 410.200 ;
        RECT 183.000 401.600 183.800 406.200 ;
        RECT 185.800 401.600 186.600 406.200 ;
        RECT 190.000 401.600 190.800 410.200 ;
        RECT 218.600 410.000 219.600 410.200 ;
        RECT 222.000 409.600 222.800 410.200 ;
        RECT 191.600 401.600 192.400 406.200 ;
        RECT 194.800 401.600 195.600 406.200 ;
        RECT 198.000 401.600 198.800 406.200 ;
        RECT 201.200 401.600 202.000 406.200 ;
        RECT 209.200 401.600 210.000 406.200 ;
        RECT 212.400 401.600 213.200 406.200 ;
        RECT 218.800 401.600 219.600 406.200 ;
        RECT 222.000 401.600 222.800 406.200 ;
        RECT 225.200 401.600 226.000 406.200 ;
        RECT 226.800 401.600 227.600 406.200 ;
        RECT 230.000 401.600 230.800 406.200 ;
        RECT 231.600 401.600 232.400 406.200 ;
        RECT 234.800 401.600 235.600 406.200 ;
        RECT 236.400 401.600 237.200 406.200 ;
        RECT 239.600 401.600 240.400 409.800 ;
        RECT 242.800 401.600 243.600 410.200 ;
        RECT 247.000 401.600 247.800 406.200 ;
        RECT 249.200 401.600 250.000 406.200 ;
        RECT 252.400 401.600 253.200 406.200 ;
        RECT 254.600 401.600 255.400 406.200 ;
        RECT 258.800 401.600 259.600 410.200 ;
        RECT 265.200 401.600 266.000 406.200 ;
        RECT 268.400 401.600 269.200 406.200 ;
        RECT 271.600 401.600 272.400 406.200 ;
        RECT 278.000 401.600 278.800 406.400 ;
        RECT 281.200 401.600 282.000 406.200 ;
        RECT 289.200 401.600 290.000 406.200 ;
        RECT 292.400 401.600 293.200 406.200 ;
        RECT 295.600 401.600 296.400 406.200 ;
        RECT 298.800 401.600 299.600 406.200 ;
        RECT 300.400 401.600 301.200 406.200 ;
        RECT 303.600 401.600 304.400 406.200 ;
        RECT 306.800 401.600 307.600 406.200 ;
        RECT 308.400 401.600 309.200 406.200 ;
        RECT 311.600 401.600 312.400 406.200 ;
        RECT 316.400 401.600 317.200 410.200 ;
        RECT 321.200 401.600 322.000 410.200 ;
        RECT 323.400 401.600 324.200 406.200 ;
        RECT 327.600 401.600 328.400 410.200 ;
        RECT 332.400 401.600 333.200 409.000 ;
        RECT 335.600 401.600 336.400 406.200 ;
        RECT 338.800 401.600 339.600 406.200 ;
        RECT 341.000 401.600 341.800 406.200 ;
        RECT 345.200 401.600 346.000 410.200 ;
        RECT 350.000 401.600 350.800 409.000 ;
        RECT 353.200 401.600 354.000 410.200 ;
        RECT 358.000 401.600 358.800 406.200 ;
        RECT 361.200 401.600 362.000 406.200 ;
        RECT 364.400 401.600 365.200 405.800 ;
        RECT 367.600 401.600 368.400 406.200 ;
        RECT 369.200 401.600 370.000 406.200 ;
        RECT 372.400 401.600 373.200 405.800 ;
        RECT 377.200 401.600 378.000 405.800 ;
        RECT 380.400 401.600 381.200 406.200 ;
        RECT 383.600 401.600 384.400 410.200 ;
        RECT 390.000 401.600 390.800 409.000 ;
        RECT 393.200 401.600 394.000 406.200 ;
        RECT 396.400 401.600 397.200 405.800 ;
        RECT 402.800 401.600 403.600 409.000 ;
        RECT 409.200 401.600 410.000 410.200 ;
        RECT 442.600 410.000 443.600 410.200 ;
        RECT 446.000 409.600 446.800 410.200 ;
        RECT 454.000 410.200 481.000 410.800 ;
        RECT 512.600 410.800 513.400 411.000 ;
        RECT 581.400 410.800 582.200 411.000 ;
        RECT 653.400 410.800 654.200 411.000 ;
        RECT 512.600 410.200 539.600 410.800 ;
        RECT 581.400 410.200 608.400 410.800 ;
        RECT 653.400 410.200 680.400 410.800 ;
        RECT 454.000 409.600 454.800 410.200 ;
        RECT 457.400 410.000 458.200 410.200 ;
        RECT 415.600 401.600 416.400 406.200 ;
        RECT 418.800 401.600 419.600 406.200 ;
        RECT 422.000 401.600 422.800 406.200 ;
        RECT 425.200 401.600 426.000 406.200 ;
        RECT 433.200 401.600 434.000 406.200 ;
        RECT 436.400 401.600 437.200 406.200 ;
        RECT 442.800 401.600 443.600 406.200 ;
        RECT 446.000 401.600 446.800 406.200 ;
        RECT 449.200 401.600 450.000 406.200 ;
        RECT 450.800 401.600 451.600 406.200 ;
        RECT 454.000 401.600 454.800 406.200 ;
        RECT 457.200 401.600 458.000 406.200 ;
        RECT 463.600 401.600 464.400 406.200 ;
        RECT 466.800 401.600 467.600 406.200 ;
        RECT 474.800 401.600 475.600 406.200 ;
        RECT 478.000 401.600 478.800 406.200 ;
        RECT 481.200 401.600 482.000 406.200 ;
        RECT 484.400 401.600 485.200 406.200 ;
        RECT 486.000 401.600 486.800 410.200 ;
        RECT 490.200 401.600 491.000 406.200 ;
        RECT 493.000 401.600 493.800 406.200 ;
        RECT 497.200 401.600 498.000 410.200 ;
        RECT 500.400 401.600 501.200 406.200 ;
        RECT 502.000 401.600 502.800 410.200 ;
        RECT 535.400 410.000 536.200 410.200 ;
        RECT 538.800 409.600 539.600 410.200 ;
        RECT 506.200 401.600 507.000 406.200 ;
        RECT 508.400 401.600 509.200 406.200 ;
        RECT 511.600 401.600 512.400 406.200 ;
        RECT 514.800 401.600 515.600 406.200 ;
        RECT 518.000 401.600 518.800 406.200 ;
        RECT 526.000 401.600 526.800 406.200 ;
        RECT 529.200 401.600 530.000 406.200 ;
        RECT 535.600 401.600 536.400 406.200 ;
        RECT 538.800 401.600 539.600 406.200 ;
        RECT 542.000 401.600 542.800 406.200 ;
        RECT 543.600 401.600 544.400 410.200 ;
        RECT 546.800 401.600 547.600 409.000 ;
        RECT 550.000 401.600 550.800 410.200 ;
        RECT 554.200 401.600 555.000 406.200 ;
        RECT 558.000 401.600 558.800 406.200 ;
        RECT 560.200 401.600 561.000 406.200 ;
        RECT 564.400 401.600 565.200 410.200 ;
        RECT 566.000 401.600 566.800 410.200 ;
        RECT 604.200 410.000 605.200 410.200 ;
        RECT 607.600 409.600 608.400 410.200 ;
        RECT 570.200 401.600 571.000 406.200 ;
        RECT 577.200 401.600 578.000 406.200 ;
        RECT 580.400 401.600 581.200 406.200 ;
        RECT 583.600 401.600 584.400 406.200 ;
        RECT 586.800 401.600 587.600 406.200 ;
        RECT 594.800 401.600 595.600 406.200 ;
        RECT 598.000 401.600 598.800 406.200 ;
        RECT 604.400 401.600 605.200 406.200 ;
        RECT 607.600 401.600 608.400 406.200 ;
        RECT 610.800 401.600 611.600 406.200 ;
        RECT 614.000 402.200 615.000 408.800 ;
        RECT 614.200 401.600 615.000 402.200 ;
        RECT 620.200 401.600 621.200 408.800 ;
        RECT 623.600 401.600 624.400 406.200 ;
        RECT 626.800 401.600 627.600 406.200 ;
        RECT 628.400 401.600 629.200 410.200 ;
        RECT 631.600 401.600 632.400 410.200 ;
        RECT 676.200 410.000 677.200 410.200 ;
        RECT 679.600 409.600 680.400 410.200 ;
        RECT 635.800 401.600 636.600 406.200 ;
        RECT 639.600 402.200 640.600 408.800 ;
        RECT 639.800 401.600 640.600 402.200 ;
        RECT 645.800 401.600 646.800 408.800 ;
        RECT 649.200 401.600 650.000 406.200 ;
        RECT 652.400 401.600 653.200 406.200 ;
        RECT 655.600 401.600 656.400 406.200 ;
        RECT 658.800 401.600 659.600 406.200 ;
        RECT 666.800 401.600 667.600 406.200 ;
        RECT 670.000 401.600 670.800 406.200 ;
        RECT 676.400 401.600 677.200 406.200 ;
        RECT 679.600 401.600 680.400 406.200 ;
        RECT 682.800 401.600 683.600 406.200 ;
        RECT 0.400 400.400 689.200 401.600 ;
        RECT 2.800 393.000 3.600 400.400 ;
        RECT 7.600 392.000 8.400 400.400 ;
        RECT 13.200 395.800 14.000 400.400 ;
        RECT 16.400 395.800 17.200 400.400 ;
        RECT 22.000 391.800 22.800 400.400 ;
        RECT 25.800 395.800 26.600 400.400 ;
        RECT 30.000 391.800 30.800 400.400 ;
        RECT 31.600 391.800 32.400 400.400 ;
        RECT 34.800 393.000 35.600 400.400 ;
        RECT 38.000 391.800 38.800 400.400 ;
        RECT 42.200 395.800 43.000 400.400 ;
        RECT 45.000 395.800 45.800 400.400 ;
        RECT 49.200 391.800 50.000 400.400 ;
        RECT 52.000 391.800 52.800 400.400 ;
        RECT 57.200 392.200 58.000 400.400 ;
        RECT 61.600 391.800 62.400 400.400 ;
        RECT 66.800 392.200 67.600 400.400 ;
        RECT 70.000 395.800 70.800 400.400 ;
        RECT 73.200 391.800 74.000 400.400 ;
        RECT 76.400 393.000 77.200 400.400 ;
        RECT 79.600 395.800 80.400 400.400 ;
        RECT 82.800 395.800 83.600 400.400 ;
        RECT 86.000 393.000 86.800 400.400 ;
        RECT 89.200 391.800 90.000 400.400 ;
        RECT 91.400 395.800 92.200 400.400 ;
        RECT 95.600 391.800 96.400 400.400 ;
        RECT 97.200 391.800 98.000 400.400 ;
        RECT 100.400 393.000 101.200 400.400 ;
        RECT 103.600 391.800 104.400 400.400 ;
        RECT 107.800 395.800 108.600 400.400 ;
        RECT 114.800 391.800 115.600 400.400 ;
        RECT 119.600 391.800 120.400 400.400 ;
        RECT 123.800 395.800 124.600 400.400 ;
        RECT 126.600 395.800 127.400 400.400 ;
        RECT 130.800 391.800 131.600 400.400 ;
        RECT 134.000 396.200 134.800 400.400 ;
        RECT 137.200 395.800 138.000 400.400 ;
        RECT 139.400 395.800 140.200 400.400 ;
        RECT 143.600 391.800 144.400 400.400 ;
        RECT 145.200 395.800 146.000 400.400 ;
        RECT 148.400 395.800 149.200 400.400 ;
        RECT 150.600 395.800 151.400 400.400 ;
        RECT 154.800 391.800 155.600 400.400 ;
        RECT 158.000 392.200 158.800 400.400 ;
        RECT 163.200 391.800 164.000 400.400 ;
        RECT 166.000 391.800 166.800 400.400 ;
        RECT 170.200 395.800 171.000 400.400 ;
        RECT 173.000 395.800 173.800 400.400 ;
        RECT 177.200 391.800 178.000 400.400 ;
        RECT 180.400 392.200 181.200 400.400 ;
        RECT 185.600 391.800 186.400 400.400 ;
        RECT 188.400 391.800 189.200 400.400 ;
        RECT 192.600 395.800 193.400 400.400 ;
        RECT 194.800 391.800 195.600 400.400 ;
        RECT 199.000 395.800 199.800 400.400 ;
        RECT 202.800 391.800 203.600 400.400 ;
        RECT 208.400 395.800 209.200 400.400 ;
        RECT 211.600 395.800 212.400 400.400 ;
        RECT 217.200 392.000 218.000 400.400 ;
        RECT 222.200 399.800 223.000 400.400 ;
        RECT 222.000 393.200 223.000 399.800 ;
        RECT 228.200 393.200 229.200 400.400 ;
        RECT 233.200 392.200 234.000 400.400 ;
        RECT 238.400 391.800 239.200 400.400 ;
        RECT 242.800 392.200 243.600 400.400 ;
        RECT 248.000 391.800 248.800 400.400 ;
        RECT 252.400 393.000 253.200 400.400 ;
        RECT 255.600 391.800 256.400 400.400 ;
        RECT 257.200 391.800 258.000 400.400 ;
        RECT 260.400 391.800 261.200 400.400 ;
        RECT 263.600 391.800 264.400 400.400 ;
        RECT 271.200 391.800 272.000 400.400 ;
        RECT 276.400 392.200 277.200 400.400 ;
        RECT 279.600 395.800 280.400 400.400 ;
        RECT 282.800 395.800 283.600 400.400 ;
        RECT 286.000 395.800 286.800 400.400 ;
        RECT 292.400 395.800 293.200 400.400 ;
        RECT 295.600 395.800 296.400 400.400 ;
        RECT 303.600 395.800 304.400 400.400 ;
        RECT 306.800 395.800 307.600 400.400 ;
        RECT 310.000 395.800 310.800 400.400 ;
        RECT 313.200 395.800 314.000 400.400 ;
        RECT 314.800 395.800 315.600 400.400 ;
        RECT 318.000 395.800 318.800 400.400 ;
        RECT 282.800 391.800 283.600 392.400 ;
        RECT 286.000 391.800 287.000 392.000 ;
        RECT 319.600 391.800 320.400 400.400 ;
        RECT 323.800 395.800 324.600 400.400 ;
        RECT 326.000 395.800 326.800 400.400 ;
        RECT 329.200 395.800 330.000 400.400 ;
        RECT 331.400 395.800 332.200 400.400 ;
        RECT 335.600 391.800 336.400 400.400 ;
        RECT 337.800 395.800 338.600 400.400 ;
        RECT 342.000 391.800 342.800 400.400 ;
        RECT 346.800 393.000 347.600 400.400 ;
        RECT 350.000 391.800 350.800 400.400 ;
        RECT 356.400 391.800 357.200 400.400 ;
        RECT 358.000 391.800 358.800 400.400 ;
        RECT 366.000 393.000 366.800 400.400 ;
        RECT 369.200 395.800 370.000 400.400 ;
        RECT 372.400 395.800 373.200 400.400 ;
        RECT 374.000 395.800 374.800 400.400 ;
        RECT 377.200 396.200 378.000 400.400 ;
        RECT 380.400 395.800 381.200 400.400 ;
        RECT 383.600 395.800 384.400 400.400 ;
        RECT 385.200 395.800 386.000 400.400 ;
        RECT 388.400 395.800 389.200 400.400 ;
        RECT 391.600 395.800 392.400 400.400 ;
        RECT 398.000 395.800 398.800 400.400 ;
        RECT 401.200 395.800 402.000 400.400 ;
        RECT 409.200 395.800 410.000 400.400 ;
        RECT 412.400 395.800 413.200 400.400 ;
        RECT 415.600 395.800 416.400 400.400 ;
        RECT 418.800 395.800 419.600 400.400 ;
        RECT 388.400 391.800 389.200 392.400 ;
        RECT 426.800 392.200 427.600 400.400 ;
        RECT 391.800 391.800 392.600 392.000 ;
        RECT 432.000 391.800 432.800 400.400 ;
        RECT 434.800 391.800 435.600 400.400 ;
        RECT 438.000 393.000 438.800 400.400 ;
        RECT 441.200 391.800 442.000 400.400 ;
        RECT 445.400 395.800 446.200 400.400 ;
        RECT 447.600 395.800 448.400 400.400 ;
        RECT 450.800 395.800 451.600 400.400 ;
        RECT 454.000 395.800 454.800 400.400 ;
        RECT 457.200 395.800 458.000 400.400 ;
        RECT 465.200 395.800 466.000 400.400 ;
        RECT 468.400 395.800 469.200 400.400 ;
        RECT 474.800 395.800 475.600 400.400 ;
        RECT 478.000 395.800 478.800 400.400 ;
        RECT 481.200 395.800 482.000 400.400 ;
        RECT 482.800 395.800 483.600 400.400 ;
        RECT 486.000 395.800 486.800 400.400 ;
        RECT 487.600 395.800 488.400 400.400 ;
        RECT 490.800 395.800 491.600 400.400 ;
        RECT 474.600 391.800 475.400 392.000 ;
        RECT 478.000 391.800 478.800 392.400 ;
        RECT 492.400 391.800 493.200 400.400 ;
        RECT 495.600 391.800 496.400 400.400 ;
        RECT 498.800 391.800 499.600 400.400 ;
        RECT 500.400 395.800 501.200 400.400 ;
        RECT 503.600 395.800 504.400 400.400 ;
        RECT 505.800 395.800 506.600 400.400 ;
        RECT 510.000 391.800 510.800 400.400 ;
        RECT 512.200 395.800 513.000 400.400 ;
        RECT 516.400 391.800 517.200 400.400 ;
        RECT 518.600 395.800 519.400 400.400 ;
        RECT 522.800 391.800 523.600 400.400 ;
        RECT 524.400 391.800 525.200 400.400 ;
        RECT 527.600 393.000 528.400 400.400 ;
        RECT 530.800 395.800 531.600 400.400 ;
        RECT 534.000 395.800 534.800 400.400 ;
        RECT 535.600 391.800 536.400 400.400 ;
        RECT 539.800 395.800 540.600 400.400 ;
        RECT 542.600 395.800 543.400 400.400 ;
        RECT 546.800 391.800 547.600 400.400 ;
        RECT 550.000 392.000 550.800 400.400 ;
        RECT 555.600 395.800 556.400 400.400 ;
        RECT 558.800 395.800 559.600 400.400 ;
        RECT 564.400 391.800 565.200 400.400 ;
        RECT 569.200 395.800 570.000 400.400 ;
        RECT 575.600 395.800 576.400 400.400 ;
        RECT 578.800 395.800 579.600 400.400 ;
        RECT 581.000 395.800 581.800 400.400 ;
        RECT 585.200 391.800 586.000 400.400 ;
        RECT 588.400 392.000 589.200 400.400 ;
        RECT 594.000 395.800 594.800 400.400 ;
        RECT 597.200 395.800 598.000 400.400 ;
        RECT 602.800 391.800 603.600 400.400 ;
        RECT 607.600 396.200 608.400 400.400 ;
        RECT 610.800 395.800 611.600 400.400 ;
        RECT 612.400 391.800 613.200 400.400 ;
        RECT 616.600 395.800 617.400 400.400 ;
        RECT 618.800 395.800 619.600 400.400 ;
        RECT 622.000 395.800 622.800 400.400 ;
        RECT 625.200 391.800 626.000 400.400 ;
        RECT 630.800 395.800 631.600 400.400 ;
        RECT 634.000 395.800 634.800 400.400 ;
        RECT 639.600 392.000 640.400 400.400 ;
        RECT 643.400 395.800 644.200 400.400 ;
        RECT 647.600 391.800 648.400 400.400 ;
        RECT 649.200 395.800 650.000 400.400 ;
        RECT 652.400 395.800 653.200 400.400 ;
        RECT 655.600 395.800 656.400 400.400 ;
        RECT 662.000 395.800 662.800 400.400 ;
        RECT 665.200 395.800 666.000 400.400 ;
        RECT 673.200 395.800 674.000 400.400 ;
        RECT 676.400 395.800 677.200 400.400 ;
        RECT 679.600 395.800 680.400 400.400 ;
        RECT 682.800 395.800 683.600 400.400 ;
        RECT 652.400 391.800 653.200 392.400 ;
        RECT 655.800 391.800 656.600 392.000 ;
        RECT 282.800 391.200 309.800 391.800 ;
        RECT 388.400 391.200 415.400 391.800 ;
        RECT 309.000 391.000 309.800 391.200 ;
        RECT 414.600 391.000 415.400 391.200 ;
        RECT 451.800 391.200 478.800 391.800 ;
        RECT 652.400 391.200 679.400 391.800 ;
        RECT 451.800 391.000 452.600 391.200 ;
        RECT 678.600 391.000 679.400 391.200 ;
        RECT 209.800 370.800 210.600 371.000 ;
        RECT 267.400 370.800 268.200 371.000 ;
        RECT 183.600 370.200 210.600 370.800 ;
        RECT 241.200 370.200 268.200 370.800 ;
        RECT 419.800 370.800 420.600 371.000 ;
        RECT 480.200 370.800 481.000 371.000 ;
        RECT 419.800 370.200 446.800 370.800 ;
        RECT 2.800 361.600 3.600 370.000 ;
        RECT 8.400 361.600 9.200 366.200 ;
        RECT 11.600 361.600 12.400 366.200 ;
        RECT 17.200 361.600 18.000 370.200 ;
        RECT 20.400 361.600 21.200 366.200 ;
        RECT 23.600 361.600 24.400 370.200 ;
        RECT 27.800 361.600 28.600 366.200 ;
        RECT 30.600 361.600 31.400 366.200 ;
        RECT 34.800 361.600 35.600 370.200 ;
        RECT 37.600 361.600 38.400 370.200 ;
        RECT 42.800 361.600 43.600 369.800 ;
        RECT 47.200 361.600 48.000 370.200 ;
        RECT 52.400 361.600 53.200 369.800 ;
        RECT 55.600 361.600 56.400 366.200 ;
        RECT 59.400 361.600 60.200 366.200 ;
        RECT 63.600 361.600 64.400 370.200 ;
        RECT 65.200 361.600 66.000 366.200 ;
        RECT 68.400 361.600 69.200 366.200 ;
        RECT 70.000 361.600 70.800 366.200 ;
        RECT 73.200 361.600 74.000 370.200 ;
        RECT 77.400 361.600 78.200 366.200 ;
        RECT 79.600 361.600 80.400 366.200 ;
        RECT 84.400 361.600 85.200 369.000 ;
        RECT 87.600 361.600 88.400 370.200 ;
        RECT 89.200 361.600 90.000 370.200 ;
        RECT 93.400 361.600 94.200 366.200 ;
        RECT 95.600 361.600 96.400 370.200 ;
        RECT 99.800 361.600 100.600 366.200 ;
        RECT 102.000 361.600 102.800 370.200 ;
        RECT 106.200 361.600 107.000 366.200 ;
        RECT 113.200 361.600 114.000 366.200 ;
        RECT 116.400 361.600 117.200 365.800 ;
        RECT 120.200 361.600 121.000 366.200 ;
        RECT 124.400 361.600 125.200 370.200 ;
        RECT 127.600 361.600 128.400 369.000 ;
        RECT 130.800 361.600 131.600 370.200 ;
        RECT 135.600 361.600 136.400 370.200 ;
        RECT 137.800 361.600 138.600 366.200 ;
        RECT 142.000 361.600 142.800 370.200 ;
        RECT 145.200 361.600 146.000 366.200 ;
        RECT 148.400 361.600 149.200 366.200 ;
        RECT 151.600 361.600 152.400 370.200 ;
        RECT 157.200 361.600 158.000 366.200 ;
        RECT 160.400 361.600 161.200 366.200 ;
        RECT 166.000 361.600 166.800 370.000 ;
        RECT 170.800 361.600 171.600 369.000 ;
        RECT 174.000 361.600 174.800 370.200 ;
        RECT 183.600 369.600 184.400 370.200 ;
        RECT 187.000 370.000 187.800 370.200 ;
        RECT 175.600 361.600 176.400 366.200 ;
        RECT 178.800 361.600 179.600 366.200 ;
        RECT 180.400 361.600 181.200 366.200 ;
        RECT 183.600 361.600 184.400 366.200 ;
        RECT 186.800 361.600 187.600 366.200 ;
        RECT 193.200 361.600 194.000 366.200 ;
        RECT 196.400 361.600 197.200 366.200 ;
        RECT 204.400 361.600 205.200 366.200 ;
        RECT 207.600 361.600 208.400 366.200 ;
        RECT 210.800 361.600 211.600 366.200 ;
        RECT 214.000 361.600 214.800 366.200 ;
        RECT 216.200 361.600 217.000 366.200 ;
        RECT 220.400 361.600 221.200 370.200 ;
        RECT 223.600 361.600 224.400 369.000 ;
        RECT 228.400 361.600 229.200 369.000 ;
        RECT 231.600 361.600 232.400 370.200 ;
        RECT 241.200 369.600 242.000 370.200 ;
        RECT 244.400 370.000 245.400 370.200 ;
        RECT 233.200 361.600 234.000 366.200 ;
        RECT 236.400 361.600 237.200 366.200 ;
        RECT 238.000 361.600 238.800 366.200 ;
        RECT 241.200 361.600 242.000 366.200 ;
        RECT 244.400 361.600 245.200 366.200 ;
        RECT 250.800 361.600 251.600 366.200 ;
        RECT 254.000 361.600 254.800 366.200 ;
        RECT 262.000 361.600 262.800 366.200 ;
        RECT 265.200 361.600 266.000 366.200 ;
        RECT 268.400 361.600 269.200 366.200 ;
        RECT 271.600 361.600 272.400 366.200 ;
        RECT 278.600 361.600 279.400 366.200 ;
        RECT 282.800 361.600 283.600 370.200 ;
        RECT 286.000 361.600 286.800 369.000 ;
        RECT 289.200 361.600 290.000 370.200 ;
        RECT 290.800 361.600 291.600 370.200 ;
        RECT 294.000 361.600 294.800 370.200 ;
        RECT 297.200 361.600 298.000 370.200 ;
        RECT 300.400 361.600 301.200 370.200 ;
        RECT 303.600 361.600 304.400 370.200 ;
        RECT 305.200 361.600 306.000 366.200 ;
        RECT 308.400 361.600 309.200 370.200 ;
        RECT 312.600 361.600 313.400 366.200 ;
        RECT 319.600 361.600 320.400 369.000 ;
        RECT 324.400 361.600 325.200 366.200 ;
        RECT 326.000 361.600 326.800 366.200 ;
        RECT 330.800 361.600 331.600 369.000 ;
        RECT 337.200 361.600 338.000 366.200 ;
        RECT 340.400 361.600 341.200 365.800 ;
        RECT 343.600 361.600 344.400 366.200 ;
        RECT 346.800 361.600 347.600 365.800 ;
        RECT 351.600 361.600 352.400 365.800 ;
        RECT 354.800 361.600 355.600 366.200 ;
        RECT 356.400 361.600 357.200 366.200 ;
        RECT 364.400 361.600 365.200 369.000 ;
        RECT 367.600 361.600 368.400 366.200 ;
        RECT 372.400 361.600 373.200 369.000 ;
        RECT 380.400 361.600 381.200 365.800 ;
        RECT 383.600 361.600 384.400 366.200 ;
        RECT 385.200 361.600 386.000 366.200 ;
        RECT 388.400 361.600 389.200 365.800 ;
        RECT 391.600 361.600 392.400 366.200 ;
        RECT 394.800 361.600 395.600 365.800 ;
        RECT 398.000 361.600 398.800 370.200 ;
        RECT 402.800 361.600 403.600 370.200 ;
        RECT 406.000 361.600 406.800 370.200 ;
        RECT 409.200 361.600 410.000 370.200 ;
        RECT 442.600 370.000 443.400 370.200 ;
        RECT 446.000 369.600 446.800 370.200 ;
        RECT 454.000 370.200 481.000 370.800 ;
        RECT 656.600 370.800 657.400 371.000 ;
        RECT 656.600 370.200 683.600 370.800 ;
        RECT 454.000 369.600 454.800 370.200 ;
        RECT 457.400 370.000 458.200 370.200 ;
        RECT 415.600 361.600 416.400 366.200 ;
        RECT 418.800 361.600 419.600 366.200 ;
        RECT 422.000 361.600 422.800 366.200 ;
        RECT 425.200 361.600 426.000 366.200 ;
        RECT 433.200 361.600 434.000 366.200 ;
        RECT 436.400 361.600 437.200 366.200 ;
        RECT 442.800 361.600 443.600 366.200 ;
        RECT 446.000 361.600 446.800 366.200 ;
        RECT 449.200 361.600 450.000 366.200 ;
        RECT 450.800 361.600 451.600 366.200 ;
        RECT 454.000 361.600 454.800 366.200 ;
        RECT 457.200 361.600 458.000 366.200 ;
        RECT 463.600 361.600 464.400 366.200 ;
        RECT 466.800 361.600 467.600 366.200 ;
        RECT 474.800 361.600 475.600 366.200 ;
        RECT 478.000 361.600 478.800 366.200 ;
        RECT 481.200 361.600 482.000 366.200 ;
        RECT 484.400 361.600 485.200 366.200 ;
        RECT 486.000 361.600 486.800 370.200 ;
        RECT 489.200 361.600 490.000 370.200 ;
        RECT 492.400 361.600 493.200 370.200 ;
        RECT 495.600 361.600 496.400 370.200 ;
        RECT 498.800 361.600 499.600 370.200 ;
        RECT 500.400 361.600 501.200 366.200 ;
        RECT 503.600 361.600 504.400 366.200 ;
        RECT 505.800 361.600 506.600 366.200 ;
        RECT 510.000 361.600 510.800 370.200 ;
        RECT 512.800 361.600 513.600 370.200 ;
        RECT 518.000 361.600 518.800 369.800 ;
        RECT 521.200 361.600 522.000 370.200 ;
        RECT 525.400 361.600 526.200 366.200 ;
        RECT 528.200 361.600 529.000 366.200 ;
        RECT 532.400 361.600 533.200 370.200 ;
        RECT 534.000 361.600 534.800 366.200 ;
        RECT 537.200 361.600 538.000 365.800 ;
        RECT 541.600 361.600 542.400 370.200 ;
        RECT 546.800 361.600 547.600 369.800 ;
        RECT 551.600 361.600 552.400 370.200 ;
        RECT 557.200 361.600 558.000 366.200 ;
        RECT 560.400 361.600 561.200 366.200 ;
        RECT 566.000 361.600 566.800 370.000 ;
        RECT 569.200 361.600 570.000 366.200 ;
        RECT 572.400 361.600 573.200 366.200 ;
        RECT 578.800 361.600 579.600 370.200 ;
        RECT 583.000 361.600 583.800 366.200 ;
        RECT 585.800 361.600 586.600 366.200 ;
        RECT 590.000 361.600 590.800 370.200 ;
        RECT 591.600 361.600 592.400 370.200 ;
        RECT 594.800 361.600 595.600 369.000 ;
        RECT 598.000 361.600 598.800 370.200 ;
        RECT 601.200 361.600 602.000 369.000 ;
        RECT 606.000 361.600 606.800 366.200 ;
        RECT 610.800 361.600 611.600 370.200 ;
        RECT 612.400 361.600 613.200 366.200 ;
        RECT 615.600 361.600 616.400 366.200 ;
        RECT 618.800 361.600 619.600 366.200 ;
        RECT 620.400 361.600 621.200 370.200 ;
        RECT 624.600 361.600 625.400 366.200 ;
        RECT 628.400 361.600 629.200 369.800 ;
        RECT 633.600 361.600 634.400 370.200 ;
        RECT 637.000 361.600 637.800 366.200 ;
        RECT 641.200 361.600 642.000 370.200 ;
        RECT 642.800 361.600 643.600 366.200 ;
        RECT 646.000 361.600 646.800 366.200 ;
        RECT 647.600 361.600 648.400 370.200 ;
        RECT 679.400 370.000 680.400 370.200 ;
        RECT 682.800 369.600 683.600 370.200 ;
        RECT 652.400 361.600 653.200 366.200 ;
        RECT 655.600 361.600 656.400 366.200 ;
        RECT 658.800 361.600 659.600 366.200 ;
        RECT 662.000 361.600 662.800 366.200 ;
        RECT 670.000 361.600 670.800 366.200 ;
        RECT 673.200 361.600 674.000 366.200 ;
        RECT 679.600 361.600 680.400 366.200 ;
        RECT 682.800 361.600 683.600 366.200 ;
        RECT 686.000 361.600 686.800 366.200 ;
        RECT 0.400 360.400 689.200 361.600 ;
        RECT 2.800 352.000 3.600 360.400 ;
        RECT 8.400 355.800 9.200 360.400 ;
        RECT 11.600 355.800 12.400 360.400 ;
        RECT 17.200 351.800 18.000 360.400 ;
        RECT 21.000 355.800 21.800 360.400 ;
        RECT 25.200 351.800 26.000 360.400 ;
        RECT 27.400 355.800 28.200 360.400 ;
        RECT 31.600 351.800 32.400 360.400 ;
        RECT 33.200 351.800 34.000 360.400 ;
        RECT 37.400 355.800 38.200 360.400 ;
        RECT 40.200 355.800 41.000 360.400 ;
        RECT 44.400 351.800 45.200 360.400 ;
        RECT 47.200 351.800 48.000 360.400 ;
        RECT 52.400 352.200 53.200 360.400 ;
        RECT 55.600 355.800 56.400 360.400 ;
        RECT 58.800 355.800 59.600 360.400 ;
        RECT 61.600 351.800 62.400 360.400 ;
        RECT 66.800 352.200 67.600 360.400 ;
        RECT 70.600 355.800 71.400 360.400 ;
        RECT 74.800 351.800 75.600 360.400 ;
        RECT 76.400 351.800 77.200 360.400 ;
        RECT 80.600 355.800 81.400 360.400 ;
        RECT 83.400 355.800 84.200 360.400 ;
        RECT 87.600 351.800 88.400 360.400 ;
        RECT 89.800 355.800 90.600 360.400 ;
        RECT 94.000 351.800 94.800 360.400 ;
        RECT 95.600 351.800 96.400 360.400 ;
        RECT 98.800 353.000 99.600 360.400 ;
        RECT 102.000 351.800 102.800 360.400 ;
        RECT 106.200 355.800 107.000 360.400 ;
        RECT 113.200 351.800 114.000 360.400 ;
        RECT 117.400 355.800 118.200 360.400 ;
        RECT 121.200 352.200 122.000 360.400 ;
        RECT 126.400 351.800 127.200 360.400 ;
        RECT 129.200 355.800 130.000 360.400 ;
        RECT 133.000 355.800 133.800 360.400 ;
        RECT 137.200 351.800 138.000 360.400 ;
        RECT 139.400 355.800 140.200 360.400 ;
        RECT 143.600 351.800 144.400 360.400 ;
        RECT 145.200 351.800 146.000 360.400 ;
        RECT 149.400 355.800 150.200 360.400 ;
        RECT 152.200 355.800 153.000 360.400 ;
        RECT 156.400 351.800 157.200 360.400 ;
        RECT 158.600 355.800 159.400 360.400 ;
        RECT 162.800 351.800 163.600 360.400 ;
        RECT 165.000 355.800 165.800 360.400 ;
        RECT 169.200 351.800 170.000 360.400 ;
        RECT 170.800 355.800 171.600 360.400 ;
        RECT 174.000 355.800 174.800 360.400 ;
        RECT 177.200 355.800 178.000 360.400 ;
        RECT 183.600 355.800 184.400 360.400 ;
        RECT 186.800 355.800 187.600 360.400 ;
        RECT 194.800 355.800 195.600 360.400 ;
        RECT 198.000 355.800 198.800 360.400 ;
        RECT 201.200 355.800 202.000 360.400 ;
        RECT 204.400 355.800 205.200 360.400 ;
        RECT 207.600 353.200 208.600 360.400 ;
        RECT 213.800 359.800 214.600 360.400 ;
        RECT 213.800 353.200 214.800 359.800 ;
        RECT 217.800 355.800 218.600 360.400 ;
        RECT 174.000 351.800 174.800 352.400 ;
        RECT 177.400 351.800 178.200 352.000 ;
        RECT 222.000 351.800 222.800 360.400 ;
        RECT 226.200 351.800 227.000 360.400 ;
        RECT 230.000 351.800 230.800 360.400 ;
        RECT 234.200 355.800 235.000 360.400 ;
        RECT 236.400 355.800 237.200 360.400 ;
        RECT 239.600 355.800 240.400 360.400 ;
        RECT 241.200 355.800 242.000 360.400 ;
        RECT 244.400 355.800 245.200 360.400 ;
        RECT 247.600 355.800 248.400 360.400 ;
        RECT 254.000 355.800 254.800 360.400 ;
        RECT 257.200 355.800 258.000 360.400 ;
        RECT 265.200 355.800 266.000 360.400 ;
        RECT 268.400 355.800 269.200 360.400 ;
        RECT 271.600 355.800 272.400 360.400 ;
        RECT 274.800 355.800 275.600 360.400 ;
        RECT 244.400 351.800 245.200 352.400 ;
        RECT 247.600 351.800 248.600 352.000 ;
        RECT 281.200 351.800 282.000 360.400 ;
        RECT 284.400 351.800 285.200 360.400 ;
        RECT 287.600 351.800 288.400 360.400 ;
        RECT 290.800 351.800 291.600 360.400 ;
        RECT 294.000 351.800 294.800 360.400 ;
        RECT 297.200 355.800 298.000 360.400 ;
        RECT 298.800 355.800 299.600 360.400 ;
        RECT 302.000 355.800 302.800 360.400 ;
        RECT 304.200 355.800 305.000 360.400 ;
        RECT 308.400 351.800 309.200 360.400 ;
        RECT 311.600 356.200 312.400 360.400 ;
        RECT 314.800 355.800 315.600 360.400 ;
        RECT 318.000 353.000 318.800 360.400 ;
        RECT 326.000 353.000 326.800 360.400 ;
        RECT 334.000 353.000 334.800 360.400 ;
        RECT 340.400 355.800 341.200 360.400 ;
        RECT 343.600 356.200 344.400 360.400 ;
        RECT 351.600 353.000 352.400 360.400 ;
        RECT 356.400 356.200 357.200 360.400 ;
        RECT 359.600 355.800 360.400 360.400 ;
        RECT 361.200 355.800 362.000 360.400 ;
        RECT 364.400 355.800 365.200 360.400 ;
        RECT 366.000 355.800 366.800 360.400 ;
        RECT 369.200 355.800 370.000 360.400 ;
        RECT 372.400 353.000 373.200 360.400 ;
        RECT 378.800 355.800 379.600 360.400 ;
        RECT 382.000 356.200 382.800 360.400 ;
        RECT 385.200 355.800 386.000 360.400 ;
        RECT 388.400 355.800 389.200 360.400 ;
        RECT 391.600 355.800 392.400 360.400 ;
        RECT 394.800 355.800 395.600 360.400 ;
        RECT 402.800 355.800 403.600 360.400 ;
        RECT 406.000 355.800 406.800 360.400 ;
        RECT 412.400 355.800 413.200 360.400 ;
        RECT 415.600 355.800 416.400 360.400 ;
        RECT 418.800 355.800 419.600 360.400 ;
        RECT 425.800 355.800 426.600 360.400 ;
        RECT 412.200 351.800 413.200 352.000 ;
        RECT 415.600 351.800 416.400 352.400 ;
        RECT 430.000 351.800 430.800 360.400 ;
        RECT 431.600 355.800 432.400 360.400 ;
        RECT 434.800 355.800 435.600 360.400 ;
        RECT 436.400 355.800 437.200 360.400 ;
        RECT 439.600 355.800 440.400 360.400 ;
        RECT 442.800 355.800 443.600 360.400 ;
        RECT 446.000 355.800 446.800 360.400 ;
        RECT 454.000 355.800 454.800 360.400 ;
        RECT 457.200 355.800 458.000 360.400 ;
        RECT 463.600 355.800 464.400 360.400 ;
        RECT 466.800 355.800 467.600 360.400 ;
        RECT 470.000 355.800 470.800 360.400 ;
        RECT 471.600 355.800 472.400 360.400 ;
        RECT 474.800 355.800 475.600 360.400 ;
        RECT 463.400 351.800 464.200 352.000 ;
        RECT 466.800 351.800 467.600 352.400 ;
        RECT 476.400 351.800 477.200 360.400 ;
        RECT 480.600 355.800 481.400 360.400 ;
        RECT 484.400 351.800 485.200 360.400 ;
        RECT 490.000 355.800 490.800 360.400 ;
        RECT 493.200 355.800 494.000 360.400 ;
        RECT 498.800 352.000 499.600 360.400 ;
        RECT 503.600 352.000 504.400 360.400 ;
        RECT 509.200 355.800 510.000 360.400 ;
        RECT 512.400 355.800 513.200 360.400 ;
        RECT 518.000 351.800 518.800 360.400 ;
        RECT 521.200 355.800 522.000 360.400 ;
        RECT 525.000 355.800 525.800 360.400 ;
        RECT 529.200 351.800 530.000 360.400 ;
        RECT 532.400 352.200 533.200 360.400 ;
        RECT 537.600 351.800 538.400 360.400 ;
        RECT 540.400 351.800 541.200 360.400 ;
        RECT 544.600 355.800 545.400 360.400 ;
        RECT 546.800 351.800 547.600 360.400 ;
        RECT 551.000 355.800 551.800 360.400 ;
        RECT 553.800 355.800 554.600 360.400 ;
        RECT 558.000 351.800 558.800 360.400 ;
        RECT 561.200 355.800 562.000 360.400 ;
        RECT 562.800 355.800 563.600 360.400 ;
        RECT 566.000 355.800 566.800 360.400 ;
        RECT 573.600 351.800 574.400 360.400 ;
        RECT 578.800 352.200 579.600 360.400 ;
        RECT 583.200 351.800 584.000 360.400 ;
        RECT 588.400 352.200 589.200 360.400 ;
        RECT 593.200 352.000 594.000 360.400 ;
        RECT 598.800 355.800 599.600 360.400 ;
        RECT 602.000 355.800 602.800 360.400 ;
        RECT 607.600 351.800 608.400 360.400 ;
        RECT 610.800 351.800 611.600 360.400 ;
        RECT 615.000 355.800 615.800 360.400 ;
        RECT 617.800 355.800 618.600 360.400 ;
        RECT 622.000 351.800 622.800 360.400 ;
        RECT 625.200 352.200 626.000 360.400 ;
        RECT 630.400 351.800 631.200 360.400 ;
        RECT 633.200 351.800 634.000 360.400 ;
        RECT 637.400 355.800 638.200 360.400 ;
        RECT 640.200 355.800 641.000 360.400 ;
        RECT 644.400 351.800 645.200 360.400 ;
        RECT 649.200 351.800 650.000 360.400 ;
        RECT 652.400 351.800 653.200 360.400 ;
        RECT 658.000 355.800 658.800 360.400 ;
        RECT 661.200 355.800 662.000 360.400 ;
        RECT 666.800 352.000 667.600 360.400 ;
        RECT 673.200 351.800 674.000 360.400 ;
        RECT 678.000 351.800 678.800 360.400 ;
        RECT 679.600 355.800 680.400 360.400 ;
        RECT 174.000 351.200 201.000 351.800 ;
        RECT 244.400 351.200 271.400 351.800 ;
        RECT 200.200 351.000 201.000 351.200 ;
        RECT 270.600 351.000 271.400 351.200 ;
        RECT 389.400 351.200 416.400 351.800 ;
        RECT 440.600 351.200 467.600 351.800 ;
        RECT 389.400 351.000 390.200 351.200 ;
        RECT 440.600 351.000 441.400 351.200 ;
        RECT 171.800 330.800 172.600 331.000 ;
        RECT 234.200 330.800 235.000 331.000 ;
        RECT 299.400 330.800 300.200 331.000 ;
        RECT 171.800 330.200 198.800 330.800 ;
        RECT 234.200 330.200 261.200 330.800 ;
        RECT 2.800 321.600 3.600 330.000 ;
        RECT 8.400 321.600 9.200 326.200 ;
        RECT 11.600 321.600 12.400 326.200 ;
        RECT 17.200 321.600 18.000 330.200 ;
        RECT 21.000 321.600 21.800 326.200 ;
        RECT 25.200 321.600 26.000 330.200 ;
        RECT 27.400 321.600 28.200 326.200 ;
        RECT 31.600 321.600 32.400 330.200 ;
        RECT 34.400 321.600 35.200 330.200 ;
        RECT 39.600 321.600 40.400 329.800 ;
        RECT 44.400 321.600 45.200 330.000 ;
        RECT 50.000 321.600 50.800 326.200 ;
        RECT 53.200 321.600 54.000 326.200 ;
        RECT 58.800 321.600 59.600 330.200 ;
        RECT 62.000 321.600 62.800 326.200 ;
        RECT 65.200 321.600 66.000 326.200 ;
        RECT 69.000 321.600 69.800 330.200 ;
        RECT 74.800 321.600 75.600 330.000 ;
        RECT 80.400 321.600 81.200 326.200 ;
        RECT 83.600 321.600 84.400 326.200 ;
        RECT 89.200 321.600 90.000 330.200 ;
        RECT 92.400 321.600 93.200 330.200 ;
        RECT 96.600 321.600 97.400 326.200 ;
        RECT 98.800 321.600 99.600 330.200 ;
        RECT 103.000 321.600 103.800 326.200 ;
        RECT 111.600 321.600 112.400 330.000 ;
        RECT 117.200 321.600 118.000 326.200 ;
        RECT 120.400 321.600 121.200 326.200 ;
        RECT 126.000 321.600 126.800 330.200 ;
        RECT 129.200 321.600 130.000 326.200 ;
        RECT 132.400 321.600 133.200 326.200 ;
        RECT 134.000 321.600 134.800 326.200 ;
        RECT 137.200 321.600 138.000 326.200 ;
        RECT 140.400 321.600 141.200 326.200 ;
        RECT 143.600 322.200 144.600 328.800 ;
        RECT 143.800 321.600 144.600 322.200 ;
        RECT 149.800 321.600 150.800 328.800 ;
        RECT 153.200 321.600 154.000 330.200 ;
        RECT 156.400 321.600 157.200 326.200 ;
        RECT 159.600 321.600 160.400 326.200 ;
        RECT 161.200 321.600 162.000 330.200 ;
        RECT 194.600 330.000 195.600 330.200 ;
        RECT 198.000 329.600 198.800 330.200 ;
        RECT 165.400 321.600 166.200 326.200 ;
        RECT 167.600 321.600 168.400 326.200 ;
        RECT 170.800 321.600 171.600 326.200 ;
        RECT 174.000 321.600 174.800 326.200 ;
        RECT 177.200 321.600 178.000 326.200 ;
        RECT 185.200 321.600 186.000 326.200 ;
        RECT 188.400 321.600 189.200 326.200 ;
        RECT 194.800 321.600 195.600 326.200 ;
        RECT 198.000 321.600 198.800 326.200 ;
        RECT 201.200 321.600 202.000 326.200 ;
        RECT 202.800 321.600 203.600 330.200 ;
        RECT 206.000 321.600 206.800 329.000 ;
        RECT 210.800 321.600 211.600 329.000 ;
        RECT 214.000 321.600 214.800 330.200 ;
        RECT 216.200 321.600 217.000 326.200 ;
        RECT 220.400 321.600 221.200 330.200 ;
        RECT 223.600 321.600 224.400 326.200 ;
        RECT 228.400 321.600 229.200 330.200 ;
        RECT 257.000 330.000 257.800 330.200 ;
        RECT 260.400 329.600 261.200 330.200 ;
        RECT 273.200 330.200 300.200 330.800 ;
        RECT 439.000 330.800 439.800 331.000 ;
        RECT 439.000 330.200 466.000 330.800 ;
        RECT 273.200 329.600 274.000 330.200 ;
        RECT 276.400 330.000 277.400 330.200 ;
        RECT 230.000 321.600 230.800 326.200 ;
        RECT 233.200 321.600 234.000 326.200 ;
        RECT 236.400 321.600 237.200 326.200 ;
        RECT 239.600 321.600 240.400 326.200 ;
        RECT 247.600 321.600 248.400 326.200 ;
        RECT 250.800 321.600 251.600 326.200 ;
        RECT 257.200 321.600 258.000 326.200 ;
        RECT 260.400 321.600 261.200 326.200 ;
        RECT 263.600 321.600 264.400 326.200 ;
        RECT 270.000 321.600 270.800 326.200 ;
        RECT 273.200 321.600 274.000 326.200 ;
        RECT 276.400 321.600 277.200 326.200 ;
        RECT 282.800 321.600 283.600 326.200 ;
        RECT 286.000 321.600 286.800 326.200 ;
        RECT 294.000 321.600 294.800 326.200 ;
        RECT 297.200 321.600 298.000 326.200 ;
        RECT 300.400 321.600 301.200 326.200 ;
        RECT 303.600 321.600 304.400 326.200 ;
        RECT 305.800 321.600 306.600 326.200 ;
        RECT 310.000 321.600 310.800 330.200 ;
        RECT 312.200 321.600 313.000 326.200 ;
        RECT 316.400 321.600 317.200 330.200 ;
        RECT 318.000 321.600 318.800 326.200 ;
        RECT 321.200 321.600 322.000 326.200 ;
        RECT 327.600 321.600 328.400 329.000 ;
        RECT 335.600 321.600 336.400 329.000 ;
        RECT 343.600 321.600 344.400 329.000 ;
        RECT 351.600 321.600 352.400 329.000 ;
        RECT 356.400 321.600 357.200 329.000 ;
        RECT 362.800 321.600 363.600 326.200 ;
        RECT 366.000 321.600 366.800 326.200 ;
        RECT 372.400 321.600 373.200 329.000 ;
        RECT 375.600 321.600 376.400 326.200 ;
        RECT 378.800 321.600 379.600 326.200 ;
        RECT 380.400 321.600 381.200 326.200 ;
        RECT 383.600 321.600 384.400 326.200 ;
        RECT 390.000 321.600 390.800 329.000 ;
        RECT 393.200 321.600 394.000 326.200 ;
        RECT 396.400 321.600 397.200 326.200 ;
        RECT 399.600 321.600 400.400 329.000 ;
        RECT 406.600 321.600 407.400 326.200 ;
        RECT 410.800 321.600 411.600 330.200 ;
        RECT 412.400 321.600 413.200 326.200 ;
        RECT 415.600 321.600 416.400 326.200 ;
        RECT 422.000 321.600 422.800 330.200 ;
        RECT 426.200 321.600 427.000 326.200 ;
        RECT 428.400 321.600 429.200 330.200 ;
        RECT 461.800 330.000 462.800 330.200 ;
        RECT 465.200 329.600 466.000 330.200 ;
        RECT 432.600 321.600 433.400 326.200 ;
        RECT 434.800 321.600 435.600 326.200 ;
        RECT 438.000 321.600 438.800 326.200 ;
        RECT 441.200 321.600 442.000 326.200 ;
        RECT 444.400 321.600 445.200 326.200 ;
        RECT 452.400 321.600 453.200 326.200 ;
        RECT 455.600 321.600 456.400 326.200 ;
        RECT 462.000 321.600 462.800 326.200 ;
        RECT 465.200 321.600 466.000 326.200 ;
        RECT 468.400 321.600 469.200 326.200 ;
        RECT 470.000 321.600 470.800 326.200 ;
        RECT 473.200 321.600 474.000 326.200 ;
        RECT 474.800 321.600 475.600 326.200 ;
        RECT 478.000 321.600 478.800 326.200 ;
        RECT 479.600 321.600 480.400 326.200 ;
        RECT 482.800 321.600 483.600 330.200 ;
        RECT 487.000 321.600 487.800 326.200 ;
        RECT 489.200 321.600 490.000 330.200 ;
        RECT 492.400 321.600 493.200 329.000 ;
        RECT 497.200 321.600 498.000 329.800 ;
        RECT 502.400 321.600 503.200 330.200 ;
        RECT 505.200 321.600 506.000 330.200 ;
        RECT 509.400 321.600 510.200 326.200 ;
        RECT 512.200 321.600 513.000 326.200 ;
        RECT 516.400 321.600 517.200 330.200 ;
        RECT 518.000 321.600 518.800 326.200 ;
        RECT 521.200 321.600 522.000 330.200 ;
        RECT 525.400 321.600 526.200 326.200 ;
        RECT 529.200 321.600 530.000 329.000 ;
        RECT 532.400 321.600 533.200 330.200 ;
        RECT 534.000 321.600 534.800 326.200 ;
        RECT 537.200 321.600 538.000 325.800 ;
        RECT 540.400 321.600 541.200 330.200 ;
        RECT 544.600 321.600 545.400 326.200 ;
        RECT 546.800 321.600 547.600 326.200 ;
        RECT 550.000 321.600 550.800 325.800 ;
        RECT 553.200 321.600 554.000 330.200 ;
        RECT 557.400 321.600 558.200 326.200 ;
        RECT 561.200 321.600 562.000 330.200 ;
        RECT 566.800 321.600 567.600 326.200 ;
        RECT 570.000 321.600 570.800 326.200 ;
        RECT 575.600 321.600 576.400 330.000 ;
        RECT 583.600 321.600 584.400 330.200 ;
        RECT 587.800 321.600 588.600 326.200 ;
        RECT 590.600 321.600 591.400 326.200 ;
        RECT 594.800 321.600 595.600 330.200 ;
        RECT 596.400 321.600 597.200 326.200 ;
        RECT 599.600 321.600 600.400 325.800 ;
        RECT 604.400 321.600 605.200 329.000 ;
        RECT 607.600 321.600 608.400 330.200 ;
        RECT 609.800 321.600 610.600 326.200 ;
        RECT 614.000 321.600 614.800 330.200 ;
        RECT 617.200 321.600 618.000 329.000 ;
        RECT 620.400 321.600 621.200 330.200 ;
        RECT 622.000 321.600 622.800 330.200 ;
        RECT 626.200 321.600 627.000 326.200 ;
        RECT 630.000 321.600 630.800 325.800 ;
        RECT 633.200 321.600 634.000 326.200 ;
        RECT 636.400 321.600 637.200 326.200 ;
        RECT 639.600 321.600 640.400 329.800 ;
        RECT 644.800 321.600 645.600 330.200 ;
        RECT 647.600 321.600 648.400 330.200 ;
        RECT 651.800 321.600 652.600 326.200 ;
        RECT 655.600 321.600 656.400 329.800 ;
        RECT 660.800 321.600 661.600 330.200 ;
        RECT 664.200 321.600 665.000 326.200 ;
        RECT 668.400 321.600 669.200 330.200 ;
        RECT 671.600 321.600 672.400 330.000 ;
        RECT 677.200 321.600 678.000 326.200 ;
        RECT 680.400 321.600 681.200 326.200 ;
        RECT 686.000 321.600 686.800 330.200 ;
        RECT 0.400 320.400 689.200 321.600 ;
        RECT 1.200 315.800 2.000 320.400 ;
        RECT 4.400 315.800 5.200 320.400 ;
        RECT 7.600 315.800 8.400 320.400 ;
        RECT 14.000 315.800 14.800 320.400 ;
        RECT 17.200 315.800 18.000 320.400 ;
        RECT 25.200 315.800 26.000 320.400 ;
        RECT 28.400 315.800 29.200 320.400 ;
        RECT 31.600 315.800 32.400 320.400 ;
        RECT 34.800 315.800 35.600 320.400 ;
        RECT 4.400 311.800 5.200 312.400 ;
        RECT 7.800 311.800 8.600 312.000 ;
        RECT 36.400 311.800 37.200 320.400 ;
        RECT 40.600 315.800 41.400 320.400 ;
        RECT 43.400 315.800 44.200 320.400 ;
        RECT 47.600 311.800 48.400 320.400 ;
        RECT 50.800 315.800 51.600 320.400 ;
        RECT 52.400 315.800 53.200 320.400 ;
        RECT 55.600 315.800 56.400 320.400 ;
        RECT 57.200 315.800 58.000 320.400 ;
        RECT 60.400 315.800 61.200 320.400 ;
        RECT 62.000 315.800 62.800 320.400 ;
        RECT 65.200 315.800 66.000 320.400 ;
        RECT 68.400 315.800 69.200 320.400 ;
        RECT 74.800 315.800 75.600 320.400 ;
        RECT 78.000 315.800 78.800 320.400 ;
        RECT 86.000 315.800 86.800 320.400 ;
        RECT 89.200 315.800 90.000 320.400 ;
        RECT 92.400 315.800 93.200 320.400 ;
        RECT 95.600 315.800 96.400 320.400 ;
        RECT 98.800 315.800 99.600 320.400 ;
        RECT 100.400 315.800 101.200 320.400 ;
        RECT 103.600 316.200 104.400 320.400 ;
        RECT 111.600 315.800 112.400 320.400 ;
        RECT 114.800 315.800 115.600 320.400 ;
        RECT 118.000 315.800 118.800 320.400 ;
        RECT 124.400 315.800 125.200 320.400 ;
        RECT 127.600 315.800 128.400 320.400 ;
        RECT 135.600 315.800 136.400 320.400 ;
        RECT 138.800 315.800 139.600 320.400 ;
        RECT 142.000 315.800 142.800 320.400 ;
        RECT 145.200 315.800 146.000 320.400 ;
        RECT 147.400 315.800 148.200 320.400 ;
        RECT 65.200 311.800 66.000 312.400 ;
        RECT 68.600 311.800 69.400 312.000 ;
        RECT 114.800 311.800 115.600 312.400 ;
        RECT 118.200 311.800 119.000 312.000 ;
        RECT 151.600 311.800 152.400 320.400 ;
        RECT 153.200 315.800 154.000 320.400 ;
        RECT 156.400 315.800 157.200 320.400 ;
        RECT 158.000 315.800 158.800 320.400 ;
        RECT 161.200 311.800 162.000 320.400 ;
        RECT 164.400 313.000 165.200 320.400 ;
        RECT 167.600 315.800 168.400 320.400 ;
        RECT 170.800 315.800 171.600 320.400 ;
        RECT 174.000 315.800 174.800 320.400 ;
        RECT 177.200 315.800 178.000 320.400 ;
        RECT 185.200 315.800 186.000 320.400 ;
        RECT 188.400 315.800 189.200 320.400 ;
        RECT 194.800 315.800 195.600 320.400 ;
        RECT 198.000 315.800 198.800 320.400 ;
        RECT 201.200 315.800 202.000 320.400 ;
        RECT 202.800 315.800 203.600 320.400 ;
        RECT 206.000 315.800 206.800 320.400 ;
        RECT 207.600 315.800 208.400 320.400 ;
        RECT 210.800 315.800 211.600 320.400 ;
        RECT 213.000 315.800 213.800 320.400 ;
        RECT 194.600 311.800 195.600 312.000 ;
        RECT 198.000 311.800 198.800 312.400 ;
        RECT 217.200 311.800 218.000 320.400 ;
        RECT 220.400 313.000 221.200 320.400 ;
        RECT 225.200 313.000 226.000 320.400 ;
        RECT 228.400 311.800 229.200 320.400 ;
        RECT 230.000 311.800 230.800 320.400 ;
        RECT 233.200 311.800 234.000 320.400 ;
        RECT 236.400 311.800 237.200 320.400 ;
        RECT 238.000 315.800 238.800 320.400 ;
        RECT 241.200 315.800 242.000 320.400 ;
        RECT 242.800 311.800 243.600 320.400 ;
        RECT 247.000 315.800 247.800 320.400 ;
        RECT 254.000 315.800 254.800 320.400 ;
        RECT 257.200 315.800 258.000 320.400 ;
        RECT 260.400 315.800 261.200 320.400 ;
        RECT 266.800 315.800 267.600 320.400 ;
        RECT 270.000 315.800 270.800 320.400 ;
        RECT 278.000 315.800 278.800 320.400 ;
        RECT 281.200 315.800 282.000 320.400 ;
        RECT 284.400 315.800 285.200 320.400 ;
        RECT 287.600 315.800 288.400 320.400 ;
        RECT 257.200 311.800 258.000 312.400 ;
        RECT 260.400 311.800 261.400 312.000 ;
        RECT 289.200 311.800 290.000 320.400 ;
        RECT 292.400 311.800 293.200 320.400 ;
        RECT 294.000 315.800 294.800 320.400 ;
        RECT 297.200 315.800 298.000 320.400 ;
        RECT 298.800 311.800 299.600 320.400 ;
        RECT 303.000 315.800 303.800 320.400 ;
        RECT 306.800 315.800 307.600 320.400 ;
        RECT 308.400 315.800 309.200 320.400 ;
        RECT 311.600 315.800 312.400 320.400 ;
        RECT 314.800 316.200 315.600 320.400 ;
        RECT 318.000 315.800 318.800 320.400 ;
        RECT 319.600 315.800 320.400 320.400 ;
        RECT 322.800 315.800 323.600 320.400 ;
        RECT 326.000 313.000 326.800 320.400 ;
        RECT 329.200 311.800 330.000 320.400 ;
        RECT 330.800 315.800 331.600 320.400 ;
        RECT 334.000 316.200 334.800 320.400 ;
        RECT 337.200 311.800 338.000 320.400 ;
        RECT 340.400 313.000 341.200 320.400 ;
        RECT 343.600 311.800 344.400 320.400 ;
        RECT 346.800 311.800 347.600 320.400 ;
        RECT 348.400 315.800 349.200 320.400 ;
        RECT 351.600 315.800 352.400 320.400 ;
        RECT 353.200 311.800 354.000 320.400 ;
        RECT 359.600 311.800 360.400 320.400 ;
        RECT 361.200 311.800 362.000 320.400 ;
        RECT 365.400 315.800 366.200 320.400 ;
        RECT 367.600 315.800 368.400 320.400 ;
        RECT 370.800 315.800 371.600 320.400 ;
        RECT 374.000 315.800 374.800 320.400 ;
        RECT 377.200 315.800 378.000 320.400 ;
        RECT 385.200 315.800 386.000 320.400 ;
        RECT 388.400 315.800 389.200 320.400 ;
        RECT 394.800 315.800 395.600 320.400 ;
        RECT 398.000 315.800 398.800 320.400 ;
        RECT 401.200 315.800 402.000 320.400 ;
        RECT 407.600 315.800 408.400 320.400 ;
        RECT 410.800 315.800 411.600 320.400 ;
        RECT 414.000 315.800 414.800 320.400 ;
        RECT 420.400 315.800 421.200 320.400 ;
        RECT 423.600 315.800 424.400 320.400 ;
        RECT 431.600 315.800 432.400 320.400 ;
        RECT 434.800 315.800 435.600 320.400 ;
        RECT 438.000 315.800 438.800 320.400 ;
        RECT 441.200 315.800 442.000 320.400 ;
        RECT 442.800 315.800 443.600 320.400 ;
        RECT 394.600 311.800 395.400 312.000 ;
        RECT 398.000 311.800 398.800 312.400 ;
        RECT 4.400 311.200 31.400 311.800 ;
        RECT 65.200 311.200 92.200 311.800 ;
        RECT 114.800 311.200 141.800 311.800 ;
        RECT 30.600 311.000 31.400 311.200 ;
        RECT 91.400 311.000 92.200 311.200 ;
        RECT 141.000 311.000 141.800 311.200 ;
        RECT 171.800 311.200 198.800 311.800 ;
        RECT 257.200 311.200 284.200 311.800 ;
        RECT 171.800 311.000 172.600 311.200 ;
        RECT 283.400 311.000 284.200 311.200 ;
        RECT 371.800 311.200 398.800 311.800 ;
        RECT 410.800 311.800 411.600 312.400 ;
        RECT 447.600 312.000 448.400 320.400 ;
        RECT 453.200 315.800 454.000 320.400 ;
        RECT 456.400 315.800 457.200 320.400 ;
        RECT 414.000 311.800 415.000 312.000 ;
        RECT 462.000 311.800 462.800 320.400 ;
        RECT 465.200 315.800 466.000 320.400 ;
        RECT 468.400 311.800 469.200 320.400 ;
        RECT 472.600 315.800 473.400 320.400 ;
        RECT 476.000 311.800 476.800 320.400 ;
        RECT 481.200 312.200 482.000 320.400 ;
        RECT 484.400 311.800 485.200 320.400 ;
        RECT 488.600 315.800 489.400 320.400 ;
        RECT 491.400 315.800 492.200 320.400 ;
        RECT 495.600 311.800 496.400 320.400 ;
        RECT 497.800 315.800 498.600 320.400 ;
        RECT 502.000 311.800 502.800 320.400 ;
        RECT 503.600 315.800 504.400 320.400 ;
        RECT 507.400 315.800 508.200 320.400 ;
        RECT 511.600 311.800 512.400 320.400 ;
        RECT 513.200 311.800 514.000 320.400 ;
        RECT 519.600 313.000 520.400 320.400 ;
        RECT 522.800 311.800 523.600 320.400 ;
        RECT 524.400 311.800 525.200 320.400 ;
        RECT 527.600 313.000 528.400 320.400 ;
        RECT 530.800 311.800 531.600 320.400 ;
        RECT 535.000 315.800 535.800 320.400 ;
        RECT 537.200 311.800 538.000 320.400 ;
        RECT 541.400 315.800 542.200 320.400 ;
        RECT 545.200 313.000 546.000 320.400 ;
        RECT 548.400 311.800 549.200 320.400 ;
        RECT 550.600 315.800 551.400 320.400 ;
        RECT 554.800 311.800 555.600 320.400 ;
        RECT 556.400 311.800 557.200 320.400 ;
        RECT 560.600 315.800 561.400 320.400 ;
        RECT 563.400 315.800 564.200 320.400 ;
        RECT 567.600 311.800 568.400 320.400 ;
        RECT 570.800 315.800 571.600 320.400 ;
        RECT 578.800 312.000 579.600 320.400 ;
        RECT 584.400 315.800 585.200 320.400 ;
        RECT 587.600 315.800 588.400 320.400 ;
        RECT 593.200 311.800 594.000 320.400 ;
        RECT 596.400 311.800 597.200 320.400 ;
        RECT 600.600 315.800 601.400 320.400 ;
        RECT 603.400 315.800 604.200 320.400 ;
        RECT 607.600 311.800 608.400 320.400 ;
        RECT 610.800 312.200 611.600 320.400 ;
        RECT 616.000 311.800 616.800 320.400 ;
        RECT 620.400 313.000 621.200 320.400 ;
        RECT 623.600 311.800 624.400 320.400 ;
        RECT 625.200 315.800 626.000 320.400 ;
        RECT 628.400 315.800 629.200 320.400 ;
        RECT 630.600 315.800 631.400 320.400 ;
        RECT 634.800 311.800 635.600 320.400 ;
        RECT 638.600 311.800 639.400 320.400 ;
        RECT 644.400 315.800 645.200 320.400 ;
        RECT 647.200 311.800 648.000 320.400 ;
        RECT 652.400 312.200 653.200 320.400 ;
        RECT 655.600 311.800 656.400 320.400 ;
        RECT 659.800 315.800 660.600 320.400 ;
        RECT 662.600 315.800 663.400 320.400 ;
        RECT 666.800 311.800 667.600 320.400 ;
        RECT 670.000 312.000 670.800 320.400 ;
        RECT 675.600 315.800 676.400 320.400 ;
        RECT 678.800 315.800 679.600 320.400 ;
        RECT 684.400 311.800 685.200 320.400 ;
        RECT 410.800 311.200 437.800 311.800 ;
        RECT 371.800 311.000 372.600 311.200 ;
        RECT 437.000 311.000 437.800 311.200 ;
        RECT 91.400 290.800 92.200 291.000 ;
        RECT 147.400 290.800 148.200 291.000 ;
        RECT 193.800 290.800 194.600 291.000 ;
        RECT 235.400 290.800 236.200 291.000 ;
        RECT 288.200 290.800 289.000 291.000 ;
        RECT 65.200 290.200 92.200 290.800 ;
        RECT 121.200 290.200 148.200 290.800 ;
        RECT 167.600 290.200 194.600 290.800 ;
        RECT 209.200 290.200 236.200 290.800 ;
        RECT 262.000 290.200 289.000 290.800 ;
        RECT 371.800 290.800 372.600 291.000 ;
        RECT 449.800 290.800 450.600 291.000 ;
        RECT 371.800 290.200 398.800 290.800 ;
        RECT 423.600 290.200 450.600 290.800 ;
        RECT 1.200 281.600 2.000 286.200 ;
        RECT 4.400 281.600 5.200 290.200 ;
        RECT 8.600 281.600 9.400 286.200 ;
        RECT 11.400 281.600 12.200 286.200 ;
        RECT 15.600 281.600 16.400 290.200 ;
        RECT 17.200 281.600 18.000 286.200 ;
        RECT 20.400 281.600 21.200 286.200 ;
        RECT 22.600 281.600 23.400 286.200 ;
        RECT 26.800 281.600 27.600 290.200 ;
        RECT 28.400 281.600 29.200 290.200 ;
        RECT 32.600 281.600 33.400 286.200 ;
        RECT 35.400 281.600 36.200 286.200 ;
        RECT 39.600 281.600 40.400 290.200 ;
        RECT 42.800 281.600 43.600 286.200 ;
        RECT 44.400 281.600 45.200 286.200 ;
        RECT 47.600 281.600 48.400 286.200 ;
        RECT 49.800 281.600 50.600 286.200 ;
        RECT 54.000 281.600 54.800 290.200 ;
        RECT 56.200 281.600 57.000 286.200 ;
        RECT 60.400 281.600 61.200 290.200 ;
        RECT 65.200 289.600 66.000 290.200 ;
        RECT 68.400 290.000 69.400 290.200 ;
        RECT 62.000 281.600 62.800 286.200 ;
        RECT 65.200 281.600 66.000 286.200 ;
        RECT 68.400 281.600 69.200 286.200 ;
        RECT 74.800 281.600 75.600 286.200 ;
        RECT 78.000 281.600 78.800 286.200 ;
        RECT 86.000 281.600 86.800 286.200 ;
        RECT 89.200 281.600 90.000 286.200 ;
        RECT 92.400 281.600 93.200 286.200 ;
        RECT 95.600 281.600 96.400 286.200 ;
        RECT 97.200 281.600 98.000 286.200 ;
        RECT 100.400 281.600 101.200 286.200 ;
        RECT 102.600 281.600 103.400 286.200 ;
        RECT 106.800 281.600 107.600 290.200 ;
        RECT 121.200 289.600 122.000 290.200 ;
        RECT 124.600 290.000 125.400 290.200 ;
        RECT 108.400 281.600 109.200 286.200 ;
        RECT 111.600 281.600 112.400 286.200 ;
        RECT 118.000 281.600 118.800 286.200 ;
        RECT 121.200 281.600 122.000 286.200 ;
        RECT 124.400 281.600 125.200 286.200 ;
        RECT 130.800 281.600 131.600 286.200 ;
        RECT 134.000 281.600 134.800 286.200 ;
        RECT 142.000 281.600 142.800 286.200 ;
        RECT 145.200 281.600 146.000 286.200 ;
        RECT 148.400 281.600 149.200 286.200 ;
        RECT 151.600 281.600 152.400 286.200 ;
        RECT 153.200 281.600 154.000 286.200 ;
        RECT 156.400 281.600 157.200 286.200 ;
        RECT 158.600 281.600 159.400 286.200 ;
        RECT 162.800 281.600 163.600 290.200 ;
        RECT 167.600 289.600 168.400 290.200 ;
        RECT 171.000 290.000 171.800 290.200 ;
        RECT 164.400 281.600 165.200 286.200 ;
        RECT 167.600 281.600 168.400 286.200 ;
        RECT 170.800 281.600 171.600 286.200 ;
        RECT 177.200 281.600 178.000 286.200 ;
        RECT 180.400 281.600 181.200 286.200 ;
        RECT 188.400 281.600 189.200 286.200 ;
        RECT 191.600 281.600 192.400 286.200 ;
        RECT 194.800 281.600 195.600 286.200 ;
        RECT 198.000 281.600 198.800 286.200 ;
        RECT 199.600 281.600 200.400 290.200 ;
        RECT 209.200 289.600 210.000 290.200 ;
        RECT 212.400 290.000 213.400 290.200 ;
        RECT 203.800 281.600 204.600 286.200 ;
        RECT 206.000 281.600 206.800 286.200 ;
        RECT 209.200 281.600 210.000 286.200 ;
        RECT 212.400 281.600 213.200 286.200 ;
        RECT 218.800 281.600 219.600 286.200 ;
        RECT 222.000 281.600 222.800 286.200 ;
        RECT 230.000 281.600 230.800 286.200 ;
        RECT 233.200 281.600 234.000 286.200 ;
        RECT 236.400 281.600 237.200 286.200 ;
        RECT 239.600 281.600 240.400 286.200 ;
        RECT 241.200 281.600 242.000 290.200 ;
        RECT 262.000 289.600 262.800 290.200 ;
        RECT 265.200 290.000 266.200 290.200 ;
        RECT 244.400 281.600 245.200 286.200 ;
        RECT 247.600 281.600 248.400 286.200 ;
        RECT 249.200 281.600 250.000 286.200 ;
        RECT 252.400 281.600 253.200 286.200 ;
        RECT 258.800 281.600 259.600 286.200 ;
        RECT 262.000 281.600 262.800 286.200 ;
        RECT 265.200 281.600 266.000 286.200 ;
        RECT 271.600 281.600 272.400 286.200 ;
        RECT 274.800 281.600 275.600 286.200 ;
        RECT 282.800 281.600 283.600 286.200 ;
        RECT 286.000 281.600 286.800 286.200 ;
        RECT 289.200 281.600 290.000 286.200 ;
        RECT 292.400 281.600 293.200 286.200 ;
        RECT 294.000 281.600 294.800 286.200 ;
        RECT 297.200 281.600 298.000 285.800 ;
        RECT 302.000 281.600 302.800 289.000 ;
        RECT 306.800 281.600 307.600 285.800 ;
        RECT 310.000 281.600 310.800 286.200 ;
        RECT 313.200 281.600 314.000 285.800 ;
        RECT 316.400 281.600 317.200 286.200 ;
        RECT 319.600 281.600 320.400 285.800 ;
        RECT 322.800 281.600 323.600 286.200 ;
        RECT 324.400 281.600 325.200 286.200 ;
        RECT 327.600 281.600 328.400 286.200 ;
        RECT 330.800 281.600 331.600 285.800 ;
        RECT 334.000 281.600 334.800 286.200 ;
        RECT 335.600 281.600 336.400 286.200 ;
        RECT 338.800 281.600 339.600 285.800 ;
        RECT 343.600 281.600 344.400 285.800 ;
        RECT 346.800 281.600 347.600 286.200 ;
        RECT 348.400 281.600 349.200 286.200 ;
        RECT 351.600 281.600 352.400 285.800 ;
        RECT 356.000 281.600 356.800 290.200 ;
        RECT 394.600 290.000 395.400 290.200 ;
        RECT 361.200 281.600 362.000 289.800 ;
        RECT 398.000 289.600 398.800 290.200 ;
        RECT 366.000 281.600 366.800 286.200 ;
        RECT 367.600 281.600 368.400 286.200 ;
        RECT 370.800 281.600 371.600 286.200 ;
        RECT 374.000 281.600 374.800 286.200 ;
        RECT 377.200 281.600 378.000 286.200 ;
        RECT 385.200 281.600 386.000 286.200 ;
        RECT 388.400 281.600 389.200 286.200 ;
        RECT 394.800 281.600 395.600 286.200 ;
        RECT 398.000 281.600 398.800 286.200 ;
        RECT 401.200 281.600 402.000 286.200 ;
        RECT 404.400 281.600 405.200 289.800 ;
        RECT 409.600 281.600 410.400 290.200 ;
        RECT 423.600 289.600 424.400 290.200 ;
        RECT 427.000 290.000 427.800 290.200 ;
        RECT 414.000 281.600 414.800 286.200 ;
        RECT 420.400 281.600 421.200 286.200 ;
        RECT 423.600 281.600 424.400 286.200 ;
        RECT 426.800 281.600 427.600 286.200 ;
        RECT 433.200 281.600 434.000 286.200 ;
        RECT 436.400 281.600 437.200 286.200 ;
        RECT 444.400 281.600 445.200 286.200 ;
        RECT 447.600 281.600 448.400 286.200 ;
        RECT 450.800 281.600 451.600 286.200 ;
        RECT 454.000 281.600 454.800 286.200 ;
        RECT 456.200 281.600 457.000 286.200 ;
        RECT 460.400 281.600 461.200 290.200 ;
        RECT 463.600 281.600 464.400 286.200 ;
        RECT 465.200 281.600 466.000 290.200 ;
        RECT 469.400 281.600 470.200 286.200 ;
        RECT 472.800 281.600 473.600 290.200 ;
        RECT 478.000 281.600 478.800 289.800 ;
        RECT 481.200 281.600 482.000 290.200 ;
        RECT 485.400 281.600 486.200 286.200 ;
        RECT 489.200 281.600 490.000 290.200 ;
        RECT 494.800 281.600 495.600 286.200 ;
        RECT 498.000 281.600 498.800 286.200 ;
        RECT 503.600 281.600 504.400 290.000 ;
        RECT 506.800 281.600 507.600 286.200 ;
        RECT 511.200 281.600 512.000 290.200 ;
        RECT 516.400 281.600 517.200 289.800 ;
        RECT 520.200 281.600 521.000 286.200 ;
        RECT 524.400 281.600 525.200 290.200 ;
        RECT 526.000 281.600 526.800 290.200 ;
        RECT 530.200 281.600 531.000 286.200 ;
        RECT 534.000 281.600 534.800 289.800 ;
        RECT 539.200 281.600 540.000 290.200 ;
        RECT 542.600 281.600 543.400 286.200 ;
        RECT 546.800 281.600 547.600 290.200 ;
        RECT 550.000 281.600 550.800 286.200 ;
        RECT 553.200 281.600 554.000 289.000 ;
        RECT 556.400 281.600 557.200 290.200 ;
        RECT 559.600 281.600 560.400 290.000 ;
        RECT 565.200 281.600 566.000 286.200 ;
        RECT 568.400 281.600 569.200 286.200 ;
        RECT 574.000 281.600 574.800 290.200 ;
        RECT 583.600 281.600 584.400 289.800 ;
        RECT 588.800 281.600 589.600 290.200 ;
        RECT 593.200 281.600 594.000 289.800 ;
        RECT 598.400 281.600 599.200 290.200 ;
        RECT 601.200 281.600 602.000 290.200 ;
        RECT 605.400 281.600 606.200 286.200 ;
        RECT 608.200 281.600 609.000 286.200 ;
        RECT 612.400 281.600 613.200 290.200 ;
        RECT 614.600 281.600 615.400 286.200 ;
        RECT 618.800 281.600 619.600 290.200 ;
        RECT 621.000 281.600 621.800 286.200 ;
        RECT 625.200 281.600 626.000 290.200 ;
        RECT 626.800 281.600 627.600 286.200 ;
        RECT 630.000 281.600 630.800 286.200 ;
        RECT 633.200 281.600 634.000 286.200 ;
        RECT 636.400 281.600 637.200 289.800 ;
        RECT 641.600 281.600 642.400 290.200 ;
        RECT 644.400 281.600 645.200 290.200 ;
        RECT 648.600 281.600 649.400 286.200 ;
        RECT 652.400 281.600 653.200 290.200 ;
        RECT 658.000 281.600 658.800 286.200 ;
        RECT 661.200 281.600 662.000 286.200 ;
        RECT 666.800 281.600 667.600 290.000 ;
        RECT 670.000 281.600 670.800 290.200 ;
        RECT 673.200 281.600 674.000 290.200 ;
        RECT 676.400 281.600 677.200 290.200 ;
        RECT 679.600 281.600 680.400 290.200 ;
        RECT 682.800 281.600 683.600 290.200 ;
        RECT 0.400 280.400 689.200 281.600 ;
        RECT 1.200 275.800 2.000 280.400 ;
        RECT 4.400 275.800 5.200 280.400 ;
        RECT 7.600 275.800 8.400 280.400 ;
        RECT 14.000 275.800 14.800 280.400 ;
        RECT 17.200 275.800 18.000 280.400 ;
        RECT 25.200 275.800 26.000 280.400 ;
        RECT 28.400 275.800 29.200 280.400 ;
        RECT 31.600 275.800 32.400 280.400 ;
        RECT 34.800 275.800 35.600 280.400 ;
        RECT 4.400 271.800 5.200 272.400 ;
        RECT 7.800 271.800 8.600 272.000 ;
        RECT 36.400 271.800 37.200 280.400 ;
        RECT 39.600 271.800 40.400 280.400 ;
        RECT 42.800 271.800 43.600 280.400 ;
        RECT 46.000 271.800 46.800 280.400 ;
        RECT 49.200 271.800 50.000 280.400 ;
        RECT 51.400 275.800 52.200 280.400 ;
        RECT 55.600 271.800 56.400 280.400 ;
        RECT 57.200 275.800 58.000 280.400 ;
        RECT 60.400 271.800 61.200 280.400 ;
        RECT 64.600 275.800 65.400 280.400 ;
        RECT 66.800 275.800 67.600 280.400 ;
        RECT 70.000 275.800 70.800 280.400 ;
        RECT 73.200 275.800 74.000 280.400 ;
        RECT 76.400 275.800 77.200 280.400 ;
        RECT 84.400 275.800 85.200 280.400 ;
        RECT 87.600 275.800 88.400 280.400 ;
        RECT 94.000 275.800 94.800 280.400 ;
        RECT 97.200 275.800 98.000 280.400 ;
        RECT 100.400 275.800 101.200 280.400 ;
        RECT 103.600 275.800 104.400 280.400 ;
        RECT 106.800 275.800 107.600 280.400 ;
        RECT 108.400 275.800 109.200 280.400 ;
        RECT 111.600 275.800 112.400 280.400 ;
        RECT 93.800 271.800 94.600 272.000 ;
        RECT 97.200 271.800 98.000 272.400 ;
        RECT 118.000 271.800 118.800 280.400 ;
        RECT 121.200 271.800 122.000 280.400 ;
        RECT 124.400 271.800 125.200 280.400 ;
        RECT 127.600 271.800 128.400 280.400 ;
        RECT 130.800 271.800 131.600 280.400 ;
        RECT 134.000 275.800 134.800 280.400 ;
        RECT 135.600 275.800 136.400 280.400 ;
        RECT 138.800 275.800 139.600 280.400 ;
        RECT 142.000 275.800 142.800 280.400 ;
        RECT 145.200 275.800 146.000 280.400 ;
        RECT 153.200 275.800 154.000 280.400 ;
        RECT 156.400 275.800 157.200 280.400 ;
        RECT 162.800 275.800 163.600 280.400 ;
        RECT 166.000 275.800 166.800 280.400 ;
        RECT 169.200 275.800 170.000 280.400 ;
        RECT 170.800 275.800 171.600 280.400 ;
        RECT 174.000 275.800 174.800 280.400 ;
        RECT 176.200 275.800 177.000 280.400 ;
        RECT 162.600 271.800 163.600 272.000 ;
        RECT 166.000 271.800 166.800 272.400 ;
        RECT 180.400 271.800 181.200 280.400 ;
        RECT 182.000 271.800 182.800 280.400 ;
        RECT 185.200 273.000 186.000 280.400 ;
        RECT 188.400 275.800 189.200 280.400 ;
        RECT 191.600 275.800 192.400 280.400 ;
        RECT 194.800 275.800 195.600 280.400 ;
        RECT 198.000 275.800 198.800 280.400 ;
        RECT 206.000 275.800 206.800 280.400 ;
        RECT 209.200 275.800 210.000 280.400 ;
        RECT 215.600 275.800 216.400 280.400 ;
        RECT 218.800 275.800 219.600 280.400 ;
        RECT 222.000 275.800 222.800 280.400 ;
        RECT 215.400 271.800 216.200 272.000 ;
        RECT 218.800 271.800 219.600 272.400 ;
        RECT 226.800 271.800 227.600 280.400 ;
        RECT 228.400 275.800 229.200 280.400 ;
        RECT 231.600 275.800 232.400 280.400 ;
        RECT 234.800 275.800 235.600 280.400 ;
        RECT 238.000 275.800 238.800 280.400 ;
        RECT 246.000 275.800 246.800 280.400 ;
        RECT 249.200 275.800 250.000 280.400 ;
        RECT 255.600 275.800 256.400 280.400 ;
        RECT 258.800 275.800 259.600 280.400 ;
        RECT 262.000 275.800 262.800 280.400 ;
        RECT 270.000 273.000 270.800 280.400 ;
        RECT 255.400 271.800 256.200 272.000 ;
        RECT 258.800 271.800 259.600 272.400 ;
        RECT 273.200 271.800 274.000 280.400 ;
        RECT 276.400 276.200 277.200 280.400 ;
        RECT 279.600 275.800 280.400 280.400 ;
        RECT 281.800 275.800 282.600 280.400 ;
        RECT 286.000 271.800 286.800 280.400 ;
        RECT 287.600 271.800 288.400 280.400 ;
        RECT 291.800 275.800 292.600 280.400 ;
        RECT 294.000 275.800 294.800 280.400 ;
        RECT 297.200 275.800 298.000 280.400 ;
        RECT 300.400 275.800 301.200 280.400 ;
        RECT 306.800 275.800 307.600 280.400 ;
        RECT 310.000 275.800 310.800 280.400 ;
        RECT 318.000 275.800 318.800 280.400 ;
        RECT 321.200 275.800 322.000 280.400 ;
        RECT 324.400 275.800 325.200 280.400 ;
        RECT 327.600 275.800 328.400 280.400 ;
        RECT 329.200 275.800 330.000 280.400 ;
        RECT 332.400 275.800 333.200 280.400 ;
        RECT 297.200 271.800 298.000 272.400 ;
        RECT 300.400 271.800 301.400 272.000 ;
        RECT 335.600 271.800 336.400 280.400 ;
        RECT 337.200 275.800 338.000 280.400 ;
        RECT 340.400 275.800 341.200 280.400 ;
        RECT 342.000 275.800 342.800 280.400 ;
        RECT 345.200 275.800 346.000 280.400 ;
        RECT 347.400 275.800 348.200 280.400 ;
        RECT 351.600 271.800 352.400 280.400 ;
        RECT 354.800 275.800 355.600 280.400 ;
        RECT 356.400 271.800 357.200 280.400 ;
        RECT 360.600 275.800 361.400 280.400 ;
        RECT 363.400 275.800 364.200 280.400 ;
        RECT 367.600 271.800 368.400 280.400 ;
        RECT 370.800 275.800 371.600 280.400 ;
        RECT 372.400 275.800 373.200 280.400 ;
        RECT 375.600 275.800 376.400 280.400 ;
        RECT 377.200 275.800 378.000 280.400 ;
        RECT 380.400 276.200 381.200 280.400 ;
        RECT 383.600 271.800 384.400 280.400 ;
        RECT 386.800 271.800 387.600 280.400 ;
        RECT 390.000 271.800 390.800 280.400 ;
        RECT 393.200 273.000 394.000 280.400 ;
        RECT 396.400 271.800 397.200 280.400 ;
        RECT 399.600 273.000 400.400 280.400 ;
        RECT 402.800 275.800 403.600 280.400 ;
        RECT 406.000 276.200 406.800 280.400 ;
        RECT 410.800 272.200 411.600 280.400 ;
        RECT 416.000 271.800 416.800 280.400 ;
        RECT 425.200 275.800 426.000 280.400 ;
        RECT 426.800 275.800 427.600 280.400 ;
        RECT 430.000 275.800 430.800 280.400 ;
        RECT 433.200 275.800 434.000 280.400 ;
        RECT 439.600 275.800 440.400 280.400 ;
        RECT 442.800 275.800 443.600 280.400 ;
        RECT 450.800 275.800 451.600 280.400 ;
        RECT 454.000 275.800 454.800 280.400 ;
        RECT 457.200 275.800 458.000 280.400 ;
        RECT 460.400 275.800 461.200 280.400 ;
        RECT 462.000 275.800 462.800 280.400 ;
        RECT 465.200 275.800 466.000 280.400 ;
        RECT 468.400 275.800 469.200 280.400 ;
        RECT 471.600 275.800 472.400 280.400 ;
        RECT 478.000 275.800 478.800 280.400 ;
        RECT 481.200 275.800 482.000 280.400 ;
        RECT 489.200 275.800 490.000 280.400 ;
        RECT 492.400 275.800 493.200 280.400 ;
        RECT 495.600 275.800 496.400 280.400 ;
        RECT 498.800 275.800 499.600 280.400 ;
        RECT 500.400 275.800 501.200 280.400 ;
        RECT 505.200 275.800 506.000 280.400 ;
        RECT 430.000 271.800 430.800 272.400 ;
        RECT 433.400 271.800 434.200 272.000 ;
        RECT 468.400 271.800 469.200 272.400 ;
        RECT 471.800 271.800 472.600 272.000 ;
        RECT 506.800 271.800 507.600 280.400 ;
        RECT 510.000 271.800 510.800 280.400 ;
        RECT 513.200 271.800 514.000 280.400 ;
        RECT 516.400 271.800 517.200 280.400 ;
        RECT 519.600 271.800 520.400 280.400 ;
        RECT 521.800 275.800 522.600 280.400 ;
        RECT 526.000 271.800 526.800 280.400 ;
        RECT 527.600 271.800 528.400 280.400 ;
        RECT 530.800 273.000 531.600 280.400 ;
        RECT 534.000 271.800 534.800 280.400 ;
        RECT 538.200 275.800 539.000 280.400 ;
        RECT 542.000 272.000 542.800 280.400 ;
        RECT 547.600 275.800 548.400 280.400 ;
        RECT 550.800 275.800 551.600 280.400 ;
        RECT 556.400 271.800 557.200 280.400 ;
        RECT 559.600 275.800 560.400 280.400 ;
        RECT 562.800 275.800 563.600 280.400 ;
        RECT 565.600 271.800 566.400 280.400 ;
        RECT 570.800 272.200 571.600 280.400 ;
        RECT 580.000 271.800 580.800 280.400 ;
        RECT 585.200 272.200 586.000 280.400 ;
        RECT 589.000 275.800 589.800 280.400 ;
        RECT 593.200 271.800 594.000 280.400 ;
        RECT 595.400 275.800 596.200 280.400 ;
        RECT 599.600 271.800 600.400 280.400 ;
        RECT 602.800 273.000 603.600 280.400 ;
        RECT 606.000 271.800 606.800 280.400 ;
        RECT 607.600 271.800 608.400 280.400 ;
        RECT 611.800 275.800 612.600 280.400 ;
        RECT 614.600 275.800 615.400 280.400 ;
        RECT 618.800 271.800 619.600 280.400 ;
        RECT 622.000 275.800 622.800 280.400 ;
        RECT 623.600 275.800 624.400 280.400 ;
        RECT 626.800 275.800 627.600 280.400 ;
        RECT 630.000 272.200 630.800 280.400 ;
        RECT 635.200 271.800 636.000 280.400 ;
        RECT 638.000 271.800 638.800 280.400 ;
        RECT 642.200 275.800 643.000 280.400 ;
        RECT 644.400 271.800 645.200 280.400 ;
        RECT 648.600 275.800 649.400 280.400 ;
        RECT 652.000 271.800 652.800 280.400 ;
        RECT 657.200 272.200 658.000 280.400 ;
        RECT 661.000 275.800 661.800 280.400 ;
        RECT 665.200 271.800 666.000 280.400 ;
        RECT 668.400 271.800 669.200 280.400 ;
        RECT 674.000 275.800 674.800 280.400 ;
        RECT 677.200 275.800 678.000 280.400 ;
        RECT 682.800 272.000 683.600 280.400 ;
        RECT 4.400 271.200 31.400 271.800 ;
        RECT 30.600 271.000 31.400 271.200 ;
        RECT 71.000 271.200 98.000 271.800 ;
        RECT 139.800 271.200 166.800 271.800 ;
        RECT 192.600 271.200 219.600 271.800 ;
        RECT 232.600 271.200 259.600 271.800 ;
        RECT 297.200 271.200 324.200 271.800 ;
        RECT 430.000 271.200 457.000 271.800 ;
        RECT 468.400 271.200 495.400 271.800 ;
        RECT 71.000 271.000 71.800 271.200 ;
        RECT 139.800 271.000 140.600 271.200 ;
        RECT 192.600 271.000 193.400 271.200 ;
        RECT 232.600 271.000 233.400 271.200 ;
        RECT 323.400 271.000 324.200 271.200 ;
        RECT 456.200 271.000 457.000 271.200 ;
        RECT 494.600 271.000 495.400 271.200 ;
        RECT 18.200 250.800 19.000 251.000 ;
        RECT 53.400 250.800 54.200 251.000 ;
        RECT 91.800 250.800 92.600 251.000 ;
        RECT 214.600 250.800 215.400 251.000 ;
        RECT 18.200 250.200 45.200 250.800 ;
        RECT 53.400 250.200 80.400 250.800 ;
        RECT 91.800 250.200 118.800 250.800 ;
        RECT 188.400 250.200 215.400 250.800 ;
        RECT 227.800 250.800 228.600 251.000 ;
        RECT 277.400 250.800 278.200 251.000 ;
        RECT 453.000 250.800 453.800 251.000 ;
        RECT 541.000 250.800 541.800 251.000 ;
        RECT 227.800 250.200 254.800 250.800 ;
        RECT 277.400 250.200 304.400 250.800 ;
        RECT 426.800 250.200 453.800 250.800 ;
        RECT 514.800 250.200 541.800 250.800 ;
        RECT 41.000 250.000 41.800 250.200 ;
        RECT 44.400 249.600 45.200 250.200 ;
        RECT 76.200 250.000 77.000 250.200 ;
        RECT 79.600 249.600 80.400 250.200 ;
        RECT 114.600 250.000 115.600 250.200 ;
        RECT 118.000 249.600 118.800 250.200 ;
        RECT 2.800 241.600 3.600 249.000 ;
        RECT 7.600 241.600 8.400 249.000 ;
        RECT 10.800 241.600 11.600 246.200 ;
        RECT 14.000 241.600 14.800 246.200 ;
        RECT 17.200 241.600 18.000 246.200 ;
        RECT 20.400 241.600 21.200 246.200 ;
        RECT 23.600 241.600 24.400 246.200 ;
        RECT 31.600 241.600 32.400 246.200 ;
        RECT 34.800 241.600 35.600 246.200 ;
        RECT 41.200 241.600 42.000 246.200 ;
        RECT 44.400 241.600 45.200 246.200 ;
        RECT 47.600 241.600 48.400 246.200 ;
        RECT 49.200 241.600 50.000 246.200 ;
        RECT 52.400 241.600 53.200 246.200 ;
        RECT 55.600 241.600 56.400 246.200 ;
        RECT 58.800 241.600 59.600 246.200 ;
        RECT 66.800 241.600 67.600 246.200 ;
        RECT 70.000 241.600 70.800 246.200 ;
        RECT 76.400 241.600 77.200 246.200 ;
        RECT 79.600 241.600 80.400 246.200 ;
        RECT 82.800 241.600 83.600 246.200 ;
        RECT 86.000 241.600 86.800 246.200 ;
        RECT 87.600 241.600 88.400 246.200 ;
        RECT 90.800 241.600 91.600 246.200 ;
        RECT 94.000 241.600 94.800 246.200 ;
        RECT 97.200 241.600 98.000 246.200 ;
        RECT 105.200 241.600 106.000 246.200 ;
        RECT 108.400 241.600 109.200 246.200 ;
        RECT 114.800 241.600 115.600 246.200 ;
        RECT 118.000 241.600 118.800 246.200 ;
        RECT 121.200 241.600 122.000 246.200 ;
        RECT 127.600 241.600 128.400 250.200 ;
        RECT 130.800 241.600 131.600 250.200 ;
        RECT 134.000 241.600 134.800 250.200 ;
        RECT 137.200 241.600 138.000 250.200 ;
        RECT 140.400 241.600 141.200 250.200 ;
        RECT 142.000 241.600 142.800 250.200 ;
        RECT 145.200 241.600 146.000 250.200 ;
        RECT 148.400 241.600 149.200 250.200 ;
        RECT 151.600 241.600 152.400 250.200 ;
        RECT 154.800 241.600 155.600 250.200 ;
        RECT 156.400 241.600 157.200 246.200 ;
        RECT 160.800 241.600 161.600 250.200 ;
        RECT 166.000 241.600 166.800 249.800 ;
        RECT 169.200 241.600 170.000 246.200 ;
        RECT 173.600 241.600 174.400 250.200 ;
        RECT 178.800 241.600 179.600 249.800 ;
        RECT 188.400 249.600 189.200 250.200 ;
        RECT 191.600 250.000 192.600 250.200 ;
        RECT 250.600 250.000 251.600 250.200 ;
        RECT 254.000 249.600 254.800 250.200 ;
        RECT 182.000 241.600 182.800 246.200 ;
        RECT 185.200 241.600 186.000 246.200 ;
        RECT 188.400 241.600 189.200 246.200 ;
        RECT 191.600 241.600 192.400 246.200 ;
        RECT 198.000 241.600 198.800 246.200 ;
        RECT 201.200 241.600 202.000 246.200 ;
        RECT 209.200 241.600 210.000 246.200 ;
        RECT 212.400 241.600 213.200 246.200 ;
        RECT 215.600 241.600 216.400 246.200 ;
        RECT 218.800 241.600 219.600 246.200 ;
        RECT 220.400 241.600 221.200 246.200 ;
        RECT 223.600 241.600 224.400 246.200 ;
        RECT 226.800 241.600 227.600 246.200 ;
        RECT 230.000 241.600 230.800 246.200 ;
        RECT 233.200 241.600 234.000 246.200 ;
        RECT 241.200 241.600 242.000 246.200 ;
        RECT 244.400 241.600 245.200 246.200 ;
        RECT 250.800 241.600 251.600 246.200 ;
        RECT 254.000 241.600 254.800 246.200 ;
        RECT 257.200 241.600 258.000 246.200 ;
        RECT 258.800 241.600 259.600 246.200 ;
        RECT 266.800 241.600 267.600 250.200 ;
        RECT 300.200 250.000 301.200 250.200 ;
        RECT 303.600 249.600 304.400 250.200 ;
        RECT 271.000 241.600 271.800 246.200 ;
        RECT 273.200 241.600 274.000 246.200 ;
        RECT 276.400 241.600 277.200 246.200 ;
        RECT 279.600 241.600 280.400 246.200 ;
        RECT 282.800 241.600 283.600 246.200 ;
        RECT 290.800 241.600 291.600 246.200 ;
        RECT 294.000 241.600 294.800 246.200 ;
        RECT 300.400 241.600 301.200 246.200 ;
        RECT 303.600 241.600 304.400 246.200 ;
        RECT 306.800 241.600 307.600 246.200 ;
        RECT 308.400 241.600 309.200 246.200 ;
        RECT 311.600 241.600 312.400 245.800 ;
        RECT 314.800 241.600 315.600 246.200 ;
        RECT 318.000 241.600 318.800 245.800 ;
        RECT 321.800 241.600 322.600 246.200 ;
        RECT 326.000 241.600 326.800 250.200 ;
        RECT 327.600 241.600 328.400 250.200 ;
        RECT 334.000 241.600 334.800 250.200 ;
        RECT 335.600 241.600 336.400 246.200 ;
        RECT 338.800 241.600 339.600 246.200 ;
        RECT 340.400 241.600 341.200 250.200 ;
        RECT 343.600 241.600 344.400 250.200 ;
        RECT 346.800 241.600 347.600 250.200 ;
        RECT 350.000 241.600 350.800 250.200 ;
        RECT 353.200 241.600 354.000 250.200 ;
        RECT 355.400 241.600 356.200 246.200 ;
        RECT 359.600 241.600 360.400 250.200 ;
        RECT 361.200 241.600 362.000 250.200 ;
        RECT 367.600 241.600 368.400 250.200 ;
        RECT 369.200 241.600 370.000 246.200 ;
        RECT 372.400 241.600 373.200 246.200 ;
        RECT 374.000 241.600 374.800 250.200 ;
        RECT 378.200 241.600 379.000 246.200 ;
        RECT 380.400 241.600 381.200 250.200 ;
        RECT 385.200 241.600 386.000 246.200 ;
        RECT 388.400 241.600 389.200 245.800 ;
        RECT 393.200 241.600 394.000 246.200 ;
        RECT 394.800 241.600 395.600 246.200 ;
        RECT 398.000 241.600 398.800 246.200 ;
        RECT 401.200 241.600 402.000 249.000 ;
        RECT 404.400 241.600 405.200 250.200 ;
        RECT 408.200 241.600 409.000 250.200 ;
        RECT 426.800 249.600 427.600 250.200 ;
        RECT 430.000 250.000 431.000 250.200 ;
        RECT 412.400 241.600 413.200 246.200 ;
        RECT 415.600 241.600 416.400 245.800 ;
        RECT 423.600 241.600 424.400 246.200 ;
        RECT 426.800 241.600 427.600 246.200 ;
        RECT 430.000 241.600 430.800 246.200 ;
        RECT 436.400 241.600 437.200 246.200 ;
        RECT 439.600 241.600 440.400 246.200 ;
        RECT 447.600 241.600 448.400 246.200 ;
        RECT 450.800 241.600 451.600 246.200 ;
        RECT 454.000 241.600 454.800 246.200 ;
        RECT 457.200 241.600 458.000 246.200 ;
        RECT 460.400 241.600 461.200 249.800 ;
        RECT 465.600 241.600 466.400 250.200 ;
        RECT 470.000 241.600 470.800 246.200 ;
        RECT 471.600 241.600 472.400 250.200 ;
        RECT 474.800 241.600 475.600 250.200 ;
        RECT 478.000 241.600 478.800 250.200 ;
        RECT 481.200 241.600 482.000 250.200 ;
        RECT 484.400 241.600 485.200 250.200 ;
        RECT 487.600 241.600 488.400 249.800 ;
        RECT 492.800 241.600 493.600 250.200 ;
        RECT 497.200 241.600 498.000 246.200 ;
        RECT 500.400 241.600 501.200 249.800 ;
        RECT 505.600 241.600 506.400 250.200 ;
        RECT 514.800 249.600 515.600 250.200 ;
        RECT 518.000 250.000 519.000 250.200 ;
        RECT 510.000 241.600 510.800 246.200 ;
        RECT 511.600 241.600 512.400 246.200 ;
        RECT 514.800 241.600 515.600 246.200 ;
        RECT 518.000 241.600 518.800 246.200 ;
        RECT 524.400 241.600 525.200 246.200 ;
        RECT 527.600 241.600 528.400 246.200 ;
        RECT 535.600 241.600 536.400 246.200 ;
        RECT 538.800 241.600 539.600 246.200 ;
        RECT 542.000 241.600 542.800 246.200 ;
        RECT 545.200 241.600 546.000 246.200 ;
        RECT 548.400 241.600 549.200 250.200 ;
        RECT 554.000 241.600 554.800 246.200 ;
        RECT 557.200 241.600 558.000 246.200 ;
        RECT 562.800 241.600 563.600 250.000 ;
        RECT 566.000 241.600 566.800 250.200 ;
        RECT 570.200 241.600 571.000 246.200 ;
        RECT 577.800 241.600 578.600 246.200 ;
        RECT 582.000 241.600 582.800 250.200 ;
        RECT 585.200 241.600 586.000 250.000 ;
        RECT 590.800 241.600 591.600 246.200 ;
        RECT 594.000 241.600 594.800 246.200 ;
        RECT 599.600 241.600 600.400 250.200 ;
        RECT 604.400 241.600 605.200 250.200 ;
        RECT 610.000 241.600 610.800 246.200 ;
        RECT 613.200 241.600 614.000 246.200 ;
        RECT 618.800 241.600 619.600 250.000 ;
        RECT 623.600 241.600 624.400 250.200 ;
        RECT 629.200 241.600 630.000 246.200 ;
        RECT 632.400 241.600 633.200 246.200 ;
        RECT 638.000 241.600 638.800 250.000 ;
        RECT 641.800 241.600 642.600 246.200 ;
        RECT 646.000 241.600 646.800 250.200 ;
        RECT 648.200 241.600 649.000 246.200 ;
        RECT 652.400 241.600 653.200 250.200 ;
        RECT 655.200 241.600 656.000 250.200 ;
        RECT 660.400 241.600 661.200 249.800 ;
        RECT 663.600 241.600 664.400 250.200 ;
        RECT 667.800 241.600 668.600 246.200 ;
        RECT 671.600 241.600 672.400 250.000 ;
        RECT 677.200 241.600 678.000 246.200 ;
        RECT 680.400 241.600 681.200 246.200 ;
        RECT 686.000 241.600 686.800 250.200 ;
        RECT 0.400 240.400 689.200 241.600 ;
        RECT 1.200 231.800 2.000 240.400 ;
        RECT 4.400 231.800 5.200 240.400 ;
        RECT 7.600 231.800 8.400 240.400 ;
        RECT 10.800 231.800 11.600 240.400 ;
        RECT 14.000 231.800 14.800 240.400 ;
        RECT 17.200 235.800 18.000 240.400 ;
        RECT 18.800 235.800 19.600 240.400 ;
        RECT 22.000 235.800 22.800 240.400 ;
        RECT 25.200 235.800 26.000 240.400 ;
        RECT 28.400 235.800 29.200 240.400 ;
        RECT 31.600 235.800 32.400 240.400 ;
        RECT 39.600 235.800 40.400 240.400 ;
        RECT 42.800 235.800 43.600 240.400 ;
        RECT 49.200 235.800 50.000 240.400 ;
        RECT 52.400 235.800 53.200 240.400 ;
        RECT 55.600 235.800 56.400 240.400 ;
        RECT 49.000 231.800 49.800 232.000 ;
        RECT 52.400 231.800 53.200 232.400 ;
        RECT 58.400 231.800 59.200 240.400 ;
        RECT 63.600 232.200 64.400 240.400 ;
        RECT 66.800 231.800 67.600 240.400 ;
        RECT 74.800 233.000 75.600 240.400 ;
        RECT 79.600 232.200 80.400 240.400 ;
        RECT 84.800 231.800 85.600 240.400 ;
        RECT 87.600 235.800 88.400 240.400 ;
        RECT 90.800 235.800 91.600 240.400 ;
        RECT 94.000 235.800 94.800 240.400 ;
        RECT 100.400 235.800 101.200 240.400 ;
        RECT 103.600 235.800 104.400 240.400 ;
        RECT 111.600 235.800 112.400 240.400 ;
        RECT 114.800 235.800 115.600 240.400 ;
        RECT 118.000 235.800 118.800 240.400 ;
        RECT 121.200 235.800 122.000 240.400 ;
        RECT 90.800 231.800 91.600 232.400 ;
        RECT 94.200 231.800 95.000 232.000 ;
        RECT 130.800 231.800 131.600 240.400 ;
        RECT 135.600 233.000 136.400 240.400 ;
        RECT 138.800 235.800 139.600 240.400 ;
        RECT 142.000 235.800 142.800 240.400 ;
        RECT 145.200 235.800 146.000 240.400 ;
        RECT 148.400 235.800 149.200 240.400 ;
        RECT 156.400 235.800 157.200 240.400 ;
        RECT 159.600 235.800 160.400 240.400 ;
        RECT 166.000 235.800 166.800 240.400 ;
        RECT 169.200 235.800 170.000 240.400 ;
        RECT 172.400 235.800 173.200 240.400 ;
        RECT 174.000 235.800 174.800 240.400 ;
        RECT 165.800 231.800 166.800 232.000 ;
        RECT 169.200 231.800 170.000 232.400 ;
        RECT 178.400 231.800 179.200 240.400 ;
        RECT 183.600 232.200 184.400 240.400 ;
        RECT 186.800 235.800 187.600 240.400 ;
        RECT 190.000 235.800 190.800 240.400 ;
        RECT 193.200 235.800 194.000 240.400 ;
        RECT 196.400 235.800 197.200 240.400 ;
        RECT 204.400 235.800 205.200 240.400 ;
        RECT 207.600 235.800 208.400 240.400 ;
        RECT 214.000 235.800 214.800 240.400 ;
        RECT 217.200 235.800 218.000 240.400 ;
        RECT 220.400 235.800 221.200 240.400 ;
        RECT 213.800 231.800 214.800 232.000 ;
        RECT 217.200 231.800 218.000 232.400 ;
        RECT 223.200 231.800 224.000 240.400 ;
        RECT 228.400 232.200 229.200 240.400 ;
        RECT 232.200 235.800 233.000 240.400 ;
        RECT 236.400 231.800 237.200 240.400 ;
        RECT 238.000 235.800 238.800 240.400 ;
        RECT 241.200 235.800 242.000 240.400 ;
        RECT 244.400 235.800 245.200 240.400 ;
        RECT 250.800 235.800 251.600 240.400 ;
        RECT 254.000 235.800 254.800 240.400 ;
        RECT 262.000 235.800 262.800 240.400 ;
        RECT 265.200 235.800 266.000 240.400 ;
        RECT 268.400 235.800 269.200 240.400 ;
        RECT 271.600 235.800 272.400 240.400 ;
        RECT 241.200 231.800 242.000 232.400 ;
        RECT 244.400 231.800 245.400 232.000 ;
        RECT 280.200 231.800 281.000 240.400 ;
        RECT 286.000 235.800 286.800 240.400 ;
        RECT 287.600 231.800 288.400 240.400 ;
        RECT 290.800 235.800 291.600 240.400 ;
        RECT 294.000 235.800 294.800 240.400 ;
        RECT 296.200 235.800 297.000 240.400 ;
        RECT 300.400 231.800 301.200 240.400 ;
        RECT 302.000 235.800 302.800 240.400 ;
        RECT 305.200 231.800 306.000 240.400 ;
        RECT 309.400 235.800 310.200 240.400 ;
        RECT 311.600 231.800 312.400 240.400 ;
        RECT 315.800 235.800 316.600 240.400 ;
        RECT 318.000 235.800 318.800 240.400 ;
        RECT 321.200 235.800 322.000 240.400 ;
        RECT 324.400 235.800 325.200 240.400 ;
        RECT 330.800 235.800 331.600 240.400 ;
        RECT 334.000 235.800 334.800 240.400 ;
        RECT 342.000 235.800 342.800 240.400 ;
        RECT 345.200 235.800 346.000 240.400 ;
        RECT 348.400 235.800 349.200 240.400 ;
        RECT 351.600 235.800 352.400 240.400 ;
        RECT 321.200 231.800 322.000 232.400 ;
        RECT 324.400 231.800 325.400 232.000 ;
        RECT 353.200 231.800 354.000 240.400 ;
        RECT 356.400 235.800 357.200 240.400 ;
        RECT 359.600 235.800 360.400 240.400 ;
        RECT 361.800 235.800 362.600 240.400 ;
        RECT 366.000 231.800 366.800 240.400 ;
        RECT 369.200 233.000 370.000 240.400 ;
        RECT 372.400 231.800 373.200 240.400 ;
        RECT 375.600 236.200 376.400 240.400 ;
        RECT 378.800 235.800 379.600 240.400 ;
        RECT 382.000 236.200 382.800 240.400 ;
        RECT 385.200 235.800 386.000 240.400 ;
        RECT 386.800 235.800 387.600 240.400 ;
        RECT 390.000 235.800 390.800 240.400 ;
        RECT 393.200 235.800 394.000 240.400 ;
        RECT 399.600 235.800 400.400 240.400 ;
        RECT 402.800 235.800 403.600 240.400 ;
        RECT 410.800 235.800 411.600 240.400 ;
        RECT 414.000 235.800 414.800 240.400 ;
        RECT 417.200 235.800 418.000 240.400 ;
        RECT 420.400 235.800 421.200 240.400 ;
        RECT 390.000 231.800 390.800 232.400 ;
        RECT 428.400 232.200 429.200 240.400 ;
        RECT 393.400 231.800 394.200 232.000 ;
        RECT 433.600 231.800 434.400 240.400 ;
        RECT 436.400 235.800 437.200 240.400 ;
        RECT 439.600 231.800 440.400 240.400 ;
        RECT 442.800 231.800 443.600 240.400 ;
        RECT 446.000 231.800 446.800 240.400 ;
        RECT 449.200 231.800 450.000 240.400 ;
        RECT 452.400 231.800 453.200 240.400 ;
        RECT 454.000 235.800 454.800 240.400 ;
        RECT 457.200 235.800 458.000 240.400 ;
        RECT 460.400 235.800 461.200 240.400 ;
        RECT 466.800 235.800 467.600 240.400 ;
        RECT 470.000 235.800 470.800 240.400 ;
        RECT 478.000 235.800 478.800 240.400 ;
        RECT 481.200 235.800 482.000 240.400 ;
        RECT 484.400 235.800 485.200 240.400 ;
        RECT 487.600 235.800 488.400 240.400 ;
        RECT 457.200 231.800 458.000 232.400 ;
        RECT 490.800 232.200 491.600 240.400 ;
        RECT 460.400 231.800 461.400 232.000 ;
        RECT 496.000 231.800 496.800 240.400 ;
        RECT 500.400 235.800 501.200 240.400 ;
        RECT 502.000 235.800 502.800 240.400 ;
        RECT 505.200 235.800 506.000 240.400 ;
        RECT 508.400 235.800 509.200 240.400 ;
        RECT 514.800 235.800 515.600 240.400 ;
        RECT 518.000 235.800 518.800 240.400 ;
        RECT 526.000 235.800 526.800 240.400 ;
        RECT 529.200 235.800 530.000 240.400 ;
        RECT 532.400 235.800 533.200 240.400 ;
        RECT 535.600 235.800 536.400 240.400 ;
        RECT 538.800 235.800 539.600 240.400 ;
        RECT 540.400 235.800 541.200 240.400 ;
        RECT 505.200 231.800 506.000 232.400 ;
        RECT 543.600 232.200 544.400 240.400 ;
        RECT 546.800 235.800 547.600 240.400 ;
        RECT 551.600 233.000 552.400 240.400 ;
        RECT 555.400 235.800 556.200 240.400 ;
        RECT 508.400 231.800 509.400 232.000 ;
        RECT 559.600 231.800 560.400 240.400 ;
        RECT 561.200 235.800 562.000 240.400 ;
        RECT 564.400 235.800 565.200 240.400 ;
        RECT 566.000 235.800 566.800 240.400 ;
        RECT 569.200 235.800 570.000 240.400 ;
        RECT 575.600 235.800 576.400 240.400 ;
        RECT 578.800 235.800 579.600 240.400 ;
        RECT 582.000 235.800 582.800 240.400 ;
        RECT 585.200 235.800 586.000 240.400 ;
        RECT 593.200 235.800 594.000 240.400 ;
        RECT 596.400 235.800 597.200 240.400 ;
        RECT 602.800 235.800 603.600 240.400 ;
        RECT 606.000 235.800 606.800 240.400 ;
        RECT 609.200 235.800 610.000 240.400 ;
        RECT 602.600 231.800 603.400 232.000 ;
        RECT 606.000 231.800 606.800 232.400 ;
        RECT 612.400 231.800 613.200 240.400 ;
        RECT 618.000 235.800 618.800 240.400 ;
        RECT 621.200 235.800 622.000 240.400 ;
        RECT 626.800 232.000 627.600 240.400 ;
        RECT 630.000 235.800 630.800 240.400 ;
        RECT 633.200 235.800 634.000 240.400 ;
        RECT 636.400 235.800 637.200 240.400 ;
        RECT 642.800 235.800 643.600 240.400 ;
        RECT 646.000 235.800 646.800 240.400 ;
        RECT 654.000 235.800 654.800 240.400 ;
        RECT 657.200 235.800 658.000 240.400 ;
        RECT 660.400 235.800 661.200 240.400 ;
        RECT 663.600 235.800 664.400 240.400 ;
        RECT 665.200 235.800 666.000 240.400 ;
        RECT 633.200 231.800 634.000 232.400 ;
        RECT 670.000 232.000 670.800 240.400 ;
        RECT 675.600 235.800 676.400 240.400 ;
        RECT 678.800 235.800 679.600 240.400 ;
        RECT 636.600 231.800 637.400 232.000 ;
        RECT 684.400 231.800 685.200 240.400 ;
        RECT 26.200 231.200 53.200 231.800 ;
        RECT 90.800 231.200 117.800 231.800 ;
        RECT 26.200 231.000 27.000 231.200 ;
        RECT 117.000 231.000 117.800 231.200 ;
        RECT 143.000 231.200 170.000 231.800 ;
        RECT 191.000 231.200 218.000 231.800 ;
        RECT 241.200 231.200 268.200 231.800 ;
        RECT 321.200 231.200 348.200 231.800 ;
        RECT 390.000 231.200 417.000 231.800 ;
        RECT 457.200 231.200 484.200 231.800 ;
        RECT 505.200 231.200 532.200 231.800 ;
        RECT 143.000 231.000 143.800 231.200 ;
        RECT 191.000 231.000 191.800 231.200 ;
        RECT 267.400 231.000 268.200 231.200 ;
        RECT 347.400 231.000 348.200 231.200 ;
        RECT 416.200 231.000 417.000 231.200 ;
        RECT 483.400 231.000 484.200 231.200 ;
        RECT 531.400 231.000 532.200 231.200 ;
        RECT 579.800 231.200 606.800 231.800 ;
        RECT 633.200 231.200 660.200 231.800 ;
        RECT 579.800 231.000 580.600 231.200 ;
        RECT 659.400 231.000 660.200 231.200 ;
        RECT 458.800 212.000 459.600 212.600 ;
        RECT 470.000 212.000 470.800 212.400 ;
        RECT 476.400 212.000 477.200 212.400 ;
        RECT 481.400 212.000 482.200 212.200 ;
        RECT 458.800 211.400 482.200 212.000 ;
        RECT 40.200 210.800 41.000 211.000 ;
        RECT 14.000 210.200 41.000 210.800 ;
        RECT 64.600 210.800 65.400 211.000 ;
        RECT 122.200 210.800 123.000 211.000 ;
        RECT 157.400 210.800 158.200 211.000 ;
        RECT 217.800 210.800 218.600 211.000 ;
        RECT 294.600 210.800 295.400 211.000 ;
        RECT 64.600 210.200 91.600 210.800 ;
        RECT 122.200 210.200 149.200 210.800 ;
        RECT 157.400 210.200 184.400 210.800 ;
        RECT 1.200 201.600 2.000 206.200 ;
        RECT 4.400 201.600 5.200 210.200 ;
        RECT 14.000 209.600 14.800 210.200 ;
        RECT 17.400 210.000 18.200 210.200 ;
        RECT 8.600 201.600 9.400 206.200 ;
        RECT 10.800 201.600 11.600 206.200 ;
        RECT 14.000 201.600 14.800 206.200 ;
        RECT 17.200 201.600 18.000 206.200 ;
        RECT 23.600 201.600 24.400 206.200 ;
        RECT 26.800 201.600 27.600 206.200 ;
        RECT 34.800 201.600 35.600 206.200 ;
        RECT 38.000 201.600 38.800 206.200 ;
        RECT 41.200 201.600 42.000 206.200 ;
        RECT 44.400 201.600 45.200 206.200 ;
        RECT 46.000 201.600 46.800 210.200 ;
        RECT 49.200 201.600 50.000 210.200 ;
        RECT 52.400 201.600 53.200 210.200 ;
        RECT 55.600 201.600 56.400 210.200 ;
        RECT 58.800 201.600 59.600 210.200 ;
        RECT 87.400 210.000 88.200 210.200 ;
        RECT 90.800 209.600 91.600 210.200 ;
        RECT 60.400 201.600 61.200 206.200 ;
        RECT 63.600 201.600 64.400 206.200 ;
        RECT 66.800 201.600 67.600 206.200 ;
        RECT 70.000 201.600 70.800 206.200 ;
        RECT 78.000 201.600 78.800 206.200 ;
        RECT 81.200 201.600 82.000 206.200 ;
        RECT 87.600 201.600 88.400 206.200 ;
        RECT 90.800 201.600 91.600 206.200 ;
        RECT 94.000 201.600 94.800 206.200 ;
        RECT 95.600 201.600 96.400 210.200 ;
        RECT 98.800 201.600 99.600 210.200 ;
        RECT 102.000 201.600 102.800 210.200 ;
        RECT 105.200 201.600 106.000 210.200 ;
        RECT 108.400 201.600 109.200 210.200 ;
        RECT 145.000 210.000 146.000 210.200 ;
        RECT 148.400 209.600 149.200 210.200 ;
        RECT 180.200 210.000 181.000 210.200 ;
        RECT 183.600 209.600 184.400 210.200 ;
        RECT 191.600 210.200 218.600 210.800 ;
        RECT 268.400 210.200 295.400 210.800 ;
        RECT 359.000 210.800 359.800 211.000 ;
        RECT 437.000 210.800 437.800 211.000 ;
        RECT 517.000 210.800 517.800 211.000 ;
        RECT 359.000 210.200 386.000 210.800 ;
        RECT 410.800 210.200 437.800 210.800 ;
        RECT 490.800 210.200 517.800 210.800 ;
        RECT 615.000 210.800 615.800 211.000 ;
        RECT 615.000 210.200 642.000 210.800 ;
        RECT 191.600 209.600 192.400 210.200 ;
        RECT 195.000 210.000 195.800 210.200 ;
        RECT 116.400 201.600 117.200 206.200 ;
        RECT 118.000 201.600 118.800 206.200 ;
        RECT 121.200 201.600 122.000 206.200 ;
        RECT 124.400 201.600 125.200 206.200 ;
        RECT 127.600 201.600 128.400 206.200 ;
        RECT 135.600 201.600 136.400 206.200 ;
        RECT 138.800 201.600 139.600 206.200 ;
        RECT 145.200 201.600 146.000 206.200 ;
        RECT 148.400 201.600 149.200 206.200 ;
        RECT 151.600 201.600 152.400 206.200 ;
        RECT 153.200 201.600 154.000 206.200 ;
        RECT 156.400 201.600 157.200 206.200 ;
        RECT 159.600 201.600 160.400 206.200 ;
        RECT 162.800 201.600 163.600 206.200 ;
        RECT 170.800 201.600 171.600 206.200 ;
        RECT 174.000 201.600 174.800 206.200 ;
        RECT 180.400 201.600 181.200 206.200 ;
        RECT 183.600 201.600 184.400 206.200 ;
        RECT 186.800 201.600 187.600 206.200 ;
        RECT 188.400 201.600 189.200 206.200 ;
        RECT 191.600 201.600 192.400 206.200 ;
        RECT 194.800 201.600 195.600 206.200 ;
        RECT 201.200 201.600 202.000 206.200 ;
        RECT 204.400 201.600 205.200 206.200 ;
        RECT 212.400 201.600 213.200 206.200 ;
        RECT 215.600 201.600 216.400 206.200 ;
        RECT 218.800 201.600 219.600 206.200 ;
        RECT 222.000 201.600 222.800 206.200 ;
        RECT 223.600 201.600 224.400 210.200 ;
        RECT 231.600 201.600 232.400 209.000 ;
        RECT 234.800 201.600 235.600 206.200 ;
        RECT 238.000 201.600 238.800 206.200 ;
        RECT 239.600 201.600 240.400 210.200 ;
        RECT 244.400 201.600 245.200 210.200 ;
        RECT 247.600 201.600 248.400 209.000 ;
        RECT 250.800 201.600 251.600 210.200 ;
        RECT 268.400 209.600 269.200 210.200 ;
        RECT 271.800 210.000 272.600 210.200 ;
        RECT 254.000 201.600 254.800 209.000 ;
        RECT 258.800 201.600 259.600 206.200 ;
        RECT 265.200 201.600 266.000 206.200 ;
        RECT 268.400 201.600 269.200 206.200 ;
        RECT 271.600 201.600 272.400 206.200 ;
        RECT 278.000 201.600 278.800 206.200 ;
        RECT 281.200 201.600 282.000 206.200 ;
        RECT 289.200 201.600 290.000 206.200 ;
        RECT 292.400 201.600 293.200 206.200 ;
        RECT 295.600 201.600 296.400 206.200 ;
        RECT 298.800 201.600 299.600 206.200 ;
        RECT 300.400 201.600 301.200 206.200 ;
        RECT 303.600 201.600 304.400 206.200 ;
        RECT 305.200 201.600 306.000 210.200 ;
        RECT 309.400 201.600 310.200 206.200 ;
        RECT 311.600 201.600 312.400 210.200 ;
        RECT 314.800 201.600 315.600 210.200 ;
        RECT 316.400 201.600 317.200 210.200 ;
        RECT 319.600 201.600 320.400 210.200 ;
        RECT 322.800 201.600 323.600 209.000 ;
        RECT 326.000 201.600 326.800 210.200 ;
        RECT 328.200 201.600 329.000 206.200 ;
        RECT 332.400 201.600 333.200 210.200 ;
        RECT 334.000 201.600 334.800 206.200 ;
        RECT 337.200 201.600 338.000 206.200 ;
        RECT 338.800 201.600 339.600 206.200 ;
        RECT 342.000 201.600 342.800 206.200 ;
        RECT 343.600 201.600 344.400 210.200 ;
        RECT 381.800 210.000 382.800 210.200 ;
        RECT 385.200 209.600 386.000 210.200 ;
        RECT 347.800 201.600 348.600 206.200 ;
        RECT 350.000 201.600 350.800 206.200 ;
        RECT 353.200 201.600 354.000 206.200 ;
        RECT 354.800 201.600 355.600 206.200 ;
        RECT 358.000 201.600 358.800 206.200 ;
        RECT 361.200 201.600 362.000 206.200 ;
        RECT 364.400 201.600 365.200 206.200 ;
        RECT 372.400 201.600 373.200 206.200 ;
        RECT 375.600 201.600 376.400 206.200 ;
        RECT 382.000 201.600 382.800 206.200 ;
        RECT 385.200 201.600 386.000 206.200 ;
        RECT 388.400 201.600 389.200 206.200 ;
        RECT 390.000 201.600 390.800 210.200 ;
        RECT 393.200 201.600 394.000 209.000 ;
        RECT 396.400 201.600 397.200 210.200 ;
        RECT 410.800 209.600 411.600 210.200 ;
        RECT 414.000 210.000 415.000 210.200 ;
        RECT 400.600 201.600 401.400 206.200 ;
        RECT 407.600 201.600 408.400 206.200 ;
        RECT 410.800 201.600 411.600 206.200 ;
        RECT 414.000 201.600 414.800 206.200 ;
        RECT 420.400 201.600 421.200 206.200 ;
        RECT 423.600 201.600 424.400 206.200 ;
        RECT 431.600 201.600 432.400 206.200 ;
        RECT 434.800 201.600 435.600 206.200 ;
        RECT 438.000 201.600 438.800 206.200 ;
        RECT 441.200 201.600 442.000 206.200 ;
        RECT 444.400 201.600 445.200 209.000 ;
        RECT 447.600 201.600 448.400 210.200 ;
        RECT 490.800 209.600 491.600 210.200 ;
        RECT 494.000 210.000 495.000 210.200 ;
        RECT 449.200 201.600 450.000 206.200 ;
        RECT 452.400 201.600 453.200 206.200 ;
        RECT 455.600 201.600 456.400 206.200 ;
        RECT 458.800 201.600 459.600 206.200 ;
        RECT 466.800 201.600 467.600 206.200 ;
        RECT 470.000 201.600 470.800 206.400 ;
        RECT 476.400 201.600 477.200 206.200 ;
        RECT 479.600 201.600 480.400 206.200 ;
        RECT 482.800 201.600 483.600 206.200 ;
        RECT 484.400 201.600 485.200 206.200 ;
        RECT 487.600 201.600 488.400 206.200 ;
        RECT 490.800 201.600 491.600 206.200 ;
        RECT 494.000 201.600 494.800 206.200 ;
        RECT 500.400 201.600 501.200 206.200 ;
        RECT 503.600 201.600 504.400 206.200 ;
        RECT 511.600 201.600 512.400 206.200 ;
        RECT 514.800 201.600 515.600 206.200 ;
        RECT 518.000 201.600 518.800 206.200 ;
        RECT 521.200 201.600 522.000 206.200 ;
        RECT 522.800 201.600 523.600 210.200 ;
        RECT 527.000 201.600 527.800 206.200 ;
        RECT 529.200 201.600 530.000 206.200 ;
        RECT 532.400 201.600 533.200 206.200 ;
        RECT 534.600 201.600 535.400 206.200 ;
        RECT 538.800 201.600 539.600 210.200 ;
        RECT 540.400 201.600 541.200 210.200 ;
        RECT 548.400 201.600 549.200 210.200 ;
        RECT 550.000 201.600 550.800 210.200 ;
        RECT 554.200 201.600 555.000 206.200 ;
        RECT 559.600 201.600 560.400 209.000 ;
        RECT 564.400 201.600 565.200 205.800 ;
        RECT 567.600 201.600 568.400 206.200 ;
        RECT 576.200 201.600 577.000 210.200 ;
        RECT 582.000 202.200 583.000 208.800 ;
        RECT 582.200 201.600 583.000 202.200 ;
        RECT 588.200 201.600 589.200 208.800 ;
        RECT 593.200 201.600 594.000 209.800 ;
        RECT 598.400 201.600 599.200 210.200 ;
        RECT 602.800 201.600 603.600 209.800 ;
        RECT 608.000 201.600 608.800 210.200 ;
        RECT 637.800 210.000 638.600 210.200 ;
        RECT 641.200 209.600 642.000 210.200 ;
        RECT 610.800 201.600 611.600 206.200 ;
        RECT 614.000 201.600 614.800 206.200 ;
        RECT 617.200 201.600 618.000 206.200 ;
        RECT 620.400 201.600 621.200 206.200 ;
        RECT 628.400 201.600 629.200 206.200 ;
        RECT 631.600 201.600 632.400 206.200 ;
        RECT 638.000 201.600 638.800 206.200 ;
        RECT 641.200 201.600 642.000 206.200 ;
        RECT 644.400 201.600 645.200 206.200 ;
        RECT 647.600 202.200 648.600 208.800 ;
        RECT 647.800 201.600 648.600 202.200 ;
        RECT 653.800 201.600 654.800 208.800 ;
        RECT 657.200 201.600 658.000 210.200 ;
        RECT 660.400 201.600 661.200 210.200 ;
        RECT 663.600 201.600 664.400 210.200 ;
        RECT 666.800 201.600 667.600 210.200 ;
        RECT 670.000 201.600 670.800 210.200 ;
        RECT 671.600 201.600 672.400 210.200 ;
        RECT 674.800 201.600 675.600 210.200 ;
        RECT 678.000 201.600 678.800 210.200 ;
        RECT 681.200 201.600 682.000 210.200 ;
        RECT 684.400 201.600 685.200 210.200 ;
        RECT 0.400 200.400 689.200 201.600 ;
        RECT 1.200 195.800 2.000 200.400 ;
        RECT 4.400 191.800 5.200 200.400 ;
        RECT 8.600 195.800 9.400 200.400 ;
        RECT 11.400 195.800 12.200 200.400 ;
        RECT 15.600 191.800 16.400 200.400 ;
        RECT 17.200 195.800 18.000 200.400 ;
        RECT 20.400 195.800 21.200 200.400 ;
        RECT 23.600 195.800 24.400 200.400 ;
        RECT 30.000 195.800 30.800 200.400 ;
        RECT 33.200 195.800 34.000 200.400 ;
        RECT 41.200 195.800 42.000 200.400 ;
        RECT 44.400 195.800 45.200 200.400 ;
        RECT 47.600 195.800 48.400 200.400 ;
        RECT 50.800 195.800 51.600 200.400 ;
        RECT 53.000 195.800 53.800 200.400 ;
        RECT 20.400 191.800 21.200 192.400 ;
        RECT 23.800 191.800 24.600 192.000 ;
        RECT 57.200 191.800 58.000 200.400 ;
        RECT 61.400 191.800 62.200 200.400 ;
        RECT 65.200 195.800 66.000 200.400 ;
        RECT 68.400 195.800 69.200 200.400 ;
        RECT 70.000 195.800 70.800 200.400 ;
        RECT 73.800 195.800 74.600 200.400 ;
        RECT 78.000 191.800 78.800 200.400 ;
        RECT 80.200 195.800 81.000 200.400 ;
        RECT 84.400 191.800 85.200 200.400 ;
        RECT 87.600 192.000 88.400 200.400 ;
        RECT 93.200 195.800 94.000 200.400 ;
        RECT 96.400 195.800 97.200 200.400 ;
        RECT 102.000 191.800 102.800 200.400 ;
        RECT 105.200 195.800 106.000 200.400 ;
        RECT 108.400 195.800 109.200 200.400 ;
        RECT 115.400 195.800 116.200 200.400 ;
        RECT 119.600 191.800 120.400 200.400 ;
        RECT 122.800 192.000 123.600 200.400 ;
        RECT 128.400 195.800 129.200 200.400 ;
        RECT 131.600 195.800 132.400 200.400 ;
        RECT 137.200 191.800 138.000 200.400 ;
        RECT 142.000 195.800 142.800 200.400 ;
        RECT 145.200 192.000 146.000 200.400 ;
        RECT 150.800 195.800 151.600 200.400 ;
        RECT 154.000 195.800 154.800 200.400 ;
        RECT 159.600 191.800 160.400 200.400 ;
        RECT 164.400 192.000 165.200 200.400 ;
        RECT 170.000 195.800 170.800 200.400 ;
        RECT 173.200 195.800 174.000 200.400 ;
        RECT 178.800 191.800 179.600 200.400 ;
        RECT 182.000 195.800 182.800 200.400 ;
        RECT 185.200 195.800 186.000 200.400 ;
        RECT 188.400 195.800 189.200 200.400 ;
        RECT 191.600 195.800 192.400 200.400 ;
        RECT 199.600 195.800 200.400 200.400 ;
        RECT 202.800 195.800 203.600 200.400 ;
        RECT 209.200 195.800 210.000 200.400 ;
        RECT 212.400 195.800 213.200 200.400 ;
        RECT 215.600 195.800 216.400 200.400 ;
        RECT 209.000 191.800 209.800 192.000 ;
        RECT 212.400 191.800 213.200 192.400 ;
        RECT 220.400 191.800 221.200 200.400 ;
        RECT 225.200 193.000 226.000 200.400 ;
        RECT 228.400 195.800 229.200 200.400 ;
        RECT 231.600 195.800 232.400 200.400 ;
        RECT 234.800 195.800 235.600 200.400 ;
        RECT 238.000 195.800 238.800 200.400 ;
        RECT 246.000 195.800 246.800 200.400 ;
        RECT 249.200 195.800 250.000 200.400 ;
        RECT 255.600 195.800 256.400 200.400 ;
        RECT 258.800 195.800 259.600 200.400 ;
        RECT 262.000 195.800 262.800 200.400 ;
        RECT 268.400 195.800 269.200 200.400 ;
        RECT 271.600 195.800 272.400 200.400 ;
        RECT 274.800 195.800 275.600 200.400 ;
        RECT 278.000 195.800 278.800 200.400 ;
        RECT 286.000 195.800 286.800 200.400 ;
        RECT 289.200 195.800 290.000 200.400 ;
        RECT 295.600 195.800 296.400 200.400 ;
        RECT 298.800 195.800 299.600 200.400 ;
        RECT 302.000 195.800 302.800 200.400 ;
        RECT 305.200 195.800 306.000 200.400 ;
        RECT 306.800 195.800 307.600 200.400 ;
        RECT 310.000 195.800 310.800 200.400 ;
        RECT 313.200 195.800 314.000 200.400 ;
        RECT 319.600 195.800 320.400 200.400 ;
        RECT 322.800 195.800 323.600 200.400 ;
        RECT 330.800 195.800 331.600 200.400 ;
        RECT 334.000 195.800 334.800 200.400 ;
        RECT 337.200 195.800 338.000 200.400 ;
        RECT 340.400 195.800 341.200 200.400 ;
        RECT 342.000 195.800 342.800 200.400 ;
        RECT 345.200 195.800 346.000 200.400 ;
        RECT 346.800 195.800 347.600 200.400 ;
        RECT 350.000 195.800 350.800 200.400 ;
        RECT 255.400 191.800 256.200 192.000 ;
        RECT 258.800 191.800 259.600 192.400 ;
        RECT 295.400 191.800 296.200 192.000 ;
        RECT 298.800 191.800 299.600 192.400 ;
        RECT 20.400 191.200 47.400 191.800 ;
        RECT 46.600 191.000 47.400 191.200 ;
        RECT 186.200 191.200 213.200 191.800 ;
        RECT 232.600 191.200 259.600 191.800 ;
        RECT 272.600 191.200 299.600 191.800 ;
        RECT 310.000 191.800 310.800 192.400 ;
        RECT 313.400 191.800 314.200 192.000 ;
        RECT 351.600 191.800 352.400 200.400 ;
        RECT 354.800 191.800 355.600 200.400 ;
        RECT 358.000 191.800 358.800 200.400 ;
        RECT 361.200 191.800 362.000 200.400 ;
        RECT 364.400 191.800 365.200 200.400 ;
        RECT 367.600 191.800 368.400 200.400 ;
        RECT 369.200 191.800 370.000 200.400 ;
        RECT 372.400 195.800 373.200 200.400 ;
        RECT 375.600 195.800 376.400 200.400 ;
        RECT 377.200 195.800 378.000 200.400 ;
        RECT 380.400 195.800 381.200 200.400 ;
        RECT 382.000 191.800 382.800 200.400 ;
        RECT 388.400 191.800 389.200 200.400 ;
        RECT 390.000 195.800 390.800 200.400 ;
        RECT 393.200 195.800 394.000 200.400 ;
        RECT 394.800 195.800 395.600 200.400 ;
        RECT 398.000 196.200 398.800 200.400 ;
        RECT 401.200 195.800 402.000 200.400 ;
        RECT 404.400 196.200 405.200 200.400 ;
        RECT 407.600 191.800 408.400 200.400 ;
        RECT 410.800 191.800 411.600 200.400 ;
        RECT 414.000 191.800 414.800 200.400 ;
        RECT 417.200 191.800 418.000 200.400 ;
        RECT 420.400 191.800 421.200 200.400 ;
        RECT 426.800 195.800 427.600 200.400 ;
        RECT 430.000 195.800 430.800 200.400 ;
        RECT 433.200 195.800 434.000 200.400 ;
        RECT 436.400 195.800 437.200 200.400 ;
        RECT 444.400 195.800 445.200 200.400 ;
        RECT 447.600 195.800 448.400 200.400 ;
        RECT 454.000 195.800 454.800 200.400 ;
        RECT 457.200 195.800 458.000 200.400 ;
        RECT 460.400 195.800 461.200 200.400 ;
        RECT 462.600 195.800 463.400 200.400 ;
        RECT 453.800 191.800 454.800 192.000 ;
        RECT 457.200 191.800 458.000 192.400 ;
        RECT 466.800 191.800 467.600 200.400 ;
        RECT 468.400 191.800 469.200 200.400 ;
        RECT 471.600 191.800 472.400 200.400 ;
        RECT 474.800 191.800 475.600 200.400 ;
        RECT 478.000 191.800 478.800 200.400 ;
        RECT 481.200 191.800 482.000 200.400 ;
        RECT 484.400 192.200 485.200 200.400 ;
        RECT 489.600 191.800 490.400 200.400 ;
        RECT 494.000 195.800 494.800 200.400 ;
        RECT 495.600 191.800 496.400 200.400 ;
        RECT 498.800 191.800 499.600 200.400 ;
        RECT 502.000 191.800 502.800 200.400 ;
        RECT 505.200 191.800 506.000 200.400 ;
        RECT 508.400 191.800 509.200 200.400 ;
        RECT 511.600 193.000 512.400 200.400 ;
        RECT 514.800 191.800 515.600 200.400 ;
        RECT 519.000 191.800 519.800 200.400 ;
        RECT 522.800 191.800 523.600 200.400 ;
        RECT 529.400 199.800 530.200 200.400 ;
        RECT 529.200 193.200 530.200 199.800 ;
        RECT 535.400 193.200 536.400 200.400 ;
        RECT 540.400 192.000 541.200 200.400 ;
        RECT 546.000 195.800 546.800 200.400 ;
        RECT 549.200 195.800 550.000 200.400 ;
        RECT 554.800 191.800 555.600 200.400 ;
        RECT 558.000 191.800 558.800 200.400 ;
        RECT 562.200 195.800 563.000 200.400 ;
        RECT 565.000 195.800 565.800 200.400 ;
        RECT 569.200 191.800 570.000 200.400 ;
        RECT 577.200 192.200 578.000 200.400 ;
        RECT 582.400 191.800 583.200 200.400 ;
        RECT 585.200 191.800 586.000 200.400 ;
        RECT 589.400 195.800 590.200 200.400 ;
        RECT 592.200 195.800 593.000 200.400 ;
        RECT 596.400 191.800 597.200 200.400 ;
        RECT 599.600 191.800 600.400 200.400 ;
        RECT 605.200 195.800 606.000 200.400 ;
        RECT 608.400 195.800 609.200 200.400 ;
        RECT 614.000 192.000 614.800 200.400 ;
        RECT 617.200 191.800 618.000 200.400 ;
        RECT 621.400 195.800 622.200 200.400 ;
        RECT 623.600 191.800 624.400 200.400 ;
        RECT 627.800 195.800 628.600 200.400 ;
        RECT 631.200 191.800 632.000 200.400 ;
        RECT 636.400 192.200 637.200 200.400 ;
        RECT 641.200 191.800 642.000 200.400 ;
        RECT 646.800 195.800 647.600 200.400 ;
        RECT 650.000 195.800 650.800 200.400 ;
        RECT 655.600 192.000 656.400 200.400 ;
        RECT 658.800 191.800 659.600 200.400 ;
        RECT 663.600 195.800 664.400 200.400 ;
        RECT 670.000 191.800 670.800 200.400 ;
        RECT 672.200 195.800 673.000 200.400 ;
        RECT 676.400 191.800 677.200 200.400 ;
        RECT 679.600 193.200 680.600 200.400 ;
        RECT 685.800 199.800 686.600 200.400 ;
        RECT 685.800 193.200 686.800 199.800 ;
        RECT 310.000 191.200 337.000 191.800 ;
        RECT 186.200 191.000 187.000 191.200 ;
        RECT 232.600 191.000 233.400 191.200 ;
        RECT 272.600 191.000 273.400 191.200 ;
        RECT 336.200 191.000 337.000 191.200 ;
        RECT 431.000 191.200 458.000 191.800 ;
        RECT 431.000 191.000 431.800 191.200 ;
        RECT 30.600 170.800 31.400 171.000 ;
        RECT 105.800 170.800 106.600 171.000 ;
        RECT 4.400 170.200 31.400 170.800 ;
        RECT 79.600 170.200 106.600 170.800 ;
        RECT 224.600 170.800 225.400 171.000 ;
        RECT 301.000 170.800 301.800 171.000 ;
        RECT 353.800 170.800 354.600 171.000 ;
        RECT 224.600 170.200 251.600 170.800 ;
        RECT 274.800 170.200 301.800 170.800 ;
        RECT 327.600 170.200 354.600 170.800 ;
        RECT 363.800 170.800 364.600 171.000 ;
        RECT 419.800 170.800 420.600 171.000 ;
        RECT 534.600 170.800 535.400 171.000 ;
        RECT 363.800 170.200 390.800 170.800 ;
        RECT 419.800 170.200 446.800 170.800 ;
        RECT 508.400 170.200 535.400 170.800 ;
        RECT 658.200 170.800 659.000 171.000 ;
        RECT 658.200 170.200 685.200 170.800 ;
        RECT 4.400 169.600 5.200 170.200 ;
        RECT 7.800 170.000 8.600 170.200 ;
        RECT 1.200 161.600 2.000 166.200 ;
        RECT 4.400 161.600 5.200 166.200 ;
        RECT 7.600 161.600 8.400 166.200 ;
        RECT 14.000 161.600 14.800 166.200 ;
        RECT 17.200 161.600 18.000 166.200 ;
        RECT 25.200 161.600 26.000 166.200 ;
        RECT 28.400 161.600 29.200 166.200 ;
        RECT 31.600 161.600 32.400 166.200 ;
        RECT 34.800 161.600 35.600 166.200 ;
        RECT 38.000 161.600 38.800 170.000 ;
        RECT 43.600 161.600 44.400 166.200 ;
        RECT 46.800 161.600 47.600 166.200 ;
        RECT 52.400 161.600 53.200 170.200 ;
        RECT 55.600 161.600 56.400 166.200 ;
        RECT 58.800 161.600 59.600 166.200 ;
        RECT 60.400 161.600 61.200 170.200 ;
        RECT 64.600 161.600 65.400 166.200 ;
        RECT 67.400 161.600 68.200 166.200 ;
        RECT 71.600 161.600 72.400 170.200 ;
        RECT 79.600 169.600 80.400 170.200 ;
        RECT 83.000 170.000 83.800 170.200 ;
        RECT 74.800 161.600 75.600 166.200 ;
        RECT 76.400 161.600 77.200 166.200 ;
        RECT 79.600 161.600 80.400 166.200 ;
        RECT 82.800 161.600 83.600 166.200 ;
        RECT 89.200 161.600 90.000 166.200 ;
        RECT 92.400 161.600 93.200 166.200 ;
        RECT 100.400 161.600 101.200 166.200 ;
        RECT 103.600 161.600 104.400 166.200 ;
        RECT 106.800 161.600 107.600 166.200 ;
        RECT 110.000 161.600 110.800 166.200 ;
        RECT 118.000 161.600 118.800 166.200 ;
        RECT 119.600 161.600 120.400 166.200 ;
        RECT 122.800 161.600 123.600 166.200 ;
        RECT 126.000 161.600 126.800 169.000 ;
        RECT 129.200 161.600 130.000 170.200 ;
        RECT 131.400 161.600 132.200 166.200 ;
        RECT 135.600 161.600 136.400 170.200 ;
        RECT 138.800 161.600 139.600 169.800 ;
        RECT 144.000 161.600 144.800 170.200 ;
        RECT 150.000 161.600 150.800 170.200 ;
        RECT 152.200 161.600 153.000 166.200 ;
        RECT 156.400 161.600 157.200 170.200 ;
        RECT 158.000 161.600 158.800 170.200 ;
        RECT 162.200 161.600 163.000 166.200 ;
        RECT 166.000 161.600 166.800 166.200 ;
        RECT 169.200 161.600 170.000 169.800 ;
        RECT 174.400 161.600 175.200 170.200 ;
        RECT 177.200 161.600 178.000 170.200 ;
        RECT 181.400 161.600 182.200 166.200 ;
        RECT 183.600 161.600 184.400 170.200 ;
        RECT 187.800 161.600 188.600 166.200 ;
        RECT 190.600 161.600 191.400 166.200 ;
        RECT 194.800 161.600 195.600 170.200 ;
        RECT 198.000 161.600 198.800 166.200 ;
        RECT 200.200 161.600 201.000 166.200 ;
        RECT 204.400 161.600 205.200 170.200 ;
        RECT 206.000 161.600 206.800 170.200 ;
        RECT 247.400 170.000 248.200 170.200 ;
        RECT 250.800 169.600 251.600 170.200 ;
        RECT 214.000 161.600 214.800 169.000 ;
        RECT 218.800 161.600 219.600 166.200 ;
        RECT 220.400 161.600 221.200 166.200 ;
        RECT 223.600 161.600 224.400 166.200 ;
        RECT 226.800 161.600 227.600 166.200 ;
        RECT 230.000 161.600 230.800 166.200 ;
        RECT 238.000 161.600 238.800 166.200 ;
        RECT 241.200 161.600 242.000 166.200 ;
        RECT 247.600 161.600 248.400 166.200 ;
        RECT 250.800 161.600 251.600 166.200 ;
        RECT 254.000 161.600 254.800 166.200 ;
        RECT 258.800 161.600 259.600 170.200 ;
        RECT 274.800 169.600 275.600 170.200 ;
        RECT 278.000 170.000 279.000 170.200 ;
        RECT 263.600 161.600 264.400 169.000 ;
        RECT 271.600 161.600 272.400 166.200 ;
        RECT 274.800 161.600 275.600 166.200 ;
        RECT 278.000 161.600 278.800 166.200 ;
        RECT 284.400 161.600 285.200 166.200 ;
        RECT 287.600 161.600 288.400 166.200 ;
        RECT 295.600 161.600 296.400 166.200 ;
        RECT 298.800 161.600 299.600 166.200 ;
        RECT 302.000 161.600 302.800 166.200 ;
        RECT 305.200 161.600 306.000 166.200 ;
        RECT 308.400 161.600 309.200 169.000 ;
        RECT 311.600 161.600 312.400 170.200 ;
        RECT 313.200 161.600 314.000 166.200 ;
        RECT 316.400 161.600 317.200 166.200 ;
        RECT 318.000 161.600 318.800 170.200 ;
        RECT 327.600 169.600 328.400 170.200 ;
        RECT 331.000 170.000 331.800 170.200 ;
        RECT 386.600 170.000 387.600 170.200 ;
        RECT 390.000 169.600 390.800 170.200 ;
        RECT 322.200 161.600 323.000 166.200 ;
        RECT 324.400 161.600 325.200 166.200 ;
        RECT 327.600 161.600 328.400 166.200 ;
        RECT 330.800 161.600 331.600 166.200 ;
        RECT 337.200 161.600 338.000 166.200 ;
        RECT 340.400 161.600 341.200 166.200 ;
        RECT 348.400 161.600 349.200 166.200 ;
        RECT 351.600 161.600 352.400 166.200 ;
        RECT 354.800 161.600 355.600 166.200 ;
        RECT 358.000 161.600 358.800 166.200 ;
        RECT 359.600 161.600 360.400 166.200 ;
        RECT 362.800 161.600 363.600 166.200 ;
        RECT 366.000 161.600 366.800 166.200 ;
        RECT 369.200 161.600 370.000 166.200 ;
        RECT 377.200 161.600 378.000 166.200 ;
        RECT 380.400 161.600 381.200 166.200 ;
        RECT 386.800 161.600 387.600 166.200 ;
        RECT 390.000 161.600 390.800 166.200 ;
        RECT 393.200 161.600 394.000 166.200 ;
        RECT 396.400 161.600 397.200 169.800 ;
        RECT 401.600 161.600 402.400 170.200 ;
        RECT 406.000 161.600 406.800 169.000 ;
        RECT 409.200 161.600 410.000 170.200 ;
        RECT 442.600 170.000 443.600 170.200 ;
        RECT 446.000 169.600 446.800 170.200 ;
        RECT 415.600 161.600 416.400 166.200 ;
        RECT 418.800 161.600 419.600 166.200 ;
        RECT 422.000 161.600 422.800 166.200 ;
        RECT 425.200 161.600 426.000 166.200 ;
        RECT 433.200 161.600 434.000 166.200 ;
        RECT 436.400 161.600 437.200 166.200 ;
        RECT 442.800 161.600 443.600 166.200 ;
        RECT 446.000 161.600 446.800 166.200 ;
        RECT 449.200 161.600 450.000 166.200 ;
        RECT 450.800 161.600 451.600 166.200 ;
        RECT 454.000 161.600 454.800 166.200 ;
        RECT 455.600 161.600 456.400 166.200 ;
        RECT 458.800 161.600 459.600 166.200 ;
        RECT 462.000 161.600 462.800 166.200 ;
        RECT 465.200 161.600 466.000 169.800 ;
        RECT 470.400 161.600 471.200 170.200 ;
        RECT 474.800 161.600 475.600 169.800 ;
        RECT 480.000 161.600 480.800 170.200 ;
        RECT 484.400 161.600 485.200 166.200 ;
        RECT 486.600 161.600 487.400 166.200 ;
        RECT 490.800 161.600 491.600 170.200 ;
        RECT 494.000 161.600 494.800 166.200 ;
        RECT 495.600 161.600 496.400 166.200 ;
        RECT 498.800 161.600 499.600 170.200 ;
        RECT 508.400 169.600 509.200 170.200 ;
        RECT 511.800 170.000 512.600 170.200 ;
        RECT 502.000 161.600 502.800 169.000 ;
        RECT 505.200 161.600 506.000 166.200 ;
        RECT 508.400 161.600 509.200 166.200 ;
        RECT 511.600 161.600 512.400 166.200 ;
        RECT 518.000 161.600 518.800 166.200 ;
        RECT 521.200 161.600 522.000 166.200 ;
        RECT 529.200 161.600 530.000 166.200 ;
        RECT 532.400 161.600 533.200 166.200 ;
        RECT 535.600 161.600 536.400 166.200 ;
        RECT 538.800 161.600 539.600 166.200 ;
        RECT 540.400 161.600 541.200 170.200 ;
        RECT 543.600 161.600 544.400 169.000 ;
        RECT 548.400 161.600 549.200 169.000 ;
        RECT 551.600 161.600 552.400 170.200 ;
        RECT 554.800 161.600 555.600 166.200 ;
        RECT 557.000 161.600 557.800 166.200 ;
        RECT 561.200 161.600 562.000 170.200 ;
        RECT 562.800 161.600 563.600 166.200 ;
        RECT 566.000 161.600 566.800 166.200 ;
        RECT 573.600 161.600 574.400 170.200 ;
        RECT 578.800 161.600 579.600 169.800 ;
        RECT 582.600 161.600 583.400 166.200 ;
        RECT 586.800 161.600 587.600 170.200 ;
        RECT 590.000 161.600 590.800 166.200 ;
        RECT 593.200 161.600 594.000 170.200 ;
        RECT 598.800 161.600 599.600 166.200 ;
        RECT 602.000 161.600 602.800 166.200 ;
        RECT 607.600 161.600 608.400 170.000 ;
        RECT 612.400 161.600 613.200 166.200 ;
        RECT 614.000 161.600 614.800 170.200 ;
        RECT 618.200 161.600 619.000 166.200 ;
        RECT 621.000 161.600 621.800 166.200 ;
        RECT 625.200 161.600 626.000 170.200 ;
        RECT 628.400 161.600 629.200 169.800 ;
        RECT 633.600 161.600 634.400 170.200 ;
        RECT 636.400 161.600 637.200 166.200 ;
        RECT 639.600 161.600 640.400 166.200 ;
        RECT 641.200 161.600 642.000 170.200 ;
        RECT 649.200 161.600 650.000 170.200 ;
        RECT 681.000 170.000 682.000 170.200 ;
        RECT 684.400 169.600 685.200 170.200 ;
        RECT 652.400 161.600 653.200 166.200 ;
        RECT 654.000 161.600 654.800 166.200 ;
        RECT 657.200 161.600 658.000 166.200 ;
        RECT 660.400 161.600 661.200 166.200 ;
        RECT 663.600 161.600 664.400 166.200 ;
        RECT 671.600 161.600 672.400 166.200 ;
        RECT 674.800 161.600 675.600 166.200 ;
        RECT 681.200 161.600 682.000 166.200 ;
        RECT 684.400 161.600 685.200 166.200 ;
        RECT 687.600 161.600 688.400 166.200 ;
        RECT 0.400 160.400 689.200 161.600 ;
        RECT 2.800 155.800 3.600 160.400 ;
        RECT 4.400 151.800 5.200 160.400 ;
        RECT 8.600 155.800 9.400 160.400 ;
        RECT 11.400 155.800 12.200 160.400 ;
        RECT 15.600 151.800 16.400 160.400 ;
        RECT 17.200 151.800 18.000 160.400 ;
        RECT 20.400 153.000 21.200 160.400 ;
        RECT 23.600 151.800 24.400 160.400 ;
        RECT 26.800 153.000 27.600 160.400 ;
        RECT 30.000 151.800 30.800 160.400 ;
        RECT 34.200 155.800 35.000 160.400 ;
        RECT 37.000 155.800 37.800 160.400 ;
        RECT 41.200 151.800 42.000 160.400 ;
        RECT 44.000 151.800 44.800 160.400 ;
        RECT 49.200 152.200 50.000 160.400 ;
        RECT 53.600 151.800 54.400 160.400 ;
        RECT 58.800 152.200 59.600 160.400 ;
        RECT 62.000 151.800 62.800 160.400 ;
        RECT 66.200 155.800 67.000 160.400 ;
        RECT 69.000 155.800 69.800 160.400 ;
        RECT 73.200 151.800 74.000 160.400 ;
        RECT 74.800 151.800 75.600 160.400 ;
        RECT 78.000 153.000 78.800 160.400 ;
        RECT 81.200 151.800 82.000 160.400 ;
        RECT 85.400 155.800 86.200 160.400 ;
        RECT 88.200 155.800 89.000 160.400 ;
        RECT 92.400 151.800 93.200 160.400 ;
        RECT 95.600 151.800 96.400 160.400 ;
        RECT 101.200 155.800 102.000 160.400 ;
        RECT 104.400 155.800 105.200 160.400 ;
        RECT 110.000 152.000 110.800 160.400 ;
        RECT 119.600 152.200 120.400 160.400 ;
        RECT 124.800 151.800 125.600 160.400 ;
        RECT 127.600 151.800 128.400 160.400 ;
        RECT 131.800 155.800 132.600 160.400 ;
        RECT 135.600 153.000 136.400 160.400 ;
        RECT 138.800 151.800 139.600 160.400 ;
        RECT 142.000 152.200 142.800 160.400 ;
        RECT 147.200 151.800 148.000 160.400 ;
        RECT 150.000 151.800 150.800 160.400 ;
        RECT 154.200 155.800 155.000 160.400 ;
        RECT 157.000 155.800 157.800 160.400 ;
        RECT 161.200 151.800 162.000 160.400 ;
        RECT 164.400 152.000 165.200 160.400 ;
        RECT 170.000 155.800 170.800 160.400 ;
        RECT 173.200 155.800 174.000 160.400 ;
        RECT 178.800 151.800 179.600 160.400 ;
        RECT 182.000 155.800 182.800 160.400 ;
        RECT 186.800 152.200 187.600 160.400 ;
        RECT 192.000 151.800 192.800 160.400 ;
        RECT 196.400 152.200 197.200 160.400 ;
        RECT 201.600 151.800 202.400 160.400 ;
        RECT 204.400 151.800 205.200 160.400 ;
        RECT 208.600 155.800 209.400 160.400 ;
        RECT 211.400 155.800 212.200 160.400 ;
        RECT 215.600 151.800 216.400 160.400 ;
        RECT 218.800 151.800 219.600 160.400 ;
        RECT 224.400 155.800 225.200 160.400 ;
        RECT 227.600 155.800 228.400 160.400 ;
        RECT 233.200 152.000 234.000 160.400 ;
        RECT 238.000 152.200 238.800 160.400 ;
        RECT 243.200 151.800 244.000 160.400 ;
        RECT 247.600 152.200 248.400 160.400 ;
        RECT 252.800 151.800 253.600 160.400 ;
        RECT 257.400 159.800 258.200 160.400 ;
        RECT 257.200 153.200 258.200 159.800 ;
        RECT 263.400 153.200 264.400 160.400 ;
        RECT 271.600 155.800 272.400 160.400 ;
        RECT 274.800 155.800 275.600 160.400 ;
        RECT 278.000 155.800 278.800 160.400 ;
        RECT 284.400 155.800 285.200 160.400 ;
        RECT 287.600 155.800 288.400 160.400 ;
        RECT 295.600 155.800 296.400 160.400 ;
        RECT 298.800 155.800 299.600 160.400 ;
        RECT 302.000 155.800 302.800 160.400 ;
        RECT 305.200 155.800 306.000 160.400 ;
        RECT 306.800 151.800 307.600 160.400 ;
        RECT 311.000 155.800 311.800 160.400 ;
        RECT 313.200 155.800 314.000 160.400 ;
        RECT 316.400 155.800 317.200 160.400 ;
        RECT 319.600 155.800 320.400 160.400 ;
        RECT 326.000 155.800 326.800 160.400 ;
        RECT 329.200 155.800 330.000 160.400 ;
        RECT 337.200 155.800 338.000 160.400 ;
        RECT 340.400 155.800 341.200 160.400 ;
        RECT 343.600 155.800 344.400 160.400 ;
        RECT 346.800 155.800 347.600 160.400 ;
        RECT 348.400 155.800 349.200 160.400 ;
        RECT 351.600 155.800 352.400 160.400 ;
        RECT 354.800 155.800 355.600 160.400 ;
        RECT 358.000 155.800 358.800 160.400 ;
        RECT 366.000 155.800 366.800 160.400 ;
        RECT 369.200 155.800 370.000 160.400 ;
        RECT 375.600 155.800 376.400 160.400 ;
        RECT 378.800 155.800 379.600 160.400 ;
        RECT 382.000 155.800 382.800 160.400 ;
        RECT 383.600 155.800 384.400 160.400 ;
        RECT 386.800 155.800 387.600 160.400 ;
        RECT 390.000 155.800 390.800 160.400 ;
        RECT 396.400 155.800 397.200 160.400 ;
        RECT 399.600 155.800 400.400 160.400 ;
        RECT 407.600 155.800 408.400 160.400 ;
        RECT 410.800 155.800 411.600 160.400 ;
        RECT 414.000 155.800 414.800 160.400 ;
        RECT 417.200 155.800 418.000 160.400 ;
        RECT 425.200 155.800 426.000 160.400 ;
        RECT 316.400 151.800 317.200 152.400 ;
        RECT 319.800 151.800 320.600 152.000 ;
        RECT 375.400 151.800 376.200 152.000 ;
        RECT 378.800 151.800 379.600 152.400 ;
        RECT 316.400 151.200 343.400 151.800 ;
        RECT 342.600 151.000 343.400 151.200 ;
        RECT 352.600 151.200 379.600 151.800 ;
        RECT 386.800 151.800 387.600 152.400 ;
        RECT 390.000 151.800 391.000 152.000 ;
        RECT 426.800 151.800 427.600 160.400 ;
        RECT 431.000 155.800 431.800 160.400 ;
        RECT 433.200 155.800 434.000 160.400 ;
        RECT 436.400 155.800 437.200 160.400 ;
        RECT 438.000 155.800 438.800 160.400 ;
        RECT 441.200 155.800 442.000 160.400 ;
        RECT 444.400 155.800 445.200 160.400 ;
        RECT 450.800 155.800 451.600 160.400 ;
        RECT 454.000 155.800 454.800 160.400 ;
        RECT 462.000 155.800 462.800 160.400 ;
        RECT 465.200 155.800 466.000 160.400 ;
        RECT 468.400 155.800 469.200 160.400 ;
        RECT 471.600 155.800 472.400 160.400 ;
        RECT 474.800 155.800 475.600 160.400 ;
        RECT 476.400 155.800 477.200 160.400 ;
        RECT 479.600 155.800 480.400 160.400 ;
        RECT 482.800 155.800 483.600 160.400 ;
        RECT 489.200 155.800 490.000 160.400 ;
        RECT 492.400 155.800 493.200 160.400 ;
        RECT 500.400 155.800 501.200 160.400 ;
        RECT 503.600 155.800 504.400 160.400 ;
        RECT 506.800 155.800 507.600 160.400 ;
        RECT 510.000 155.800 510.800 160.400 ;
        RECT 511.600 155.800 512.400 160.400 ;
        RECT 515.400 155.800 516.200 160.400 ;
        RECT 441.200 151.800 442.000 152.400 ;
        RECT 444.400 151.800 445.400 152.000 ;
        RECT 479.600 151.800 480.400 152.400 ;
        RECT 483.000 151.800 483.800 152.000 ;
        RECT 519.600 151.800 520.400 160.400 ;
        RECT 521.200 151.800 522.000 160.400 ;
        RECT 525.400 155.800 526.200 160.400 ;
        RECT 528.200 155.800 529.000 160.400 ;
        RECT 532.400 151.800 533.200 160.400 ;
        RECT 534.000 151.800 534.800 160.400 ;
        RECT 538.800 155.800 539.600 160.400 ;
        RECT 542.000 151.800 542.800 160.400 ;
        RECT 546.200 155.800 547.000 160.400 ;
        RECT 550.000 151.800 550.800 160.400 ;
        RECT 551.600 155.800 552.400 160.400 ;
        RECT 554.800 155.800 555.600 160.400 ;
        RECT 556.400 151.800 557.200 160.400 ;
        RECT 559.600 153.000 560.400 160.400 ;
        RECT 563.400 155.800 564.200 160.400 ;
        RECT 567.600 151.800 568.400 160.400 ;
        RECT 574.600 155.800 575.400 160.400 ;
        RECT 578.800 151.800 579.600 160.400 ;
        RECT 580.400 151.800 581.200 160.400 ;
        RECT 584.600 155.800 585.400 160.400 ;
        RECT 587.400 155.800 588.200 160.400 ;
        RECT 591.600 151.800 592.400 160.400 ;
        RECT 594.800 152.200 595.600 160.400 ;
        RECT 600.000 151.800 600.800 160.400 ;
        RECT 604.400 153.000 605.200 160.400 ;
        RECT 607.600 151.800 608.400 160.400 ;
        RECT 609.200 151.800 610.000 160.400 ;
        RECT 613.400 155.800 614.200 160.400 ;
        RECT 615.600 151.800 616.400 160.400 ;
        RECT 618.800 153.000 619.600 160.400 ;
        RECT 623.600 156.200 624.400 160.400 ;
        RECT 626.800 155.800 627.600 160.400 ;
        RECT 630.000 153.000 630.800 160.400 ;
        RECT 633.200 151.800 634.000 160.400 ;
        RECT 636.400 153.000 637.200 160.400 ;
        RECT 639.600 151.800 640.400 160.400 ;
        RECT 642.800 155.800 643.600 160.400 ;
        RECT 646.000 152.200 646.800 160.400 ;
        RECT 651.200 151.800 652.000 160.400 ;
        RECT 655.600 152.200 656.400 160.400 ;
        RECT 660.800 151.800 661.600 160.400 ;
        RECT 663.600 151.800 664.400 160.400 ;
        RECT 667.800 155.800 668.600 160.400 ;
        RECT 671.600 151.800 672.400 160.400 ;
        RECT 677.200 155.800 678.000 160.400 ;
        RECT 680.400 155.800 681.200 160.400 ;
        RECT 686.000 152.000 686.800 160.400 ;
        RECT 386.800 151.200 413.800 151.800 ;
        RECT 441.200 151.200 468.200 151.800 ;
        RECT 479.600 151.200 506.600 151.800 ;
        RECT 352.600 151.000 353.400 151.200 ;
        RECT 413.000 151.000 413.800 151.200 ;
        RECT 467.400 151.000 468.200 151.200 ;
        RECT 505.800 151.000 506.600 151.200 ;
        RECT 273.000 150.000 296.400 150.600 ;
        RECT 273.000 149.800 273.800 150.000 ;
        RECT 278.000 149.600 278.800 150.000 ;
        RECT 295.600 149.400 296.400 150.000 ;
        RECT 205.400 130.800 206.200 131.000 ;
        RECT 311.000 130.800 311.800 131.000 ;
        RECT 381.000 130.800 381.800 131.000 ;
        RECT 205.400 130.200 232.400 130.800 ;
        RECT 311.000 130.200 338.000 130.800 ;
        RECT 354.800 130.200 381.800 130.800 ;
        RECT 397.400 130.800 398.200 131.000 ;
        RECT 470.600 130.800 471.400 131.000 ;
        RECT 505.800 130.800 506.600 131.000 ;
        RECT 397.400 130.200 424.400 130.800 ;
        RECT 2.800 121.600 3.600 130.000 ;
        RECT 8.400 121.600 9.200 126.200 ;
        RECT 11.600 121.600 12.400 126.200 ;
        RECT 17.200 121.600 18.000 130.200 ;
        RECT 21.000 121.600 21.800 126.200 ;
        RECT 25.200 121.600 26.000 130.200 ;
        RECT 27.400 121.600 28.200 126.200 ;
        RECT 31.600 121.600 32.400 130.200 ;
        RECT 34.800 121.600 35.600 130.000 ;
        RECT 40.400 121.600 41.200 126.200 ;
        RECT 43.600 121.600 44.400 126.200 ;
        RECT 49.200 121.600 50.000 130.200 ;
        RECT 52.400 121.600 53.200 130.200 ;
        RECT 56.600 121.600 57.400 126.200 ;
        RECT 59.400 121.600 60.200 126.200 ;
        RECT 63.600 121.600 64.400 130.200 ;
        RECT 66.400 121.600 67.200 130.200 ;
        RECT 71.600 121.600 72.400 129.800 ;
        RECT 74.800 121.600 75.600 130.200 ;
        RECT 79.000 121.600 79.800 126.200 ;
        RECT 81.800 121.600 82.600 126.200 ;
        RECT 86.000 121.600 86.800 130.200 ;
        RECT 87.600 121.600 88.400 126.200 ;
        RECT 92.000 121.600 92.800 130.200 ;
        RECT 97.200 121.600 98.000 129.800 ;
        RECT 100.400 121.600 101.200 126.200 ;
        RECT 103.600 121.600 104.400 125.800 ;
        RECT 107.400 121.600 108.200 126.200 ;
        RECT 111.600 121.600 112.400 130.200 ;
        RECT 118.000 121.600 118.800 126.200 ;
        RECT 121.200 121.600 122.000 126.200 ;
        RECT 123.400 121.600 124.200 126.200 ;
        RECT 127.600 121.600 128.400 130.200 ;
        RECT 130.800 121.600 131.600 126.200 ;
        RECT 132.400 121.600 133.200 126.200 ;
        RECT 135.600 121.600 136.400 125.800 ;
        RECT 138.800 121.600 139.600 126.200 ;
        RECT 142.000 121.600 142.800 130.200 ;
        RECT 146.200 121.600 147.000 126.200 ;
        RECT 149.000 121.600 149.800 126.200 ;
        RECT 153.200 121.600 154.000 130.200 ;
        RECT 154.800 121.600 155.600 130.200 ;
        RECT 159.000 121.600 159.800 126.200 ;
        RECT 162.800 121.600 163.600 126.200 ;
        RECT 166.000 121.600 166.800 129.000 ;
        RECT 169.200 121.600 170.000 130.200 ;
        RECT 172.400 121.600 173.200 125.800 ;
        RECT 175.600 121.600 176.400 126.200 ;
        RECT 177.800 121.600 178.600 126.200 ;
        RECT 182.000 121.600 182.800 130.200 ;
        RECT 183.600 121.600 184.400 126.200 ;
        RECT 186.800 121.600 187.600 126.200 ;
        RECT 189.000 121.600 189.800 126.200 ;
        RECT 193.200 121.600 194.000 130.200 ;
        RECT 194.800 121.600 195.600 130.200 ;
        RECT 228.200 130.000 229.200 130.200 ;
        RECT 231.600 129.600 232.400 130.200 ;
        RECT 199.000 121.600 199.800 126.200 ;
        RECT 201.200 121.600 202.000 126.200 ;
        RECT 204.400 121.600 205.200 126.200 ;
        RECT 207.600 121.600 208.400 126.200 ;
        RECT 210.800 121.600 211.600 126.200 ;
        RECT 218.800 121.600 219.600 126.200 ;
        RECT 222.000 121.600 222.800 126.200 ;
        RECT 228.400 121.600 229.200 126.200 ;
        RECT 231.600 121.600 232.400 126.200 ;
        RECT 234.800 121.600 235.600 126.200 ;
        RECT 238.000 121.600 238.800 125.800 ;
        RECT 241.200 121.600 242.000 126.200 ;
        RECT 245.000 121.600 245.800 130.200 ;
        RECT 252.400 121.600 253.200 130.200 ;
        RECT 254.000 121.600 254.800 130.200 ;
        RECT 257.200 121.600 258.000 130.200 ;
        RECT 260.400 121.600 261.200 130.200 ;
        RECT 266.800 121.600 267.600 130.200 ;
        RECT 270.000 121.600 270.800 129.000 ;
        RECT 273.200 121.600 274.000 130.200 ;
        RECT 276.400 121.600 277.200 129.000 ;
        RECT 279.600 121.600 280.400 126.200 ;
        RECT 282.800 121.600 283.600 126.200 ;
        RECT 285.000 121.600 285.800 126.200 ;
        RECT 289.200 121.600 290.000 130.200 ;
        RECT 290.800 121.600 291.600 126.200 ;
        RECT 294.000 121.600 294.800 126.200 ;
        RECT 295.600 121.600 296.400 130.200 ;
        RECT 333.800 130.000 334.800 130.200 ;
        RECT 337.200 129.600 338.000 130.200 ;
        RECT 299.800 121.600 300.600 126.200 ;
        RECT 302.000 121.600 302.800 126.200 ;
        RECT 305.200 121.600 306.000 126.200 ;
        RECT 306.800 121.600 307.600 126.200 ;
        RECT 310.000 121.600 310.800 126.200 ;
        RECT 313.200 121.600 314.000 126.200 ;
        RECT 316.400 121.600 317.200 126.200 ;
        RECT 324.400 121.600 325.200 126.200 ;
        RECT 327.600 121.600 328.400 126.200 ;
        RECT 334.000 121.600 334.800 126.200 ;
        RECT 337.200 121.600 338.000 126.200 ;
        RECT 340.400 121.600 341.200 126.200 ;
        RECT 345.200 121.600 346.000 130.200 ;
        RECT 346.800 121.600 347.600 130.200 ;
        RECT 354.800 129.600 355.600 130.200 ;
        RECT 358.000 130.000 359.000 130.200 ;
        RECT 351.600 121.600 352.400 126.200 ;
        RECT 354.800 121.600 355.600 126.200 ;
        RECT 358.000 121.600 358.800 126.200 ;
        RECT 364.400 121.600 365.200 126.200 ;
        RECT 367.600 121.600 368.400 126.200 ;
        RECT 375.600 121.600 376.400 126.200 ;
        RECT 378.800 121.600 379.600 126.200 ;
        RECT 382.000 121.600 382.800 126.200 ;
        RECT 385.200 121.600 386.000 126.200 ;
        RECT 386.800 121.600 387.600 130.200 ;
        RECT 420.200 130.000 421.200 130.200 ;
        RECT 423.600 129.600 424.400 130.200 ;
        RECT 444.400 130.200 471.400 130.800 ;
        RECT 479.600 130.200 506.600 130.800 ;
        RECT 444.400 129.600 445.200 130.200 ;
        RECT 447.600 130.000 448.600 130.200 ;
        RECT 479.600 129.600 480.400 130.200 ;
        RECT 483.000 130.000 483.800 130.200 ;
        RECT 390.000 121.600 390.800 129.000 ;
        RECT 393.200 121.600 394.000 126.200 ;
        RECT 396.400 121.600 397.200 126.200 ;
        RECT 399.600 121.600 400.400 126.200 ;
        RECT 402.800 121.600 403.600 126.200 ;
        RECT 410.800 121.600 411.600 126.200 ;
        RECT 414.000 121.600 414.800 126.200 ;
        RECT 420.400 121.600 421.200 126.200 ;
        RECT 423.600 121.600 424.400 126.200 ;
        RECT 426.800 121.600 427.600 126.200 ;
        RECT 434.800 121.600 435.600 129.000 ;
        RECT 438.000 121.600 438.800 126.200 ;
        RECT 441.200 121.600 442.000 126.200 ;
        RECT 444.400 121.600 445.200 126.200 ;
        RECT 447.600 121.600 448.400 126.200 ;
        RECT 454.000 121.600 454.800 126.200 ;
        RECT 457.200 121.600 458.000 126.200 ;
        RECT 465.200 121.600 466.000 126.200 ;
        RECT 468.400 121.600 469.200 126.200 ;
        RECT 471.600 121.600 472.400 126.200 ;
        RECT 474.800 121.600 475.600 126.200 ;
        RECT 476.400 121.600 477.200 126.200 ;
        RECT 479.600 121.600 480.400 126.200 ;
        RECT 482.800 121.600 483.600 126.200 ;
        RECT 489.200 121.600 490.000 126.200 ;
        RECT 492.400 121.600 493.200 126.200 ;
        RECT 500.400 121.600 501.200 126.200 ;
        RECT 503.600 121.600 504.400 126.200 ;
        RECT 506.800 121.600 507.600 126.200 ;
        RECT 510.000 121.600 510.800 126.200 ;
        RECT 512.200 121.600 513.000 126.200 ;
        RECT 516.400 121.600 517.200 130.200 ;
        RECT 519.600 121.600 520.400 130.200 ;
        RECT 525.200 121.600 526.000 126.200 ;
        RECT 528.400 121.600 529.200 126.200 ;
        RECT 534.000 121.600 534.800 130.000 ;
        RECT 538.800 121.600 539.600 129.000 ;
        RECT 542.000 121.600 542.800 130.200 ;
        RECT 543.600 121.600 544.400 130.200 ;
        RECT 547.800 121.600 548.600 126.200 ;
        RECT 550.600 121.600 551.400 126.200 ;
        RECT 554.800 121.600 555.600 130.200 ;
        RECT 556.400 121.600 557.200 130.200 ;
        RECT 562.800 121.600 563.600 130.000 ;
        RECT 568.400 121.600 569.200 126.200 ;
        RECT 571.600 121.600 572.400 126.200 ;
        RECT 577.200 121.600 578.000 130.200 ;
        RECT 585.200 121.600 586.000 126.200 ;
        RECT 588.400 121.600 589.200 126.200 ;
        RECT 591.600 121.600 592.400 125.800 ;
        RECT 594.800 121.600 595.600 126.200 ;
        RECT 597.000 121.600 597.800 126.200 ;
        RECT 601.200 121.600 602.000 130.200 ;
        RECT 604.400 121.600 605.200 129.800 ;
        RECT 609.600 121.600 610.400 130.200 ;
        RECT 612.400 121.600 613.200 130.200 ;
        RECT 616.600 121.600 617.400 126.200 ;
        RECT 618.800 121.600 619.600 130.200 ;
        RECT 623.000 121.600 623.800 126.200 ;
        RECT 626.800 121.600 627.600 130.200 ;
        RECT 632.400 121.600 633.200 126.200 ;
        RECT 635.600 121.600 636.400 126.200 ;
        RECT 641.200 121.600 642.000 130.000 ;
        RECT 646.000 121.600 646.800 126.200 ;
        RECT 649.200 121.600 650.000 129.800 ;
        RECT 654.400 121.600 655.200 130.200 ;
        RECT 658.800 121.600 659.600 129.000 ;
        RECT 662.000 121.600 662.800 130.200 ;
        RECT 663.600 121.600 664.400 130.200 ;
        RECT 667.800 121.600 668.600 126.200 ;
        RECT 671.600 121.600 672.400 130.200 ;
        RECT 677.200 121.600 678.000 126.200 ;
        RECT 680.400 121.600 681.200 126.200 ;
        RECT 686.000 121.600 686.800 130.000 ;
        RECT 0.400 120.400 689.200 121.600 ;
        RECT 2.800 112.000 3.600 120.400 ;
        RECT 8.400 115.800 9.200 120.400 ;
        RECT 11.600 115.800 12.400 120.400 ;
        RECT 17.200 111.800 18.000 120.400 ;
        RECT 20.400 111.800 21.200 120.400 ;
        RECT 23.600 113.000 24.400 120.400 ;
        RECT 28.400 112.200 29.200 120.400 ;
        RECT 33.600 111.800 34.400 120.400 ;
        RECT 38.000 113.000 38.800 120.400 ;
        RECT 41.200 111.800 42.000 120.400 ;
        RECT 44.400 113.000 45.200 120.400 ;
        RECT 47.600 111.800 48.400 120.400 ;
        RECT 50.800 112.000 51.600 120.400 ;
        RECT 56.400 115.800 57.200 120.400 ;
        RECT 59.600 115.800 60.400 120.400 ;
        RECT 65.200 111.800 66.000 120.400 ;
        RECT 70.000 112.200 70.800 120.400 ;
        RECT 75.200 111.800 76.000 120.400 ;
        RECT 78.000 115.800 78.800 120.400 ;
        RECT 82.800 112.000 83.600 120.400 ;
        RECT 88.400 115.800 89.200 120.400 ;
        RECT 91.600 115.800 92.400 120.400 ;
        RECT 97.200 111.800 98.000 120.400 ;
        RECT 100.400 111.800 101.200 120.400 ;
        RECT 104.600 115.800 105.400 120.400 ;
        RECT 107.400 115.800 108.200 120.400 ;
        RECT 111.600 111.800 112.400 120.400 ;
        RECT 119.600 113.000 120.400 120.400 ;
        RECT 122.800 111.800 123.600 120.400 ;
        RECT 124.400 115.800 125.200 120.400 ;
        RECT 127.600 115.800 128.400 120.400 ;
        RECT 129.200 111.800 130.000 120.400 ;
        RECT 133.400 115.800 134.200 120.400 ;
        RECT 136.800 111.800 137.600 120.400 ;
        RECT 142.000 112.200 142.800 120.400 ;
        RECT 145.200 111.800 146.000 120.400 ;
        RECT 149.400 115.800 150.200 120.400 ;
        RECT 153.200 112.000 154.000 120.400 ;
        RECT 158.800 115.800 159.600 120.400 ;
        RECT 162.000 115.800 162.800 120.400 ;
        RECT 167.600 111.800 168.400 120.400 ;
        RECT 170.800 115.800 171.600 120.400 ;
        RECT 174.000 111.800 174.800 120.400 ;
        RECT 178.200 115.800 179.000 120.400 ;
        RECT 180.400 111.800 181.200 120.400 ;
        RECT 184.600 115.800 185.400 120.400 ;
        RECT 188.400 111.800 189.200 120.400 ;
        RECT 190.600 115.800 191.400 120.400 ;
        RECT 194.800 111.800 195.600 120.400 ;
        RECT 197.000 115.800 197.800 120.400 ;
        RECT 201.200 111.800 202.000 120.400 ;
        RECT 202.800 111.800 203.600 120.400 ;
        RECT 209.800 111.800 210.600 120.400 ;
        RECT 214.000 115.800 214.800 120.400 ;
        RECT 217.200 115.800 218.000 120.400 ;
        RECT 220.400 115.800 221.200 120.400 ;
        RECT 225.200 111.800 226.000 120.400 ;
        RECT 228.400 113.000 229.200 120.400 ;
        RECT 233.200 111.800 234.000 120.400 ;
        RECT 237.400 115.800 238.200 120.400 ;
        RECT 239.600 111.800 240.400 120.400 ;
        RECT 243.800 115.800 244.600 120.400 ;
        RECT 246.000 115.800 246.800 120.400 ;
        RECT 249.200 115.800 250.000 120.400 ;
        RECT 250.800 111.800 251.600 120.400 ;
        RECT 255.000 115.800 255.800 120.400 ;
        RECT 257.200 115.800 258.000 120.400 ;
        RECT 260.400 115.800 261.200 120.400 ;
        RECT 266.800 115.800 267.600 120.400 ;
        RECT 270.000 115.800 270.800 120.400 ;
        RECT 273.200 115.800 274.000 120.400 ;
        RECT 276.400 115.800 277.200 120.400 ;
        RECT 284.400 115.800 285.200 120.400 ;
        RECT 287.600 115.800 288.400 120.400 ;
        RECT 294.000 115.800 294.800 120.400 ;
        RECT 297.200 115.800 298.000 120.400 ;
        RECT 300.400 115.800 301.200 120.400 ;
        RECT 303.600 113.000 304.400 120.400 ;
        RECT 293.800 111.800 294.800 112.000 ;
        RECT 297.200 111.800 298.000 112.400 ;
        RECT 306.800 111.800 307.600 120.400 ;
        RECT 310.000 113.000 310.800 120.400 ;
        RECT 314.800 115.800 315.600 120.400 ;
        RECT 316.400 111.800 317.200 120.400 ;
        RECT 320.600 115.800 321.400 120.400 ;
        RECT 322.800 115.800 323.600 120.400 ;
        RECT 326.000 115.800 326.800 120.400 ;
        RECT 327.600 115.800 328.400 120.400 ;
        RECT 330.800 115.800 331.600 120.400 ;
        RECT 334.000 115.800 334.800 120.400 ;
        RECT 337.200 115.800 338.000 120.400 ;
        RECT 345.200 115.800 346.000 120.400 ;
        RECT 348.400 115.800 349.200 120.400 ;
        RECT 354.800 115.800 355.600 120.400 ;
        RECT 358.000 115.800 358.800 120.400 ;
        RECT 361.200 115.800 362.000 120.400 ;
        RECT 362.800 115.800 363.600 120.400 ;
        RECT 366.000 115.800 366.800 120.400 ;
        RECT 369.200 115.800 370.000 120.400 ;
        RECT 372.400 115.800 373.200 120.400 ;
        RECT 380.400 115.800 381.200 120.400 ;
        RECT 383.600 115.800 384.400 120.400 ;
        RECT 390.000 115.800 390.800 120.400 ;
        RECT 393.200 115.800 394.000 120.400 ;
        RECT 396.400 115.800 397.200 120.400 ;
        RECT 399.600 115.800 400.400 120.400 ;
        RECT 401.800 115.800 402.600 120.400 ;
        RECT 354.600 111.800 355.400 112.000 ;
        RECT 358.000 111.800 358.800 112.400 ;
        RECT 389.800 111.800 390.800 112.000 ;
        RECT 393.200 111.800 394.000 112.400 ;
        RECT 406.000 111.800 406.800 120.400 ;
        RECT 407.600 115.800 408.400 120.400 ;
        RECT 410.800 115.800 411.600 120.400 ;
        RECT 413.000 115.800 413.800 120.400 ;
        RECT 417.200 111.800 418.000 120.400 ;
        RECT 423.600 115.800 424.400 120.400 ;
        RECT 426.800 115.800 427.600 120.400 ;
        RECT 430.000 115.800 430.800 120.400 ;
        RECT 433.200 115.800 434.000 120.400 ;
        RECT 441.200 115.800 442.000 120.400 ;
        RECT 444.400 115.800 445.200 120.400 ;
        RECT 450.800 115.800 451.600 120.400 ;
        RECT 454.000 115.800 454.800 120.400 ;
        RECT 457.200 115.800 458.000 120.400 ;
        RECT 450.600 111.800 451.400 112.000 ;
        RECT 454.000 111.800 454.800 112.400 ;
        RECT 458.800 111.800 459.600 120.400 ;
        RECT 462.000 113.000 462.800 120.400 ;
        RECT 465.200 111.800 466.000 120.400 ;
        RECT 469.400 115.800 470.200 120.400 ;
        RECT 471.600 115.800 472.400 120.400 ;
        RECT 474.800 115.800 475.600 120.400 ;
        RECT 476.400 115.800 477.200 120.400 ;
        RECT 479.600 115.800 480.400 120.400 ;
        RECT 481.200 115.800 482.000 120.400 ;
        RECT 484.400 115.800 485.200 120.400 ;
        RECT 487.600 115.800 488.400 120.400 ;
        RECT 490.800 115.800 491.600 120.400 ;
        RECT 498.800 115.800 499.600 120.400 ;
        RECT 502.000 115.800 502.800 120.400 ;
        RECT 508.400 115.800 509.200 120.400 ;
        RECT 511.600 115.800 512.400 120.400 ;
        RECT 514.800 115.800 515.600 120.400 ;
        RECT 508.200 111.800 509.200 112.000 ;
        RECT 511.600 111.800 512.400 112.400 ;
        RECT 516.400 111.800 517.200 120.400 ;
        RECT 519.600 113.000 520.400 120.400 ;
        RECT 523.400 115.800 524.200 120.400 ;
        RECT 527.600 111.800 528.400 120.400 ;
        RECT 529.200 111.800 530.000 120.400 ;
        RECT 532.400 111.800 533.200 120.400 ;
        RECT 535.600 111.800 536.400 120.400 ;
        RECT 538.800 111.800 539.600 120.400 ;
        RECT 542.000 111.800 542.800 120.400 ;
        RECT 544.200 115.800 545.000 120.400 ;
        RECT 548.400 111.800 549.200 120.400 ;
        RECT 550.000 115.800 550.800 120.400 ;
        RECT 553.200 115.800 554.000 120.400 ;
        RECT 556.000 111.800 556.800 120.400 ;
        RECT 561.200 112.200 562.000 120.400 ;
        RECT 566.000 113.000 566.800 120.400 ;
        RECT 569.200 111.800 570.000 120.400 ;
        RECT 575.600 115.800 576.400 120.400 ;
        RECT 578.800 115.800 579.600 120.400 ;
        RECT 582.000 115.800 582.800 120.400 ;
        RECT 584.200 115.800 585.000 120.400 ;
        RECT 588.400 111.800 589.200 120.400 ;
        RECT 590.000 111.800 590.800 120.400 ;
        RECT 594.200 115.800 595.000 120.400 ;
        RECT 596.400 115.800 597.200 120.400 ;
        RECT 599.600 115.800 600.400 120.400 ;
        RECT 602.800 115.800 603.600 120.400 ;
        RECT 606.000 111.800 606.800 120.400 ;
        RECT 611.600 115.800 612.400 120.400 ;
        RECT 614.800 115.800 615.600 120.400 ;
        RECT 620.400 112.000 621.200 120.400 ;
        RECT 623.600 111.800 624.400 120.400 ;
        RECT 627.800 115.800 628.600 120.400 ;
        RECT 630.600 115.800 631.400 120.400 ;
        RECT 634.800 111.800 635.600 120.400 ;
        RECT 638.000 112.200 638.800 120.400 ;
        RECT 643.200 111.800 644.000 120.400 ;
        RECT 646.000 111.800 646.800 120.400 ;
        RECT 649.200 113.000 650.000 120.400 ;
        RECT 652.400 111.800 653.200 120.400 ;
        RECT 655.600 113.000 656.400 120.400 ;
        RECT 658.800 111.800 659.600 120.400 ;
        RECT 662.000 111.800 662.800 120.400 ;
        RECT 665.200 111.800 666.000 120.400 ;
        RECT 668.400 111.800 669.200 120.400 ;
        RECT 671.600 111.800 672.400 120.400 ;
        RECT 673.200 111.800 674.000 120.400 ;
        RECT 677.400 115.800 678.200 120.400 ;
        RECT 681.200 112.200 682.000 120.400 ;
        RECT 686.400 111.800 687.200 120.400 ;
        RECT 271.000 111.200 298.000 111.800 ;
        RECT 331.800 111.200 358.800 111.800 ;
        RECT 367.000 111.200 394.000 111.800 ;
        RECT 427.800 111.200 454.800 111.800 ;
        RECT 485.400 111.200 512.400 111.800 ;
        RECT 271.000 111.000 271.800 111.200 ;
        RECT 331.800 111.000 332.600 111.200 ;
        RECT 367.000 111.000 367.800 111.200 ;
        RECT 427.800 111.000 428.600 111.200 ;
        RECT 485.400 111.000 486.200 111.200 ;
        RECT 179.800 90.800 180.600 91.000 ;
        RECT 258.200 90.800 259.000 91.000 ;
        RECT 311.000 90.800 311.800 91.000 ;
        RECT 374.600 90.800 375.400 91.000 ;
        RECT 179.800 90.200 206.800 90.800 ;
        RECT 258.200 90.200 285.200 90.800 ;
        RECT 311.000 90.200 338.000 90.800 ;
        RECT 1.800 81.600 2.600 86.200 ;
        RECT 6.000 81.600 6.800 90.200 ;
        RECT 8.800 81.600 9.600 90.200 ;
        RECT 14.000 81.600 14.800 89.800 ;
        RECT 17.800 81.600 18.600 86.200 ;
        RECT 22.000 81.600 22.800 90.200 ;
        RECT 24.200 81.600 25.000 86.200 ;
        RECT 28.400 81.600 29.200 90.200 ;
        RECT 30.000 81.600 30.800 90.200 ;
        RECT 34.200 81.600 35.000 86.200 ;
        RECT 36.400 81.600 37.200 90.200 ;
        RECT 40.600 81.600 41.400 86.200 ;
        RECT 42.800 81.600 43.600 90.200 ;
        RECT 47.000 81.600 47.800 86.200 ;
        RECT 49.800 81.600 50.600 86.200 ;
        RECT 54.000 81.600 54.800 90.200 ;
        RECT 57.200 81.600 58.000 89.800 ;
        RECT 62.400 81.600 63.200 90.200 ;
        RECT 65.200 81.600 66.000 90.200 ;
        RECT 68.400 81.600 69.200 89.000 ;
        RECT 73.200 81.600 74.000 90.200 ;
        RECT 78.800 81.600 79.600 86.200 ;
        RECT 82.000 81.600 82.800 86.200 ;
        RECT 87.600 81.600 88.400 90.000 ;
        RECT 90.800 81.600 91.600 86.200 ;
        RECT 95.600 81.600 96.400 89.000 ;
        RECT 98.800 81.600 99.600 90.200 ;
        RECT 100.400 81.600 101.200 86.200 ;
        RECT 103.600 81.600 104.400 85.800 ;
        RECT 107.400 81.600 108.200 86.200 ;
        RECT 111.600 81.600 112.400 90.200 ;
        RECT 119.600 81.600 120.400 89.000 ;
        RECT 122.800 81.600 123.600 90.200 ;
        RECT 125.600 81.600 126.400 90.200 ;
        RECT 130.800 81.600 131.600 89.800 ;
        RECT 134.000 81.600 134.800 90.200 ;
        RECT 138.200 81.600 139.000 86.200 ;
        RECT 141.000 81.600 141.800 86.200 ;
        RECT 145.200 81.600 146.000 90.200 ;
        RECT 150.000 81.600 150.800 90.200 ;
        RECT 153.200 81.600 154.000 90.000 ;
        RECT 158.800 81.600 159.600 86.200 ;
        RECT 162.000 81.600 162.800 86.200 ;
        RECT 167.600 81.600 168.400 90.200 ;
        RECT 202.600 90.000 203.600 90.200 ;
        RECT 206.000 89.600 206.800 90.200 ;
        RECT 170.800 81.600 171.600 86.200 ;
        RECT 174.000 81.600 174.800 86.200 ;
        RECT 175.600 81.600 176.400 86.200 ;
        RECT 178.800 81.600 179.600 86.200 ;
        RECT 182.000 81.600 182.800 86.200 ;
        RECT 185.200 81.600 186.000 86.200 ;
        RECT 193.200 81.600 194.000 86.200 ;
        RECT 196.400 81.600 197.200 86.200 ;
        RECT 202.800 81.600 203.600 86.200 ;
        RECT 206.000 81.600 206.800 86.200 ;
        RECT 209.200 81.600 210.000 86.200 ;
        RECT 210.800 81.600 211.600 86.200 ;
        RECT 214.000 81.600 214.800 86.200 ;
        RECT 215.600 81.600 216.400 90.200 ;
        RECT 219.800 81.600 220.600 86.200 ;
        RECT 222.000 81.600 222.800 86.200 ;
        RECT 225.200 81.600 226.000 86.200 ;
        RECT 228.400 81.600 229.200 89.800 ;
        RECT 233.200 81.600 234.200 88.800 ;
        RECT 239.400 82.200 240.400 88.800 ;
        RECT 239.400 81.600 240.200 82.200 ;
        RECT 243.400 81.600 244.200 86.200 ;
        RECT 247.600 81.600 248.400 90.200 ;
        RECT 281.000 90.000 281.800 90.200 ;
        RECT 284.400 89.600 285.200 90.200 ;
        RECT 254.000 81.600 254.800 86.200 ;
        RECT 257.200 81.600 258.000 86.200 ;
        RECT 260.400 81.600 261.200 86.200 ;
        RECT 263.600 81.600 264.400 86.200 ;
        RECT 271.600 81.600 272.400 86.200 ;
        RECT 274.800 81.600 275.600 86.200 ;
        RECT 281.200 81.600 282.000 86.200 ;
        RECT 284.400 81.600 285.200 86.200 ;
        RECT 287.600 81.600 288.400 86.200 ;
        RECT 290.800 81.600 291.600 89.000 ;
        RECT 294.000 81.600 294.800 90.200 ;
        RECT 295.600 81.600 296.400 90.200 ;
        RECT 333.800 90.000 334.800 90.200 ;
        RECT 337.200 89.600 338.000 90.200 ;
        RECT 348.400 90.200 375.400 90.800 ;
        RECT 411.800 90.800 412.600 91.000 ;
        RECT 471.000 90.800 471.800 91.000 ;
        RECT 411.800 90.200 438.800 90.800 ;
        RECT 471.000 90.200 498.000 90.800 ;
        RECT 348.400 89.600 349.200 90.200 ;
        RECT 351.600 90.000 352.600 90.200 ;
        RECT 299.800 81.600 300.600 86.200 ;
        RECT 302.000 81.600 302.800 86.200 ;
        RECT 305.200 81.600 306.000 86.200 ;
        RECT 306.800 81.600 307.600 86.200 ;
        RECT 310.000 81.600 310.800 86.200 ;
        RECT 313.200 81.600 314.000 86.200 ;
        RECT 316.400 81.600 317.200 86.200 ;
        RECT 324.400 81.600 325.200 86.200 ;
        RECT 327.600 81.600 328.400 86.200 ;
        RECT 334.000 81.600 334.800 86.200 ;
        RECT 337.200 81.600 338.000 86.200 ;
        RECT 340.400 81.600 341.200 86.200 ;
        RECT 342.000 81.600 342.800 86.200 ;
        RECT 345.200 81.600 346.000 86.200 ;
        RECT 348.400 81.600 349.200 86.200 ;
        RECT 351.600 81.600 352.400 86.200 ;
        RECT 358.000 81.600 358.800 86.200 ;
        RECT 361.200 81.600 362.000 86.200 ;
        RECT 369.200 81.600 370.000 86.200 ;
        RECT 372.400 81.600 373.200 86.200 ;
        RECT 375.600 81.600 376.400 86.200 ;
        RECT 378.800 81.600 379.600 86.200 ;
        RECT 380.400 81.600 381.200 90.200 ;
        RECT 384.600 81.600 385.400 86.200 ;
        RECT 386.800 81.600 387.600 86.200 ;
        RECT 390.000 81.600 390.800 86.200 ;
        RECT 391.600 81.600 392.400 90.200 ;
        RECT 434.600 90.000 435.600 90.200 ;
        RECT 438.000 89.600 438.800 90.200 ;
        RECT 395.800 81.600 396.600 86.200 ;
        RECT 398.000 81.600 398.800 86.200 ;
        RECT 401.200 81.600 402.000 86.200 ;
        RECT 407.600 81.600 408.400 86.200 ;
        RECT 410.800 81.600 411.600 86.200 ;
        RECT 414.000 81.600 414.800 86.200 ;
        RECT 417.200 81.600 418.000 86.200 ;
        RECT 425.200 81.600 426.000 86.200 ;
        RECT 428.400 81.600 429.200 86.200 ;
        RECT 434.800 81.600 435.600 86.200 ;
        RECT 438.000 81.600 438.800 86.200 ;
        RECT 441.200 81.600 442.000 86.200 ;
        RECT 442.800 81.600 443.600 86.200 ;
        RECT 446.000 81.600 446.800 86.200 ;
        RECT 448.200 81.600 449.000 86.200 ;
        RECT 452.400 81.600 453.200 90.200 ;
        RECT 454.600 81.600 455.400 86.200 ;
        RECT 458.800 81.600 459.600 90.200 ;
        RECT 460.400 81.600 461.200 90.200 ;
        RECT 493.800 90.000 494.800 90.200 ;
        RECT 497.200 89.600 498.000 90.200 ;
        RECT 464.600 81.600 465.400 86.200 ;
        RECT 466.800 81.600 467.600 86.200 ;
        RECT 470.000 81.600 470.800 86.200 ;
        RECT 473.200 81.600 474.000 86.200 ;
        RECT 476.400 81.600 477.200 86.200 ;
        RECT 484.400 81.600 485.200 86.200 ;
        RECT 487.600 81.600 488.400 86.200 ;
        RECT 494.000 81.600 494.800 86.200 ;
        RECT 497.200 81.600 498.000 86.200 ;
        RECT 500.400 81.600 501.200 86.200 ;
        RECT 502.000 81.600 502.800 90.200 ;
        RECT 506.200 81.600 507.000 86.200 ;
        RECT 508.400 81.600 509.200 86.200 ;
        RECT 511.600 81.600 512.400 86.200 ;
        RECT 513.200 81.600 514.000 86.200 ;
        RECT 516.400 81.600 517.200 86.200 ;
        RECT 518.000 81.600 518.800 86.200 ;
        RECT 521.200 81.600 522.000 90.200 ;
        RECT 525.400 81.600 526.200 86.200 ;
        RECT 528.200 81.600 529.000 86.200 ;
        RECT 532.400 81.600 533.200 90.200 ;
        RECT 535.600 81.600 536.400 86.200 ;
        RECT 537.800 81.600 538.600 86.200 ;
        RECT 542.000 81.600 542.800 90.200 ;
        RECT 544.200 81.600 545.000 86.200 ;
        RECT 548.400 81.600 549.200 90.200 ;
        RECT 551.600 81.600 552.400 86.200 ;
        RECT 553.800 81.600 554.600 86.200 ;
        RECT 558.000 81.600 558.800 90.200 ;
        RECT 560.200 81.600 561.000 86.200 ;
        RECT 564.400 81.600 565.200 90.200 ;
        RECT 567.200 81.600 568.000 90.200 ;
        RECT 572.400 81.600 573.200 89.800 ;
        RECT 582.000 81.600 582.800 86.200 ;
        RECT 585.200 81.600 586.000 90.200 ;
        RECT 590.800 81.600 591.600 86.200 ;
        RECT 594.000 81.600 594.800 86.200 ;
        RECT 599.600 81.600 600.400 90.000 ;
        RECT 604.400 81.600 605.200 89.800 ;
        RECT 609.600 81.600 610.400 90.200 ;
        RECT 613.000 81.600 613.800 86.200 ;
        RECT 617.200 81.600 618.000 90.200 ;
        RECT 618.800 81.600 619.600 90.200 ;
        RECT 623.000 81.600 623.800 86.200 ;
        RECT 625.800 81.600 626.600 86.200 ;
        RECT 630.000 81.600 630.800 90.200 ;
        RECT 633.200 81.600 634.000 89.000 ;
        RECT 636.400 81.600 637.200 90.200 ;
        RECT 638.000 81.600 638.800 90.200 ;
        RECT 642.200 81.600 643.000 86.200 ;
        RECT 644.400 81.600 645.200 90.200 ;
        RECT 648.600 81.600 649.400 86.200 ;
        RECT 652.400 81.600 653.200 90.200 ;
        RECT 658.000 81.600 658.800 86.200 ;
        RECT 661.200 81.600 662.000 86.200 ;
        RECT 666.800 81.600 667.600 90.000 ;
        RECT 671.600 81.600 672.400 90.000 ;
        RECT 677.200 81.600 678.000 86.200 ;
        RECT 680.400 81.600 681.200 86.200 ;
        RECT 686.000 81.600 686.800 90.200 ;
        RECT 0.400 80.400 689.200 81.600 ;
        RECT 2.800 72.000 3.600 80.400 ;
        RECT 8.400 75.800 9.200 80.400 ;
        RECT 11.600 75.800 12.400 80.400 ;
        RECT 17.200 71.800 18.000 80.400 ;
        RECT 20.400 71.800 21.200 80.400 ;
        RECT 24.600 75.800 25.400 80.400 ;
        RECT 27.400 75.800 28.200 80.400 ;
        RECT 31.600 71.800 32.400 80.400 ;
        RECT 34.800 72.200 35.600 80.400 ;
        RECT 40.000 71.800 40.800 80.400 ;
        RECT 43.400 75.800 44.200 80.400 ;
        RECT 47.600 71.800 48.400 80.400 ;
        RECT 50.400 71.800 51.200 80.400 ;
        RECT 55.600 72.200 56.400 80.400 ;
        RECT 60.000 71.800 60.800 80.400 ;
        RECT 65.200 72.200 66.000 80.400 ;
        RECT 70.000 72.000 70.800 80.400 ;
        RECT 75.600 75.800 76.400 80.400 ;
        RECT 78.800 75.800 79.600 80.400 ;
        RECT 84.400 71.800 85.200 80.400 ;
        RECT 87.600 75.800 88.400 80.400 ;
        RECT 90.800 75.800 91.600 80.400 ;
        RECT 94.000 75.800 94.800 80.400 ;
        RECT 97.200 72.000 98.000 80.400 ;
        RECT 102.800 75.800 103.600 80.400 ;
        RECT 106.000 75.800 106.800 80.400 ;
        RECT 111.600 71.800 112.400 80.400 ;
        RECT 120.200 75.800 121.000 80.400 ;
        RECT 124.400 71.800 125.200 80.400 ;
        RECT 126.000 71.800 126.800 80.400 ;
        RECT 130.200 75.800 131.000 80.400 ;
        RECT 132.400 75.800 133.200 80.400 ;
        RECT 135.600 71.800 136.400 80.400 ;
        RECT 139.800 75.800 140.600 80.400 ;
        RECT 142.000 75.800 142.800 80.400 ;
        RECT 145.200 76.200 146.000 80.400 ;
        RECT 148.400 71.800 149.200 80.400 ;
        RECT 152.600 75.800 153.400 80.400 ;
        RECT 154.800 71.800 155.600 80.400 ;
        RECT 159.000 75.800 159.800 80.400 ;
        RECT 161.200 71.800 162.000 80.400 ;
        RECT 165.400 75.800 166.200 80.400 ;
        RECT 167.600 71.800 168.400 80.400 ;
        RECT 171.800 75.800 172.600 80.400 ;
        RECT 175.600 73.000 176.400 80.400 ;
        RECT 178.800 71.800 179.600 80.400 ;
        RECT 180.400 75.800 181.200 80.400 ;
        RECT 183.600 75.800 184.400 80.400 ;
        RECT 185.200 75.800 186.000 80.400 ;
        RECT 188.400 75.800 189.200 80.400 ;
        RECT 191.600 75.800 192.400 80.400 ;
        RECT 194.800 73.200 195.800 80.400 ;
        RECT 201.000 79.800 201.800 80.400 ;
        RECT 201.000 73.200 202.000 79.800 ;
        RECT 204.400 71.800 205.200 80.400 ;
        RECT 207.600 71.800 208.400 80.400 ;
        RECT 210.800 71.800 211.600 80.400 ;
        RECT 214.000 71.800 214.800 80.400 ;
        RECT 217.200 71.800 218.000 80.400 ;
        RECT 218.800 71.800 219.600 80.400 ;
        RECT 222.000 73.000 222.800 80.400 ;
        RECT 225.200 71.800 226.000 80.400 ;
        RECT 228.400 73.000 229.200 80.400 ;
        RECT 231.600 75.800 232.400 80.400 ;
        RECT 234.800 75.800 235.600 80.400 ;
        RECT 236.400 75.800 237.200 80.400 ;
        RECT 239.600 75.800 240.400 80.400 ;
        RECT 242.800 75.800 243.600 80.400 ;
        RECT 249.200 75.800 250.000 80.400 ;
        RECT 252.400 75.800 253.200 80.400 ;
        RECT 260.400 75.800 261.200 80.400 ;
        RECT 263.600 75.800 264.400 80.400 ;
        RECT 266.800 75.800 267.600 80.400 ;
        RECT 270.000 75.800 270.800 80.400 ;
        RECT 239.600 71.800 240.400 72.400 ;
        RECT 243.000 71.800 243.800 72.000 ;
        RECT 276.400 71.800 277.200 80.400 ;
        RECT 279.600 71.800 280.400 80.400 ;
        RECT 282.800 71.800 283.600 80.400 ;
        RECT 286.000 71.800 286.800 80.400 ;
        RECT 289.200 71.800 290.000 80.400 ;
        RECT 290.800 75.800 291.600 80.400 ;
        RECT 294.000 75.800 294.800 80.400 ;
        RECT 295.600 71.800 296.400 80.400 ;
        RECT 299.800 75.800 300.600 80.400 ;
        RECT 302.000 75.800 302.800 80.400 ;
        RECT 305.200 75.800 306.000 80.400 ;
        RECT 308.400 75.800 309.200 80.400 ;
        RECT 314.800 75.800 315.600 80.400 ;
        RECT 318.000 75.800 318.800 80.400 ;
        RECT 326.000 75.800 326.800 80.400 ;
        RECT 329.200 75.800 330.000 80.400 ;
        RECT 332.400 75.800 333.200 80.400 ;
        RECT 335.600 75.800 336.400 80.400 ;
        RECT 337.200 75.800 338.000 80.400 ;
        RECT 340.400 75.800 341.200 80.400 ;
        RECT 343.600 75.800 344.400 80.400 ;
        RECT 350.000 75.800 350.800 80.400 ;
        RECT 353.200 75.800 354.000 80.400 ;
        RECT 361.200 75.800 362.000 80.400 ;
        RECT 364.400 75.800 365.200 80.400 ;
        RECT 367.600 75.800 368.400 80.400 ;
        RECT 370.800 75.800 371.600 80.400 ;
        RECT 305.200 71.800 306.000 72.400 ;
        RECT 308.400 71.800 309.400 72.000 ;
        RECT 340.400 71.800 341.200 72.400 ;
        RECT 343.800 71.800 344.600 72.000 ;
        RECT 372.400 71.800 373.200 80.400 ;
        RECT 375.600 71.800 376.400 80.400 ;
        RECT 378.800 71.800 379.600 80.400 ;
        RECT 382.000 71.800 382.800 80.400 ;
        RECT 385.200 71.800 386.000 80.400 ;
        RECT 386.800 75.800 387.600 80.400 ;
        RECT 390.000 71.800 390.800 80.400 ;
        RECT 394.200 75.800 395.000 80.400 ;
        RECT 396.400 75.800 397.200 80.400 ;
        RECT 399.600 75.800 400.400 80.400 ;
        RECT 401.200 75.800 402.000 80.400 ;
        RECT 404.400 75.800 405.200 80.400 ;
        RECT 410.800 75.800 411.600 80.400 ;
        RECT 414.000 75.800 414.800 80.400 ;
        RECT 417.200 75.800 418.000 80.400 ;
        RECT 420.400 75.800 421.200 80.400 ;
        RECT 428.400 75.800 429.200 80.400 ;
        RECT 431.600 75.800 432.400 80.400 ;
        RECT 438.000 75.800 438.800 80.400 ;
        RECT 441.200 75.800 442.000 80.400 ;
        RECT 444.400 75.800 445.200 80.400 ;
        RECT 446.000 75.800 446.800 80.400 ;
        RECT 449.200 75.800 450.000 80.400 ;
        RECT 451.400 75.800 452.200 80.400 ;
        RECT 437.800 71.800 438.800 72.000 ;
        RECT 441.200 71.800 442.000 72.400 ;
        RECT 455.600 71.800 456.400 80.400 ;
        RECT 457.200 71.800 458.000 80.400 ;
        RECT 460.400 71.800 461.200 80.400 ;
        RECT 463.600 71.800 464.400 80.400 ;
        RECT 465.200 75.800 466.000 80.400 ;
        RECT 468.400 75.800 469.200 80.400 ;
        RECT 471.600 75.800 472.400 80.400 ;
        RECT 478.000 75.800 478.800 80.400 ;
        RECT 481.200 75.800 482.000 80.400 ;
        RECT 489.200 75.800 490.000 80.400 ;
        RECT 492.400 75.800 493.200 80.400 ;
        RECT 495.600 75.800 496.400 80.400 ;
        RECT 498.800 75.800 499.600 80.400 ;
        RECT 502.000 75.800 502.800 80.400 ;
        RECT 503.600 75.800 504.400 80.400 ;
        RECT 468.400 71.800 469.200 72.400 ;
        RECT 471.800 71.800 472.600 72.000 ;
        RECT 506.800 71.800 507.600 80.400 ;
        RECT 511.000 75.800 511.800 80.400 ;
        RECT 513.800 75.800 514.600 80.400 ;
        RECT 518.000 71.800 518.800 80.400 ;
        RECT 519.600 71.800 520.400 80.400 ;
        RECT 522.800 71.800 523.600 80.400 ;
        RECT 526.000 71.800 526.800 80.400 ;
        RECT 529.200 71.800 530.000 80.400 ;
        RECT 532.400 71.800 533.200 80.400 ;
        RECT 535.600 72.000 536.400 80.400 ;
        RECT 541.200 75.800 542.000 80.400 ;
        RECT 544.400 75.800 545.200 80.400 ;
        RECT 550.000 71.800 550.800 80.400 ;
        RECT 554.800 76.200 555.600 80.400 ;
        RECT 558.000 75.800 558.800 80.400 ;
        RECT 559.600 71.800 560.400 80.400 ;
        RECT 563.800 75.800 564.600 80.400 ;
        RECT 566.600 75.800 567.400 80.400 ;
        RECT 570.800 71.800 571.600 80.400 ;
        RECT 577.800 75.800 578.600 80.400 ;
        RECT 582.000 71.800 582.800 80.400 ;
        RECT 585.200 76.200 586.000 80.400 ;
        RECT 588.400 75.800 589.200 80.400 ;
        RECT 591.600 71.800 592.400 80.400 ;
        RECT 597.200 75.800 598.000 80.400 ;
        RECT 600.400 75.800 601.200 80.400 ;
        RECT 606.000 72.000 606.800 80.400 ;
        RECT 610.800 76.200 611.600 80.400 ;
        RECT 614.000 75.800 614.800 80.400 ;
        RECT 615.600 71.800 616.400 80.400 ;
        RECT 619.800 75.800 620.600 80.400 ;
        RECT 623.600 76.200 624.400 80.400 ;
        RECT 626.800 75.800 627.600 80.400 ;
        RECT 630.000 72.200 630.800 80.400 ;
        RECT 635.200 71.800 636.000 80.400 ;
        RECT 638.000 71.800 638.800 80.400 ;
        RECT 642.200 75.800 643.000 80.400 ;
        RECT 646.000 71.800 646.800 80.400 ;
        RECT 651.600 75.800 652.400 80.400 ;
        RECT 654.800 75.800 655.600 80.400 ;
        RECT 660.400 72.000 661.200 80.400 ;
        RECT 664.200 75.800 665.000 80.400 ;
        RECT 668.400 71.800 669.200 80.400 ;
        RECT 671.600 75.800 672.400 80.400 ;
        RECT 673.200 71.800 674.000 80.400 ;
        RECT 676.400 71.800 677.200 80.400 ;
        RECT 679.600 71.800 680.400 80.400 ;
        RECT 682.800 71.800 683.600 80.400 ;
        RECT 686.000 71.800 686.800 80.400 ;
        RECT 239.600 71.200 266.600 71.800 ;
        RECT 305.200 71.200 332.200 71.800 ;
        RECT 340.400 71.200 367.400 71.800 ;
        RECT 265.800 71.000 266.600 71.200 ;
        RECT 331.400 71.000 332.200 71.200 ;
        RECT 366.600 71.000 367.400 71.200 ;
        RECT 415.000 71.200 442.000 71.800 ;
        RECT 468.400 71.200 495.400 71.800 ;
        RECT 415.000 71.000 415.800 71.200 ;
        RECT 494.600 71.000 495.400 71.200 ;
        RECT 179.800 50.800 180.600 51.000 ;
        RECT 246.600 50.800 247.400 51.000 ;
        RECT 293.000 50.800 293.800 51.000 ;
        RECT 179.800 50.200 206.800 50.800 ;
        RECT 220.400 50.200 247.400 50.800 ;
        RECT 266.800 50.200 293.800 50.800 ;
        RECT 319.000 50.800 319.800 51.000 ;
        RECT 362.200 50.800 363.000 51.000 ;
        RECT 402.200 50.800 403.000 51.000 ;
        RECT 488.200 50.800 489.000 51.000 ;
        RECT 319.000 50.200 346.000 50.800 ;
        RECT 362.200 50.200 389.200 50.800 ;
        RECT 402.200 50.200 429.200 50.800 ;
        RECT 462.000 50.200 489.000 50.800 ;
        RECT 2.800 41.600 3.600 50.000 ;
        RECT 8.400 41.600 9.200 46.200 ;
        RECT 11.600 41.600 12.400 46.200 ;
        RECT 17.200 41.600 18.000 50.200 ;
        RECT 20.400 41.600 21.200 50.200 ;
        RECT 24.600 41.600 25.400 46.200 ;
        RECT 27.400 41.600 28.200 46.200 ;
        RECT 31.600 41.600 32.400 50.200 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 38.000 41.600 38.800 46.200 ;
        RECT 41.200 41.600 42.000 46.200 ;
        RECT 44.000 41.600 44.800 50.200 ;
        RECT 49.200 41.600 50.000 49.800 ;
        RECT 52.400 41.600 53.200 50.200 ;
        RECT 56.600 41.600 57.400 46.200 ;
        RECT 59.400 41.600 60.200 46.200 ;
        RECT 63.600 41.600 64.400 50.200 ;
        RECT 66.800 41.600 67.600 50.000 ;
        RECT 72.400 41.600 73.200 46.200 ;
        RECT 75.600 41.600 76.400 46.200 ;
        RECT 81.200 41.600 82.000 50.200 ;
        RECT 84.400 41.600 85.200 46.200 ;
        RECT 87.600 41.600 88.400 46.200 ;
        RECT 89.200 41.600 90.000 46.200 ;
        RECT 92.400 41.600 93.200 46.200 ;
        RECT 95.600 41.600 96.400 49.800 ;
        RECT 100.800 41.600 101.600 50.200 ;
        RECT 104.800 41.600 105.600 50.200 ;
        RECT 110.000 41.600 110.800 49.800 ;
        RECT 118.000 41.600 118.800 50.200 ;
        RECT 122.200 41.600 123.000 46.200 ;
        RECT 124.400 41.600 125.200 50.200 ;
        RECT 128.600 41.600 129.400 46.200 ;
        RECT 130.800 41.600 131.600 50.200 ;
        RECT 135.000 41.600 135.800 46.200 ;
        RECT 138.800 41.600 139.600 49.800 ;
        RECT 144.000 41.600 144.800 50.200 ;
        RECT 146.800 41.600 147.600 46.200 ;
        RECT 151.200 41.600 152.000 50.200 ;
        RECT 156.400 41.600 157.200 49.800 ;
        RECT 159.600 41.600 160.400 46.200 ;
        RECT 162.800 41.600 163.600 50.200 ;
        RECT 202.600 50.000 203.600 50.200 ;
        RECT 206.000 49.600 206.800 50.200 ;
        RECT 167.000 41.600 167.800 46.200 ;
        RECT 169.200 41.600 170.000 46.200 ;
        RECT 172.400 41.600 173.200 45.800 ;
        RECT 175.600 41.600 176.400 46.200 ;
        RECT 178.800 41.600 179.600 46.200 ;
        RECT 182.000 41.600 182.800 46.200 ;
        RECT 185.200 41.600 186.000 46.200 ;
        RECT 193.200 41.600 194.000 46.200 ;
        RECT 196.400 41.600 197.200 46.200 ;
        RECT 202.800 41.600 203.600 46.200 ;
        RECT 206.000 41.600 206.800 46.200 ;
        RECT 209.200 41.600 210.000 46.200 ;
        RECT 210.800 41.600 211.600 50.200 ;
        RECT 220.400 49.600 221.200 50.200 ;
        RECT 223.600 50.000 224.600 50.200 ;
        RECT 214.000 41.600 214.800 49.000 ;
        RECT 217.200 41.600 218.000 46.200 ;
        RECT 220.400 41.600 221.200 46.200 ;
        RECT 223.600 41.600 224.400 46.200 ;
        RECT 230.000 41.600 230.800 46.200 ;
        RECT 233.200 41.600 234.000 46.200 ;
        RECT 241.200 41.600 242.000 46.200 ;
        RECT 244.400 41.600 245.200 46.200 ;
        RECT 247.600 41.600 248.400 46.200 ;
        RECT 250.800 41.600 251.600 46.200 ;
        RECT 253.000 41.600 253.800 46.200 ;
        RECT 257.200 41.600 258.000 50.200 ;
        RECT 266.800 49.600 267.600 50.200 ;
        RECT 270.000 50.000 271.000 50.200 ;
        RECT 263.600 41.600 264.400 46.200 ;
        RECT 266.800 41.600 267.600 46.200 ;
        RECT 270.000 41.600 270.800 46.200 ;
        RECT 276.400 41.600 277.200 46.200 ;
        RECT 279.600 41.600 280.400 46.200 ;
        RECT 287.600 41.600 288.400 46.200 ;
        RECT 290.800 41.600 291.600 46.200 ;
        RECT 294.000 41.600 294.800 46.200 ;
        RECT 297.200 41.600 298.000 46.200 ;
        RECT 298.800 41.600 299.600 46.200 ;
        RECT 302.000 41.600 302.800 46.200 ;
        RECT 304.200 41.600 305.000 46.200 ;
        RECT 308.400 41.600 309.200 50.200 ;
        RECT 341.800 50.000 342.800 50.200 ;
        RECT 345.200 49.600 346.000 50.200 ;
        RECT 310.000 41.600 310.800 46.200 ;
        RECT 313.200 41.600 314.000 46.200 ;
        RECT 314.800 41.600 315.600 46.200 ;
        RECT 318.000 41.600 318.800 46.200 ;
        RECT 321.200 41.600 322.000 46.200 ;
        RECT 324.400 41.600 325.200 46.200 ;
        RECT 332.400 41.600 333.200 46.200 ;
        RECT 335.600 41.600 336.400 46.200 ;
        RECT 342.000 41.600 342.800 46.200 ;
        RECT 345.200 41.600 346.000 46.200 ;
        RECT 348.400 41.600 349.200 46.200 ;
        RECT 350.000 41.600 350.800 50.200 ;
        RECT 353.200 41.600 354.000 50.200 ;
        RECT 356.400 41.600 357.200 50.200 ;
        RECT 385.000 50.000 385.800 50.200 ;
        RECT 388.400 49.600 389.200 50.200 ;
        RECT 425.000 50.000 426.000 50.200 ;
        RECT 428.400 49.600 429.200 50.200 ;
        RECT 358.000 41.600 358.800 46.200 ;
        RECT 361.200 41.600 362.000 46.200 ;
        RECT 364.400 41.600 365.200 46.200 ;
        RECT 367.600 41.600 368.400 46.200 ;
        RECT 375.600 41.600 376.400 46.200 ;
        RECT 378.800 41.600 379.600 46.200 ;
        RECT 385.200 41.600 386.000 46.200 ;
        RECT 388.400 41.600 389.200 46.200 ;
        RECT 391.600 41.600 392.400 46.200 ;
        RECT 393.200 41.600 394.000 46.200 ;
        RECT 396.400 41.600 397.200 46.200 ;
        RECT 398.000 41.600 398.800 46.200 ;
        RECT 401.200 41.600 402.000 46.200 ;
        RECT 404.400 41.600 405.200 46.200 ;
        RECT 407.600 41.600 408.400 46.200 ;
        RECT 415.600 41.600 416.400 46.200 ;
        RECT 418.800 41.600 419.600 46.200 ;
        RECT 425.200 41.600 426.000 46.200 ;
        RECT 428.400 41.600 429.200 46.200 ;
        RECT 431.600 41.600 432.400 46.200 ;
        RECT 438.000 41.600 438.800 46.200 ;
        RECT 441.200 41.600 442.000 46.200 ;
        RECT 445.400 41.600 446.200 50.200 ;
        RECT 462.000 49.600 462.800 50.200 ;
        RECT 465.200 50.000 466.200 50.200 ;
        RECT 449.200 41.600 450.000 46.200 ;
        RECT 452.400 41.600 453.200 46.200 ;
        RECT 454.000 41.600 454.800 46.200 ;
        RECT 457.200 41.600 458.000 46.200 ;
        RECT 458.800 41.600 459.600 46.200 ;
        RECT 462.000 41.600 462.800 46.200 ;
        RECT 465.200 41.600 466.000 46.200 ;
        RECT 471.600 41.600 472.400 46.200 ;
        RECT 474.800 41.600 475.600 46.200 ;
        RECT 482.800 41.600 483.600 46.200 ;
        RECT 486.000 41.600 486.800 46.200 ;
        RECT 489.200 41.600 490.000 46.200 ;
        RECT 492.400 41.600 493.200 46.200 ;
        RECT 494.600 41.600 495.400 46.200 ;
        RECT 498.800 41.600 499.600 50.200 ;
        RECT 501.000 41.600 501.800 46.200 ;
        RECT 505.200 41.600 506.000 50.200 ;
        RECT 506.800 41.600 507.600 46.200 ;
        RECT 510.000 41.600 510.800 46.200 ;
        RECT 512.200 41.600 513.000 46.200 ;
        RECT 516.400 41.600 517.200 50.200 ;
        RECT 518.000 41.600 518.800 50.200 ;
        RECT 521.200 41.600 522.000 49.000 ;
        RECT 524.400 41.600 525.200 46.200 ;
        RECT 527.600 41.600 528.400 46.200 ;
        RECT 529.200 41.600 530.000 50.200 ;
        RECT 533.400 41.600 534.200 46.200 ;
        RECT 536.200 41.600 537.000 46.200 ;
        RECT 540.400 41.600 541.200 50.200 ;
        RECT 543.200 41.600 544.000 50.200 ;
        RECT 548.400 41.600 549.200 49.800 ;
        RECT 551.600 41.600 552.400 50.200 ;
        RECT 555.800 41.600 556.600 46.200 ;
        RECT 558.000 41.600 558.800 46.200 ;
        RECT 561.200 41.600 562.000 46.200 ;
        RECT 563.400 41.600 564.200 46.200 ;
        RECT 567.600 41.600 568.400 50.200 ;
        RECT 575.600 41.600 576.600 48.800 ;
        RECT 581.800 42.200 582.800 48.800 ;
        RECT 581.800 41.600 582.600 42.200 ;
        RECT 585.200 41.600 586.000 46.200 ;
        RECT 588.400 41.600 589.200 46.200 ;
        RECT 591.200 41.600 592.000 50.200 ;
        RECT 596.400 41.600 597.200 49.800 ;
        RECT 601.200 41.600 602.000 50.200 ;
        RECT 606.800 41.600 607.600 46.200 ;
        RECT 610.000 41.600 610.800 46.200 ;
        RECT 615.600 41.600 616.400 50.000 ;
        RECT 620.400 41.600 621.200 49.800 ;
        RECT 625.600 41.600 626.400 50.200 ;
        RECT 628.400 41.600 629.200 50.200 ;
        RECT 631.600 41.600 632.400 49.000 ;
        RECT 636.400 41.600 637.200 49.800 ;
        RECT 641.600 41.600 642.400 50.200 ;
        RECT 645.000 41.600 645.800 46.200 ;
        RECT 649.200 41.600 650.000 50.200 ;
        RECT 651.400 41.600 652.200 46.200 ;
        RECT 655.600 41.600 656.400 50.200 ;
        RECT 658.400 41.600 659.200 50.200 ;
        RECT 663.600 41.600 664.400 49.800 ;
        RECT 668.400 41.600 669.200 49.800 ;
        RECT 673.600 41.600 674.400 50.200 ;
        RECT 676.400 41.600 677.200 50.200 ;
        RECT 680.600 41.600 681.400 46.200 ;
        RECT 683.400 41.600 684.200 46.200 ;
        RECT 687.600 41.600 688.400 50.200 ;
        RECT 0.400 40.400 689.200 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 4.400 35.800 5.200 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 14.000 35.800 14.800 40.400 ;
        RECT 17.200 35.800 18.000 40.400 ;
        RECT 25.200 35.800 26.000 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 36.400 35.800 37.200 40.400 ;
        RECT 4.400 31.800 5.200 32.400 ;
        RECT 7.800 31.800 8.600 32.000 ;
        RECT 39.600 31.800 40.400 40.400 ;
        RECT 43.800 35.800 44.600 40.400 ;
        RECT 46.600 35.800 47.400 40.400 ;
        RECT 50.800 31.800 51.600 40.400 ;
        RECT 52.400 31.800 53.200 40.400 ;
        RECT 56.600 35.800 57.400 40.400 ;
        RECT 58.800 31.800 59.600 40.400 ;
        RECT 63.000 35.800 63.800 40.400 ;
        RECT 65.200 31.800 66.000 40.400 ;
        RECT 68.400 31.800 69.200 40.400 ;
        RECT 71.600 31.800 72.400 40.400 ;
        RECT 74.800 31.800 75.600 40.400 ;
        RECT 78.000 31.800 78.800 40.400 ;
        RECT 79.600 31.800 80.400 40.400 ;
        RECT 82.800 31.800 83.600 40.400 ;
        RECT 86.000 31.800 86.800 40.400 ;
        RECT 89.200 31.800 90.000 40.400 ;
        RECT 92.400 31.800 93.200 40.400 ;
        RECT 94.600 35.800 95.400 40.400 ;
        RECT 98.800 31.800 99.600 40.400 ;
        RECT 101.000 35.800 101.800 40.400 ;
        RECT 105.200 31.800 106.000 40.400 ;
        RECT 107.400 35.800 108.200 40.400 ;
        RECT 111.600 31.800 112.400 40.400 ;
        RECT 119.600 32.000 120.400 40.400 ;
        RECT 125.200 35.800 126.000 40.400 ;
        RECT 128.400 35.800 129.200 40.400 ;
        RECT 134.000 31.800 134.800 40.400 ;
        RECT 137.200 31.800 138.000 40.400 ;
        RECT 141.400 35.800 142.200 40.400 ;
        RECT 143.600 35.800 144.400 40.400 ;
        RECT 146.800 35.800 147.600 40.400 ;
        RECT 149.000 35.800 149.800 40.400 ;
        RECT 153.200 31.800 154.000 40.400 ;
        RECT 156.400 32.000 157.200 40.400 ;
        RECT 162.000 35.800 162.800 40.400 ;
        RECT 165.200 35.800 166.000 40.400 ;
        RECT 170.800 31.800 171.600 40.400 ;
        RECT 174.000 31.800 174.800 40.400 ;
        RECT 180.400 35.800 181.200 40.400 ;
        RECT 182.000 31.800 182.800 40.400 ;
        RECT 188.600 39.800 189.400 40.400 ;
        RECT 188.400 33.200 189.400 39.800 ;
        RECT 194.600 33.200 195.600 40.400 ;
        RECT 198.000 35.800 198.800 40.400 ;
        RECT 201.200 35.800 202.000 40.400 ;
        RECT 204.400 35.800 205.200 40.400 ;
        RECT 207.600 35.800 208.400 40.400 ;
        RECT 215.600 35.800 216.400 40.400 ;
        RECT 218.800 35.800 219.600 40.400 ;
        RECT 225.200 35.800 226.000 40.400 ;
        RECT 228.400 35.800 229.200 40.400 ;
        RECT 231.600 35.800 232.400 40.400 ;
        RECT 233.200 35.800 234.000 40.400 ;
        RECT 236.400 35.800 237.200 40.400 ;
        RECT 239.600 35.800 240.400 40.400 ;
        RECT 246.000 35.800 246.800 40.400 ;
        RECT 249.200 35.800 250.000 40.400 ;
        RECT 257.200 35.800 258.000 40.400 ;
        RECT 260.400 35.800 261.200 40.400 ;
        RECT 263.600 35.800 264.400 40.400 ;
        RECT 266.800 35.800 267.600 40.400 ;
        RECT 225.000 31.800 225.800 32.000 ;
        RECT 228.400 31.800 229.200 32.400 ;
        RECT 4.400 31.200 31.400 31.800 ;
        RECT 30.600 31.000 31.400 31.200 ;
        RECT 202.200 31.200 229.200 31.800 ;
        RECT 236.400 31.800 237.200 32.400 ;
        RECT 239.600 31.800 240.600 32.000 ;
        RECT 273.200 31.800 274.000 40.400 ;
        RECT 277.400 35.800 278.200 40.400 ;
        RECT 279.600 35.800 280.400 40.400 ;
        RECT 282.800 35.800 283.600 40.400 ;
        RECT 284.400 35.800 285.200 40.400 ;
        RECT 287.600 35.800 288.400 40.400 ;
        RECT 289.200 31.800 290.000 40.400 ;
        RECT 292.400 31.800 293.200 40.400 ;
        RECT 295.600 31.800 296.400 40.400 ;
        RECT 298.800 31.800 299.600 40.400 ;
        RECT 302.000 31.800 302.800 40.400 ;
        RECT 303.600 31.800 304.400 40.400 ;
        RECT 307.800 35.800 308.600 40.400 ;
        RECT 311.600 35.800 312.400 40.400 ;
        RECT 313.200 35.800 314.000 40.400 ;
        RECT 316.400 35.800 317.200 40.400 ;
        RECT 319.600 35.800 320.400 40.400 ;
        RECT 322.800 35.800 323.600 40.400 ;
        RECT 330.800 35.800 331.600 40.400 ;
        RECT 334.000 35.800 334.800 40.400 ;
        RECT 340.400 35.800 341.200 40.400 ;
        RECT 343.600 35.800 344.400 40.400 ;
        RECT 346.800 35.800 347.600 40.400 ;
        RECT 340.200 31.800 341.200 32.000 ;
        RECT 343.600 31.800 344.400 32.400 ;
        RECT 348.400 31.800 349.200 40.400 ;
        RECT 351.600 31.800 352.400 40.400 ;
        RECT 354.800 31.800 355.600 40.400 ;
        RECT 358.000 31.800 358.800 40.400 ;
        RECT 361.200 31.800 362.000 40.400 ;
        RECT 362.800 35.800 363.600 40.400 ;
        RECT 366.000 31.800 366.800 40.400 ;
        RECT 370.200 35.800 371.000 40.400 ;
        RECT 372.400 35.800 373.200 40.400 ;
        RECT 375.600 35.800 376.400 40.400 ;
        RECT 378.800 35.800 379.600 40.400 ;
        RECT 385.200 35.800 386.000 40.400 ;
        RECT 388.400 35.800 389.200 40.400 ;
        RECT 396.400 35.800 397.200 40.400 ;
        RECT 399.600 35.800 400.400 40.400 ;
        RECT 402.800 35.800 403.600 40.400 ;
        RECT 406.000 35.800 406.800 40.400 ;
        RECT 407.600 35.800 408.400 40.400 ;
        RECT 411.400 35.800 412.200 40.400 ;
        RECT 375.600 31.800 376.400 32.400 ;
        RECT 379.000 31.800 379.800 32.000 ;
        RECT 415.600 31.800 416.400 40.400 ;
        RECT 422.600 35.800 423.400 40.400 ;
        RECT 426.800 31.800 427.600 40.400 ;
        RECT 430.000 35.800 430.800 40.400 ;
        RECT 431.600 35.800 432.400 40.400 ;
        RECT 434.800 35.800 435.600 40.400 ;
        RECT 438.000 35.800 438.800 40.400 ;
        RECT 444.400 35.800 445.200 40.400 ;
        RECT 447.600 35.800 448.400 40.400 ;
        RECT 455.600 35.800 456.400 40.400 ;
        RECT 458.800 35.800 459.600 40.400 ;
        RECT 462.000 35.800 462.800 40.400 ;
        RECT 465.200 35.800 466.000 40.400 ;
        RECT 434.800 31.800 435.600 32.400 ;
        RECT 438.000 31.800 439.000 32.000 ;
        RECT 466.800 31.800 467.600 40.400 ;
        RECT 471.000 35.800 471.800 40.400 ;
        RECT 473.800 35.800 474.600 40.400 ;
        RECT 478.000 31.800 478.800 40.400 ;
        RECT 480.200 35.800 481.000 40.400 ;
        RECT 484.400 31.800 485.200 40.400 ;
        RECT 486.600 35.800 487.400 40.400 ;
        RECT 490.800 31.800 491.600 40.400 ;
        RECT 494.000 35.800 494.800 40.400 ;
        RECT 495.600 35.800 496.400 40.400 ;
        RECT 498.800 35.800 499.600 40.400 ;
        RECT 502.000 35.800 502.800 40.400 ;
        RECT 505.200 35.800 506.000 40.400 ;
        RECT 513.200 35.800 514.000 40.400 ;
        RECT 516.400 35.800 517.200 40.400 ;
        RECT 522.800 35.800 523.600 40.400 ;
        RECT 526.000 35.800 526.800 40.400 ;
        RECT 529.200 35.800 530.000 40.400 ;
        RECT 531.400 35.800 532.200 40.400 ;
        RECT 522.600 31.800 523.400 32.000 ;
        RECT 526.000 31.800 526.800 32.400 ;
        RECT 535.600 31.800 536.400 40.400 ;
        RECT 537.200 31.800 538.000 40.400 ;
        RECT 541.400 35.800 542.200 40.400 ;
        RECT 544.200 35.800 545.000 40.400 ;
        RECT 548.400 31.800 549.200 40.400 ;
        RECT 550.000 31.800 550.800 40.400 ;
        RECT 554.200 35.800 555.000 40.400 ;
        RECT 556.400 35.800 557.200 40.400 ;
        RECT 559.600 35.800 560.400 40.400 ;
        RECT 562.400 31.800 563.200 40.400 ;
        RECT 567.600 32.200 568.400 40.400 ;
        RECT 577.200 31.800 578.000 40.400 ;
        RECT 582.800 35.800 583.600 40.400 ;
        RECT 586.000 35.800 586.800 40.400 ;
        RECT 591.600 32.000 592.400 40.400 ;
        RECT 596.400 35.800 597.200 40.400 ;
        RECT 599.600 31.800 600.400 40.400 ;
        RECT 605.200 35.800 606.000 40.400 ;
        RECT 608.400 35.800 609.200 40.400 ;
        RECT 614.000 32.000 614.800 40.400 ;
        RECT 617.200 31.800 618.000 40.400 ;
        RECT 621.400 35.800 622.200 40.400 ;
        RECT 624.200 35.800 625.000 40.400 ;
        RECT 628.400 31.800 629.200 40.400 ;
        RECT 631.200 31.800 632.000 40.400 ;
        RECT 636.400 32.200 637.200 40.400 ;
        RECT 641.200 32.200 642.000 40.400 ;
        RECT 646.400 31.800 647.200 40.400 ;
        RECT 649.200 31.800 650.000 40.400 ;
        RECT 653.400 35.800 654.200 40.400 ;
        RECT 656.200 35.800 657.000 40.400 ;
        RECT 660.400 31.800 661.200 40.400 ;
        RECT 662.000 31.800 662.800 40.400 ;
        RECT 666.200 35.800 667.000 40.400 ;
        RECT 669.000 35.800 669.800 40.400 ;
        RECT 673.200 31.800 674.000 40.400 ;
        RECT 676.400 33.200 677.400 40.400 ;
        RECT 682.600 39.800 683.400 40.400 ;
        RECT 682.600 33.200 683.600 39.800 ;
        RECT 236.400 31.200 263.400 31.800 ;
        RECT 202.200 31.000 203.000 31.200 ;
        RECT 262.600 31.000 263.400 31.200 ;
        RECT 317.400 31.200 344.400 31.800 ;
        RECT 375.600 31.200 402.600 31.800 ;
        RECT 434.800 31.200 461.800 31.800 ;
        RECT 317.400 31.000 318.200 31.200 ;
        RECT 401.800 31.000 402.600 31.200 ;
        RECT 461.000 31.000 461.800 31.200 ;
        RECT 499.800 31.200 526.800 31.800 ;
        RECT 499.800 31.000 500.600 31.200 ;
        RECT 33.800 10.800 34.600 11.000 ;
        RECT 7.600 10.200 34.600 10.800 ;
        RECT 51.800 10.800 52.600 11.000 ;
        RECT 87.000 10.800 87.800 11.000 ;
        RECT 170.200 10.800 171.000 11.000 ;
        RECT 230.600 10.800 231.400 11.000 ;
        RECT 51.800 10.200 78.800 10.800 ;
        RECT 87.000 10.200 114.000 10.800 ;
        RECT 170.200 10.200 197.200 10.800 ;
        RECT 7.600 9.600 8.400 10.200 ;
        RECT 10.800 10.000 11.800 10.200 ;
        RECT 74.600 10.000 75.400 10.200 ;
        RECT 78.000 9.600 78.800 10.200 ;
        RECT 109.800 10.000 110.600 10.200 ;
        RECT 113.200 9.600 114.000 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 10.800 1.600 11.600 6.200 ;
        RECT 17.200 1.600 18.000 6.200 ;
        RECT 20.400 1.600 21.200 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 38.000 1.600 38.800 6.200 ;
        RECT 41.200 1.600 42.000 9.000 ;
        RECT 44.400 1.600 45.200 6.200 ;
        RECT 47.600 1.600 48.400 6.200 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 54.000 1.600 54.800 6.200 ;
        RECT 57.200 1.600 58.000 6.200 ;
        RECT 65.200 1.600 66.000 6.200 ;
        RECT 68.400 1.600 69.200 6.200 ;
        RECT 74.800 1.600 75.600 6.200 ;
        RECT 78.000 1.600 78.800 6.200 ;
        RECT 81.200 1.600 82.000 6.200 ;
        RECT 82.800 1.600 83.600 6.200 ;
        RECT 86.000 1.600 86.800 6.200 ;
        RECT 89.200 1.600 90.000 6.200 ;
        RECT 92.400 1.600 93.200 6.200 ;
        RECT 100.400 1.600 101.200 6.200 ;
        RECT 103.600 1.600 104.400 6.200 ;
        RECT 110.000 1.600 110.800 6.200 ;
        RECT 113.200 1.600 114.000 6.200 ;
        RECT 116.400 1.600 117.200 6.200 ;
        RECT 124.400 1.600 125.200 10.000 ;
        RECT 130.000 1.600 130.800 6.200 ;
        RECT 133.200 1.600 134.000 6.200 ;
        RECT 138.800 1.600 139.600 10.200 ;
        RECT 145.200 1.600 146.000 10.200 ;
        RECT 148.400 2.200 149.400 8.800 ;
        RECT 148.600 1.600 149.400 2.200 ;
        RECT 154.600 1.600 155.600 8.800 ;
        RECT 159.600 1.600 160.400 6.200 ;
        RECT 161.200 1.600 162.000 10.200 ;
        RECT 193.000 10.000 193.800 10.200 ;
        RECT 196.400 9.600 197.200 10.200 ;
        RECT 204.400 10.200 231.400 10.800 ;
        RECT 287.000 10.800 287.800 11.000 ;
        RECT 339.800 10.800 340.600 11.000 ;
        RECT 409.800 10.800 410.600 11.000 ;
        RECT 454.600 10.800 455.400 11.000 ;
        RECT 287.000 10.200 314.000 10.800 ;
        RECT 339.800 10.200 366.800 10.800 ;
        RECT 204.400 9.600 205.200 10.200 ;
        RECT 207.600 10.000 208.600 10.200 ;
        RECT 166.000 1.600 166.800 6.200 ;
        RECT 169.200 1.600 170.000 6.200 ;
        RECT 172.400 1.600 173.200 6.200 ;
        RECT 175.600 1.600 176.400 6.200 ;
        RECT 183.600 1.600 184.400 6.200 ;
        RECT 186.800 1.600 187.600 6.200 ;
        RECT 193.200 1.600 194.000 6.200 ;
        RECT 196.400 1.600 197.200 6.200 ;
        RECT 199.600 1.600 200.400 6.200 ;
        RECT 201.200 1.600 202.000 6.200 ;
        RECT 204.400 1.600 205.200 6.200 ;
        RECT 207.600 1.600 208.400 6.200 ;
        RECT 214.000 1.600 214.800 6.200 ;
        RECT 217.200 1.600 218.000 6.200 ;
        RECT 225.200 1.600 226.000 6.200 ;
        RECT 228.400 1.600 229.200 6.200 ;
        RECT 231.600 1.600 232.400 6.200 ;
        RECT 234.800 1.600 235.600 6.200 ;
        RECT 236.400 1.600 237.200 6.200 ;
        RECT 241.200 1.600 242.000 9.000 ;
        RECT 245.000 1.600 245.800 6.200 ;
        RECT 249.200 1.600 250.000 10.200 ;
        RECT 250.800 1.600 251.600 6.200 ;
        RECT 254.000 1.600 254.800 6.200 ;
        RECT 257.200 1.600 258.000 9.000 ;
        RECT 260.400 1.600 261.200 6.200 ;
        RECT 270.000 1.600 270.800 9.000 ;
        RECT 273.200 1.600 274.000 6.200 ;
        RECT 276.400 1.600 277.200 10.200 ;
        RECT 309.800 10.000 310.800 10.200 ;
        RECT 313.200 9.600 314.000 10.200 ;
        RECT 280.600 1.600 281.400 6.200 ;
        RECT 282.800 1.600 283.600 6.200 ;
        RECT 286.000 1.600 286.800 6.200 ;
        RECT 289.200 1.600 290.000 6.200 ;
        RECT 292.400 1.600 293.200 6.200 ;
        RECT 300.400 1.600 301.200 6.200 ;
        RECT 303.600 1.600 304.400 6.200 ;
        RECT 310.000 1.600 310.800 6.200 ;
        RECT 313.200 1.600 314.000 6.200 ;
        RECT 316.400 1.600 317.200 6.200 ;
        RECT 319.600 1.600 320.400 9.000 ;
        RECT 322.800 1.600 323.600 10.200 ;
        RECT 326.000 1.600 326.800 10.200 ;
        RECT 329.200 1.600 330.000 10.200 ;
        RECT 362.600 10.000 363.400 10.200 ;
        RECT 366.000 9.600 366.800 10.200 ;
        RECT 383.600 10.200 410.600 10.800 ;
        RECT 428.400 10.200 455.400 10.800 ;
        RECT 471.000 10.800 471.800 11.000 ;
        RECT 534.600 10.800 535.400 11.000 ;
        RECT 573.000 10.800 573.800 11.000 ;
        RECT 471.000 10.200 498.000 10.800 ;
        RECT 383.600 9.600 384.400 10.200 ;
        RECT 387.000 10.000 387.800 10.200 ;
        RECT 428.400 9.600 429.200 10.200 ;
        RECT 431.800 10.000 432.600 10.200 ;
        RECT 493.800 10.000 494.800 10.200 ;
        RECT 497.200 9.600 498.000 10.200 ;
        RECT 508.400 10.200 535.400 10.800 ;
        RECT 546.800 10.200 573.800 10.800 ;
        RECT 508.400 9.600 509.200 10.200 ;
        RECT 511.800 10.000 512.600 10.200 ;
        RECT 546.800 9.600 547.600 10.200 ;
        RECT 550.000 10.000 551.000 10.200 ;
        RECT 332.400 1.600 333.200 9.000 ;
        RECT 335.600 1.600 336.400 6.200 ;
        RECT 338.800 1.600 339.600 6.200 ;
        RECT 342.000 1.600 342.800 6.200 ;
        RECT 345.200 1.600 346.000 6.200 ;
        RECT 353.200 1.600 354.000 6.200 ;
        RECT 356.400 1.600 357.200 6.200 ;
        RECT 362.800 1.600 363.600 6.200 ;
        RECT 366.000 1.600 366.800 6.200 ;
        RECT 369.200 1.600 370.000 6.200 ;
        RECT 372.400 1.600 373.200 9.000 ;
        RECT 377.200 1.600 378.000 9.000 ;
        RECT 380.400 1.600 381.200 6.200 ;
        RECT 383.600 1.600 384.400 6.200 ;
        RECT 386.800 1.600 387.600 6.200 ;
        RECT 393.200 1.600 394.000 6.200 ;
        RECT 396.400 1.600 397.200 6.200 ;
        RECT 404.400 1.600 405.200 6.200 ;
        RECT 407.600 1.600 408.400 6.200 ;
        RECT 410.800 1.600 411.600 6.200 ;
        RECT 414.000 1.600 414.800 6.200 ;
        RECT 417.200 1.600 418.000 9.000 ;
        RECT 425.200 1.600 426.000 6.200 ;
        RECT 428.400 1.600 429.200 6.200 ;
        RECT 431.600 1.600 432.400 6.200 ;
        RECT 438.000 1.600 438.800 6.200 ;
        RECT 441.200 1.600 442.000 6.200 ;
        RECT 449.200 1.600 450.000 6.200 ;
        RECT 452.400 1.600 453.200 6.200 ;
        RECT 455.600 1.600 456.400 6.200 ;
        RECT 458.800 1.600 459.600 6.200 ;
        RECT 462.000 1.600 462.800 6.200 ;
        RECT 463.600 1.600 464.400 6.200 ;
        RECT 466.800 1.600 467.600 6.200 ;
        RECT 470.000 1.600 470.800 6.200 ;
        RECT 473.200 1.600 474.000 6.200 ;
        RECT 476.400 1.600 477.200 6.200 ;
        RECT 484.400 1.600 485.200 6.200 ;
        RECT 487.600 1.600 488.400 6.200 ;
        RECT 494.000 1.600 494.800 6.200 ;
        RECT 497.200 1.600 498.000 6.200 ;
        RECT 500.400 1.600 501.200 6.200 ;
        RECT 502.000 1.600 502.800 6.200 ;
        RECT 505.200 1.600 506.000 6.200 ;
        RECT 508.400 1.600 509.200 6.200 ;
        RECT 511.600 1.600 512.400 6.200 ;
        RECT 518.000 1.600 518.800 6.200 ;
        RECT 521.200 1.600 522.000 6.200 ;
        RECT 529.200 1.600 530.000 6.200 ;
        RECT 532.400 1.600 533.200 6.200 ;
        RECT 535.600 1.600 536.400 6.200 ;
        RECT 538.800 1.600 539.600 6.200 ;
        RECT 542.000 1.600 542.800 6.200 ;
        RECT 543.600 1.600 544.400 6.200 ;
        RECT 546.800 1.600 547.600 6.200 ;
        RECT 550.000 1.600 550.800 6.200 ;
        RECT 556.400 1.600 557.200 6.200 ;
        RECT 559.600 1.600 560.400 6.200 ;
        RECT 567.600 1.600 568.400 6.200 ;
        RECT 570.800 1.600 571.600 6.200 ;
        RECT 574.000 1.600 574.800 6.200 ;
        RECT 577.200 1.600 578.000 6.200 ;
        RECT 585.200 1.600 586.000 9.000 ;
        RECT 590.000 1.600 590.800 10.200 ;
        RECT 595.600 1.600 596.400 6.200 ;
        RECT 598.800 1.600 599.600 6.200 ;
        RECT 604.400 1.600 605.200 10.000 ;
        RECT 607.600 1.600 608.400 10.200 ;
        RECT 611.800 1.600 612.600 6.200 ;
        RECT 614.600 1.600 615.400 6.200 ;
        RECT 618.800 1.600 619.600 10.200 ;
        RECT 620.400 1.600 621.200 10.200 ;
        RECT 624.600 1.600 625.400 6.200 ;
        RECT 627.400 1.600 628.200 6.200 ;
        RECT 631.600 1.600 632.400 10.200 ;
        RECT 634.800 1.600 635.600 6.200 ;
        RECT 637.000 1.600 637.800 6.200 ;
        RECT 641.200 1.600 642.000 10.200 ;
        RECT 644.400 1.600 645.200 10.200 ;
        RECT 650.000 1.600 650.800 6.200 ;
        RECT 653.200 1.600 654.000 6.200 ;
        RECT 658.800 1.600 659.600 10.000 ;
        RECT 663.600 1.600 664.400 10.200 ;
        RECT 669.200 1.600 670.000 6.200 ;
        RECT 672.400 1.600 673.200 6.200 ;
        RECT 678.000 1.600 678.800 10.000 ;
        RECT 681.800 1.600 682.600 6.200 ;
        RECT 686.000 1.600 686.800 10.200 ;
        RECT 0.400 0.400 689.200 1.600 ;
      LAYER via1 ;
        RECT 4.400 483.600 5.200 484.400 ;
        RECT 52.400 483.600 53.200 484.400 ;
        RECT 196.400 483.600 197.200 484.400 ;
        RECT 234.800 483.600 235.600 484.400 ;
        RECT 372.400 490.000 373.200 490.800 ;
        RECT 412.400 490.000 413.200 490.800 ;
        RECT 262.000 483.600 262.800 484.400 ;
        RECT 302.000 483.600 302.800 484.400 ;
        RECT 372.400 485.400 373.200 486.200 ;
        RECT 412.400 485.400 413.200 486.200 ;
        RECT 518.000 490.000 518.800 490.800 ;
        RECT 474.800 483.600 475.600 484.400 ;
        RECT 518.000 485.400 518.800 486.200 ;
        RECT 577.200 490.000 578.000 490.800 ;
        RECT 577.200 485.400 578.000 486.200 ;
        RECT 593.200 483.600 594.000 484.400 ;
        RECT 681.200 483.600 682.000 484.400 ;
        RECT 111.800 480.600 112.600 481.400 ;
        RECT 113.200 480.600 114.000 481.400 ;
        RECT 114.600 480.600 115.400 481.400 ;
        RECT 415.800 480.600 416.600 481.400 ;
        RECT 417.200 480.600 418.000 481.400 ;
        RECT 418.600 480.600 419.400 481.400 ;
        RECT 31.600 477.600 32.400 478.400 ;
        RECT 31.600 471.600 32.400 472.400 ;
        RECT 215.600 477.600 216.400 478.400 ;
        RECT 215.600 471.600 216.400 472.400 ;
        RECT 258.800 471.200 259.600 472.000 ;
        RECT 380.400 477.600 381.200 478.400 ;
        RECT 380.400 471.600 381.200 472.400 ;
        RECT 474.800 477.600 475.600 478.400 ;
        RECT 474.800 471.600 475.600 472.400 ;
        RECT 486.000 471.200 486.800 472.000 ;
        RECT 562.800 477.600 563.600 478.400 ;
        RECT 562.800 471.600 563.600 472.400 ;
        RECT 254.000 450.000 254.800 450.800 ;
        RECT 254.000 445.400 254.800 446.200 ;
        RECT 273.200 443.600 274.000 444.400 ;
        RECT 420.400 450.000 421.200 450.800 ;
        RECT 420.400 445.400 421.200 446.200 ;
        RECT 444.400 445.400 445.200 446.200 ;
        RECT 500.400 443.600 501.200 444.400 ;
        RECT 588.400 450.000 589.200 450.800 ;
        RECT 588.400 445.400 589.200 446.200 ;
        RECT 665.200 443.600 666.000 444.400 ;
        RECT 111.800 440.600 112.600 441.400 ;
        RECT 113.200 440.600 114.000 441.400 ;
        RECT 114.600 440.600 115.400 441.400 ;
        RECT 415.800 440.600 416.600 441.400 ;
        RECT 417.200 440.600 418.000 441.400 ;
        RECT 418.600 440.600 419.400 441.400 ;
        RECT 266.800 431.200 267.600 432.000 ;
        RECT 412.400 431.200 413.200 432.000 ;
        RECT 468.400 437.600 469.200 438.400 ;
        RECT 468.400 431.600 469.200 432.400 ;
        RECT 630.000 437.600 630.800 438.400 ;
        RECT 630.000 431.600 630.800 432.400 ;
        RECT 676.400 431.200 677.200 432.000 ;
        RECT 562.800 429.600 563.600 430.400 ;
        RECT 278.000 411.600 278.800 412.400 ;
        RECT 218.800 410.000 219.600 410.800 ;
        RECT 218.800 405.400 219.600 406.200 ;
        RECT 278.000 405.600 278.800 406.400 ;
        RECT 442.800 410.000 443.600 410.800 ;
        RECT 442.800 403.600 443.600 404.400 ;
        RECT 454.000 403.600 454.800 404.400 ;
        RECT 538.800 403.600 539.600 404.400 ;
        RECT 604.400 410.000 605.200 410.800 ;
        RECT 604.400 405.400 605.200 406.200 ;
        RECT 676.400 410.000 677.200 410.800 ;
        RECT 676.400 405.400 677.200 406.200 ;
        RECT 111.800 400.600 112.600 401.400 ;
        RECT 113.200 400.600 114.000 401.400 ;
        RECT 114.600 400.600 115.400 401.400 ;
        RECT 415.800 400.600 416.600 401.400 ;
        RECT 417.200 400.600 418.000 401.400 ;
        RECT 418.600 400.600 419.400 401.400 ;
        RECT 286.000 391.200 286.800 392.000 ;
        RECT 388.400 397.600 389.200 398.400 ;
        RECT 388.400 391.600 389.200 392.400 ;
        RECT 478.000 397.600 478.800 398.400 ;
        RECT 478.000 391.600 478.800 392.400 ;
        RECT 652.400 397.600 653.200 398.400 ;
        RECT 652.400 391.600 653.200 392.400 ;
        RECT 183.600 363.600 184.400 364.400 ;
        RECT 244.400 365.400 245.200 366.200 ;
        RECT 446.000 363.600 446.800 364.400 ;
        RECT 454.000 363.600 454.800 364.400 ;
        RECT 679.600 370.000 680.400 370.800 ;
        RECT 679.600 363.600 680.400 364.400 ;
        RECT 111.800 360.600 112.600 361.400 ;
        RECT 113.200 360.600 114.000 361.400 ;
        RECT 114.600 360.600 115.400 361.400 ;
        RECT 415.800 360.600 416.600 361.400 ;
        RECT 417.200 360.600 418.000 361.400 ;
        RECT 418.600 360.600 419.400 361.400 ;
        RECT 174.000 357.600 174.800 358.400 ;
        RECT 174.000 351.600 174.800 352.400 ;
        RECT 247.600 351.200 248.400 352.000 ;
        RECT 412.400 351.200 413.200 352.000 ;
        RECT 466.800 357.600 467.600 358.400 ;
        RECT 466.800 351.600 467.600 352.400 ;
        RECT 194.800 330.000 195.600 330.800 ;
        RECT 194.800 325.400 195.600 326.200 ;
        RECT 260.400 323.600 261.200 324.400 ;
        RECT 276.400 325.400 277.200 326.200 ;
        RECT 462.000 330.000 462.800 330.800 ;
        RECT 462.000 325.400 462.800 326.200 ;
        RECT 111.800 320.600 112.600 321.400 ;
        RECT 113.200 320.600 114.000 321.400 ;
        RECT 114.600 320.600 115.400 321.400 ;
        RECT 415.800 320.600 416.600 321.400 ;
        RECT 417.200 320.600 418.000 321.400 ;
        RECT 418.600 320.600 419.400 321.400 ;
        RECT 4.400 317.600 5.200 318.400 ;
        RECT 4.400 311.600 5.200 312.400 ;
        RECT 65.200 317.600 66.000 318.400 ;
        RECT 114.800 317.600 115.600 318.400 ;
        RECT 65.200 311.600 66.000 312.400 ;
        RECT 114.800 311.600 115.600 312.400 ;
        RECT 194.800 311.200 195.600 312.000 ;
        RECT 260.400 311.200 261.200 312.000 ;
        RECT 398.000 317.600 398.800 318.400 ;
        RECT 398.000 311.600 398.800 312.400 ;
        RECT 414.000 311.200 414.800 312.000 ;
        RECT 68.400 283.600 69.200 284.400 ;
        RECT 121.200 283.600 122.000 284.400 ;
        RECT 167.600 283.600 168.400 284.400 ;
        RECT 212.400 285.400 213.200 286.200 ;
        RECT 265.200 283.600 266.000 284.400 ;
        RECT 398.000 283.600 398.800 284.400 ;
        RECT 423.600 283.600 424.400 284.400 ;
        RECT 111.800 280.600 112.600 281.400 ;
        RECT 113.200 280.600 114.000 281.400 ;
        RECT 114.600 280.600 115.400 281.400 ;
        RECT 415.800 280.600 416.600 281.400 ;
        RECT 417.200 280.600 418.000 281.400 ;
        RECT 418.600 280.600 419.400 281.400 ;
        RECT 4.400 277.600 5.200 278.400 ;
        RECT 4.400 271.600 5.200 272.400 ;
        RECT 97.200 277.600 98.000 278.400 ;
        RECT 97.200 271.600 98.000 272.400 ;
        RECT 162.800 271.200 163.600 272.000 ;
        RECT 218.800 277.600 219.600 278.400 ;
        RECT 218.800 271.600 219.600 272.400 ;
        RECT 258.800 277.600 259.600 278.400 ;
        RECT 258.800 271.600 259.600 272.400 ;
        RECT 300.400 271.200 301.200 272.000 ;
        RECT 430.000 277.600 430.800 278.400 ;
        RECT 468.400 277.600 469.200 278.400 ;
        RECT 430.000 271.600 430.800 272.400 ;
        RECT 468.400 271.600 469.200 272.400 ;
        RECT 114.800 250.000 115.600 250.800 ;
        RECT 44.400 243.600 45.200 244.400 ;
        RECT 79.600 243.600 80.400 244.400 ;
        RECT 114.800 245.400 115.600 246.200 ;
        RECT 250.800 250.000 251.600 250.800 ;
        RECT 191.600 245.400 192.400 246.200 ;
        RECT 250.800 245.400 251.600 246.200 ;
        RECT 300.400 250.000 301.200 250.800 ;
        RECT 300.400 245.400 301.200 246.200 ;
        RECT 430.000 245.400 430.800 246.200 ;
        RECT 518.000 245.400 518.800 246.200 ;
        RECT 111.800 240.600 112.600 241.400 ;
        RECT 113.200 240.600 114.000 241.400 ;
        RECT 114.600 240.600 115.400 241.400 ;
        RECT 415.800 240.600 416.600 241.400 ;
        RECT 417.200 240.600 418.000 241.400 ;
        RECT 418.600 240.600 419.400 241.400 ;
        RECT 52.400 237.600 53.200 238.400 ;
        RECT 52.400 231.600 53.200 232.400 ;
        RECT 90.800 237.600 91.600 238.400 ;
        RECT 90.800 231.600 91.600 232.400 ;
        RECT 166.000 231.200 166.800 232.000 ;
        RECT 214.000 231.200 214.800 232.000 ;
        RECT 244.400 231.200 245.200 232.000 ;
        RECT 324.400 231.200 325.200 232.000 ;
        RECT 390.000 237.600 390.800 238.400 ;
        RECT 390.000 231.600 390.800 232.400 ;
        RECT 460.400 231.200 461.200 232.000 ;
        RECT 508.400 231.200 509.200 232.000 ;
        RECT 606.000 237.600 606.800 238.400 ;
        RECT 606.000 231.600 606.800 232.400 ;
        RECT 633.200 237.600 634.000 238.400 ;
        RECT 633.200 231.600 634.000 232.400 ;
        RECT 470.000 211.600 470.800 212.400 ;
        RECT 14.000 203.600 14.800 204.400 ;
        RECT 90.800 203.600 91.600 204.400 ;
        RECT 145.200 210.000 146.000 210.800 ;
        RECT 145.200 205.400 146.000 206.200 ;
        RECT 183.600 203.600 184.400 204.400 ;
        RECT 191.600 203.600 192.400 204.400 ;
        RECT 268.400 203.600 269.200 204.400 ;
        RECT 382.000 210.000 382.800 210.800 ;
        RECT 382.000 205.400 382.800 206.200 ;
        RECT 414.000 205.400 414.800 206.200 ;
        RECT 470.000 205.600 470.800 206.400 ;
        RECT 494.000 205.400 494.800 206.200 ;
        RECT 641.200 203.600 642.000 204.400 ;
        RECT 111.800 200.600 112.600 201.400 ;
        RECT 113.200 200.600 114.000 201.400 ;
        RECT 114.600 200.600 115.400 201.400 ;
        RECT 415.800 200.600 416.600 201.400 ;
        RECT 417.200 200.600 418.000 201.400 ;
        RECT 418.600 200.600 419.400 201.400 ;
        RECT 20.400 197.600 21.200 198.400 ;
        RECT 20.400 191.600 21.200 192.400 ;
        RECT 212.400 197.600 213.200 198.400 ;
        RECT 212.400 191.600 213.200 192.400 ;
        RECT 258.800 197.600 259.600 198.400 ;
        RECT 298.800 197.600 299.600 198.400 ;
        RECT 310.000 197.600 310.800 198.400 ;
        RECT 258.800 191.600 259.600 192.400 ;
        RECT 298.800 191.600 299.600 192.400 ;
        RECT 310.000 191.600 310.800 192.400 ;
        RECT 454.000 191.200 454.800 192.000 ;
        RECT 4.400 163.600 5.200 164.400 ;
        RECT 79.600 163.600 80.400 164.400 ;
        RECT 250.800 163.600 251.600 164.400 ;
        RECT 278.000 165.400 278.800 166.200 ;
        RECT 386.800 170.000 387.600 170.800 ;
        RECT 327.600 163.600 328.400 164.400 ;
        RECT 386.800 163.600 387.600 164.400 ;
        RECT 442.800 170.000 443.600 170.800 ;
        RECT 442.800 163.600 443.600 164.400 ;
        RECT 508.400 163.600 509.200 164.400 ;
        RECT 681.200 170.000 682.000 170.800 ;
        RECT 681.200 165.400 682.000 166.200 ;
        RECT 111.800 160.600 112.600 161.400 ;
        RECT 113.200 160.600 114.000 161.400 ;
        RECT 114.600 160.600 115.400 161.400 ;
        RECT 415.800 160.600 416.600 161.400 ;
        RECT 417.200 160.600 418.000 161.400 ;
        RECT 418.600 160.600 419.400 161.400 ;
        RECT 316.400 157.600 317.200 158.400 ;
        RECT 378.800 157.600 379.600 158.400 ;
        RECT 316.400 151.600 317.200 152.400 ;
        RECT 378.800 151.600 379.600 152.400 ;
        RECT 390.000 151.200 390.800 152.000 ;
        RECT 479.600 157.600 480.400 158.400 ;
        RECT 444.400 151.200 445.200 152.000 ;
        RECT 479.600 151.600 480.400 152.400 ;
        RECT 295.600 149.600 296.400 150.400 ;
        RECT 228.400 130.000 229.200 130.800 ;
        RECT 228.400 123.600 229.200 124.400 ;
        RECT 334.000 130.000 334.800 130.800 ;
        RECT 334.000 125.400 334.800 126.200 ;
        RECT 358.000 125.400 358.800 126.200 ;
        RECT 420.400 130.000 421.200 130.800 ;
        RECT 420.400 125.400 421.200 126.200 ;
        RECT 447.600 123.600 448.400 124.400 ;
        RECT 479.600 123.600 480.400 124.400 ;
        RECT 111.800 120.600 112.600 121.400 ;
        RECT 113.200 120.600 114.000 121.400 ;
        RECT 114.600 120.600 115.400 121.400 ;
        RECT 415.800 120.600 416.600 121.400 ;
        RECT 417.200 120.600 418.000 121.400 ;
        RECT 418.600 120.600 419.400 121.400 ;
        RECT 294.000 111.200 294.800 112.000 ;
        RECT 358.000 117.600 358.800 118.400 ;
        RECT 358.000 111.600 358.800 112.400 ;
        RECT 390.000 111.200 390.800 112.000 ;
        RECT 454.000 117.600 454.800 118.400 ;
        RECT 454.000 111.600 454.800 112.400 ;
        RECT 508.400 111.200 509.200 112.000 ;
        RECT 202.800 90.000 203.600 90.800 ;
        RECT 202.800 85.400 203.600 86.200 ;
        RECT 284.400 83.600 285.200 84.400 ;
        RECT 334.000 90.000 334.800 90.800 ;
        RECT 334.000 85.400 334.800 86.200 ;
        RECT 351.600 83.600 352.400 84.400 ;
        RECT 434.800 90.000 435.600 90.800 ;
        RECT 434.800 83.600 435.600 84.400 ;
        RECT 494.000 90.000 494.800 90.800 ;
        RECT 494.000 85.400 494.800 86.200 ;
        RECT 111.800 80.600 112.600 81.400 ;
        RECT 113.200 80.600 114.000 81.400 ;
        RECT 114.600 80.600 115.400 81.400 ;
        RECT 415.800 80.600 416.600 81.400 ;
        RECT 417.200 80.600 418.000 81.400 ;
        RECT 418.600 80.600 419.400 81.400 ;
        RECT 239.600 77.600 240.400 78.400 ;
        RECT 239.600 71.600 240.400 72.400 ;
        RECT 340.400 77.600 341.200 78.400 ;
        RECT 308.400 71.200 309.200 72.000 ;
        RECT 340.400 71.600 341.200 72.400 ;
        RECT 438.000 71.200 438.800 72.000 ;
        RECT 468.400 77.600 469.200 78.400 ;
        RECT 468.400 71.600 469.200 72.400 ;
        RECT 202.800 50.000 203.600 50.800 ;
        RECT 202.800 45.400 203.600 46.200 ;
        RECT 223.600 45.400 224.400 46.200 ;
        RECT 270.000 45.400 270.800 46.200 ;
        RECT 342.000 50.000 342.800 50.800 ;
        RECT 342.000 45.400 342.800 46.200 ;
        RECT 425.200 50.000 426.000 50.800 ;
        RECT 388.400 43.600 389.200 44.400 ;
        RECT 425.200 43.600 426.000 44.400 ;
        RECT 465.200 43.600 466.000 44.400 ;
        RECT 111.800 40.600 112.600 41.400 ;
        RECT 113.200 40.600 114.000 41.400 ;
        RECT 114.600 40.600 115.400 41.400 ;
        RECT 415.800 40.600 416.600 41.400 ;
        RECT 417.200 40.600 418.000 41.400 ;
        RECT 418.600 40.600 419.400 41.400 ;
        RECT 4.400 37.600 5.200 38.400 ;
        RECT 4.400 31.600 5.200 32.400 ;
        RECT 228.400 37.600 229.200 38.400 ;
        RECT 228.400 31.600 229.200 32.400 ;
        RECT 239.600 31.200 240.400 32.000 ;
        RECT 340.400 31.200 341.200 32.000 ;
        RECT 375.600 37.600 376.400 38.400 ;
        RECT 375.600 31.600 376.400 32.400 ;
        RECT 438.000 31.200 438.800 32.000 ;
        RECT 526.000 37.600 526.800 38.400 ;
        RECT 526.000 31.600 526.800 32.400 ;
        RECT 10.800 3.600 11.600 4.400 ;
        RECT 78.000 3.600 78.800 4.400 ;
        RECT 113.200 3.600 114.000 4.400 ;
        RECT 196.400 3.600 197.200 4.400 ;
        RECT 207.600 5.400 208.400 6.200 ;
        RECT 310.000 10.000 310.800 10.800 ;
        RECT 310.000 5.400 310.800 6.200 ;
        RECT 494.000 10.000 494.800 10.800 ;
        RECT 366.000 3.600 366.800 4.400 ;
        RECT 383.600 3.600 384.400 4.400 ;
        RECT 428.400 3.600 429.200 4.400 ;
        RECT 494.000 5.400 494.800 6.200 ;
        RECT 508.400 3.600 509.200 4.400 ;
        RECT 550.000 5.400 550.800 6.200 ;
        RECT 111.800 0.600 112.600 1.400 ;
        RECT 113.200 0.600 114.000 1.400 ;
        RECT 114.600 0.600 115.400 1.400 ;
        RECT 415.800 0.600 416.600 1.400 ;
        RECT 417.200 0.600 418.000 1.400 ;
        RECT 418.600 0.600 419.400 1.400 ;
      LAYER metal2 ;
        RECT 4.400 489.600 5.200 490.400 ;
        RECT 52.400 490.000 53.200 490.800 ;
        RECT 4.500 484.400 5.100 489.600 ;
        RECT 52.500 484.400 53.100 490.000 ;
        RECT 196.400 489.600 197.200 490.400 ;
        RECT 234.800 489.600 235.600 490.400 ;
        RECT 262.000 489.600 262.800 490.400 ;
        RECT 302.000 489.600 302.800 490.400 ;
        RECT 372.400 490.000 373.200 490.800 ;
        RECT 412.400 490.000 413.200 490.800 ;
        RECT 196.500 484.400 197.100 489.600 ;
        RECT 234.900 484.400 235.500 489.600 ;
        RECT 262.100 484.400 262.700 489.600 ;
        RECT 302.100 484.400 302.700 489.600 ;
        RECT 372.500 486.200 373.100 490.000 ;
        RECT 412.500 486.200 413.100 490.000 ;
        RECT 474.800 489.600 475.600 490.400 ;
        RECT 518.000 490.000 518.800 490.800 ;
        RECT 577.200 490.000 578.000 490.800 ;
        RECT 372.400 485.400 373.200 486.200 ;
        RECT 412.400 485.400 413.200 486.200 ;
        RECT 474.900 484.400 475.500 489.600 ;
        RECT 518.100 486.200 518.700 490.000 ;
        RECT 577.300 486.200 577.900 490.000 ;
        RECT 593.200 489.600 594.000 490.400 ;
        RECT 681.200 489.600 682.000 490.400 ;
        RECT 518.000 485.400 518.800 486.200 ;
        RECT 577.200 485.400 578.000 486.200 ;
        RECT 593.300 484.400 593.900 489.600 ;
        RECT 681.300 484.400 681.900 489.600 ;
        RECT 4.400 483.600 5.200 484.400 ;
        RECT 52.400 483.600 53.200 484.400 ;
        RECT 196.400 483.600 197.200 484.400 ;
        RECT 234.800 483.600 235.600 484.400 ;
        RECT 262.000 483.600 262.800 484.400 ;
        RECT 302.000 483.600 302.800 484.400 ;
        RECT 474.800 483.600 475.600 484.400 ;
        RECT 593.200 483.600 594.000 484.400 ;
        RECT 681.200 483.600 682.000 484.400 ;
        RECT 111.200 480.600 116.000 481.400 ;
        RECT 415.200 480.600 420.000 481.400 ;
        RECT 31.600 477.600 32.400 478.400 ;
        RECT 215.600 477.600 216.400 478.400 ;
        RECT 380.400 477.600 381.200 478.400 ;
        RECT 474.800 477.600 475.600 478.400 ;
        RECT 562.800 477.600 563.600 478.400 ;
        RECT 31.700 472.400 32.300 477.600 ;
        RECT 215.700 472.400 216.300 477.600 ;
        RECT 258.800 475.800 259.600 476.600 ;
        RECT 31.600 471.600 32.400 472.400 ;
        RECT 215.600 471.600 216.400 472.400 ;
        RECT 258.900 472.000 259.500 475.800 ;
        RECT 380.500 472.400 381.100 477.600 ;
        RECT 474.900 472.400 475.500 477.600 ;
        RECT 486.000 475.800 486.800 476.600 ;
        RECT 258.800 471.200 259.600 472.000 ;
        RECT 380.400 471.600 381.200 472.400 ;
        RECT 474.800 471.600 475.600 472.400 ;
        RECT 486.100 472.000 486.700 475.800 ;
        RECT 562.900 472.400 563.500 477.600 ;
        RECT 486.000 471.200 486.800 472.000 ;
        RECT 562.800 471.600 563.600 472.400 ;
        RECT 254.000 450.000 254.800 450.800 ;
        RECT 273.200 450.000 274.000 450.800 ;
        RECT 420.400 450.000 421.200 450.800 ;
        RECT 444.400 450.000 445.200 450.800 ;
        RECT 254.100 446.200 254.700 450.000 ;
        RECT 254.000 445.400 254.800 446.200 ;
        RECT 273.300 444.400 273.900 450.000 ;
        RECT 420.500 446.200 421.100 450.000 ;
        RECT 444.500 446.200 445.100 450.000 ;
        RECT 500.400 449.600 501.200 450.400 ;
        RECT 588.400 450.000 589.200 450.800 ;
        RECT 420.400 445.400 421.200 446.200 ;
        RECT 444.400 445.400 445.200 446.200 ;
        RECT 500.500 444.400 501.100 449.600 ;
        RECT 588.500 446.200 589.100 450.000 ;
        RECT 665.200 449.600 666.000 450.400 ;
        RECT 588.400 445.400 589.200 446.200 ;
        RECT 665.300 444.400 665.900 449.600 ;
        RECT 273.200 443.600 274.000 444.400 ;
        RECT 500.400 443.600 501.200 444.400 ;
        RECT 665.200 443.600 666.000 444.400 ;
        RECT 111.200 440.600 116.000 441.400 ;
        RECT 415.200 440.600 420.000 441.400 ;
        RECT 468.400 437.600 469.200 438.400 ;
        RECT 630.000 437.600 630.800 438.400 ;
        RECT 266.800 435.800 267.600 436.600 ;
        RECT 412.400 435.800 413.200 436.600 ;
        RECT 266.900 432.000 267.500 435.800 ;
        RECT 412.500 432.000 413.100 435.800 ;
        RECT 468.500 432.400 469.100 437.600 ;
        RECT 562.800 435.800 563.600 436.600 ;
        RECT 266.800 431.200 267.600 432.000 ;
        RECT 412.400 431.200 413.200 432.000 ;
        RECT 468.400 431.600 469.200 432.400 ;
        RECT 562.900 430.400 563.500 435.800 ;
        RECT 630.100 432.400 630.700 437.600 ;
        RECT 676.400 435.800 677.200 436.600 ;
        RECT 630.000 431.600 630.800 432.400 ;
        RECT 676.500 432.000 677.100 435.800 ;
        RECT 676.400 431.200 677.200 432.000 ;
        RECT 562.800 429.600 563.600 430.400 ;
        RECT 278.000 411.600 278.800 412.400 ;
        RECT 218.800 410.000 219.600 410.800 ;
        RECT 218.900 406.200 219.500 410.000 ;
        RECT 278.100 406.400 278.700 411.600 ;
        RECT 442.800 410.000 443.600 410.800 ;
        RECT 218.800 405.400 219.600 406.200 ;
        RECT 278.000 405.600 278.800 406.400 ;
        RECT 442.900 404.400 443.500 410.000 ;
        RECT 454.000 409.600 454.800 410.400 ;
        RECT 538.800 409.600 539.600 410.400 ;
        RECT 604.400 410.000 605.200 410.800 ;
        RECT 676.400 410.000 677.200 410.800 ;
        RECT 454.100 404.400 454.700 409.600 ;
        RECT 538.900 404.400 539.500 409.600 ;
        RECT 604.500 406.200 605.100 410.000 ;
        RECT 676.500 406.200 677.100 410.000 ;
        RECT 604.400 405.400 605.200 406.200 ;
        RECT 676.400 405.400 677.200 406.200 ;
        RECT 442.800 403.600 443.600 404.400 ;
        RECT 454.000 403.600 454.800 404.400 ;
        RECT 538.800 403.600 539.600 404.400 ;
        RECT 111.200 400.600 116.000 401.400 ;
        RECT 415.200 400.600 420.000 401.400 ;
        RECT 388.400 397.600 389.200 398.400 ;
        RECT 478.000 397.600 478.800 398.400 ;
        RECT 652.400 397.600 653.200 398.400 ;
        RECT 286.000 395.800 286.800 396.600 ;
        RECT 286.100 392.000 286.700 395.800 ;
        RECT 388.500 392.400 389.100 397.600 ;
        RECT 478.100 392.400 478.700 397.600 ;
        RECT 652.500 392.400 653.100 397.600 ;
        RECT 286.000 391.200 286.800 392.000 ;
        RECT 388.400 391.600 389.200 392.400 ;
        RECT 478.000 391.600 478.800 392.400 ;
        RECT 652.400 391.600 653.200 392.400 ;
        RECT 183.600 369.600 184.400 370.400 ;
        RECT 244.400 370.000 245.200 370.800 ;
        RECT 183.700 364.400 184.300 369.600 ;
        RECT 244.500 366.200 245.100 370.000 ;
        RECT 446.000 369.600 446.800 370.400 ;
        RECT 454.000 369.600 454.800 370.400 ;
        RECT 679.600 370.000 680.400 370.800 ;
        RECT 244.400 365.400 245.200 366.200 ;
        RECT 446.100 364.400 446.700 369.600 ;
        RECT 454.100 364.400 454.700 369.600 ;
        RECT 679.700 364.400 680.300 370.000 ;
        RECT 183.600 363.600 184.400 364.400 ;
        RECT 446.000 363.600 446.800 364.400 ;
        RECT 454.000 363.600 454.800 364.400 ;
        RECT 679.600 363.600 680.400 364.400 ;
        RECT 111.200 360.600 116.000 361.400 ;
        RECT 415.200 360.600 420.000 361.400 ;
        RECT 174.000 357.600 174.800 358.400 ;
        RECT 466.800 357.600 467.600 358.400 ;
        RECT 174.100 352.400 174.700 357.600 ;
        RECT 247.600 355.800 248.400 356.600 ;
        RECT 412.400 355.800 413.200 356.600 ;
        RECT 174.000 351.600 174.800 352.400 ;
        RECT 247.700 352.000 248.300 355.800 ;
        RECT 412.500 352.000 413.100 355.800 ;
        RECT 466.900 352.400 467.500 357.600 ;
        RECT 247.600 351.200 248.400 352.000 ;
        RECT 412.400 351.200 413.200 352.000 ;
        RECT 466.800 351.600 467.600 352.400 ;
        RECT 194.800 330.000 195.600 330.800 ;
        RECT 194.900 326.200 195.500 330.000 ;
        RECT 260.400 329.600 261.200 330.400 ;
        RECT 276.400 330.000 277.200 330.800 ;
        RECT 462.000 330.000 462.800 330.800 ;
        RECT 194.800 325.400 195.600 326.200 ;
        RECT 260.500 324.400 261.100 329.600 ;
        RECT 276.500 326.200 277.100 330.000 ;
        RECT 462.100 326.200 462.700 330.000 ;
        RECT 276.400 325.400 277.200 326.200 ;
        RECT 462.000 325.400 462.800 326.200 ;
        RECT 260.400 323.600 261.200 324.400 ;
        RECT 111.200 320.600 116.000 321.400 ;
        RECT 415.200 320.600 420.000 321.400 ;
        RECT 4.400 317.600 5.200 318.400 ;
        RECT 65.200 317.600 66.000 318.400 ;
        RECT 114.800 317.600 115.600 318.400 ;
        RECT 398.000 317.600 398.800 318.400 ;
        RECT 4.500 312.400 5.100 317.600 ;
        RECT 65.300 312.400 65.900 317.600 ;
        RECT 114.900 312.400 115.500 317.600 ;
        RECT 194.800 315.800 195.600 316.600 ;
        RECT 260.400 315.800 261.200 316.600 ;
        RECT 4.400 311.600 5.200 312.400 ;
        RECT 65.200 311.600 66.000 312.400 ;
        RECT 114.800 311.600 115.600 312.400 ;
        RECT 194.900 312.000 195.500 315.800 ;
        RECT 260.500 312.000 261.100 315.800 ;
        RECT 398.100 312.400 398.700 317.600 ;
        RECT 414.000 315.800 414.800 316.600 ;
        RECT 194.800 311.200 195.600 312.000 ;
        RECT 260.400 311.200 261.200 312.000 ;
        RECT 398.000 311.600 398.800 312.400 ;
        RECT 414.100 312.000 414.700 315.800 ;
        RECT 414.000 311.200 414.800 312.000 ;
        RECT 68.400 290.000 69.200 290.800 ;
        RECT 68.500 284.400 69.100 290.000 ;
        RECT 121.200 289.600 122.000 290.400 ;
        RECT 167.600 289.600 168.400 290.400 ;
        RECT 212.400 290.000 213.200 290.800 ;
        RECT 265.200 290.000 266.000 290.800 ;
        RECT 121.300 284.400 121.900 289.600 ;
        RECT 167.700 284.400 168.300 289.600 ;
        RECT 212.500 286.200 213.100 290.000 ;
        RECT 212.400 285.400 213.200 286.200 ;
        RECT 265.300 284.400 265.900 290.000 ;
        RECT 398.000 289.600 398.800 290.400 ;
        RECT 423.600 289.600 424.400 290.400 ;
        RECT 398.100 284.400 398.700 289.600 ;
        RECT 423.700 284.400 424.300 289.600 ;
        RECT 68.400 283.600 69.200 284.400 ;
        RECT 121.200 283.600 122.000 284.400 ;
        RECT 167.600 283.600 168.400 284.400 ;
        RECT 265.200 283.600 266.000 284.400 ;
        RECT 398.000 283.600 398.800 284.400 ;
        RECT 423.600 283.600 424.400 284.400 ;
        RECT 111.200 280.600 116.000 281.400 ;
        RECT 415.200 280.600 420.000 281.400 ;
        RECT 4.400 277.600 5.200 278.400 ;
        RECT 97.200 277.600 98.000 278.400 ;
        RECT 218.800 277.600 219.600 278.400 ;
        RECT 258.800 277.600 259.600 278.400 ;
        RECT 430.000 277.600 430.800 278.400 ;
        RECT 468.400 277.600 469.200 278.400 ;
        RECT 4.500 272.400 5.100 277.600 ;
        RECT 97.300 272.400 97.900 277.600 ;
        RECT 162.800 275.800 163.600 276.600 ;
        RECT 4.400 271.600 5.200 272.400 ;
        RECT 97.200 271.600 98.000 272.400 ;
        RECT 162.900 272.000 163.500 275.800 ;
        RECT 218.900 272.400 219.500 277.600 ;
        RECT 258.900 272.400 259.500 277.600 ;
        RECT 300.400 275.800 301.200 276.600 ;
        RECT 162.800 271.200 163.600 272.000 ;
        RECT 218.800 271.600 219.600 272.400 ;
        RECT 258.800 271.600 259.600 272.400 ;
        RECT 300.500 272.000 301.100 275.800 ;
        RECT 430.100 272.400 430.700 277.600 ;
        RECT 468.500 272.400 469.100 277.600 ;
        RECT 300.400 271.200 301.200 272.000 ;
        RECT 430.000 271.600 430.800 272.400 ;
        RECT 468.400 271.600 469.200 272.400 ;
        RECT 44.400 249.600 45.200 250.400 ;
        RECT 79.600 249.600 80.400 250.400 ;
        RECT 114.800 250.000 115.600 250.800 ;
        RECT 191.600 250.000 192.400 250.800 ;
        RECT 250.800 250.000 251.600 250.800 ;
        RECT 300.400 250.000 301.200 250.800 ;
        RECT 430.000 250.000 430.800 250.800 ;
        RECT 518.000 250.000 518.800 250.800 ;
        RECT 44.500 244.400 45.100 249.600 ;
        RECT 79.700 244.400 80.300 249.600 ;
        RECT 114.900 246.200 115.500 250.000 ;
        RECT 191.700 246.200 192.300 250.000 ;
        RECT 250.900 246.200 251.500 250.000 ;
        RECT 300.500 246.200 301.100 250.000 ;
        RECT 430.100 246.200 430.700 250.000 ;
        RECT 518.100 246.200 518.700 250.000 ;
        RECT 114.800 245.400 115.600 246.200 ;
        RECT 191.600 245.400 192.400 246.200 ;
        RECT 250.800 245.400 251.600 246.200 ;
        RECT 300.400 245.400 301.200 246.200 ;
        RECT 430.000 245.400 430.800 246.200 ;
        RECT 518.000 245.400 518.800 246.200 ;
        RECT 44.400 243.600 45.200 244.400 ;
        RECT 79.600 243.600 80.400 244.400 ;
        RECT 111.200 240.600 116.000 241.400 ;
        RECT 415.200 240.600 420.000 241.400 ;
        RECT 52.400 237.600 53.200 238.400 ;
        RECT 90.800 237.600 91.600 238.400 ;
        RECT 390.000 237.600 390.800 238.400 ;
        RECT 606.000 237.600 606.800 238.400 ;
        RECT 633.200 237.600 634.000 238.400 ;
        RECT 52.500 232.400 53.100 237.600 ;
        RECT 90.900 232.400 91.500 237.600 ;
        RECT 166.000 235.800 166.800 236.600 ;
        RECT 214.000 235.800 214.800 236.600 ;
        RECT 244.400 235.800 245.200 236.600 ;
        RECT 324.400 235.800 325.200 236.600 ;
        RECT 52.400 231.600 53.200 232.400 ;
        RECT 90.800 231.600 91.600 232.400 ;
        RECT 166.100 232.000 166.700 235.800 ;
        RECT 214.100 232.000 214.700 235.800 ;
        RECT 244.500 232.000 245.100 235.800 ;
        RECT 324.500 232.000 325.100 235.800 ;
        RECT 390.100 232.400 390.700 237.600 ;
        RECT 460.400 235.800 461.200 236.600 ;
        RECT 508.400 235.800 509.200 236.600 ;
        RECT 166.000 231.200 166.800 232.000 ;
        RECT 214.000 231.200 214.800 232.000 ;
        RECT 244.400 231.200 245.200 232.000 ;
        RECT 324.400 231.200 325.200 232.000 ;
        RECT 390.000 231.600 390.800 232.400 ;
        RECT 460.500 232.000 461.100 235.800 ;
        RECT 508.500 232.000 509.100 235.800 ;
        RECT 606.100 232.400 606.700 237.600 ;
        RECT 633.300 232.400 633.900 237.600 ;
        RECT 460.400 231.200 461.200 232.000 ;
        RECT 508.400 231.200 509.200 232.000 ;
        RECT 606.000 231.600 606.800 232.400 ;
        RECT 633.200 231.600 634.000 232.400 ;
        RECT 470.000 211.600 470.800 212.400 ;
        RECT 14.000 209.600 14.800 210.400 ;
        RECT 90.800 209.600 91.600 210.400 ;
        RECT 145.200 210.000 146.000 210.800 ;
        RECT 14.100 204.400 14.700 209.600 ;
        RECT 90.900 204.400 91.500 209.600 ;
        RECT 145.300 206.200 145.900 210.000 ;
        RECT 183.600 209.600 184.400 210.400 ;
        RECT 191.600 209.600 192.400 210.400 ;
        RECT 268.400 209.600 269.200 210.400 ;
        RECT 382.000 210.000 382.800 210.800 ;
        RECT 414.000 210.000 414.800 210.800 ;
        RECT 145.200 205.400 146.000 206.200 ;
        RECT 183.700 204.400 184.300 209.600 ;
        RECT 191.700 204.400 192.300 209.600 ;
        RECT 268.500 204.400 269.100 209.600 ;
        RECT 382.100 206.200 382.700 210.000 ;
        RECT 414.100 206.200 414.700 210.000 ;
        RECT 470.100 206.400 470.700 211.600 ;
        RECT 494.000 210.000 494.800 210.800 ;
        RECT 382.000 205.400 382.800 206.200 ;
        RECT 414.000 205.400 414.800 206.200 ;
        RECT 470.000 205.600 470.800 206.400 ;
        RECT 494.100 206.200 494.700 210.000 ;
        RECT 641.200 209.600 642.000 210.400 ;
        RECT 494.000 205.400 494.800 206.200 ;
        RECT 641.300 204.400 641.900 209.600 ;
        RECT 14.000 203.600 14.800 204.400 ;
        RECT 90.800 203.600 91.600 204.400 ;
        RECT 183.600 203.600 184.400 204.400 ;
        RECT 191.600 203.600 192.400 204.400 ;
        RECT 268.400 203.600 269.200 204.400 ;
        RECT 641.200 203.600 642.000 204.400 ;
        RECT 111.200 200.600 116.000 201.400 ;
        RECT 415.200 200.600 420.000 201.400 ;
        RECT 20.400 197.600 21.200 198.400 ;
        RECT 212.400 197.600 213.200 198.400 ;
        RECT 258.800 197.600 259.600 198.400 ;
        RECT 298.800 197.600 299.600 198.400 ;
        RECT 310.000 197.600 310.800 198.400 ;
        RECT 20.500 192.400 21.100 197.600 ;
        RECT 212.500 192.400 213.100 197.600 ;
        RECT 258.900 192.400 259.500 197.600 ;
        RECT 298.900 192.400 299.500 197.600 ;
        RECT 310.100 192.400 310.700 197.600 ;
        RECT 454.000 195.800 454.800 196.600 ;
        RECT 20.400 191.600 21.200 192.400 ;
        RECT 212.400 191.600 213.200 192.400 ;
        RECT 258.800 191.600 259.600 192.400 ;
        RECT 298.800 191.600 299.600 192.400 ;
        RECT 310.000 191.600 310.800 192.400 ;
        RECT 454.100 192.000 454.700 195.800 ;
        RECT 454.000 191.200 454.800 192.000 ;
        RECT 4.400 169.600 5.200 170.400 ;
        RECT 79.600 169.600 80.400 170.400 ;
        RECT 250.800 169.600 251.600 170.400 ;
        RECT 278.000 170.000 278.800 170.800 ;
        RECT 4.500 164.400 5.100 169.600 ;
        RECT 79.700 164.400 80.300 169.600 ;
        RECT 250.900 164.400 251.500 169.600 ;
        RECT 278.100 166.200 278.700 170.000 ;
        RECT 327.600 169.600 328.400 170.400 ;
        RECT 386.800 170.000 387.600 170.800 ;
        RECT 442.800 170.000 443.600 170.800 ;
        RECT 278.000 165.400 278.800 166.200 ;
        RECT 327.700 164.400 328.300 169.600 ;
        RECT 386.900 164.400 387.500 170.000 ;
        RECT 442.900 164.400 443.500 170.000 ;
        RECT 508.400 169.600 509.200 170.400 ;
        RECT 681.200 170.000 682.000 170.800 ;
        RECT 508.500 164.400 509.100 169.600 ;
        RECT 681.300 166.200 681.900 170.000 ;
        RECT 681.200 165.400 682.000 166.200 ;
        RECT 4.400 163.600 5.200 164.400 ;
        RECT 79.600 163.600 80.400 164.400 ;
        RECT 250.800 163.600 251.600 164.400 ;
        RECT 327.600 163.600 328.400 164.400 ;
        RECT 386.800 163.600 387.600 164.400 ;
        RECT 442.800 163.600 443.600 164.400 ;
        RECT 508.400 163.600 509.200 164.400 ;
        RECT 111.200 160.600 116.000 161.400 ;
        RECT 415.200 160.600 420.000 161.400 ;
        RECT 316.400 157.600 317.200 158.400 ;
        RECT 378.800 157.600 379.600 158.400 ;
        RECT 479.600 157.600 480.400 158.400 ;
        RECT 295.600 155.800 296.400 156.600 ;
        RECT 295.700 150.400 296.300 155.800 ;
        RECT 316.500 152.400 317.100 157.600 ;
        RECT 378.900 152.400 379.500 157.600 ;
        RECT 390.000 155.800 390.800 156.600 ;
        RECT 444.400 155.800 445.200 156.600 ;
        RECT 316.400 151.600 317.200 152.400 ;
        RECT 378.800 151.600 379.600 152.400 ;
        RECT 390.100 152.000 390.700 155.800 ;
        RECT 444.500 152.000 445.100 155.800 ;
        RECT 479.700 152.400 480.300 157.600 ;
        RECT 390.000 151.200 390.800 152.000 ;
        RECT 444.400 151.200 445.200 152.000 ;
        RECT 479.600 151.600 480.400 152.400 ;
        RECT 295.600 149.600 296.400 150.400 ;
        RECT 228.400 130.000 229.200 130.800 ;
        RECT 334.000 130.000 334.800 130.800 ;
        RECT 358.000 130.000 358.800 130.800 ;
        RECT 420.400 130.000 421.200 130.800 ;
        RECT 447.600 130.000 448.400 130.800 ;
        RECT 228.500 124.400 229.100 130.000 ;
        RECT 334.100 126.200 334.700 130.000 ;
        RECT 358.100 126.200 358.700 130.000 ;
        RECT 420.500 126.200 421.100 130.000 ;
        RECT 334.000 125.400 334.800 126.200 ;
        RECT 358.000 125.400 358.800 126.200 ;
        RECT 420.400 125.400 421.200 126.200 ;
        RECT 447.700 124.400 448.300 130.000 ;
        RECT 479.600 129.600 480.400 130.400 ;
        RECT 479.700 124.400 480.300 129.600 ;
        RECT 228.400 123.600 229.200 124.400 ;
        RECT 447.600 123.600 448.400 124.400 ;
        RECT 479.600 123.600 480.400 124.400 ;
        RECT 111.200 120.600 116.000 121.400 ;
        RECT 415.200 120.600 420.000 121.400 ;
        RECT 358.000 117.600 358.800 118.400 ;
        RECT 454.000 117.600 454.800 118.400 ;
        RECT 294.000 115.800 294.800 116.600 ;
        RECT 294.100 112.000 294.700 115.800 ;
        RECT 358.100 112.400 358.700 117.600 ;
        RECT 390.000 115.800 390.800 116.600 ;
        RECT 294.000 111.200 294.800 112.000 ;
        RECT 358.000 111.600 358.800 112.400 ;
        RECT 390.100 112.000 390.700 115.800 ;
        RECT 454.100 112.400 454.700 117.600 ;
        RECT 508.400 115.800 509.200 116.600 ;
        RECT 390.000 111.200 390.800 112.000 ;
        RECT 454.000 111.600 454.800 112.400 ;
        RECT 508.500 112.000 509.100 115.800 ;
        RECT 508.400 111.200 509.200 112.000 ;
        RECT 202.800 90.000 203.600 90.800 ;
        RECT 202.900 86.200 203.500 90.000 ;
        RECT 284.400 89.600 285.200 90.400 ;
        RECT 334.000 90.000 334.800 90.800 ;
        RECT 351.600 90.000 352.400 90.800 ;
        RECT 434.800 90.000 435.600 90.800 ;
        RECT 494.000 90.000 494.800 90.800 ;
        RECT 202.800 85.400 203.600 86.200 ;
        RECT 284.500 84.400 285.100 89.600 ;
        RECT 334.100 86.200 334.700 90.000 ;
        RECT 334.000 85.400 334.800 86.200 ;
        RECT 351.700 84.400 352.300 90.000 ;
        RECT 434.900 84.400 435.500 90.000 ;
        RECT 494.100 86.200 494.700 90.000 ;
        RECT 494.000 85.400 494.800 86.200 ;
        RECT 284.400 83.600 285.200 84.400 ;
        RECT 351.600 83.600 352.400 84.400 ;
        RECT 434.800 83.600 435.600 84.400 ;
        RECT 111.200 80.600 116.000 81.400 ;
        RECT 415.200 80.600 420.000 81.400 ;
        RECT 239.600 77.600 240.400 78.400 ;
        RECT 340.400 77.600 341.200 78.400 ;
        RECT 468.400 77.600 469.200 78.400 ;
        RECT 239.700 72.400 240.300 77.600 ;
        RECT 308.400 75.800 309.200 76.600 ;
        RECT 239.600 71.600 240.400 72.400 ;
        RECT 308.500 72.000 309.100 75.800 ;
        RECT 340.500 72.400 341.100 77.600 ;
        RECT 438.000 75.800 438.800 76.600 ;
        RECT 308.400 71.200 309.200 72.000 ;
        RECT 340.400 71.600 341.200 72.400 ;
        RECT 438.100 72.000 438.700 75.800 ;
        RECT 468.500 72.400 469.100 77.600 ;
        RECT 438.000 71.200 438.800 72.000 ;
        RECT 468.400 71.600 469.200 72.400 ;
        RECT 202.800 50.000 203.600 50.800 ;
        RECT 223.600 50.000 224.400 50.800 ;
        RECT 270.000 50.000 270.800 50.800 ;
        RECT 342.000 50.000 342.800 50.800 ;
        RECT 202.900 46.200 203.500 50.000 ;
        RECT 223.700 46.200 224.300 50.000 ;
        RECT 270.100 46.200 270.700 50.000 ;
        RECT 342.100 46.200 342.700 50.000 ;
        RECT 388.400 49.600 389.200 50.400 ;
        RECT 425.200 50.000 426.000 50.800 ;
        RECT 465.200 50.000 466.000 50.800 ;
        RECT 202.800 45.400 203.600 46.200 ;
        RECT 223.600 45.400 224.400 46.200 ;
        RECT 270.000 45.400 270.800 46.200 ;
        RECT 342.000 45.400 342.800 46.200 ;
        RECT 388.500 44.400 389.100 49.600 ;
        RECT 425.300 44.400 425.900 50.000 ;
        RECT 465.300 44.400 465.900 50.000 ;
        RECT 388.400 43.600 389.200 44.400 ;
        RECT 425.200 43.600 426.000 44.400 ;
        RECT 465.200 43.600 466.000 44.400 ;
        RECT 111.200 40.600 116.000 41.400 ;
        RECT 415.200 40.600 420.000 41.400 ;
        RECT 4.400 37.600 5.200 38.400 ;
        RECT 228.400 37.600 229.200 38.400 ;
        RECT 375.600 37.600 376.400 38.400 ;
        RECT 526.000 37.600 526.800 38.400 ;
        RECT 4.500 32.400 5.100 37.600 ;
        RECT 228.500 32.400 229.100 37.600 ;
        RECT 239.600 35.800 240.400 36.600 ;
        RECT 340.400 35.800 341.200 36.600 ;
        RECT 4.400 31.600 5.200 32.400 ;
        RECT 228.400 31.600 229.200 32.400 ;
        RECT 239.700 32.000 240.300 35.800 ;
        RECT 340.500 32.000 341.100 35.800 ;
        RECT 375.700 32.400 376.300 37.600 ;
        RECT 438.000 35.800 438.800 36.600 ;
        RECT 239.600 31.200 240.400 32.000 ;
        RECT 340.400 31.200 341.200 32.000 ;
        RECT 375.600 31.600 376.400 32.400 ;
        RECT 438.100 32.000 438.700 35.800 ;
        RECT 526.100 32.400 526.700 37.600 ;
        RECT 438.000 31.200 438.800 32.000 ;
        RECT 526.000 31.600 526.800 32.400 ;
        RECT 10.800 10.000 11.600 10.800 ;
        RECT 10.900 4.400 11.500 10.000 ;
        RECT 78.000 9.600 78.800 10.400 ;
        RECT 113.200 9.600 114.000 10.400 ;
        RECT 196.400 9.600 197.200 10.400 ;
        RECT 207.600 10.000 208.400 10.800 ;
        RECT 310.000 10.000 310.800 10.800 ;
        RECT 78.100 4.400 78.700 9.600 ;
        RECT 113.300 4.400 113.900 9.600 ;
        RECT 196.500 4.400 197.100 9.600 ;
        RECT 207.700 6.200 208.300 10.000 ;
        RECT 310.100 6.200 310.700 10.000 ;
        RECT 366.000 9.600 366.800 10.400 ;
        RECT 383.600 9.600 384.400 10.400 ;
        RECT 428.400 9.600 429.200 10.400 ;
        RECT 494.000 10.000 494.800 10.800 ;
        RECT 207.600 5.400 208.400 6.200 ;
        RECT 310.000 5.400 310.800 6.200 ;
        RECT 366.100 4.400 366.700 9.600 ;
        RECT 383.700 4.400 384.300 9.600 ;
        RECT 428.500 4.400 429.100 9.600 ;
        RECT 494.100 6.200 494.700 10.000 ;
        RECT 508.400 9.600 509.200 10.400 ;
        RECT 550.000 10.000 550.800 10.800 ;
        RECT 494.000 5.400 494.800 6.200 ;
        RECT 508.500 4.400 509.100 9.600 ;
        RECT 550.100 6.200 550.700 10.000 ;
        RECT 550.000 5.400 550.800 6.200 ;
        RECT 10.800 3.600 11.600 4.400 ;
        RECT 78.000 3.600 78.800 4.400 ;
        RECT 113.200 3.600 114.000 4.400 ;
        RECT 196.400 3.600 197.200 4.400 ;
        RECT 366.000 3.600 366.800 4.400 ;
        RECT 383.600 3.600 384.400 4.400 ;
        RECT 428.400 3.600 429.200 4.400 ;
        RECT 508.400 3.600 509.200 4.400 ;
        RECT 111.200 0.600 116.000 1.400 ;
        RECT 415.200 0.600 420.000 1.400 ;
      LAYER via2 ;
        RECT 111.800 480.600 112.600 481.400 ;
        RECT 113.200 480.600 114.000 481.400 ;
        RECT 114.600 480.600 115.400 481.400 ;
        RECT 415.800 480.600 416.600 481.400 ;
        RECT 417.200 480.600 418.000 481.400 ;
        RECT 418.600 480.600 419.400 481.400 ;
        RECT 111.800 440.600 112.600 441.400 ;
        RECT 113.200 440.600 114.000 441.400 ;
        RECT 114.600 440.600 115.400 441.400 ;
        RECT 415.800 440.600 416.600 441.400 ;
        RECT 417.200 440.600 418.000 441.400 ;
        RECT 418.600 440.600 419.400 441.400 ;
        RECT 111.800 400.600 112.600 401.400 ;
        RECT 113.200 400.600 114.000 401.400 ;
        RECT 114.600 400.600 115.400 401.400 ;
        RECT 415.800 400.600 416.600 401.400 ;
        RECT 417.200 400.600 418.000 401.400 ;
        RECT 418.600 400.600 419.400 401.400 ;
        RECT 111.800 360.600 112.600 361.400 ;
        RECT 113.200 360.600 114.000 361.400 ;
        RECT 114.600 360.600 115.400 361.400 ;
        RECT 415.800 360.600 416.600 361.400 ;
        RECT 417.200 360.600 418.000 361.400 ;
        RECT 418.600 360.600 419.400 361.400 ;
        RECT 111.800 320.600 112.600 321.400 ;
        RECT 113.200 320.600 114.000 321.400 ;
        RECT 114.600 320.600 115.400 321.400 ;
        RECT 415.800 320.600 416.600 321.400 ;
        RECT 417.200 320.600 418.000 321.400 ;
        RECT 418.600 320.600 419.400 321.400 ;
        RECT 111.800 280.600 112.600 281.400 ;
        RECT 113.200 280.600 114.000 281.400 ;
        RECT 114.600 280.600 115.400 281.400 ;
        RECT 415.800 280.600 416.600 281.400 ;
        RECT 417.200 280.600 418.000 281.400 ;
        RECT 418.600 280.600 419.400 281.400 ;
        RECT 111.800 240.600 112.600 241.400 ;
        RECT 113.200 240.600 114.000 241.400 ;
        RECT 114.600 240.600 115.400 241.400 ;
        RECT 415.800 240.600 416.600 241.400 ;
        RECT 417.200 240.600 418.000 241.400 ;
        RECT 418.600 240.600 419.400 241.400 ;
        RECT 111.800 200.600 112.600 201.400 ;
        RECT 113.200 200.600 114.000 201.400 ;
        RECT 114.600 200.600 115.400 201.400 ;
        RECT 415.800 200.600 416.600 201.400 ;
        RECT 417.200 200.600 418.000 201.400 ;
        RECT 418.600 200.600 419.400 201.400 ;
        RECT 111.800 160.600 112.600 161.400 ;
        RECT 113.200 160.600 114.000 161.400 ;
        RECT 114.600 160.600 115.400 161.400 ;
        RECT 415.800 160.600 416.600 161.400 ;
        RECT 417.200 160.600 418.000 161.400 ;
        RECT 418.600 160.600 419.400 161.400 ;
        RECT 111.800 120.600 112.600 121.400 ;
        RECT 113.200 120.600 114.000 121.400 ;
        RECT 114.600 120.600 115.400 121.400 ;
        RECT 415.800 120.600 416.600 121.400 ;
        RECT 417.200 120.600 418.000 121.400 ;
        RECT 418.600 120.600 419.400 121.400 ;
        RECT 111.800 80.600 112.600 81.400 ;
        RECT 113.200 80.600 114.000 81.400 ;
        RECT 114.600 80.600 115.400 81.400 ;
        RECT 415.800 80.600 416.600 81.400 ;
        RECT 417.200 80.600 418.000 81.400 ;
        RECT 418.600 80.600 419.400 81.400 ;
        RECT 111.800 40.600 112.600 41.400 ;
        RECT 113.200 40.600 114.000 41.400 ;
        RECT 114.600 40.600 115.400 41.400 ;
        RECT 415.800 40.600 416.600 41.400 ;
        RECT 417.200 40.600 418.000 41.400 ;
        RECT 418.600 40.600 419.400 41.400 ;
        RECT 111.800 0.600 112.600 1.400 ;
        RECT 113.200 0.600 114.000 1.400 ;
        RECT 114.600 0.600 115.400 1.400 ;
        RECT 415.800 0.600 416.600 1.400 ;
        RECT 417.200 0.600 418.000 1.400 ;
        RECT 418.600 0.600 419.400 1.400 ;
      LAYER metal3 ;
        RECT 111.200 480.400 116.000 481.600 ;
        RECT 415.200 480.400 420.000 481.600 ;
        RECT 111.200 440.400 116.000 441.600 ;
        RECT 415.200 440.400 420.000 441.600 ;
        RECT 111.200 400.400 116.000 401.600 ;
        RECT 415.200 400.400 420.000 401.600 ;
        RECT 111.200 360.400 116.000 361.600 ;
        RECT 415.200 360.400 420.000 361.600 ;
        RECT 111.200 320.400 116.000 321.600 ;
        RECT 415.200 320.400 420.000 321.600 ;
        RECT 111.200 280.400 116.000 281.600 ;
        RECT 415.200 280.400 420.000 281.600 ;
        RECT 111.200 240.400 116.000 241.600 ;
        RECT 415.200 240.400 420.000 241.600 ;
        RECT 111.200 200.400 116.000 201.600 ;
        RECT 415.200 200.400 420.000 201.600 ;
        RECT 111.200 160.400 116.000 161.600 ;
        RECT 415.200 160.400 420.000 161.600 ;
        RECT 111.200 120.400 116.000 121.600 ;
        RECT 415.200 120.400 420.000 121.600 ;
        RECT 111.200 80.400 116.000 81.600 ;
        RECT 415.200 80.400 420.000 81.600 ;
        RECT 111.200 40.400 116.000 41.600 ;
        RECT 415.200 40.400 420.000 41.600 ;
        RECT 111.200 0.400 116.000 1.600 ;
        RECT 415.200 0.400 420.000 1.600 ;
      LAYER via3 ;
        RECT 111.600 480.600 112.400 481.400 ;
        RECT 113.200 480.600 114.000 481.400 ;
        RECT 114.800 480.600 115.600 481.400 ;
        RECT 415.600 480.600 416.400 481.400 ;
        RECT 417.200 480.600 418.000 481.400 ;
        RECT 418.800 480.600 419.600 481.400 ;
        RECT 111.600 440.600 112.400 441.400 ;
        RECT 113.200 440.600 114.000 441.400 ;
        RECT 114.800 440.600 115.600 441.400 ;
        RECT 415.600 440.600 416.400 441.400 ;
        RECT 417.200 440.600 418.000 441.400 ;
        RECT 418.800 440.600 419.600 441.400 ;
        RECT 111.600 400.600 112.400 401.400 ;
        RECT 113.200 400.600 114.000 401.400 ;
        RECT 114.800 400.600 115.600 401.400 ;
        RECT 415.600 400.600 416.400 401.400 ;
        RECT 417.200 400.600 418.000 401.400 ;
        RECT 418.800 400.600 419.600 401.400 ;
        RECT 111.600 360.600 112.400 361.400 ;
        RECT 113.200 360.600 114.000 361.400 ;
        RECT 114.800 360.600 115.600 361.400 ;
        RECT 415.600 360.600 416.400 361.400 ;
        RECT 417.200 360.600 418.000 361.400 ;
        RECT 418.800 360.600 419.600 361.400 ;
        RECT 111.600 320.600 112.400 321.400 ;
        RECT 113.200 320.600 114.000 321.400 ;
        RECT 114.800 320.600 115.600 321.400 ;
        RECT 415.600 320.600 416.400 321.400 ;
        RECT 417.200 320.600 418.000 321.400 ;
        RECT 418.800 320.600 419.600 321.400 ;
        RECT 111.600 280.600 112.400 281.400 ;
        RECT 113.200 280.600 114.000 281.400 ;
        RECT 114.800 280.600 115.600 281.400 ;
        RECT 415.600 280.600 416.400 281.400 ;
        RECT 417.200 280.600 418.000 281.400 ;
        RECT 418.800 280.600 419.600 281.400 ;
        RECT 111.600 240.600 112.400 241.400 ;
        RECT 113.200 240.600 114.000 241.400 ;
        RECT 114.800 240.600 115.600 241.400 ;
        RECT 415.600 240.600 416.400 241.400 ;
        RECT 417.200 240.600 418.000 241.400 ;
        RECT 418.800 240.600 419.600 241.400 ;
        RECT 111.600 200.600 112.400 201.400 ;
        RECT 113.200 200.600 114.000 201.400 ;
        RECT 114.800 200.600 115.600 201.400 ;
        RECT 415.600 200.600 416.400 201.400 ;
        RECT 417.200 200.600 418.000 201.400 ;
        RECT 418.800 200.600 419.600 201.400 ;
        RECT 111.600 160.600 112.400 161.400 ;
        RECT 113.200 160.600 114.000 161.400 ;
        RECT 114.800 160.600 115.600 161.400 ;
        RECT 415.600 160.600 416.400 161.400 ;
        RECT 417.200 160.600 418.000 161.400 ;
        RECT 418.800 160.600 419.600 161.400 ;
        RECT 111.600 120.600 112.400 121.400 ;
        RECT 113.200 120.600 114.000 121.400 ;
        RECT 114.800 120.600 115.600 121.400 ;
        RECT 415.600 120.600 416.400 121.400 ;
        RECT 417.200 120.600 418.000 121.400 ;
        RECT 418.800 120.600 419.600 121.400 ;
        RECT 111.600 80.600 112.400 81.400 ;
        RECT 113.200 80.600 114.000 81.400 ;
        RECT 114.800 80.600 115.600 81.400 ;
        RECT 415.600 80.600 416.400 81.400 ;
        RECT 417.200 80.600 418.000 81.400 ;
        RECT 418.800 80.600 419.600 81.400 ;
        RECT 111.600 40.600 112.400 41.400 ;
        RECT 113.200 40.600 114.000 41.400 ;
        RECT 114.800 40.600 115.600 41.400 ;
        RECT 415.600 40.600 416.400 41.400 ;
        RECT 417.200 40.600 418.000 41.400 ;
        RECT 418.800 40.600 419.600 41.400 ;
        RECT 111.600 0.600 112.400 1.400 ;
        RECT 113.200 0.600 114.000 1.400 ;
        RECT 114.800 0.600 115.600 1.400 ;
        RECT 415.600 0.600 416.400 1.400 ;
        RECT 417.200 0.600 418.000 1.400 ;
        RECT 418.800 0.600 419.600 1.400 ;
      LAYER metal4 ;
        RECT 111.200 -4.000 116.000 504.000 ;
        RECT 415.200 -4.000 420.000 504.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 500.400 689.200 501.600 ;
        RECT 4.400 495.800 5.200 500.400 ;
        RECT 14.000 497.800 14.800 500.400 ;
        RECT 17.200 497.800 18.000 500.400 ;
        RECT 28.400 495.800 29.200 500.400 ;
        RECT 34.800 497.800 35.600 500.400 ;
        RECT 39.600 496.600 40.400 500.400 ;
        RECT 44.400 497.800 45.200 500.400 ;
        RECT 49.200 495.800 50.000 500.400 ;
        RECT 58.800 497.800 59.600 500.400 ;
        RECT 62.000 497.800 62.800 500.400 ;
        RECT 73.200 495.800 74.000 500.400 ;
        RECT 79.600 497.800 80.400 500.400 ;
        RECT 81.200 497.800 82.000 500.400 ;
        RECT 86.000 496.600 86.800 500.400 ;
        RECT 94.000 496.600 94.800 500.400 ;
        RECT 97.200 495.800 98.000 500.400 ;
        RECT 100.400 495.800 101.200 500.400 ;
        RECT 103.600 495.800 104.400 500.400 ;
        RECT 106.800 495.800 107.600 500.400 ;
        RECT 110.000 495.800 110.800 500.400 ;
        RECT 118.000 495.800 118.800 500.400 ;
        RECT 123.400 497.800 124.400 500.400 ;
        RECT 126.800 497.800 127.600 500.400 ;
        RECT 132.400 496.000 133.200 500.400 ;
        RECT 135.600 495.800 136.400 500.400 ;
        RECT 138.800 495.800 139.600 500.400 ;
        RECT 142.000 495.800 142.800 500.400 ;
        RECT 145.200 495.800 146.000 500.400 ;
        RECT 148.400 495.800 149.200 500.400 ;
        RECT 151.600 496.600 152.400 500.400 ;
        RECT 156.400 497.800 157.200 500.400 ;
        RECT 161.200 496.600 162.000 500.400 ;
        RECT 166.000 497.800 166.800 500.400 ;
        RECT 172.400 495.800 173.200 500.400 ;
        RECT 183.600 497.800 184.400 500.400 ;
        RECT 186.800 497.800 187.600 500.400 ;
        RECT 196.400 495.800 197.200 500.400 ;
        RECT 201.200 497.800 202.000 500.400 ;
        RECT 204.400 497.800 205.200 500.400 ;
        RECT 210.800 495.800 211.600 500.400 ;
        RECT 222.000 497.800 222.800 500.400 ;
        RECT 225.200 497.800 226.000 500.400 ;
        RECT 234.800 495.800 235.600 500.400 ;
        RECT 239.600 495.800 240.400 500.400 ;
        RECT 242.800 495.800 243.600 500.400 ;
        RECT 246.000 495.800 246.800 500.400 ;
        RECT 249.200 495.800 250.000 500.400 ;
        RECT 252.400 495.800 253.200 500.400 ;
        RECT 262.000 495.800 262.800 500.400 ;
        RECT 271.600 497.800 272.400 500.400 ;
        RECT 274.800 497.800 275.600 500.400 ;
        RECT 286.000 495.800 286.800 500.400 ;
        RECT 292.400 497.800 293.200 500.400 ;
        RECT 295.600 495.800 296.400 500.400 ;
        RECT 302.000 495.800 302.800 500.400 ;
        RECT 311.600 497.800 312.400 500.400 ;
        RECT 314.800 497.800 315.600 500.400 ;
        RECT 326.000 495.800 326.800 500.400 ;
        RECT 332.400 497.800 333.200 500.400 ;
        RECT 335.800 499.800 336.600 500.400 ;
        RECT 335.600 496.400 336.600 499.800 ;
        RECT 341.800 496.400 342.800 500.400 ;
        RECT 345.200 497.800 346.000 500.400 ;
        RECT 351.600 495.800 352.400 500.400 ;
        RECT 362.800 497.800 363.600 500.400 ;
        RECT 366.000 497.800 366.800 500.400 ;
        RECT 375.600 495.800 376.400 500.400 ;
        RECT 382.000 495.800 382.800 500.400 ;
        RECT 385.200 497.800 386.000 500.400 ;
        RECT 391.600 495.800 392.400 500.400 ;
        RECT 402.800 497.800 403.600 500.400 ;
        RECT 406.000 497.800 406.800 500.400 ;
        RECT 415.600 495.800 416.400 500.400 ;
        RECT 426.800 495.800 427.600 500.400 ;
        RECT 430.000 497.800 430.800 500.400 ;
        RECT 434.800 496.600 435.600 500.400 ;
        RECT 439.600 495.800 440.400 500.400 ;
        RECT 444.400 497.800 445.200 500.400 ;
        RECT 450.800 495.800 451.600 500.400 ;
        RECT 462.000 497.800 462.800 500.400 ;
        RECT 465.200 497.800 466.000 500.400 ;
        RECT 474.800 495.800 475.600 500.400 ;
        RECT 479.600 497.800 480.400 500.400 ;
        RECT 484.400 497.800 485.200 500.400 ;
        RECT 487.600 495.800 488.400 500.400 ;
        RECT 490.800 497.800 491.600 500.400 ;
        RECT 497.200 495.800 498.000 500.400 ;
        RECT 508.400 497.800 509.200 500.400 ;
        RECT 511.600 497.800 512.400 500.400 ;
        RECT 521.200 495.800 522.000 500.400 ;
        RECT 526.000 497.800 526.800 500.400 ;
        RECT 530.800 496.600 531.600 500.400 ;
        RECT 538.800 495.800 539.600 500.400 ;
        RECT 543.600 496.600 544.400 500.400 ;
        RECT 548.400 497.800 549.200 500.400 ;
        RECT 550.000 497.800 550.800 500.400 ;
        RECT 556.400 495.800 557.200 500.400 ;
        RECT 567.600 497.800 568.400 500.400 ;
        RECT 570.800 497.800 571.600 500.400 ;
        RECT 580.400 495.800 581.200 500.400 ;
        RECT 593.200 495.800 594.000 500.400 ;
        RECT 602.800 497.800 603.600 500.400 ;
        RECT 606.000 497.800 606.800 500.400 ;
        RECT 617.200 495.800 618.000 500.400 ;
        RECT 623.600 497.800 624.400 500.400 ;
        RECT 627.000 499.800 627.800 500.400 ;
        RECT 626.800 496.400 627.800 499.800 ;
        RECT 633.000 496.400 634.000 500.400 ;
        RECT 636.400 495.800 637.200 500.400 ;
        RECT 639.600 495.800 640.400 500.400 ;
        RECT 642.800 495.800 643.600 500.400 ;
        RECT 646.000 495.800 646.800 500.400 ;
        RECT 649.200 495.800 650.000 500.400 ;
        RECT 650.800 497.800 651.600 500.400 ;
        RECT 657.200 495.800 658.000 500.400 ;
        RECT 668.400 497.800 669.200 500.400 ;
        RECT 671.600 497.800 672.400 500.400 ;
        RECT 681.200 495.800 682.000 500.400 ;
        RECT 1.200 461.600 2.000 464.200 ;
        RECT 7.600 461.600 8.400 466.200 ;
        RECT 18.800 461.600 19.600 464.200 ;
        RECT 22.000 461.600 22.800 464.200 ;
        RECT 31.600 461.600 32.400 466.200 ;
        RECT 39.600 461.600 40.400 465.400 ;
        RECT 46.000 461.600 46.800 466.200 ;
        RECT 49.200 461.600 50.000 466.200 ;
        RECT 54.600 461.600 55.600 464.200 ;
        RECT 58.000 461.600 58.800 464.200 ;
        RECT 63.600 461.600 64.400 466.000 ;
        RECT 68.000 461.600 68.800 467.000 ;
        RECT 73.200 461.600 74.000 466.600 ;
        RECT 78.000 461.600 78.800 465.400 ;
        RECT 86.000 461.600 86.800 465.400 ;
        RECT 92.400 461.600 93.200 466.200 ;
        RECT 95.600 461.600 96.400 466.200 ;
        RECT 101.000 461.600 102.000 464.200 ;
        RECT 104.400 461.600 105.200 464.200 ;
        RECT 110.000 461.600 110.800 466.000 ;
        RECT 119.600 461.600 120.400 465.400 ;
        RECT 127.600 461.600 128.400 465.400 ;
        RECT 132.400 461.600 133.200 466.600 ;
        RECT 137.600 461.600 138.400 467.000 ;
        RECT 142.000 461.600 142.800 466.000 ;
        RECT 147.600 461.600 148.400 464.200 ;
        RECT 150.800 461.600 151.800 464.200 ;
        RECT 156.400 461.600 157.200 466.200 ;
        RECT 159.600 461.600 160.400 466.200 ;
        RECT 164.400 461.600 165.200 466.200 ;
        RECT 169.200 461.600 170.000 464.200 ;
        RECT 172.400 461.600 173.200 464.200 ;
        RECT 174.000 461.600 174.800 464.200 ;
        RECT 177.200 461.600 178.000 464.200 ;
        RECT 180.400 461.600 181.200 464.200 ;
        RECT 183.600 461.600 184.400 464.200 ;
        RECT 185.200 461.600 186.000 464.200 ;
        RECT 191.600 461.600 192.400 466.200 ;
        RECT 202.800 461.600 203.600 464.200 ;
        RECT 206.000 461.600 206.800 464.200 ;
        RECT 215.600 461.600 216.400 466.200 ;
        RECT 222.000 462.200 223.000 465.600 ;
        RECT 222.200 461.600 223.000 462.200 ;
        RECT 228.200 461.600 229.200 465.600 ;
        RECT 231.600 461.600 232.400 464.200 ;
        RECT 238.000 461.600 238.800 466.200 ;
        RECT 249.200 461.600 250.000 464.200 ;
        RECT 252.400 461.600 253.200 464.200 ;
        RECT 262.000 461.600 262.800 466.200 ;
        RECT 273.200 461.600 274.000 465.400 ;
        RECT 279.600 461.600 280.400 464.200 ;
        RECT 281.200 461.600 282.000 466.200 ;
        RECT 284.400 461.600 285.200 466.200 ;
        RECT 287.600 461.600 288.400 466.200 ;
        RECT 290.800 461.600 291.600 466.200 ;
        RECT 294.000 461.600 294.800 466.200 ;
        RECT 295.600 461.600 296.400 464.200 ;
        RECT 298.800 461.600 299.600 464.200 ;
        RECT 303.600 461.600 304.400 465.400 ;
        RECT 306.800 461.600 307.600 464.200 ;
        RECT 310.000 461.600 310.800 464.200 ;
        RECT 311.600 461.600 312.400 464.200 ;
        RECT 314.800 461.600 315.600 464.200 ;
        RECT 319.600 461.600 320.400 466.200 ;
        RECT 321.200 461.600 322.000 464.200 ;
        RECT 325.400 461.600 326.200 466.200 ;
        RECT 327.600 461.600 328.400 466.200 ;
        RECT 332.400 461.600 333.200 466.200 ;
        RECT 338.800 461.600 339.600 465.400 ;
        RECT 343.600 461.600 344.400 466.200 ;
        RECT 348.400 461.600 349.200 466.200 ;
        RECT 351.600 461.600 352.400 466.200 ;
        RECT 356.400 461.600 357.200 466.200 ;
        RECT 359.600 461.600 360.400 466.200 ;
        RECT 361.200 461.600 362.000 466.200 ;
        RECT 369.200 461.600 370.000 465.400 ;
        RECT 372.400 461.600 373.200 466.200 ;
        RECT 380.400 461.600 381.200 466.200 ;
        RECT 390.000 461.600 390.800 464.200 ;
        RECT 393.200 461.600 394.000 464.200 ;
        RECT 404.400 461.600 405.200 466.200 ;
        RECT 410.800 461.600 411.600 464.200 ;
        RECT 412.400 461.600 413.200 464.200 ;
        RECT 423.600 461.600 424.400 465.400 ;
        RECT 430.000 461.600 430.800 466.200 ;
        RECT 434.800 461.600 435.600 465.400 ;
        RECT 439.600 461.600 440.400 465.400 ;
        RECT 444.400 461.600 445.200 464.200 ;
        RECT 450.800 461.600 451.600 466.200 ;
        RECT 462.000 461.600 462.800 464.200 ;
        RECT 465.200 461.600 466.000 464.200 ;
        RECT 474.800 461.600 475.600 466.200 ;
        RECT 482.800 461.600 483.600 466.200 ;
        RECT 492.400 461.600 493.200 464.200 ;
        RECT 495.600 461.600 496.400 464.200 ;
        RECT 506.800 461.600 507.600 466.200 ;
        RECT 513.200 461.600 514.000 464.200 ;
        RECT 518.000 461.600 518.800 465.400 ;
        RECT 522.800 461.600 523.600 465.400 ;
        RECT 527.600 461.600 528.400 466.200 ;
        RECT 532.400 461.600 533.200 464.200 ;
        RECT 538.800 461.600 539.600 466.200 ;
        RECT 550.000 461.600 550.800 464.200 ;
        RECT 553.200 461.600 554.000 464.200 ;
        RECT 562.800 461.600 563.600 466.200 ;
        RECT 567.600 461.600 568.400 464.200 ;
        RECT 570.800 461.600 571.600 465.800 ;
        RECT 580.400 461.600 581.200 465.400 ;
        RECT 585.200 461.600 586.000 466.200 ;
        RECT 593.200 461.600 594.000 465.400 ;
        RECT 598.600 461.600 599.400 466.000 ;
        RECT 604.400 461.600 605.200 464.200 ;
        RECT 609.200 461.600 610.000 465.400 ;
        RECT 612.400 461.600 613.200 466.200 ;
        RECT 620.400 461.600 621.200 466.200 ;
        RECT 623.600 461.600 624.600 465.600 ;
        RECT 629.800 462.200 630.800 465.600 ;
        RECT 629.800 461.600 630.600 462.200 ;
        RECT 634.800 461.600 635.600 466.600 ;
        RECT 640.000 461.600 640.800 467.000 ;
        RECT 644.400 461.600 645.200 466.600 ;
        RECT 649.600 461.600 650.400 467.000 ;
        RECT 655.600 461.600 656.400 465.400 ;
        RECT 660.400 461.600 661.200 466.000 ;
        RECT 666.000 461.600 666.800 464.200 ;
        RECT 669.200 461.600 670.200 464.200 ;
        RECT 674.800 461.600 675.600 466.200 ;
        RECT 679.600 461.600 680.400 466.200 ;
        RECT 0.400 460.400 689.200 461.600 ;
        RECT 2.800 456.000 3.600 460.400 ;
        RECT 8.400 457.800 9.200 460.400 ;
        RECT 11.600 457.800 12.600 460.400 ;
        RECT 17.200 455.800 18.000 460.400 ;
        RECT 22.000 456.600 22.800 460.400 ;
        RECT 30.000 456.600 30.800 460.400 ;
        RECT 34.800 456.600 35.600 460.400 ;
        RECT 42.800 455.800 43.600 460.400 ;
        RECT 46.000 456.600 46.800 460.400 ;
        RECT 54.000 456.600 54.800 460.400 ;
        RECT 58.400 455.000 59.200 460.400 ;
        RECT 63.600 455.400 64.400 460.400 ;
        RECT 70.000 456.600 70.800 460.400 ;
        RECT 76.400 456.600 77.200 460.400 ;
        RECT 81.200 455.800 82.000 460.400 ;
        RECT 86.600 457.800 87.600 460.400 ;
        RECT 90.000 457.800 90.800 460.400 ;
        RECT 95.600 456.000 96.400 460.400 ;
        RECT 100.400 456.600 101.200 460.400 ;
        RECT 108.400 456.600 109.200 460.400 ;
        RECT 118.000 456.000 118.800 460.400 ;
        RECT 123.600 457.800 124.400 460.400 ;
        RECT 126.800 457.800 127.800 460.400 ;
        RECT 132.400 455.800 133.200 460.400 ;
        RECT 137.200 457.800 138.000 460.400 ;
        RECT 140.400 455.400 141.200 460.400 ;
        RECT 145.600 455.000 146.400 460.400 ;
        RECT 150.000 456.600 150.800 460.400 ;
        RECT 156.400 455.400 157.200 460.400 ;
        RECT 161.600 455.000 162.400 460.400 ;
        RECT 164.400 457.800 165.200 460.400 ;
        RECT 167.600 457.800 168.400 460.400 ;
        RECT 170.800 456.600 171.600 460.400 ;
        RECT 177.200 455.800 178.000 460.400 ;
        RECT 182.600 457.800 183.600 460.400 ;
        RECT 186.000 457.800 186.800 460.400 ;
        RECT 191.600 456.000 192.400 460.400 ;
        RECT 194.800 457.800 195.600 460.400 ;
        RECT 198.000 457.800 198.800 460.400 ;
        RECT 201.200 456.400 202.200 460.400 ;
        RECT 207.400 459.800 208.200 460.400 ;
        RECT 207.400 456.400 208.400 459.800 ;
        RECT 215.600 453.800 216.400 460.400 ;
        RECT 218.800 456.600 219.600 460.400 ;
        RECT 223.600 457.800 224.400 460.400 ;
        RECT 226.800 457.800 227.600 460.400 ;
        RECT 233.200 455.800 234.000 460.400 ;
        RECT 244.400 457.800 245.200 460.400 ;
        RECT 247.600 457.800 248.400 460.400 ;
        RECT 257.200 455.800 258.000 460.400 ;
        RECT 270.000 455.800 270.800 460.400 ;
        RECT 279.600 457.800 280.400 460.400 ;
        RECT 282.800 457.800 283.600 460.400 ;
        RECT 294.000 455.800 294.800 460.400 ;
        RECT 300.400 457.800 301.200 460.400 ;
        RECT 305.200 456.600 306.000 460.400 ;
        RECT 308.400 457.800 309.200 460.400 ;
        RECT 312.600 455.800 313.400 460.400 ;
        RECT 314.800 457.800 315.600 460.400 ;
        RECT 318.000 457.800 318.800 460.400 ;
        RECT 324.400 453.800 325.200 460.400 ;
        RECT 329.200 456.600 330.000 460.400 ;
        RECT 335.600 456.600 336.400 460.400 ;
        RECT 338.800 457.800 339.600 460.400 ;
        RECT 342.000 457.800 342.800 460.400 ;
        RECT 345.200 456.600 346.000 460.400 ;
        RECT 353.200 456.600 354.000 460.400 ;
        RECT 361.200 457.800 362.000 460.400 ;
        RECT 367.600 453.800 368.400 460.400 ;
        RECT 374.000 453.800 374.800 460.400 ;
        RECT 375.600 457.800 376.400 460.400 ;
        RECT 378.800 457.800 379.600 460.400 ;
        RECT 380.400 453.800 381.200 460.400 ;
        RECT 386.800 453.800 387.600 460.400 ;
        RECT 393.200 457.800 394.000 460.400 ;
        RECT 399.600 455.800 400.400 460.400 ;
        RECT 410.800 457.800 411.600 460.400 ;
        RECT 414.000 457.800 414.800 460.400 ;
        RECT 423.600 455.800 424.400 460.400 ;
        RECT 433.200 455.800 434.000 460.400 ;
        RECT 441.200 455.800 442.000 460.400 ;
        RECT 450.800 457.800 451.600 460.400 ;
        RECT 454.000 457.800 454.800 460.400 ;
        RECT 465.200 455.800 466.000 460.400 ;
        RECT 471.600 457.800 472.400 460.400 ;
        RECT 473.200 455.800 474.000 460.400 ;
        RECT 479.600 457.800 480.400 460.400 ;
        RECT 482.800 456.600 483.600 460.400 ;
        RECT 489.200 457.800 490.000 460.400 ;
        RECT 490.800 455.800 491.600 460.400 ;
        RECT 494.000 455.800 494.800 460.400 ;
        RECT 500.400 455.800 501.200 460.400 ;
        RECT 510.000 457.800 510.800 460.400 ;
        RECT 513.200 457.800 514.000 460.400 ;
        RECT 524.400 455.800 525.200 460.400 ;
        RECT 530.800 457.800 531.600 460.400 ;
        RECT 535.600 456.600 536.400 460.400 ;
        RECT 540.400 457.800 541.200 460.400 ;
        RECT 542.000 455.800 542.800 460.400 ;
        RECT 546.800 455.800 547.600 460.400 ;
        RECT 551.600 457.800 552.400 460.400 ;
        RECT 554.800 457.800 555.600 460.400 ;
        RECT 561.200 457.800 562.000 460.400 ;
        RECT 567.600 455.800 568.400 460.400 ;
        RECT 578.800 457.800 579.600 460.400 ;
        RECT 582.000 457.800 582.800 460.400 ;
        RECT 591.600 455.800 592.400 460.400 ;
        RECT 599.600 456.600 600.400 460.400 ;
        RECT 604.400 455.800 605.200 460.400 ;
        RECT 607.600 455.800 608.400 460.400 ;
        RECT 609.200 457.800 610.000 460.400 ;
        RECT 613.400 455.800 614.200 460.400 ;
        RECT 615.600 457.800 616.400 460.400 ;
        RECT 618.800 457.800 619.600 460.400 ;
        RECT 620.400 457.800 621.200 460.400 ;
        RECT 623.600 457.800 624.400 460.400 ;
        RECT 625.200 457.800 626.000 460.400 ;
        RECT 633.200 453.800 634.000 460.400 ;
        RECT 634.800 457.800 635.600 460.400 ;
        RECT 641.200 455.800 642.000 460.400 ;
        RECT 652.400 457.800 653.200 460.400 ;
        RECT 655.600 457.800 656.400 460.400 ;
        RECT 665.200 455.800 666.000 460.400 ;
        RECT 670.000 455.800 670.800 460.400 ;
        RECT 673.200 455.800 674.000 460.400 ;
        RECT 676.400 455.800 677.200 460.400 ;
        RECT 679.600 455.800 680.400 460.400 ;
        RECT 682.800 455.800 683.600 460.400 ;
        RECT 2.800 421.600 3.600 426.000 ;
        RECT 8.400 421.600 9.200 424.200 ;
        RECT 11.600 421.600 12.600 424.200 ;
        RECT 17.200 421.600 18.000 426.200 ;
        RECT 22.000 421.600 22.800 425.400 ;
        RECT 30.000 421.600 30.800 425.400 ;
        RECT 34.400 421.600 35.200 427.000 ;
        RECT 39.600 421.600 40.400 426.600 ;
        RECT 46.000 421.600 46.800 425.400 ;
        RECT 49.200 421.600 50.000 426.200 ;
        RECT 52.400 421.600 53.200 426.200 ;
        RECT 57.200 421.600 58.000 426.600 ;
        RECT 62.400 421.600 63.200 427.000 ;
        RECT 66.400 421.600 67.200 427.000 ;
        RECT 71.600 421.600 72.400 426.600 ;
        RECT 76.400 421.600 77.200 425.400 ;
        RECT 84.400 421.600 85.200 425.400 ;
        RECT 89.200 421.600 90.000 426.000 ;
        RECT 94.800 421.600 95.600 424.200 ;
        RECT 98.000 421.600 99.000 424.200 ;
        RECT 103.600 421.600 104.400 426.200 ;
        RECT 112.800 421.600 113.600 427.000 ;
        RECT 118.000 421.600 118.800 426.600 ;
        RECT 122.800 421.600 123.600 426.200 ;
        RECT 126.000 421.600 126.800 426.200 ;
        RECT 127.600 421.600 128.400 426.200 ;
        RECT 130.800 421.600 131.600 426.200 ;
        RECT 135.600 421.600 136.400 426.200 ;
        RECT 138.800 421.600 139.600 426.200 ;
        RECT 142.000 421.600 142.800 426.000 ;
        RECT 147.600 421.600 148.400 424.200 ;
        RECT 150.800 421.600 151.800 424.200 ;
        RECT 156.400 421.600 157.200 426.200 ;
        RECT 162.800 421.600 163.600 425.400 ;
        RECT 169.200 421.600 170.000 425.400 ;
        RECT 174.000 421.600 174.800 426.600 ;
        RECT 179.200 421.600 180.000 427.000 ;
        RECT 185.200 421.600 186.000 425.400 ;
        RECT 190.000 421.600 190.800 426.200 ;
        RECT 193.200 421.600 194.000 426.200 ;
        RECT 196.400 421.600 197.200 426.000 ;
        RECT 202.000 421.600 202.800 424.200 ;
        RECT 205.200 421.600 206.200 424.200 ;
        RECT 210.800 421.600 211.600 426.200 ;
        RECT 214.000 421.600 214.800 424.200 ;
        RECT 217.200 421.600 218.000 424.200 ;
        RECT 220.400 421.600 221.200 424.200 ;
        RECT 222.000 421.600 222.800 424.200 ;
        RECT 226.200 421.600 227.000 426.200 ;
        RECT 230.000 421.600 230.800 425.800 ;
        RECT 233.200 421.600 234.000 424.200 ;
        RECT 234.800 421.600 235.600 424.200 ;
        RECT 238.000 421.600 238.800 424.200 ;
        RECT 239.600 421.600 240.400 424.200 ;
        RECT 246.000 421.600 246.800 426.200 ;
        RECT 257.200 421.600 258.000 424.200 ;
        RECT 260.400 421.600 261.200 424.200 ;
        RECT 270.000 421.600 270.800 426.200 ;
        RECT 282.800 421.600 283.600 426.200 ;
        RECT 284.400 421.600 285.200 426.200 ;
        RECT 287.600 421.600 288.400 426.200 ;
        RECT 290.800 421.600 291.600 426.200 ;
        RECT 294.000 421.600 294.800 426.200 ;
        RECT 297.200 421.600 298.000 426.200 ;
        RECT 300.400 421.600 301.200 425.400 ;
        RECT 308.400 421.600 309.200 425.400 ;
        RECT 313.200 421.600 314.000 424.200 ;
        RECT 314.800 421.600 315.600 424.200 ;
        RECT 318.000 421.600 318.800 424.200 ;
        RECT 319.600 421.600 320.400 424.200 ;
        RECT 322.800 421.600 323.600 424.200 ;
        RECT 324.400 421.600 325.200 426.200 ;
        RECT 329.200 421.600 330.000 426.200 ;
        RECT 334.000 421.600 334.800 426.200 ;
        RECT 338.800 421.600 339.600 425.400 ;
        RECT 348.400 421.600 349.200 425.400 ;
        RECT 353.200 421.600 354.000 424.200 ;
        RECT 359.600 421.600 360.400 425.400 ;
        RECT 367.600 421.600 368.400 428.200 ;
        RECT 370.800 421.600 371.600 424.200 ;
        RECT 377.200 421.600 378.000 428.200 ;
        RECT 381.000 421.600 381.800 426.000 ;
        RECT 386.800 421.600 387.600 426.200 ;
        RECT 393.200 421.600 394.000 425.400 ;
        RECT 396.400 421.600 397.200 426.200 ;
        RECT 409.200 421.600 410.000 426.200 ;
        RECT 418.800 421.600 419.600 424.200 ;
        RECT 422.000 421.600 422.800 424.200 ;
        RECT 433.200 421.600 434.000 426.200 ;
        RECT 439.600 421.600 440.400 424.200 ;
        RECT 442.800 421.600 443.600 424.200 ;
        RECT 444.400 421.600 445.200 426.200 ;
        RECT 447.600 421.600 448.400 426.200 ;
        RECT 450.800 421.600 451.600 426.200 ;
        RECT 454.000 421.600 454.800 426.200 ;
        RECT 457.200 421.600 458.000 426.200 ;
        RECT 460.400 421.600 461.200 426.200 ;
        RECT 463.600 421.600 464.400 426.200 ;
        RECT 468.400 421.600 469.200 426.200 ;
        RECT 478.000 421.600 478.800 424.200 ;
        RECT 481.200 421.600 482.000 424.200 ;
        RECT 492.400 421.600 493.200 426.200 ;
        RECT 498.800 421.600 499.600 424.200 ;
        RECT 503.600 421.600 504.400 425.400 ;
        RECT 506.800 421.600 507.600 426.200 ;
        RECT 510.000 421.600 510.800 426.200 ;
        RECT 513.200 421.600 514.000 426.200 ;
        RECT 516.400 421.600 517.200 426.200 ;
        RECT 519.600 421.600 520.400 426.200 ;
        RECT 521.200 421.600 522.000 426.200 ;
        RECT 524.400 421.600 525.200 426.200 ;
        RECT 529.200 421.600 530.000 425.400 ;
        RECT 534.000 421.600 534.800 424.200 ;
        RECT 537.200 421.600 538.000 425.800 ;
        RECT 542.000 421.600 542.800 426.200 ;
        RECT 545.200 421.600 546.000 426.200 ;
        RECT 550.000 421.600 550.800 425.400 ;
        RECT 553.200 421.600 554.000 424.200 ;
        RECT 559.600 421.600 560.400 426.200 ;
        RECT 570.800 421.600 571.600 424.200 ;
        RECT 574.000 421.600 574.800 424.200 ;
        RECT 583.600 421.600 584.400 426.200 ;
        RECT 594.800 421.600 595.600 426.200 ;
        RECT 598.000 421.600 598.800 426.200 ;
        RECT 599.600 421.600 600.400 424.200 ;
        RECT 606.000 421.600 606.800 426.200 ;
        RECT 617.200 421.600 618.000 424.200 ;
        RECT 620.400 421.600 621.200 424.200 ;
        RECT 630.000 421.600 630.800 426.200 ;
        RECT 634.800 421.600 635.600 426.200 ;
        RECT 638.000 421.600 638.800 426.200 ;
        RECT 641.200 421.600 642.000 426.200 ;
        RECT 644.400 421.600 645.200 426.200 ;
        RECT 647.600 421.600 648.400 426.200 ;
        RECT 649.200 421.600 650.000 424.200 ;
        RECT 655.600 421.600 656.400 426.200 ;
        RECT 666.800 421.600 667.600 424.200 ;
        RECT 670.000 421.600 670.800 424.200 ;
        RECT 679.600 421.600 680.400 426.200 ;
        RECT 0.400 420.400 689.200 421.600 ;
        RECT 2.800 415.800 3.600 420.400 ;
        RECT 8.200 417.800 9.200 420.400 ;
        RECT 11.600 417.800 12.400 420.400 ;
        RECT 17.200 416.000 18.000 420.400 ;
        RECT 22.000 416.600 22.800 420.400 ;
        RECT 28.000 415.000 28.800 420.400 ;
        RECT 33.200 415.400 34.000 420.400 ;
        RECT 38.000 415.800 38.800 420.400 ;
        RECT 41.200 415.800 42.000 420.400 ;
        RECT 44.400 416.600 45.200 420.400 ;
        RECT 52.400 416.600 53.200 420.400 ;
        RECT 56.800 415.000 57.600 420.400 ;
        RECT 62.000 415.400 62.800 420.400 ;
        RECT 65.200 417.800 66.000 420.400 ;
        RECT 70.000 416.000 70.800 420.400 ;
        RECT 75.600 417.800 76.400 420.400 ;
        RECT 78.800 417.800 79.800 420.400 ;
        RECT 84.400 415.800 85.200 420.400 ;
        RECT 87.600 417.800 88.400 420.400 ;
        RECT 90.800 413.800 91.600 420.400 ;
        RECT 98.800 415.800 99.600 420.400 ;
        RECT 104.200 417.800 105.200 420.400 ;
        RECT 107.600 417.800 108.400 420.400 ;
        RECT 113.200 416.000 114.000 420.400 ;
        RECT 124.400 416.600 125.200 420.400 ;
        RECT 127.600 413.800 128.400 420.400 ;
        RECT 135.600 415.400 136.400 420.400 ;
        RECT 140.800 415.000 141.600 420.400 ;
        RECT 145.200 417.800 146.000 420.400 ;
        RECT 151.600 413.800 152.400 420.400 ;
        RECT 154.800 417.800 155.600 420.400 ;
        RECT 158.000 415.800 158.800 420.400 ;
        RECT 161.200 415.800 162.000 420.400 ;
        RECT 164.400 416.600 165.200 420.400 ;
        RECT 170.800 415.400 171.600 420.400 ;
        RECT 176.000 415.000 176.800 420.400 ;
        RECT 180.400 416.600 181.200 420.400 ;
        RECT 188.400 416.600 189.200 420.400 ;
        RECT 191.600 417.800 192.400 420.400 ;
        RECT 198.000 415.800 198.800 420.400 ;
        RECT 209.200 417.800 210.000 420.400 ;
        RECT 212.400 417.800 213.200 420.400 ;
        RECT 222.000 415.800 222.800 420.400 ;
        RECT 226.800 415.800 227.600 420.400 ;
        RECT 234.800 415.800 235.600 420.400 ;
        RECT 239.000 416.000 239.800 420.400 ;
        RECT 244.400 416.600 245.200 420.400 ;
        RECT 252.400 415.800 253.200 420.400 ;
        RECT 257.200 416.600 258.000 420.400 ;
        RECT 268.400 415.800 269.200 420.400 ;
        RECT 278.000 417.800 278.800 420.400 ;
        RECT 281.200 417.800 282.000 420.400 ;
        RECT 292.400 415.800 293.200 420.400 ;
        RECT 298.800 417.800 299.600 420.400 ;
        RECT 303.600 415.800 304.400 420.400 ;
        RECT 306.800 417.800 307.600 420.400 ;
        RECT 308.400 415.800 309.200 420.400 ;
        RECT 313.200 417.800 314.000 420.400 ;
        RECT 316.400 417.800 317.200 420.400 ;
        RECT 318.000 417.800 318.800 420.400 ;
        RECT 321.200 417.800 322.000 420.400 ;
        RECT 326.000 416.600 326.800 420.400 ;
        RECT 329.200 417.800 330.000 420.400 ;
        RECT 333.400 415.800 334.200 420.400 ;
        RECT 338.800 415.800 339.600 420.400 ;
        RECT 343.600 416.600 344.400 420.400 ;
        RECT 346.800 417.800 347.600 420.400 ;
        RECT 351.000 415.800 351.800 420.400 ;
        RECT 353.200 417.800 354.000 420.400 ;
        RECT 356.400 417.800 357.200 420.400 ;
        RECT 358.000 415.800 358.800 420.400 ;
        RECT 367.600 413.800 368.400 420.400 ;
        RECT 369.200 413.800 370.000 420.400 ;
        RECT 380.400 413.800 381.200 420.400 ;
        RECT 383.600 415.800 384.400 420.400 ;
        RECT 385.200 415.800 386.000 420.400 ;
        RECT 391.200 415.800 392.000 420.400 ;
        RECT 393.200 413.800 394.000 420.400 ;
        RECT 399.600 417.800 400.400 420.400 ;
        RECT 403.800 415.800 404.600 420.400 ;
        RECT 406.000 417.800 406.800 420.400 ;
        RECT 409.200 417.800 410.000 420.400 ;
        RECT 415.600 417.800 416.400 420.400 ;
        RECT 422.000 415.800 422.800 420.400 ;
        RECT 433.200 417.800 434.000 420.400 ;
        RECT 436.400 417.800 437.200 420.400 ;
        RECT 446.000 415.800 446.800 420.400 ;
        RECT 454.000 415.800 454.800 420.400 ;
        RECT 463.600 417.800 464.400 420.400 ;
        RECT 466.800 417.800 467.600 420.400 ;
        RECT 478.000 415.800 478.800 420.400 ;
        RECT 484.400 417.800 485.200 420.400 ;
        RECT 487.600 416.600 488.400 420.400 ;
        RECT 495.600 416.600 496.400 420.400 ;
        RECT 500.400 417.800 501.200 420.400 ;
        RECT 503.600 416.600 504.400 420.400 ;
        RECT 508.400 417.800 509.200 420.400 ;
        RECT 514.800 415.800 515.600 420.400 ;
        RECT 526.000 417.800 526.800 420.400 ;
        RECT 529.200 417.800 530.000 420.400 ;
        RECT 538.800 415.800 539.600 420.400 ;
        RECT 543.600 415.800 544.400 420.400 ;
        RECT 546.800 415.800 547.600 420.400 ;
        RECT 551.600 416.600 552.400 420.400 ;
        RECT 558.000 417.800 558.800 420.400 ;
        RECT 562.800 416.600 563.600 420.400 ;
        RECT 567.600 416.600 568.400 420.400 ;
        RECT 577.200 417.800 578.000 420.400 ;
        RECT 583.600 415.800 584.400 420.400 ;
        RECT 594.800 417.800 595.600 420.400 ;
        RECT 598.000 417.800 598.800 420.400 ;
        RECT 607.600 415.800 608.400 420.400 ;
        RECT 614.200 419.800 615.000 420.400 ;
        RECT 614.000 416.400 615.000 419.800 ;
        RECT 620.200 416.400 621.200 420.400 ;
        RECT 626.800 415.800 627.600 420.400 ;
        RECT 628.400 415.800 629.200 420.400 ;
        RECT 633.200 416.600 634.000 420.400 ;
        RECT 639.800 419.800 640.600 420.400 ;
        RECT 639.600 416.400 640.600 419.800 ;
        RECT 645.800 416.400 646.800 420.400 ;
        RECT 649.200 417.800 650.000 420.400 ;
        RECT 655.600 415.800 656.400 420.400 ;
        RECT 666.800 417.800 667.600 420.400 ;
        RECT 670.000 417.800 670.800 420.400 ;
        RECT 679.600 415.800 680.400 420.400 ;
        RECT 2.800 381.600 3.600 386.200 ;
        RECT 7.600 381.600 8.400 386.200 ;
        RECT 13.000 381.600 14.000 384.200 ;
        RECT 16.400 381.600 17.200 384.200 ;
        RECT 22.000 381.600 22.800 386.000 ;
        RECT 28.400 381.600 29.200 385.400 ;
        RECT 31.600 381.600 32.400 386.200 ;
        RECT 34.800 381.600 35.600 386.200 ;
        RECT 39.600 381.600 40.400 385.400 ;
        RECT 47.600 381.600 48.400 385.400 ;
        RECT 52.000 381.600 52.800 387.000 ;
        RECT 57.200 381.600 58.000 386.600 ;
        RECT 61.600 381.600 62.400 387.000 ;
        RECT 66.800 381.600 67.600 386.600 ;
        RECT 70.000 381.600 70.800 384.200 ;
        RECT 73.200 381.600 74.000 386.200 ;
        RECT 76.400 381.600 77.200 386.200 ;
        RECT 79.600 381.600 80.400 386.200 ;
        RECT 86.000 381.600 86.800 386.200 ;
        RECT 89.200 381.600 90.000 386.200 ;
        RECT 94.000 381.600 94.800 385.400 ;
        RECT 97.200 381.600 98.000 386.200 ;
        RECT 100.400 381.600 101.200 386.200 ;
        RECT 105.200 381.600 106.000 385.400 ;
        RECT 114.800 381.600 115.600 384.200 ;
        RECT 118.000 381.600 118.800 384.200 ;
        RECT 121.200 381.600 122.000 385.400 ;
        RECT 129.200 381.600 130.000 385.400 ;
        RECT 137.200 381.600 138.000 388.200 ;
        RECT 142.000 381.600 142.800 385.400 ;
        RECT 148.400 381.600 149.200 386.200 ;
        RECT 153.200 381.600 154.000 385.400 ;
        RECT 158.000 381.600 158.800 386.600 ;
        RECT 163.200 381.600 164.000 387.000 ;
        RECT 167.600 381.600 168.400 385.400 ;
        RECT 175.600 381.600 176.400 385.400 ;
        RECT 180.400 381.600 181.200 386.600 ;
        RECT 185.600 381.600 186.400 387.000 ;
        RECT 190.000 381.600 190.800 385.400 ;
        RECT 196.400 381.600 197.200 385.400 ;
        RECT 202.800 381.600 203.600 386.000 ;
        RECT 208.400 381.600 209.200 384.200 ;
        RECT 211.600 381.600 212.600 384.200 ;
        RECT 217.200 381.600 218.000 386.200 ;
        RECT 222.000 382.200 223.000 385.600 ;
        RECT 222.200 381.600 223.000 382.200 ;
        RECT 228.200 381.600 229.200 385.600 ;
        RECT 233.200 381.600 234.000 386.600 ;
        RECT 238.400 381.600 239.200 387.000 ;
        RECT 242.800 381.600 243.600 386.600 ;
        RECT 248.000 381.600 248.800 387.000 ;
        RECT 252.400 381.600 253.200 386.200 ;
        RECT 255.600 381.600 256.400 386.200 ;
        RECT 257.200 381.600 258.000 386.200 ;
        RECT 260.400 381.600 261.200 386.200 ;
        RECT 263.600 381.600 264.400 386.200 ;
        RECT 271.200 381.600 272.000 387.000 ;
        RECT 276.400 381.600 277.200 386.600 ;
        RECT 282.800 381.600 283.600 386.200 ;
        RECT 292.400 381.600 293.200 384.200 ;
        RECT 295.600 381.600 296.400 384.200 ;
        RECT 306.800 381.600 307.600 386.200 ;
        RECT 313.200 381.600 314.000 384.200 ;
        RECT 318.000 381.600 318.800 386.200 ;
        RECT 321.200 381.600 322.000 385.400 ;
        RECT 329.200 381.600 330.000 386.200 ;
        RECT 334.000 381.600 334.800 385.400 ;
        RECT 340.400 381.600 341.200 385.400 ;
        RECT 343.600 381.600 344.400 384.200 ;
        RECT 347.800 381.600 348.600 386.200 ;
        RECT 354.800 381.600 355.600 385.400 ;
        RECT 358.000 381.600 358.800 384.200 ;
        RECT 361.200 381.600 362.000 384.200 ;
        RECT 362.800 381.600 363.600 384.200 ;
        RECT 367.000 381.600 367.800 386.200 ;
        RECT 372.400 381.600 373.200 386.200 ;
        RECT 374.000 381.600 374.800 388.200 ;
        RECT 380.400 381.600 381.200 386.200 ;
        RECT 388.400 381.600 389.200 386.200 ;
        RECT 398.000 381.600 398.800 384.200 ;
        RECT 401.200 381.600 402.000 384.200 ;
        RECT 412.400 381.600 413.200 386.200 ;
        RECT 418.800 381.600 419.600 384.200 ;
        RECT 426.800 381.600 427.600 386.600 ;
        RECT 432.000 381.600 432.800 387.000 ;
        RECT 434.800 381.600 435.600 386.200 ;
        RECT 438.000 381.600 438.800 386.200 ;
        RECT 442.800 381.600 443.600 385.400 ;
        RECT 447.600 381.600 448.400 384.200 ;
        RECT 454.000 381.600 454.800 386.200 ;
        RECT 465.200 381.600 466.000 384.200 ;
        RECT 468.400 381.600 469.200 384.200 ;
        RECT 478.000 381.600 478.800 386.200 ;
        RECT 482.800 381.600 483.600 386.200 ;
        RECT 490.800 381.600 491.600 386.200 ;
        RECT 492.400 381.600 493.200 386.200 ;
        RECT 495.600 381.600 496.400 386.200 ;
        RECT 498.800 381.600 499.600 386.200 ;
        RECT 503.600 381.600 504.400 386.200 ;
        RECT 508.400 381.600 509.200 385.400 ;
        RECT 514.800 381.600 515.600 385.400 ;
        RECT 521.200 381.600 522.000 385.400 ;
        RECT 524.400 381.600 525.200 386.200 ;
        RECT 527.600 381.600 528.400 386.200 ;
        RECT 534.000 381.600 534.800 386.200 ;
        RECT 537.200 381.600 538.000 385.400 ;
        RECT 545.200 381.600 546.000 385.400 ;
        RECT 550.000 381.600 550.800 386.200 ;
        RECT 555.400 381.600 556.400 384.200 ;
        RECT 558.800 381.600 559.600 384.200 ;
        RECT 564.400 381.600 565.200 386.000 ;
        RECT 569.200 381.600 570.000 384.200 ;
        RECT 578.800 381.600 579.600 386.200 ;
        RECT 583.600 381.600 584.400 385.400 ;
        RECT 588.400 381.600 589.200 386.200 ;
        RECT 593.800 381.600 594.800 384.200 ;
        RECT 597.200 381.600 598.000 384.200 ;
        RECT 602.800 381.600 603.600 386.000 ;
        RECT 610.800 381.600 611.600 388.200 ;
        RECT 614.000 381.600 614.800 385.400 ;
        RECT 622.000 381.600 622.800 386.200 ;
        RECT 625.200 381.600 626.000 386.000 ;
        RECT 630.800 381.600 631.600 384.200 ;
        RECT 634.000 381.600 635.000 384.200 ;
        RECT 639.600 381.600 640.400 386.200 ;
        RECT 646.000 381.600 646.800 385.400 ;
        RECT 652.400 381.600 653.200 386.200 ;
        RECT 662.000 381.600 662.800 384.200 ;
        RECT 665.200 381.600 666.000 384.200 ;
        RECT 676.400 381.600 677.200 386.200 ;
        RECT 682.800 381.600 683.600 384.200 ;
        RECT 0.400 380.400 689.200 381.600 ;
        RECT 2.800 375.800 3.600 380.400 ;
        RECT 8.200 377.800 9.200 380.400 ;
        RECT 11.600 377.800 12.400 380.400 ;
        RECT 17.200 376.000 18.000 380.400 ;
        RECT 20.400 377.800 21.200 380.400 ;
        RECT 25.200 376.600 26.000 380.400 ;
        RECT 33.200 376.600 34.000 380.400 ;
        RECT 37.600 375.000 38.400 380.400 ;
        RECT 42.800 375.400 43.600 380.400 ;
        RECT 47.200 375.000 48.000 380.400 ;
        RECT 52.400 375.400 53.200 380.400 ;
        RECT 55.600 377.800 56.400 380.400 ;
        RECT 62.000 376.600 62.800 380.400 ;
        RECT 65.200 375.800 66.000 380.400 ;
        RECT 70.000 377.800 70.800 380.400 ;
        RECT 74.800 376.600 75.600 380.400 ;
        RECT 79.600 377.800 80.400 380.400 ;
        RECT 84.400 375.800 85.200 380.400 ;
        RECT 87.600 375.800 88.400 380.400 ;
        RECT 90.800 376.600 91.600 380.400 ;
        RECT 97.200 376.600 98.000 380.400 ;
        RECT 103.600 376.600 104.400 380.400 ;
        RECT 113.200 373.800 114.000 380.400 ;
        RECT 122.800 376.600 123.600 380.400 ;
        RECT 127.600 375.800 128.400 380.400 ;
        RECT 130.800 375.800 131.600 380.400 ;
        RECT 132.400 377.800 133.200 380.400 ;
        RECT 135.600 377.800 136.400 380.400 ;
        RECT 140.400 376.600 141.200 380.400 ;
        RECT 145.200 377.800 146.000 380.400 ;
        RECT 148.400 377.800 149.200 380.400 ;
        RECT 151.600 376.000 152.400 380.400 ;
        RECT 157.200 377.800 158.000 380.400 ;
        RECT 160.400 377.800 161.400 380.400 ;
        RECT 166.000 375.800 166.800 380.400 ;
        RECT 170.800 375.800 171.600 380.400 ;
        RECT 174.000 375.800 174.800 380.400 ;
        RECT 178.800 375.800 179.600 380.400 ;
        RECT 183.600 375.800 184.400 380.400 ;
        RECT 193.200 377.800 194.000 380.400 ;
        RECT 196.400 377.800 197.200 380.400 ;
        RECT 207.600 375.800 208.400 380.400 ;
        RECT 214.000 377.800 214.800 380.400 ;
        RECT 218.800 376.600 219.600 380.400 ;
        RECT 223.600 375.800 224.400 380.400 ;
        RECT 228.400 375.800 229.200 380.400 ;
        RECT 231.600 375.800 232.400 380.400 ;
        RECT 236.400 375.800 237.200 380.400 ;
        RECT 241.200 375.800 242.000 380.400 ;
        RECT 250.800 377.800 251.600 380.400 ;
        RECT 254.000 377.800 254.800 380.400 ;
        RECT 265.200 375.800 266.000 380.400 ;
        RECT 271.600 377.800 272.400 380.400 ;
        RECT 281.200 376.600 282.000 380.400 ;
        RECT 286.000 375.800 286.800 380.400 ;
        RECT 289.200 375.800 290.000 380.400 ;
        RECT 290.800 375.800 291.600 380.400 ;
        RECT 294.000 375.800 294.800 380.400 ;
        RECT 297.200 375.800 298.000 380.400 ;
        RECT 300.400 375.800 301.200 380.400 ;
        RECT 303.600 375.800 304.400 380.400 ;
        RECT 305.200 377.800 306.000 380.400 ;
        RECT 310.000 376.600 310.800 380.400 ;
        RECT 314.800 375.800 315.600 380.400 ;
        RECT 320.800 375.800 321.600 380.400 ;
        RECT 324.400 377.800 325.200 380.400 ;
        RECT 326.000 377.800 326.800 380.400 ;
        RECT 329.600 375.800 330.400 380.400 ;
        RECT 335.600 375.800 336.400 380.400 ;
        RECT 337.200 373.800 338.000 380.400 ;
        RECT 343.600 373.800 344.400 380.400 ;
        RECT 354.800 373.800 355.600 380.400 ;
        RECT 356.400 377.800 357.200 380.400 ;
        RECT 359.600 375.800 360.400 380.400 ;
        RECT 365.600 375.800 366.400 380.400 ;
        RECT 367.600 377.800 368.400 380.400 ;
        RECT 371.200 375.800 372.000 380.400 ;
        RECT 377.200 375.800 378.000 380.400 ;
        RECT 383.600 373.800 384.400 380.400 ;
        RECT 385.200 373.800 386.000 380.400 ;
        RECT 391.600 373.800 392.400 380.400 ;
        RECT 398.000 377.800 398.800 380.400 ;
        RECT 401.200 377.800 402.000 380.400 ;
        RECT 402.800 375.800 403.600 380.400 ;
        RECT 406.000 375.800 406.800 380.400 ;
        RECT 409.200 375.800 410.000 380.400 ;
        RECT 415.600 377.800 416.400 380.400 ;
        RECT 422.000 375.800 422.800 380.400 ;
        RECT 433.200 377.800 434.000 380.400 ;
        RECT 436.400 377.800 437.200 380.400 ;
        RECT 446.000 375.800 446.800 380.400 ;
        RECT 454.000 375.800 454.800 380.400 ;
        RECT 463.600 377.800 464.400 380.400 ;
        RECT 466.800 377.800 467.600 380.400 ;
        RECT 478.000 375.800 478.800 380.400 ;
        RECT 484.400 377.800 485.200 380.400 ;
        RECT 486.000 375.800 486.800 380.400 ;
        RECT 489.200 375.800 490.000 380.400 ;
        RECT 492.400 375.800 493.200 380.400 ;
        RECT 495.600 375.800 496.400 380.400 ;
        RECT 498.800 375.800 499.600 380.400 ;
        RECT 500.400 375.800 501.200 380.400 ;
        RECT 508.400 376.600 509.200 380.400 ;
        RECT 512.800 375.000 513.600 380.400 ;
        RECT 518.000 375.400 518.800 380.400 ;
        RECT 522.800 376.600 523.600 380.400 ;
        RECT 530.800 376.600 531.600 380.400 ;
        RECT 534.000 373.800 534.800 380.400 ;
        RECT 541.600 375.000 542.400 380.400 ;
        RECT 546.800 375.400 547.600 380.400 ;
        RECT 551.600 376.000 552.400 380.400 ;
        RECT 557.200 377.800 558.000 380.400 ;
        RECT 560.400 377.800 561.400 380.400 ;
        RECT 566.000 375.800 566.800 380.400 ;
        RECT 569.200 375.800 570.000 380.400 ;
        RECT 580.400 376.600 581.200 380.400 ;
        RECT 588.400 376.600 589.200 380.400 ;
        RECT 591.600 375.800 592.400 380.400 ;
        RECT 594.800 375.800 595.600 380.400 ;
        RECT 598.000 375.800 598.800 380.400 ;
        RECT 601.200 375.800 602.000 380.400 ;
        RECT 606.000 377.800 606.800 380.400 ;
        RECT 607.600 377.800 608.400 380.400 ;
        RECT 610.800 377.800 611.600 380.400 ;
        RECT 612.400 377.800 613.200 380.400 ;
        RECT 618.800 375.800 619.600 380.400 ;
        RECT 622.000 376.600 622.800 380.400 ;
        RECT 628.400 375.400 629.200 380.400 ;
        RECT 633.600 375.000 634.400 380.400 ;
        RECT 639.600 376.600 640.400 380.400 ;
        RECT 642.800 375.800 643.600 380.400 ;
        RECT 647.600 377.800 648.400 380.400 ;
        RECT 650.800 377.800 651.600 380.400 ;
        RECT 652.400 377.800 653.200 380.400 ;
        RECT 658.800 375.800 659.600 380.400 ;
        RECT 670.000 377.800 670.800 380.400 ;
        RECT 673.200 377.800 674.000 380.400 ;
        RECT 682.800 375.800 683.600 380.400 ;
        RECT 2.800 341.600 3.600 346.200 ;
        RECT 8.200 341.600 9.200 344.200 ;
        RECT 11.600 341.600 12.400 344.200 ;
        RECT 17.200 341.600 18.000 346.000 ;
        RECT 23.600 341.600 24.400 345.400 ;
        RECT 30.000 341.600 30.800 345.400 ;
        RECT 34.800 341.600 35.600 345.400 ;
        RECT 42.800 341.600 43.600 345.400 ;
        RECT 47.200 341.600 48.000 347.000 ;
        RECT 52.400 341.600 53.200 346.600 ;
        RECT 55.600 341.600 56.400 346.200 ;
        RECT 61.600 341.600 62.400 347.000 ;
        RECT 66.800 341.600 67.600 346.600 ;
        RECT 73.200 341.600 74.000 345.400 ;
        RECT 78.000 341.600 78.800 345.400 ;
        RECT 86.000 341.600 86.800 345.400 ;
        RECT 92.400 341.600 93.200 345.400 ;
        RECT 95.600 341.600 96.400 346.200 ;
        RECT 98.800 341.600 99.600 346.200 ;
        RECT 103.600 341.600 104.400 345.400 ;
        RECT 114.800 341.600 115.600 345.400 ;
        RECT 121.200 341.600 122.000 346.600 ;
        RECT 126.400 341.600 127.200 347.000 ;
        RECT 129.200 341.600 130.000 344.200 ;
        RECT 135.600 341.600 136.400 345.400 ;
        RECT 142.000 341.600 142.800 345.400 ;
        RECT 146.800 341.600 147.600 345.400 ;
        RECT 154.800 341.600 155.600 345.400 ;
        RECT 161.200 341.600 162.000 345.400 ;
        RECT 167.600 341.600 168.400 345.400 ;
        RECT 174.000 341.600 174.800 346.200 ;
        RECT 183.600 341.600 184.400 344.200 ;
        RECT 186.800 341.600 187.600 344.200 ;
        RECT 198.000 341.600 198.800 346.200 ;
        RECT 204.400 341.600 205.200 344.200 ;
        RECT 207.600 341.600 208.600 345.600 ;
        RECT 213.800 342.200 214.800 345.600 ;
        RECT 213.800 341.600 214.600 342.200 ;
        RECT 220.400 341.600 221.200 345.400 ;
        RECT 223.600 341.600 224.400 344.200 ;
        RECT 226.800 341.600 227.600 345.800 ;
        RECT 231.600 341.600 232.400 345.400 ;
        RECT 236.400 341.600 237.200 346.200 ;
        RECT 244.400 341.600 245.200 346.200 ;
        RECT 254.000 341.600 254.800 344.200 ;
        RECT 257.200 341.600 258.000 344.200 ;
        RECT 268.400 341.600 269.200 346.200 ;
        RECT 274.800 341.600 275.600 344.200 ;
        RECT 281.200 341.600 282.000 346.200 ;
        RECT 284.400 341.600 285.200 346.200 ;
        RECT 287.600 341.600 288.400 346.200 ;
        RECT 290.800 341.600 291.600 346.200 ;
        RECT 294.000 341.600 294.800 346.200 ;
        RECT 297.200 341.600 298.000 344.200 ;
        RECT 298.800 341.600 299.600 346.200 ;
        RECT 306.800 341.600 307.600 345.400 ;
        RECT 314.800 341.600 315.600 348.200 ;
        RECT 316.800 341.600 317.600 346.200 ;
        RECT 322.800 341.600 323.600 346.200 ;
        RECT 324.800 341.600 325.600 346.200 ;
        RECT 330.800 341.600 331.600 346.200 ;
        RECT 332.800 341.600 333.600 346.200 ;
        RECT 338.800 341.600 339.600 346.200 ;
        RECT 340.400 341.600 341.200 348.200 ;
        RECT 346.800 341.600 347.600 346.200 ;
        RECT 352.800 341.600 353.600 346.200 ;
        RECT 359.600 341.600 360.400 348.200 ;
        RECT 364.400 341.600 365.200 346.200 ;
        RECT 369.200 341.600 370.000 346.200 ;
        RECT 371.200 341.600 372.000 346.200 ;
        RECT 377.200 341.600 378.000 346.200 ;
        RECT 378.800 341.600 379.600 348.200 ;
        RECT 385.200 341.600 386.000 344.200 ;
        RECT 391.600 341.600 392.400 346.200 ;
        RECT 402.800 341.600 403.600 344.200 ;
        RECT 406.000 341.600 406.800 344.200 ;
        RECT 415.600 341.600 416.400 346.200 ;
        RECT 428.400 341.600 429.200 345.400 ;
        RECT 431.600 341.600 432.400 346.200 ;
        RECT 436.400 341.600 437.200 344.200 ;
        RECT 442.800 341.600 443.600 346.200 ;
        RECT 454.000 341.600 454.800 344.200 ;
        RECT 457.200 341.600 458.000 344.200 ;
        RECT 466.800 341.600 467.600 346.200 ;
        RECT 471.600 341.600 472.400 346.200 ;
        RECT 478.000 341.600 478.800 345.400 ;
        RECT 484.400 341.600 485.200 346.000 ;
        RECT 490.000 341.600 490.800 344.200 ;
        RECT 493.200 341.600 494.200 344.200 ;
        RECT 498.800 341.600 499.600 346.200 ;
        RECT 503.600 341.600 504.400 346.200 ;
        RECT 509.000 341.600 510.000 344.200 ;
        RECT 512.400 341.600 513.200 344.200 ;
        RECT 518.000 341.600 518.800 346.000 ;
        RECT 521.200 341.600 522.000 344.200 ;
        RECT 527.600 341.600 528.400 345.400 ;
        RECT 532.400 341.600 533.200 346.600 ;
        RECT 537.600 341.600 538.400 347.000 ;
        RECT 542.000 341.600 542.800 345.400 ;
        RECT 548.400 341.600 549.200 345.400 ;
        RECT 556.400 341.600 557.200 345.400 ;
        RECT 561.200 341.600 562.000 344.200 ;
        RECT 566.000 341.600 566.800 346.200 ;
        RECT 573.600 341.600 574.400 347.000 ;
        RECT 578.800 341.600 579.600 346.600 ;
        RECT 583.200 341.600 584.000 347.000 ;
        RECT 588.400 341.600 589.200 346.600 ;
        RECT 593.200 341.600 594.000 346.200 ;
        RECT 598.600 341.600 599.600 344.200 ;
        RECT 602.000 341.600 602.800 344.200 ;
        RECT 607.600 341.600 608.400 346.000 ;
        RECT 612.400 341.600 613.200 345.400 ;
        RECT 620.400 341.600 621.200 345.400 ;
        RECT 625.200 341.600 626.000 346.600 ;
        RECT 630.400 341.600 631.200 347.000 ;
        RECT 634.800 341.600 635.600 345.400 ;
        RECT 642.800 341.600 643.600 345.400 ;
        RECT 646.000 341.600 646.800 344.200 ;
        RECT 649.200 341.600 650.000 344.200 ;
        RECT 652.400 341.600 653.200 346.000 ;
        RECT 658.000 341.600 658.800 344.200 ;
        RECT 661.200 341.600 662.200 344.200 ;
        RECT 666.800 341.600 667.600 346.200 ;
        RECT 670.000 341.600 670.800 344.200 ;
        RECT 673.200 341.600 674.000 344.200 ;
        RECT 674.800 341.600 675.600 344.200 ;
        RECT 678.000 341.600 678.800 344.200 ;
        RECT 679.600 341.600 680.400 344.200 ;
        RECT 0.400 340.400 689.200 341.600 ;
        RECT 2.800 335.800 3.600 340.400 ;
        RECT 8.200 337.800 9.200 340.400 ;
        RECT 11.600 337.800 12.400 340.400 ;
        RECT 17.200 336.000 18.000 340.400 ;
        RECT 23.600 336.600 24.400 340.400 ;
        RECT 30.000 336.600 30.800 340.400 ;
        RECT 34.400 335.000 35.200 340.400 ;
        RECT 39.600 335.400 40.400 340.400 ;
        RECT 44.400 335.800 45.200 340.400 ;
        RECT 49.800 337.800 50.800 340.400 ;
        RECT 53.200 337.800 54.000 340.400 ;
        RECT 58.800 336.000 59.600 340.400 ;
        RECT 62.000 335.800 62.800 340.400 ;
        RECT 68.400 336.200 69.200 340.400 ;
        RECT 71.600 337.800 72.400 340.400 ;
        RECT 74.800 335.800 75.600 340.400 ;
        RECT 80.200 337.800 81.200 340.400 ;
        RECT 83.600 337.800 84.400 340.400 ;
        RECT 89.200 336.000 90.000 340.400 ;
        RECT 94.000 336.600 94.800 340.400 ;
        RECT 100.400 336.600 101.200 340.400 ;
        RECT 111.600 335.800 112.400 340.400 ;
        RECT 117.000 337.800 118.000 340.400 ;
        RECT 120.400 337.800 121.200 340.400 ;
        RECT 126.000 336.000 126.800 340.400 ;
        RECT 129.200 335.800 130.000 340.400 ;
        RECT 134.000 335.800 134.800 340.400 ;
        RECT 140.400 337.800 141.200 340.400 ;
        RECT 143.800 339.800 144.600 340.400 ;
        RECT 143.600 336.400 144.600 339.800 ;
        RECT 149.800 336.400 150.800 340.400 ;
        RECT 153.200 335.800 154.000 340.400 ;
        RECT 159.600 335.800 160.400 340.400 ;
        RECT 162.800 336.600 163.600 340.400 ;
        RECT 167.600 337.800 168.400 340.400 ;
        RECT 174.000 335.800 174.800 340.400 ;
        RECT 185.200 337.800 186.000 340.400 ;
        RECT 188.400 337.800 189.200 340.400 ;
        RECT 198.000 335.800 198.800 340.400 ;
        RECT 202.800 335.800 203.600 340.400 ;
        RECT 206.000 335.800 206.800 340.400 ;
        RECT 210.800 335.800 211.600 340.400 ;
        RECT 214.000 335.800 214.800 340.400 ;
        RECT 218.800 336.600 219.600 340.400 ;
        RECT 223.600 337.800 224.400 340.400 ;
        RECT 225.200 337.800 226.000 340.400 ;
        RECT 228.400 337.800 229.200 340.400 ;
        RECT 230.000 337.800 230.800 340.400 ;
        RECT 236.400 335.800 237.200 340.400 ;
        RECT 247.600 337.800 248.400 340.400 ;
        RECT 250.800 337.800 251.600 340.400 ;
        RECT 260.400 335.800 261.200 340.400 ;
        RECT 273.200 335.800 274.000 340.400 ;
        RECT 282.800 337.800 283.600 340.400 ;
        RECT 286.000 337.800 286.800 340.400 ;
        RECT 297.200 335.800 298.000 340.400 ;
        RECT 303.600 337.800 304.400 340.400 ;
        RECT 308.400 336.600 309.200 340.400 ;
        RECT 314.800 336.600 315.600 340.400 ;
        RECT 321.200 335.800 322.000 340.400 ;
        RECT 322.800 335.800 323.600 340.400 ;
        RECT 328.800 335.800 329.600 340.400 ;
        RECT 330.800 335.800 331.600 340.400 ;
        RECT 336.800 335.800 337.600 340.400 ;
        RECT 338.800 335.800 339.600 340.400 ;
        RECT 344.800 335.800 345.600 340.400 ;
        RECT 346.800 335.800 347.600 340.400 ;
        RECT 352.800 335.800 353.600 340.400 ;
        RECT 355.200 335.800 356.000 340.400 ;
        RECT 361.200 335.800 362.000 340.400 ;
        RECT 362.800 335.800 363.600 340.400 ;
        RECT 367.600 335.800 368.400 340.400 ;
        RECT 373.600 335.800 374.400 340.400 ;
        RECT 375.600 335.800 376.400 340.400 ;
        RECT 383.600 335.800 384.400 340.400 ;
        RECT 385.200 335.800 386.000 340.400 ;
        RECT 391.200 335.800 392.000 340.400 ;
        RECT 396.400 335.800 397.200 340.400 ;
        RECT 398.400 335.800 399.200 340.400 ;
        RECT 404.400 335.800 405.200 340.400 ;
        RECT 409.200 336.600 410.000 340.400 ;
        RECT 412.400 335.800 413.200 340.400 ;
        RECT 423.600 336.600 424.400 340.400 ;
        RECT 430.000 336.600 430.800 340.400 ;
        RECT 434.800 337.800 435.600 340.400 ;
        RECT 441.200 335.800 442.000 340.400 ;
        RECT 452.400 337.800 453.200 340.400 ;
        RECT 455.600 337.800 456.400 340.400 ;
        RECT 465.200 335.800 466.000 340.400 ;
        RECT 470.000 335.800 470.800 340.400 ;
        RECT 474.800 335.800 475.600 340.400 ;
        RECT 479.600 337.800 480.400 340.400 ;
        RECT 484.400 336.600 485.200 340.400 ;
        RECT 489.200 335.800 490.000 340.400 ;
        RECT 492.400 335.800 493.200 340.400 ;
        RECT 497.200 335.400 498.000 340.400 ;
        RECT 502.400 335.000 503.200 340.400 ;
        RECT 506.800 336.600 507.600 340.400 ;
        RECT 514.800 336.600 515.600 340.400 ;
        RECT 518.000 337.800 518.800 340.400 ;
        RECT 522.800 336.600 523.600 340.400 ;
        RECT 529.200 335.800 530.000 340.400 ;
        RECT 532.400 335.800 533.200 340.400 ;
        RECT 534.000 333.800 534.800 340.400 ;
        RECT 542.000 336.600 542.800 340.400 ;
        RECT 546.800 333.800 547.600 340.400 ;
        RECT 554.800 336.600 555.600 340.400 ;
        RECT 561.200 336.000 562.000 340.400 ;
        RECT 566.800 337.800 567.600 340.400 ;
        RECT 570.000 337.800 571.000 340.400 ;
        RECT 575.600 335.800 576.400 340.400 ;
        RECT 585.200 336.600 586.000 340.400 ;
        RECT 593.200 336.600 594.000 340.400 ;
        RECT 596.400 333.800 597.200 340.400 ;
        RECT 604.400 335.800 605.200 340.400 ;
        RECT 607.600 335.800 608.400 340.400 ;
        RECT 612.400 336.600 613.200 340.400 ;
        RECT 617.200 335.800 618.000 340.400 ;
        RECT 620.400 335.800 621.200 340.400 ;
        RECT 623.600 336.600 624.400 340.400 ;
        RECT 633.200 333.800 634.000 340.400 ;
        RECT 636.400 337.800 637.200 340.400 ;
        RECT 639.600 335.400 640.400 340.400 ;
        RECT 644.800 335.000 645.600 340.400 ;
        RECT 649.200 336.600 650.000 340.400 ;
        RECT 655.600 335.400 656.400 340.400 ;
        RECT 660.800 335.000 661.600 340.400 ;
        RECT 666.800 336.600 667.600 340.400 ;
        RECT 671.600 335.800 672.400 340.400 ;
        RECT 677.000 337.800 678.000 340.400 ;
        RECT 680.400 337.800 681.200 340.400 ;
        RECT 686.000 336.000 686.800 340.400 ;
        RECT 351.600 311.600 352.400 313.200 ;
        RECT 332.400 309.600 334.000 310.400 ;
        RECT 332.500 308.300 333.100 309.600 ;
        RECT 330.900 308.200 333.100 308.300 ;
        RECT 4.400 301.600 5.200 306.200 ;
        RECT 14.000 301.600 14.800 304.200 ;
        RECT 17.200 301.600 18.000 304.200 ;
        RECT 28.400 301.600 29.200 306.200 ;
        RECT 34.800 301.600 35.600 304.200 ;
        RECT 38.000 301.600 38.800 305.400 ;
        RECT 46.000 301.600 46.800 305.400 ;
        RECT 50.800 301.600 51.600 304.200 ;
        RECT 55.600 301.600 56.400 306.200 ;
        RECT 57.200 301.600 58.000 306.200 ;
        RECT 65.200 301.600 66.000 306.200 ;
        RECT 74.800 301.600 75.600 304.200 ;
        RECT 78.000 301.600 78.800 304.200 ;
        RECT 89.200 301.600 90.000 306.200 ;
        RECT 95.600 301.600 96.400 304.200 ;
        RECT 98.800 301.600 99.600 304.200 ;
        RECT 100.400 301.600 101.200 308.200 ;
        RECT 114.800 301.600 115.600 306.200 ;
        RECT 124.400 301.600 125.200 304.200 ;
        RECT 127.600 301.600 128.400 304.200 ;
        RECT 138.800 301.600 139.600 306.200 ;
        RECT 145.200 301.600 146.000 304.200 ;
        RECT 150.000 301.600 150.800 305.400 ;
        RECT 156.400 301.600 157.200 306.200 ;
        RECT 158.000 301.600 158.800 304.200 ;
        RECT 161.200 301.600 162.000 306.200 ;
        RECT 164.400 301.600 165.200 306.200 ;
        RECT 167.600 301.600 168.400 304.200 ;
        RECT 174.000 301.600 174.800 306.200 ;
        RECT 185.200 301.600 186.000 304.200 ;
        RECT 188.400 301.600 189.200 304.200 ;
        RECT 198.000 301.600 198.800 306.200 ;
        RECT 202.800 301.600 203.600 306.200 ;
        RECT 210.800 301.600 211.600 306.200 ;
        RECT 215.600 301.600 216.400 305.400 ;
        RECT 220.400 301.600 221.200 306.200 ;
        RECT 225.200 301.600 226.000 306.200 ;
        RECT 228.400 301.600 229.200 306.200 ;
        RECT 230.000 301.600 230.800 306.200 ;
        RECT 233.200 301.600 234.000 306.200 ;
        RECT 236.400 301.600 237.200 306.200 ;
        RECT 241.200 301.600 242.000 306.200 ;
        RECT 244.400 301.600 245.200 305.400 ;
        RECT 257.200 301.600 258.000 306.200 ;
        RECT 266.800 301.600 267.600 304.200 ;
        RECT 270.000 301.600 270.800 304.200 ;
        RECT 281.200 301.600 282.000 306.200 ;
        RECT 287.600 301.600 288.400 304.200 ;
        RECT 289.200 301.600 290.000 306.200 ;
        RECT 292.400 301.600 293.200 306.200 ;
        RECT 297.200 301.600 298.000 306.200 ;
        RECT 300.400 301.600 301.200 305.400 ;
        RECT 306.800 301.600 307.600 304.200 ;
        RECT 308.400 301.600 309.200 306.200 ;
        RECT 318.000 301.600 318.800 308.200 ;
        RECT 330.800 307.700 333.100 308.200 ;
        RECT 322.800 301.600 323.600 306.200 ;
        RECT 326.000 301.600 326.800 306.200 ;
        RECT 329.200 301.600 330.000 306.200 ;
        RECT 330.800 301.600 331.600 307.700 ;
        RECT 337.200 301.600 338.000 306.200 ;
        RECT 340.400 301.600 341.200 306.200 ;
        RECT 343.600 301.600 344.400 306.200 ;
        RECT 346.800 301.600 347.600 306.200 ;
        RECT 348.400 301.600 349.200 306.200 ;
        RECT 354.800 301.600 355.600 305.400 ;
        RECT 362.800 301.600 363.600 305.400 ;
        RECT 367.600 301.600 368.400 304.200 ;
        RECT 374.000 301.600 374.800 306.200 ;
        RECT 385.200 301.600 386.000 304.200 ;
        RECT 388.400 301.600 389.200 304.200 ;
        RECT 398.000 301.600 398.800 306.200 ;
        RECT 410.800 301.600 411.600 306.200 ;
        RECT 420.400 301.600 421.200 304.200 ;
        RECT 423.600 301.600 424.400 304.200 ;
        RECT 434.800 301.600 435.600 306.200 ;
        RECT 441.200 301.600 442.000 304.200 ;
        RECT 442.800 301.600 443.600 304.200 ;
        RECT 447.600 301.600 448.400 306.200 ;
        RECT 453.000 301.600 454.000 304.200 ;
        RECT 456.400 301.600 457.200 304.200 ;
        RECT 462.000 301.600 462.800 306.000 ;
        RECT 465.200 301.600 466.000 304.200 ;
        RECT 470.000 301.600 470.800 305.400 ;
        RECT 476.000 301.600 476.800 307.000 ;
        RECT 481.200 301.600 482.000 306.600 ;
        RECT 486.000 301.600 486.800 305.400 ;
        RECT 494.000 301.600 494.800 305.400 ;
        RECT 500.400 301.600 501.200 305.400 ;
        RECT 503.600 301.600 504.400 304.200 ;
        RECT 510.000 301.600 510.800 305.400 ;
        RECT 513.200 301.600 514.000 304.200 ;
        RECT 516.400 301.600 517.200 304.200 ;
        RECT 519.600 301.600 520.400 306.200 ;
        RECT 522.800 301.600 523.600 306.200 ;
        RECT 524.400 301.600 525.200 306.200 ;
        RECT 527.600 301.600 528.400 306.200 ;
        RECT 532.400 301.600 533.200 305.400 ;
        RECT 538.800 301.600 539.600 305.400 ;
        RECT 545.200 301.600 546.000 306.200 ;
        RECT 548.400 301.600 549.200 306.200 ;
        RECT 553.200 301.600 554.000 305.400 ;
        RECT 558.000 301.600 558.800 305.400 ;
        RECT 566.000 301.600 566.800 305.400 ;
        RECT 570.800 301.600 571.600 304.200 ;
        RECT 578.800 301.600 579.600 306.200 ;
        RECT 584.200 301.600 585.200 304.200 ;
        RECT 587.600 301.600 588.400 304.200 ;
        RECT 593.200 301.600 594.000 306.000 ;
        RECT 598.000 301.600 598.800 305.400 ;
        RECT 606.000 301.600 606.800 305.400 ;
        RECT 610.800 301.600 611.600 306.600 ;
        RECT 616.000 301.600 616.800 307.000 ;
        RECT 620.400 301.600 621.200 306.200 ;
        RECT 623.600 301.600 624.400 306.200 ;
        RECT 625.200 301.600 626.000 306.200 ;
        RECT 633.200 301.600 634.000 305.400 ;
        RECT 638.000 301.600 638.800 305.800 ;
        RECT 641.200 301.600 642.000 304.200 ;
        RECT 644.400 301.600 645.200 304.200 ;
        RECT 647.200 301.600 648.000 307.000 ;
        RECT 652.400 301.600 653.200 306.600 ;
        RECT 657.200 301.600 658.000 305.400 ;
        RECT 665.200 301.600 666.000 305.400 ;
        RECT 670.000 301.600 670.800 306.200 ;
        RECT 675.400 301.600 676.400 304.200 ;
        RECT 678.800 301.600 679.600 304.200 ;
        RECT 684.400 301.600 685.200 306.000 ;
        RECT 0.400 300.400 689.200 301.600 ;
        RECT 1.200 297.800 2.000 300.400 ;
        RECT 6.000 296.600 6.800 300.400 ;
        RECT 14.000 296.600 14.800 300.400 ;
        RECT 20.400 295.800 21.200 300.400 ;
        RECT 25.200 296.600 26.000 300.400 ;
        RECT 30.000 296.600 30.800 300.400 ;
        RECT 38.000 296.600 38.800 300.400 ;
        RECT 42.800 297.800 43.600 300.400 ;
        RECT 44.400 295.800 45.200 300.400 ;
        RECT 52.400 296.600 53.200 300.400 ;
        RECT 58.800 296.600 59.600 300.400 ;
        RECT 65.200 295.800 66.000 300.400 ;
        RECT 74.800 297.800 75.600 300.400 ;
        RECT 78.000 297.800 78.800 300.400 ;
        RECT 89.200 295.800 90.000 300.400 ;
        RECT 95.600 297.800 96.400 300.400 ;
        RECT 100.400 295.800 101.200 300.400 ;
        RECT 105.200 296.600 106.000 300.400 ;
        RECT 111.600 295.800 112.400 300.400 ;
        RECT 121.200 295.800 122.000 300.400 ;
        RECT 130.800 297.800 131.600 300.400 ;
        RECT 134.000 297.800 134.800 300.400 ;
        RECT 145.200 295.800 146.000 300.400 ;
        RECT 151.600 297.800 152.400 300.400 ;
        RECT 156.400 295.800 157.200 300.400 ;
        RECT 161.200 296.600 162.000 300.400 ;
        RECT 167.600 295.800 168.400 300.400 ;
        RECT 177.200 297.800 178.000 300.400 ;
        RECT 180.400 297.800 181.200 300.400 ;
        RECT 191.600 295.800 192.400 300.400 ;
        RECT 198.000 297.800 198.800 300.400 ;
        RECT 201.200 296.600 202.000 300.400 ;
        RECT 209.200 295.800 210.000 300.400 ;
        RECT 218.800 297.800 219.600 300.400 ;
        RECT 222.000 297.800 222.800 300.400 ;
        RECT 233.200 295.800 234.000 300.400 ;
        RECT 239.600 297.800 240.400 300.400 ;
        RECT 241.200 295.800 242.000 300.400 ;
        RECT 244.400 295.800 245.200 300.400 ;
        RECT 249.200 295.800 250.000 300.400 ;
        RECT 262.000 295.800 262.800 300.400 ;
        RECT 271.600 297.800 272.400 300.400 ;
        RECT 274.800 297.800 275.600 300.400 ;
        RECT 286.000 295.800 286.800 300.400 ;
        RECT 292.400 297.800 293.200 300.400 ;
        RECT 294.000 293.800 294.800 300.400 ;
        RECT 302.000 295.800 302.800 300.400 ;
        RECT 310.000 293.800 310.800 300.400 ;
        RECT 316.400 293.800 317.200 300.400 ;
        RECT 322.800 293.800 323.600 300.400 ;
        RECT 327.600 295.800 328.400 300.400 ;
        RECT 334.000 294.300 334.800 300.400 ;
        RECT 332.500 293.800 334.800 294.300 ;
        RECT 335.600 294.300 336.400 300.400 ;
        RECT 335.600 293.800 337.900 294.300 ;
        RECT 346.800 293.800 347.600 300.400 ;
        RECT 348.400 294.300 349.200 300.400 ;
        RECT 356.000 295.000 356.800 300.400 ;
        RECT 361.200 295.400 362.000 300.400 ;
        RECT 366.000 297.800 366.800 300.400 ;
        RECT 367.600 297.800 368.400 300.400 ;
        RECT 374.000 295.800 374.800 300.400 ;
        RECT 385.200 297.800 386.000 300.400 ;
        RECT 388.400 297.800 389.200 300.400 ;
        RECT 398.000 295.800 398.800 300.400 ;
        RECT 404.400 295.400 405.200 300.400 ;
        RECT 409.600 295.000 410.400 300.400 ;
        RECT 414.000 297.800 414.800 300.400 ;
        RECT 423.600 295.800 424.400 300.400 ;
        RECT 433.200 297.800 434.000 300.400 ;
        RECT 436.400 297.800 437.200 300.400 ;
        RECT 447.600 295.800 448.400 300.400 ;
        RECT 454.000 297.800 454.800 300.400 ;
        RECT 458.800 296.600 459.600 300.400 ;
        RECT 463.600 297.800 464.400 300.400 ;
        RECT 466.800 296.600 467.600 300.400 ;
        RECT 472.800 295.000 473.600 300.400 ;
        RECT 478.000 295.400 478.800 300.400 ;
        RECT 482.800 296.600 483.600 300.400 ;
        RECT 489.200 296.000 490.000 300.400 ;
        RECT 494.800 297.800 495.600 300.400 ;
        RECT 498.000 297.800 499.000 300.400 ;
        RECT 503.600 295.800 504.400 300.400 ;
        RECT 506.800 297.800 507.600 300.400 ;
        RECT 511.200 295.000 512.000 300.400 ;
        RECT 516.400 295.400 517.200 300.400 ;
        RECT 522.800 296.600 523.600 300.400 ;
        RECT 527.600 296.600 528.400 300.400 ;
        RECT 534.000 295.400 534.800 300.400 ;
        RECT 539.200 295.000 540.000 300.400 ;
        RECT 545.200 296.600 546.000 300.400 ;
        RECT 550.000 297.800 550.800 300.400 ;
        RECT 553.200 295.800 554.000 300.400 ;
        RECT 556.400 295.800 557.200 300.400 ;
        RECT 559.600 295.800 560.400 300.400 ;
        RECT 565.000 297.800 566.000 300.400 ;
        RECT 568.400 297.800 569.200 300.400 ;
        RECT 574.000 296.000 574.800 300.400 ;
        RECT 583.600 295.400 584.400 300.400 ;
        RECT 588.800 295.000 589.600 300.400 ;
        RECT 593.200 295.400 594.000 300.400 ;
        RECT 598.400 295.000 599.200 300.400 ;
        RECT 602.800 296.600 603.600 300.400 ;
        RECT 610.800 296.600 611.600 300.400 ;
        RECT 617.200 296.600 618.000 300.400 ;
        RECT 623.600 296.600 624.400 300.400 ;
        RECT 630.000 295.800 630.800 300.400 ;
        RECT 633.200 297.800 634.000 300.400 ;
        RECT 636.400 295.400 637.200 300.400 ;
        RECT 641.600 295.000 642.400 300.400 ;
        RECT 646.000 296.600 646.800 300.400 ;
        RECT 652.400 296.000 653.200 300.400 ;
        RECT 658.000 297.800 658.800 300.400 ;
        RECT 661.200 297.800 662.200 300.400 ;
        RECT 666.800 295.800 667.600 300.400 ;
        RECT 670.000 295.800 670.800 300.400 ;
        RECT 673.200 295.800 674.000 300.400 ;
        RECT 676.400 295.800 677.200 300.400 ;
        RECT 679.600 295.800 680.400 300.400 ;
        RECT 682.800 295.800 683.600 300.400 ;
        RECT 348.400 293.800 350.700 294.300 ;
        RECT 294.100 291.200 294.700 293.800 ;
        RECT 310.100 291.200 310.700 293.800 ;
        RECT 316.500 291.200 317.100 293.800 ;
        RECT 332.500 293.700 334.700 293.800 ;
        RECT 335.700 293.700 337.900 293.800 ;
        RECT 348.500 293.700 350.700 293.800 ;
        RECT 332.500 292.400 333.100 293.700 ;
        RECT 337.300 292.400 337.900 293.700 ;
        RECT 350.100 292.400 350.700 293.700 ;
        RECT 331.600 291.600 333.200 292.400 ;
        RECT 337.200 291.600 338.800 292.400 ;
        RECT 350.000 291.600 351.600 292.400 ;
        RECT 294.000 289.600 294.800 291.200 ;
        RECT 310.000 289.600 310.800 291.200 ;
        RECT 316.400 289.600 317.200 291.200 ;
        RECT 279.600 270.800 280.400 272.400 ;
        RECT 380.400 271.600 381.200 274.400 ;
        RECT 279.700 268.200 280.300 270.800 ;
        RECT 404.400 269.600 406.000 270.400 ;
        RECT 4.400 261.600 5.200 266.200 ;
        RECT 14.000 261.600 14.800 264.200 ;
        RECT 17.200 261.600 18.000 264.200 ;
        RECT 28.400 261.600 29.200 266.200 ;
        RECT 34.800 261.600 35.600 264.200 ;
        RECT 36.400 261.600 37.200 266.200 ;
        RECT 39.600 261.600 40.400 266.200 ;
        RECT 42.800 261.600 43.600 266.200 ;
        RECT 46.000 261.600 46.800 266.200 ;
        RECT 49.200 261.600 50.000 266.200 ;
        RECT 54.000 261.600 54.800 265.400 ;
        RECT 57.200 261.600 58.000 264.200 ;
        RECT 62.000 261.600 62.800 265.400 ;
        RECT 66.800 261.600 67.600 264.200 ;
        RECT 73.200 261.600 74.000 266.200 ;
        RECT 84.400 261.600 85.200 264.200 ;
        RECT 87.600 261.600 88.400 264.200 ;
        RECT 97.200 261.600 98.000 266.200 ;
        RECT 103.600 261.600 104.400 264.200 ;
        RECT 106.800 261.600 107.600 264.200 ;
        RECT 111.600 261.600 112.400 266.200 ;
        RECT 118.000 261.600 118.800 266.200 ;
        RECT 121.200 261.600 122.000 266.200 ;
        RECT 124.400 261.600 125.200 266.200 ;
        RECT 127.600 261.600 128.400 266.200 ;
        RECT 130.800 261.600 131.600 266.200 ;
        RECT 134.000 261.600 134.800 264.200 ;
        RECT 135.600 261.600 136.400 264.200 ;
        RECT 142.000 261.600 142.800 266.200 ;
        RECT 153.200 261.600 154.000 264.200 ;
        RECT 156.400 261.600 157.200 264.200 ;
        RECT 166.000 261.600 166.800 266.200 ;
        RECT 174.000 261.600 174.800 266.200 ;
        RECT 178.800 261.600 179.600 265.400 ;
        RECT 182.000 261.600 182.800 266.200 ;
        RECT 185.200 261.600 186.000 266.200 ;
        RECT 188.400 261.600 189.200 264.200 ;
        RECT 194.800 261.600 195.600 266.200 ;
        RECT 206.000 261.600 206.800 264.200 ;
        RECT 209.200 261.600 210.000 264.200 ;
        RECT 218.800 261.600 219.600 266.200 ;
        RECT 223.600 261.600 224.400 264.200 ;
        RECT 226.800 261.600 227.600 264.200 ;
        RECT 228.400 261.600 229.200 264.200 ;
        RECT 234.800 261.600 235.600 266.200 ;
        RECT 246.000 261.600 246.800 264.200 ;
        RECT 249.200 261.600 250.000 264.200 ;
        RECT 258.800 261.600 259.600 266.200 ;
        RECT 270.000 261.600 270.800 266.200 ;
        RECT 273.200 261.600 274.000 266.200 ;
        RECT 279.600 261.600 280.400 268.200 ;
        RECT 329.200 266.800 330.000 268.400 ;
        RECT 404.500 268.300 405.100 269.600 ;
        RECT 402.900 268.200 405.100 268.300 ;
        RECT 284.400 261.600 285.200 265.400 ;
        RECT 289.200 261.600 290.000 265.400 ;
        RECT 297.200 261.600 298.000 266.200 ;
        RECT 306.800 261.600 307.600 264.200 ;
        RECT 310.000 261.600 310.800 264.200 ;
        RECT 321.200 261.600 322.000 266.200 ;
        RECT 327.600 261.600 328.400 264.200 ;
        RECT 329.200 261.600 330.000 266.200 ;
        RECT 335.600 261.600 336.400 266.200 ;
        RECT 337.200 261.600 338.000 266.200 ;
        RECT 342.000 261.600 342.800 266.200 ;
        RECT 350.000 261.600 350.800 265.400 ;
        RECT 354.800 261.600 355.600 264.200 ;
        RECT 358.000 261.600 358.800 265.400 ;
        RECT 366.000 261.600 366.800 265.400 ;
        RECT 370.800 261.600 371.600 264.200 ;
        RECT 372.400 261.600 373.200 266.200 ;
        RECT 377.200 261.600 378.000 268.200 ;
        RECT 402.800 267.700 405.100 268.200 ;
        RECT 383.600 261.600 384.400 266.200 ;
        RECT 386.800 261.600 387.600 266.200 ;
        RECT 390.000 261.600 390.800 266.200 ;
        RECT 393.200 261.600 394.000 266.200 ;
        RECT 396.400 261.600 397.200 266.200 ;
        RECT 399.600 261.600 400.400 266.200 ;
        RECT 402.800 261.600 403.600 267.700 ;
        RECT 410.800 261.600 411.600 266.600 ;
        RECT 416.000 261.600 416.800 267.000 ;
        RECT 425.200 261.600 426.000 264.200 ;
        RECT 430.000 261.600 430.800 266.200 ;
        RECT 439.600 261.600 440.400 264.200 ;
        RECT 442.800 261.600 443.600 264.200 ;
        RECT 454.000 261.600 454.800 266.200 ;
        RECT 460.400 261.600 461.200 264.200 ;
        RECT 462.000 261.600 462.800 264.200 ;
        RECT 468.400 261.600 469.200 266.200 ;
        RECT 478.000 261.600 478.800 264.200 ;
        RECT 481.200 261.600 482.000 264.200 ;
        RECT 492.400 261.600 493.200 266.200 ;
        RECT 498.800 261.600 499.600 264.200 ;
        RECT 500.400 261.600 501.200 264.200 ;
        RECT 505.200 261.600 506.000 264.200 ;
        RECT 506.800 261.600 507.600 266.200 ;
        RECT 510.000 261.600 510.800 266.200 ;
        RECT 513.200 261.600 514.000 266.200 ;
        RECT 516.400 261.600 517.200 266.200 ;
        RECT 519.600 261.600 520.400 266.200 ;
        RECT 524.400 261.600 525.200 265.400 ;
        RECT 527.600 261.600 528.400 266.200 ;
        RECT 530.800 261.600 531.600 266.200 ;
        RECT 535.600 261.600 536.400 265.400 ;
        RECT 542.000 261.600 542.800 266.200 ;
        RECT 547.400 261.600 548.400 264.200 ;
        RECT 550.800 261.600 551.600 264.200 ;
        RECT 556.400 261.600 557.200 266.000 ;
        RECT 562.800 261.600 563.600 266.200 ;
        RECT 565.600 261.600 566.400 267.000 ;
        RECT 570.800 261.600 571.600 266.600 ;
        RECT 580.000 261.600 580.800 267.000 ;
        RECT 585.200 261.600 586.000 266.600 ;
        RECT 591.600 261.600 592.400 265.400 ;
        RECT 598.000 261.600 598.800 265.400 ;
        RECT 602.800 261.600 603.600 266.200 ;
        RECT 606.000 261.600 606.800 266.200 ;
        RECT 609.200 261.600 610.000 265.400 ;
        RECT 617.200 261.600 618.000 265.400 ;
        RECT 622.000 261.600 622.800 264.200 ;
        RECT 626.800 261.600 627.600 266.200 ;
        RECT 630.000 261.600 630.800 266.600 ;
        RECT 635.200 261.600 636.000 267.000 ;
        RECT 639.600 261.600 640.400 265.400 ;
        RECT 646.000 261.600 646.800 265.400 ;
        RECT 652.000 261.600 652.800 267.000 ;
        RECT 657.200 261.600 658.000 266.600 ;
        RECT 663.600 261.600 664.400 265.400 ;
        RECT 668.400 261.600 669.200 266.000 ;
        RECT 674.000 261.600 674.800 264.200 ;
        RECT 677.200 261.600 678.200 264.200 ;
        RECT 682.800 261.600 683.600 266.200 ;
        RECT 0.400 260.400 689.200 261.600 ;
        RECT 2.800 255.800 3.600 260.400 ;
        RECT 7.600 255.800 8.400 260.400 ;
        RECT 10.800 257.800 11.600 260.400 ;
        RECT 14.000 257.800 14.800 260.400 ;
        RECT 20.400 255.800 21.200 260.400 ;
        RECT 31.600 257.800 32.400 260.400 ;
        RECT 34.800 257.800 35.600 260.400 ;
        RECT 44.400 255.800 45.200 260.400 ;
        RECT 49.200 257.800 50.000 260.400 ;
        RECT 55.600 255.800 56.400 260.400 ;
        RECT 66.800 257.800 67.600 260.400 ;
        RECT 70.000 257.800 70.800 260.400 ;
        RECT 79.600 255.800 80.400 260.400 ;
        RECT 86.000 257.800 86.800 260.400 ;
        RECT 87.600 257.800 88.400 260.400 ;
        RECT 94.000 255.800 94.800 260.400 ;
        RECT 105.200 257.800 106.000 260.400 ;
        RECT 108.400 257.800 109.200 260.400 ;
        RECT 118.000 255.800 118.800 260.400 ;
        RECT 127.600 255.800 128.400 260.400 ;
        RECT 130.800 255.800 131.600 260.400 ;
        RECT 134.000 255.800 134.800 260.400 ;
        RECT 137.200 255.800 138.000 260.400 ;
        RECT 140.400 255.800 141.200 260.400 ;
        RECT 142.000 255.800 142.800 260.400 ;
        RECT 145.200 255.800 146.000 260.400 ;
        RECT 148.400 255.800 149.200 260.400 ;
        RECT 151.600 255.800 152.400 260.400 ;
        RECT 154.800 255.800 155.600 260.400 ;
        RECT 156.400 257.800 157.200 260.400 ;
        RECT 160.800 255.000 161.600 260.400 ;
        RECT 166.000 255.400 166.800 260.400 ;
        RECT 169.200 257.800 170.000 260.400 ;
        RECT 173.600 255.000 174.400 260.400 ;
        RECT 178.800 255.400 179.600 260.400 ;
        RECT 182.000 257.800 182.800 260.400 ;
        RECT 188.400 255.800 189.200 260.400 ;
        RECT 198.000 257.800 198.800 260.400 ;
        RECT 201.200 257.800 202.000 260.400 ;
        RECT 212.400 255.800 213.200 260.400 ;
        RECT 218.800 257.800 219.600 260.400 ;
        RECT 220.400 257.800 221.200 260.400 ;
        RECT 223.600 257.800 224.400 260.400 ;
        RECT 230.000 255.800 230.800 260.400 ;
        RECT 241.200 257.800 242.000 260.400 ;
        RECT 244.400 257.800 245.200 260.400 ;
        RECT 254.000 255.800 254.800 260.400 ;
        RECT 258.800 257.800 259.600 260.400 ;
        RECT 268.400 256.600 269.200 260.400 ;
        RECT 273.200 257.800 274.000 260.400 ;
        RECT 279.600 255.800 280.400 260.400 ;
        RECT 290.800 257.800 291.600 260.400 ;
        RECT 294.000 257.800 294.800 260.400 ;
        RECT 303.600 255.800 304.400 260.400 ;
        RECT 308.400 253.800 309.200 260.400 ;
        RECT 314.800 253.800 315.600 260.400 ;
        RECT 324.400 256.600 325.200 260.400 ;
        RECT 332.400 256.600 333.200 260.400 ;
        RECT 335.600 255.800 336.400 260.400 ;
        RECT 340.400 255.800 341.200 260.400 ;
        RECT 343.600 255.800 344.400 260.400 ;
        RECT 346.800 255.800 347.600 260.400 ;
        RECT 350.000 255.800 350.800 260.400 ;
        RECT 353.200 255.800 354.000 260.400 ;
        RECT 358.000 256.600 358.800 260.400 ;
        RECT 362.800 256.600 363.600 260.400 ;
        RECT 369.200 255.800 370.000 260.400 ;
        RECT 375.600 256.600 376.400 260.400 ;
        RECT 380.400 257.800 381.200 260.400 ;
        RECT 383.600 257.800 384.400 260.400 ;
        RECT 385.200 253.800 386.000 260.400 ;
        RECT 393.200 257.800 394.000 260.400 ;
        RECT 393.200 255.600 394.000 257.200 ;
        RECT 398.000 255.800 398.800 260.400 ;
        RECT 401.200 255.800 402.000 260.400 ;
        RECT 404.400 255.800 405.200 260.400 ;
        RECT 407.600 256.200 408.400 260.400 ;
        RECT 410.800 257.800 411.600 260.400 ;
        RECT 409.000 254.300 410.000 254.400 ;
        RECT 412.400 254.300 413.200 260.400 ;
        RECT 426.800 255.800 427.600 260.400 ;
        RECT 436.400 257.800 437.200 260.400 ;
        RECT 439.600 257.800 440.400 260.400 ;
        RECT 450.800 255.800 451.600 260.400 ;
        RECT 457.200 257.800 458.000 260.400 ;
        RECT 460.400 255.400 461.200 260.400 ;
        RECT 465.600 255.000 466.400 260.400 ;
        RECT 470.000 257.800 470.800 260.400 ;
        RECT 471.600 255.800 472.400 260.400 ;
        RECT 474.800 255.800 475.600 260.400 ;
        RECT 478.000 255.800 478.800 260.400 ;
        RECT 481.200 255.800 482.000 260.400 ;
        RECT 484.400 255.800 485.200 260.400 ;
        RECT 487.600 255.400 488.400 260.400 ;
        RECT 492.800 255.000 493.600 260.400 ;
        RECT 497.200 257.800 498.000 260.400 ;
        RECT 500.400 255.400 501.200 260.400 ;
        RECT 505.600 255.000 506.400 260.400 ;
        RECT 510.000 257.800 510.800 260.400 ;
        RECT 514.800 255.800 515.600 260.400 ;
        RECT 524.400 257.800 525.200 260.400 ;
        RECT 527.600 257.800 528.400 260.400 ;
        RECT 538.800 255.800 539.600 260.400 ;
        RECT 545.200 257.800 546.000 260.400 ;
        RECT 548.400 256.000 549.200 260.400 ;
        RECT 554.000 257.800 554.800 260.400 ;
        RECT 557.200 257.800 558.200 260.400 ;
        RECT 562.800 255.800 563.600 260.400 ;
        RECT 567.600 256.600 568.400 260.400 ;
        RECT 580.400 256.600 581.200 260.400 ;
        RECT 585.200 255.800 586.000 260.400 ;
        RECT 590.600 257.800 591.600 260.400 ;
        RECT 594.000 257.800 594.800 260.400 ;
        RECT 599.600 256.000 600.400 260.400 ;
        RECT 604.400 256.000 605.200 260.400 ;
        RECT 610.000 257.800 610.800 260.400 ;
        RECT 613.200 257.800 614.200 260.400 ;
        RECT 618.800 255.800 619.600 260.400 ;
        RECT 623.600 256.000 624.400 260.400 ;
        RECT 629.200 257.800 630.000 260.400 ;
        RECT 632.400 257.800 633.400 260.400 ;
        RECT 638.000 255.800 638.800 260.400 ;
        RECT 644.400 256.600 645.200 260.400 ;
        RECT 650.800 256.600 651.600 260.400 ;
        RECT 655.200 255.000 656.000 260.400 ;
        RECT 660.400 255.400 661.200 260.400 ;
        RECT 665.200 256.600 666.000 260.400 ;
        RECT 671.600 255.800 672.400 260.400 ;
        RECT 677.000 257.800 678.000 260.400 ;
        RECT 680.400 257.800 681.200 260.400 ;
        RECT 686.000 256.000 686.800 260.400 ;
        RECT 308.500 251.200 309.100 253.800 ;
        RECT 314.900 251.200 315.500 253.800 ;
        RECT 409.000 253.700 414.700 254.300 ;
        RECT 409.000 253.600 410.000 253.700 ;
        RECT 358.000 251.600 358.800 253.200 ;
        RECT 408.800 252.800 409.600 253.600 ;
        RECT 414.100 252.400 414.700 253.700 ;
        RECT 414.000 251.600 415.600 252.400 ;
        RECT 308.400 249.600 309.200 251.200 ;
        RECT 314.800 249.600 315.600 251.200 ;
        RECT 280.800 228.400 281.600 229.200 ;
        RECT 281.000 227.600 282.000 228.400 ;
        RECT 1.200 221.600 2.000 226.200 ;
        RECT 4.400 221.600 5.200 226.200 ;
        RECT 7.600 221.600 8.400 226.200 ;
        RECT 10.800 221.600 11.600 226.200 ;
        RECT 14.000 221.600 14.800 226.200 ;
        RECT 17.200 221.600 18.000 224.200 ;
        RECT 18.800 221.600 19.600 224.200 ;
        RECT 22.000 221.600 22.800 224.200 ;
        RECT 28.400 221.600 29.200 226.200 ;
        RECT 39.600 221.600 40.400 224.200 ;
        RECT 42.800 221.600 43.600 224.200 ;
        RECT 52.400 221.600 53.200 226.200 ;
        RECT 58.400 221.600 59.200 227.000 ;
        RECT 63.600 221.600 64.400 226.600 ;
        RECT 66.800 221.600 67.600 224.200 ;
        RECT 70.000 221.600 70.800 224.200 ;
        RECT 71.600 221.600 72.400 224.200 ;
        RECT 75.800 221.600 76.600 226.200 ;
        RECT 79.600 221.600 80.400 226.600 ;
        RECT 84.800 221.600 85.600 227.000 ;
        RECT 90.800 221.600 91.600 226.200 ;
        RECT 100.400 221.600 101.200 224.200 ;
        RECT 103.600 221.600 104.400 224.200 ;
        RECT 114.800 221.600 115.600 226.200 ;
        RECT 121.200 221.600 122.000 224.200 ;
        RECT 127.600 221.600 128.400 224.200 ;
        RECT 130.800 221.600 131.600 224.200 ;
        RECT 132.400 221.600 133.200 224.200 ;
        RECT 136.600 221.600 137.400 226.200 ;
        RECT 138.800 221.600 139.600 224.200 ;
        RECT 145.200 221.600 146.000 226.200 ;
        RECT 156.400 221.600 157.200 224.200 ;
        RECT 159.600 221.600 160.400 224.200 ;
        RECT 169.200 221.600 170.000 226.200 ;
        RECT 174.000 221.600 174.800 224.200 ;
        RECT 178.400 221.600 179.200 227.000 ;
        RECT 183.600 221.600 184.400 226.600 ;
        RECT 186.800 221.600 187.600 224.200 ;
        RECT 193.200 221.600 194.000 226.200 ;
        RECT 204.400 221.600 205.200 224.200 ;
        RECT 207.600 221.600 208.400 224.200 ;
        RECT 217.200 221.600 218.000 226.200 ;
        RECT 223.200 221.600 224.000 227.000 ;
        RECT 228.400 221.600 229.200 226.600 ;
        RECT 234.800 221.600 235.600 225.400 ;
        RECT 241.200 221.600 242.000 226.200 ;
        RECT 250.800 221.600 251.600 224.200 ;
        RECT 254.000 221.600 254.800 224.200 ;
        RECT 265.200 221.600 266.000 226.200 ;
        RECT 271.600 221.600 272.400 224.200 ;
        RECT 279.600 221.600 280.400 225.800 ;
        RECT 282.800 221.600 283.600 224.200 ;
        RECT 286.000 221.600 286.800 224.200 ;
        RECT 287.600 221.600 288.400 226.200 ;
        RECT 290.800 221.600 291.600 226.200 ;
        RECT 298.800 221.600 299.600 225.400 ;
        RECT 302.000 221.600 302.800 224.200 ;
        RECT 306.800 221.600 307.600 225.400 ;
        RECT 313.200 221.600 314.000 225.400 ;
        RECT 321.200 221.600 322.000 226.200 ;
        RECT 343.600 224.300 344.400 224.400 ;
        RECT 345.200 224.300 346.000 226.200 ;
        RECT 330.800 221.600 331.600 224.200 ;
        RECT 334.000 221.600 334.800 224.200 ;
        RECT 343.600 223.700 346.000 224.300 ;
        RECT 343.600 223.600 344.400 223.700 ;
        RECT 345.200 221.600 346.000 223.700 ;
        RECT 351.600 221.600 352.400 224.200 ;
        RECT 353.200 221.600 354.000 226.200 ;
        RECT 356.400 221.600 357.200 226.200 ;
        RECT 364.400 221.600 365.200 225.400 ;
        RECT 369.200 221.600 370.000 226.200 ;
        RECT 372.400 221.600 373.200 226.200 ;
        RECT 378.800 221.600 379.600 228.200 ;
        RECT 385.200 221.600 386.000 228.200 ;
        RECT 390.000 221.600 390.800 226.200 ;
        RECT 399.600 221.600 400.400 224.200 ;
        RECT 402.800 221.600 403.600 224.200 ;
        RECT 414.000 221.600 414.800 226.200 ;
        RECT 420.400 221.600 421.200 224.200 ;
        RECT 428.400 221.600 429.200 226.600 ;
        RECT 433.600 221.600 434.400 227.000 ;
        RECT 436.400 221.600 437.200 224.200 ;
        RECT 439.600 221.600 440.400 226.200 ;
        RECT 442.800 221.600 443.600 226.200 ;
        RECT 446.000 221.600 446.800 226.200 ;
        RECT 449.200 221.600 450.000 226.200 ;
        RECT 452.400 221.600 453.200 226.200 ;
        RECT 457.200 221.600 458.000 226.200 ;
        RECT 466.800 221.600 467.600 224.200 ;
        RECT 470.000 221.600 470.800 224.200 ;
        RECT 481.200 221.600 482.000 226.200 ;
        RECT 487.600 221.600 488.400 224.200 ;
        RECT 490.800 221.600 491.600 226.600 ;
        RECT 496.000 221.600 496.800 227.000 ;
        RECT 500.400 221.600 501.200 224.200 ;
        RECT 505.200 221.600 506.000 226.200 ;
        RECT 514.800 221.600 515.600 224.200 ;
        RECT 518.000 221.600 518.800 224.200 ;
        RECT 529.200 221.600 530.000 226.200 ;
        RECT 535.600 221.600 536.400 224.200 ;
        RECT 538.800 221.600 539.600 224.200 ;
        RECT 543.000 221.600 543.800 226.000 ;
        RECT 546.800 221.600 547.600 224.200 ;
        RECT 551.600 221.600 552.400 226.200 ;
        RECT 558.000 221.600 558.800 225.400 ;
        RECT 561.200 221.600 562.000 226.200 ;
        RECT 569.200 221.600 570.000 226.200 ;
        RECT 575.600 221.600 576.400 224.200 ;
        RECT 582.000 221.600 582.800 226.200 ;
        RECT 593.200 221.600 594.000 224.200 ;
        RECT 596.400 221.600 597.200 224.200 ;
        RECT 606.000 221.600 606.800 226.200 ;
        RECT 612.400 221.600 613.200 226.000 ;
        RECT 618.000 221.600 618.800 224.200 ;
        RECT 621.200 221.600 622.200 224.200 ;
        RECT 626.800 221.600 627.600 226.200 ;
        RECT 633.200 221.600 634.000 226.200 ;
        RECT 642.800 221.600 643.600 224.200 ;
        RECT 646.000 221.600 646.800 224.200 ;
        RECT 657.200 221.600 658.000 226.200 ;
        RECT 663.600 221.600 664.400 224.200 ;
        RECT 665.200 221.600 666.000 224.200 ;
        RECT 670.000 221.600 670.800 226.200 ;
        RECT 675.400 221.600 676.400 224.200 ;
        RECT 678.800 221.600 679.600 224.200 ;
        RECT 684.400 221.600 685.200 226.000 ;
        RECT 0.400 220.400 689.200 221.600 ;
        RECT 1.200 217.800 2.000 220.400 ;
        RECT 6.000 216.600 6.800 220.400 ;
        RECT 14.000 215.800 14.800 220.400 ;
        RECT 23.600 217.800 24.400 220.400 ;
        RECT 26.800 217.800 27.600 220.400 ;
        RECT 38.000 215.800 38.800 220.400 ;
        RECT 44.400 217.800 45.200 220.400 ;
        RECT 46.000 215.800 46.800 220.400 ;
        RECT 49.200 215.800 50.000 220.400 ;
        RECT 52.400 215.800 53.200 220.400 ;
        RECT 55.600 215.800 56.400 220.400 ;
        RECT 58.800 215.800 59.600 220.400 ;
        RECT 60.400 217.800 61.200 220.400 ;
        RECT 66.800 215.800 67.600 220.400 ;
        RECT 78.000 217.800 78.800 220.400 ;
        RECT 81.200 217.800 82.000 220.400 ;
        RECT 90.800 215.800 91.600 220.400 ;
        RECT 95.600 215.800 96.400 220.400 ;
        RECT 98.800 215.800 99.600 220.400 ;
        RECT 102.000 215.800 102.800 220.400 ;
        RECT 105.200 215.800 106.000 220.400 ;
        RECT 108.400 215.800 109.200 220.400 ;
        RECT 116.400 217.800 117.200 220.400 ;
        RECT 118.000 217.800 118.800 220.400 ;
        RECT 124.400 215.800 125.200 220.400 ;
        RECT 135.600 217.800 136.400 220.400 ;
        RECT 138.800 217.800 139.600 220.400 ;
        RECT 148.400 215.800 149.200 220.400 ;
        RECT 153.200 217.800 154.000 220.400 ;
        RECT 159.600 215.800 160.400 220.400 ;
        RECT 170.800 217.800 171.600 220.400 ;
        RECT 174.000 217.800 174.800 220.400 ;
        RECT 183.600 215.800 184.400 220.400 ;
        RECT 191.600 215.800 192.400 220.400 ;
        RECT 201.200 217.800 202.000 220.400 ;
        RECT 204.400 217.800 205.200 220.400 ;
        RECT 215.600 215.800 216.400 220.400 ;
        RECT 222.000 217.800 222.800 220.400 ;
        RECT 223.600 217.800 224.400 220.400 ;
        RECT 226.800 217.800 227.600 220.400 ;
        RECT 228.400 217.800 229.200 220.400 ;
        RECT 232.600 215.800 233.400 220.400 ;
        RECT 234.800 215.800 235.600 220.400 ;
        RECT 239.600 217.800 240.400 220.400 ;
        RECT 242.800 217.800 243.600 220.400 ;
        RECT 244.400 215.800 245.200 220.400 ;
        RECT 247.600 215.800 248.400 220.400 ;
        RECT 250.800 215.800 251.600 220.400 ;
        RECT 254.000 215.800 254.800 220.400 ;
        RECT 258.800 217.800 259.600 220.400 ;
        RECT 268.400 215.800 269.200 220.400 ;
        RECT 278.000 217.800 278.800 220.400 ;
        RECT 281.200 217.800 282.000 220.400 ;
        RECT 292.400 215.800 293.200 220.400 ;
        RECT 298.800 217.800 299.600 220.400 ;
        RECT 300.400 215.800 301.200 220.400 ;
        RECT 306.800 216.600 307.600 220.400 ;
        RECT 311.600 215.800 312.400 220.400 ;
        RECT 314.800 215.800 315.600 220.400 ;
        RECT 316.400 215.800 317.200 220.400 ;
        RECT 319.600 215.800 320.400 220.400 ;
        RECT 322.800 215.800 323.600 220.400 ;
        RECT 326.000 215.800 326.800 220.400 ;
        RECT 330.800 216.600 331.600 220.400 ;
        RECT 337.200 215.800 338.000 220.400 ;
        RECT 342.000 215.800 342.800 220.400 ;
        RECT 345.200 216.600 346.000 220.400 ;
        RECT 353.200 215.800 354.000 220.400 ;
        RECT 354.800 217.800 355.600 220.400 ;
        RECT 361.200 215.800 362.000 220.400 ;
        RECT 372.400 217.800 373.200 220.400 ;
        RECT 375.600 217.800 376.400 220.400 ;
        RECT 385.200 215.800 386.000 220.400 ;
        RECT 390.000 215.800 390.800 220.400 ;
        RECT 393.200 215.800 394.000 220.400 ;
        RECT 398.000 216.600 398.800 220.400 ;
        RECT 410.800 215.800 411.600 220.400 ;
        RECT 420.400 217.800 421.200 220.400 ;
        RECT 423.600 217.800 424.400 220.400 ;
        RECT 434.800 215.800 435.600 220.400 ;
        RECT 441.200 217.800 442.000 220.400 ;
        RECT 444.400 215.800 445.200 220.400 ;
        RECT 447.600 215.800 448.400 220.400 ;
        RECT 449.200 217.800 450.000 220.400 ;
        RECT 455.600 215.800 456.400 220.400 ;
        RECT 466.800 217.800 467.600 220.400 ;
        RECT 470.000 217.800 470.800 220.400 ;
        RECT 479.600 215.800 480.400 220.400 ;
        RECT 484.400 217.800 485.200 220.400 ;
        RECT 490.800 215.800 491.600 220.400 ;
        RECT 500.400 217.800 501.200 220.400 ;
        RECT 503.600 217.800 504.400 220.400 ;
        RECT 514.800 215.800 515.600 220.400 ;
        RECT 521.200 217.800 522.000 220.400 ;
        RECT 524.400 216.600 525.200 220.400 ;
        RECT 532.400 215.800 533.200 220.400 ;
        RECT 537.200 216.600 538.000 220.400 ;
        RECT 540.400 217.800 541.200 220.400 ;
        RECT 543.600 217.800 544.400 220.400 ;
        RECT 545.200 217.800 546.000 220.400 ;
        RECT 548.400 217.800 549.200 220.400 ;
        RECT 551.600 216.600 552.400 220.400 ;
        RECT 556.400 217.800 557.200 220.400 ;
        RECT 560.600 215.800 561.400 220.400 ;
        RECT 319.600 213.600 320.400 215.200 ;
        RECT 344.400 214.400 345.200 214.800 ;
        RECT 343.600 213.800 345.200 214.400 ;
        RECT 567.600 213.800 568.400 220.400 ;
        RECT 575.600 216.200 576.400 220.400 ;
        RECT 578.800 217.800 579.600 220.400 ;
        RECT 582.200 219.800 583.000 220.400 ;
        RECT 582.000 216.400 583.000 219.800 ;
        RECT 588.200 216.400 589.200 220.400 ;
        RECT 593.200 215.400 594.000 220.400 ;
        RECT 598.400 215.000 599.200 220.400 ;
        RECT 602.800 215.400 603.600 220.400 ;
        RECT 608.000 215.000 608.800 220.400 ;
        RECT 610.800 217.800 611.600 220.400 ;
        RECT 617.200 215.800 618.000 220.400 ;
        RECT 628.400 217.800 629.200 220.400 ;
        RECT 631.600 217.800 632.400 220.400 ;
        RECT 641.200 215.800 642.000 220.400 ;
        RECT 647.800 219.800 648.600 220.400 ;
        RECT 647.600 216.400 648.600 219.800 ;
        RECT 653.800 216.400 654.800 220.400 ;
        RECT 657.200 215.800 658.000 220.400 ;
        RECT 660.400 215.800 661.200 220.400 ;
        RECT 663.600 215.800 664.400 220.400 ;
        RECT 666.800 215.800 667.600 220.400 ;
        RECT 670.000 215.800 670.800 220.400 ;
        RECT 671.600 215.800 672.400 220.400 ;
        RECT 674.800 215.800 675.600 220.400 ;
        RECT 678.000 215.800 678.800 220.400 ;
        RECT 681.200 215.800 682.000 220.400 ;
        RECT 684.400 215.800 685.200 220.400 ;
        RECT 343.600 213.600 344.400 213.800 ;
        RECT 1.200 181.600 2.000 184.200 ;
        RECT 6.000 181.600 6.800 185.400 ;
        RECT 14.000 181.600 14.800 185.400 ;
        RECT 20.400 181.600 21.200 186.200 ;
        RECT 30.000 181.600 30.800 184.200 ;
        RECT 33.200 181.600 34.000 184.200 ;
        RECT 44.400 181.600 45.200 186.200 ;
        RECT 50.800 181.600 51.600 184.200 ;
        RECT 55.600 181.600 56.400 185.400 ;
        RECT 58.800 181.600 59.600 184.200 ;
        RECT 62.000 181.600 62.800 185.800 ;
        RECT 65.200 181.600 66.000 186.200 ;
        RECT 70.000 181.600 70.800 184.200 ;
        RECT 76.400 181.600 77.200 185.400 ;
        RECT 82.800 181.600 83.600 185.400 ;
        RECT 87.600 181.600 88.400 186.200 ;
        RECT 93.000 181.600 94.000 184.200 ;
        RECT 96.400 181.600 97.200 184.200 ;
        RECT 102.000 181.600 102.800 186.000 ;
        RECT 108.400 181.600 109.200 186.200 ;
        RECT 118.000 181.600 118.800 185.400 ;
        RECT 122.800 181.600 123.600 186.200 ;
        RECT 128.200 181.600 129.200 184.200 ;
        RECT 131.600 181.600 132.400 184.200 ;
        RECT 137.200 181.600 138.000 186.000 ;
        RECT 142.000 181.600 142.800 184.200 ;
        RECT 145.200 181.600 146.000 186.200 ;
        RECT 150.600 181.600 151.600 184.200 ;
        RECT 154.000 181.600 154.800 184.200 ;
        RECT 159.600 181.600 160.400 186.000 ;
        RECT 164.400 181.600 165.200 186.200 ;
        RECT 169.800 181.600 170.800 184.200 ;
        RECT 173.200 181.600 174.000 184.200 ;
        RECT 178.800 181.600 179.600 186.000 ;
        RECT 182.000 181.600 182.800 184.200 ;
        RECT 188.400 181.600 189.200 186.200 ;
        RECT 199.600 181.600 200.400 184.200 ;
        RECT 202.800 181.600 203.600 184.200 ;
        RECT 212.400 181.600 213.200 186.200 ;
        RECT 217.200 181.600 218.000 184.200 ;
        RECT 220.400 181.600 221.200 184.200 ;
        RECT 222.000 181.600 222.800 184.200 ;
        RECT 226.200 181.600 227.000 186.200 ;
        RECT 228.400 181.600 229.200 184.200 ;
        RECT 234.800 181.600 235.600 186.200 ;
        RECT 246.000 181.600 246.800 184.200 ;
        RECT 249.200 181.600 250.000 184.200 ;
        RECT 258.800 181.600 259.600 186.200 ;
        RECT 268.400 181.600 269.200 184.200 ;
        RECT 274.800 181.600 275.600 186.200 ;
        RECT 286.000 181.600 286.800 184.200 ;
        RECT 289.200 181.600 290.000 184.200 ;
        RECT 298.800 181.600 299.600 186.200 ;
        RECT 305.200 181.600 306.000 184.200 ;
        RECT 310.000 181.600 310.800 186.200 ;
        RECT 319.600 181.600 320.400 184.200 ;
        RECT 322.800 181.600 323.600 184.200 ;
        RECT 334.000 181.600 334.800 186.200 ;
        RECT 340.400 181.600 341.200 184.200 ;
        RECT 345.200 181.600 346.000 186.200 ;
        RECT 350.000 181.600 350.800 186.200 ;
        RECT 351.600 181.600 352.400 186.200 ;
        RECT 354.800 181.600 355.600 186.200 ;
        RECT 358.000 181.600 358.800 186.200 ;
        RECT 361.200 181.600 362.000 186.200 ;
        RECT 364.400 181.600 365.200 186.200 ;
        RECT 367.600 181.600 368.400 186.200 ;
        RECT 369.200 181.600 370.000 186.200 ;
        RECT 372.400 181.600 373.200 186.200 ;
        RECT 377.200 181.600 378.000 186.200 ;
        RECT 386.800 181.600 387.600 185.400 ;
        RECT 393.200 181.600 394.000 186.200 ;
        RECT 394.800 181.600 395.600 188.200 ;
        RECT 401.200 181.600 402.000 188.200 ;
        RECT 407.600 181.600 408.400 186.200 ;
        RECT 410.800 181.600 411.600 186.200 ;
        RECT 414.000 181.600 414.800 186.200 ;
        RECT 417.200 181.600 418.000 186.200 ;
        RECT 420.400 181.600 421.200 186.200 ;
        RECT 426.800 181.600 427.600 184.200 ;
        RECT 433.200 181.600 434.000 186.200 ;
        RECT 444.400 181.600 445.200 184.200 ;
        RECT 447.600 181.600 448.400 184.200 ;
        RECT 457.200 181.600 458.000 186.200 ;
        RECT 465.200 181.600 466.000 185.400 ;
        RECT 468.400 181.600 469.200 186.200 ;
        RECT 471.600 181.600 472.400 186.200 ;
        RECT 474.800 181.600 475.600 186.200 ;
        RECT 478.000 181.600 478.800 186.200 ;
        RECT 481.200 181.600 482.000 186.200 ;
        RECT 484.400 181.600 485.200 186.600 ;
        RECT 489.600 181.600 490.400 187.000 ;
        RECT 494.000 181.600 494.800 184.200 ;
        RECT 495.600 181.600 496.400 186.200 ;
        RECT 498.800 181.600 499.600 186.200 ;
        RECT 502.000 181.600 502.800 186.200 ;
        RECT 505.200 181.600 506.000 186.200 ;
        RECT 508.400 181.600 509.200 186.200 ;
        RECT 511.600 181.600 512.400 186.200 ;
        RECT 514.800 181.600 515.600 186.200 ;
        RECT 516.400 181.600 517.200 184.200 ;
        RECT 519.600 181.600 520.400 185.800 ;
        RECT 522.800 181.600 523.600 184.200 ;
        RECT 526.000 181.600 526.800 184.200 ;
        RECT 529.200 182.200 530.200 185.600 ;
        RECT 529.400 181.600 530.200 182.200 ;
        RECT 535.400 181.600 536.400 185.600 ;
        RECT 540.400 181.600 541.200 186.200 ;
        RECT 545.800 181.600 546.800 184.200 ;
        RECT 549.200 181.600 550.000 184.200 ;
        RECT 554.800 181.600 555.600 186.000 ;
        RECT 559.600 181.600 560.400 185.400 ;
        RECT 567.600 181.600 568.400 185.400 ;
        RECT 577.200 181.600 578.000 186.600 ;
        RECT 582.400 181.600 583.200 187.000 ;
        RECT 586.800 181.600 587.600 185.400 ;
        RECT 594.800 181.600 595.600 185.400 ;
        RECT 599.600 181.600 600.400 186.000 ;
        RECT 605.200 181.600 606.000 184.200 ;
        RECT 608.400 181.600 609.400 184.200 ;
        RECT 614.000 181.600 614.800 186.200 ;
        RECT 618.800 181.600 619.600 185.400 ;
        RECT 625.200 181.600 626.000 185.400 ;
        RECT 631.200 181.600 632.000 187.000 ;
        RECT 636.400 181.600 637.200 186.600 ;
        RECT 641.200 181.600 642.000 186.000 ;
        RECT 646.800 181.600 647.600 184.200 ;
        RECT 650.000 181.600 651.000 184.200 ;
        RECT 655.600 181.600 656.400 186.200 ;
        RECT 658.800 181.600 659.600 184.200 ;
        RECT 662.000 181.600 662.800 184.200 ;
        RECT 663.600 181.600 664.400 184.200 ;
        RECT 666.800 181.600 667.600 184.200 ;
        RECT 670.000 181.600 670.800 184.200 ;
        RECT 674.800 181.600 675.600 185.400 ;
        RECT 679.600 181.600 680.600 185.600 ;
        RECT 685.800 182.200 686.800 185.600 ;
        RECT 685.800 181.600 686.600 182.200 ;
        RECT 0.400 180.400 689.200 181.600 ;
        RECT 4.400 175.800 5.200 180.400 ;
        RECT 14.000 177.800 14.800 180.400 ;
        RECT 17.200 177.800 18.000 180.400 ;
        RECT 28.400 175.800 29.200 180.400 ;
        RECT 34.800 177.800 35.600 180.400 ;
        RECT 38.000 175.800 38.800 180.400 ;
        RECT 43.400 177.800 44.400 180.400 ;
        RECT 46.800 177.800 47.600 180.400 ;
        RECT 52.400 176.000 53.200 180.400 ;
        RECT 58.800 175.800 59.600 180.400 ;
        RECT 62.000 176.600 62.800 180.400 ;
        RECT 70.000 176.600 70.800 180.400 ;
        RECT 74.800 177.800 75.600 180.400 ;
        RECT 79.600 175.800 80.400 180.400 ;
        RECT 89.200 177.800 90.000 180.400 ;
        RECT 92.400 177.800 93.200 180.400 ;
        RECT 103.600 175.800 104.400 180.400 ;
        RECT 110.000 177.800 110.800 180.400 ;
        RECT 118.000 177.800 118.800 180.400 ;
        RECT 122.800 175.800 123.600 180.400 ;
        RECT 126.000 175.800 126.800 180.400 ;
        RECT 129.200 175.800 130.000 180.400 ;
        RECT 134.000 176.600 134.800 180.400 ;
        RECT 138.800 175.400 139.600 180.400 ;
        RECT 144.000 175.000 144.800 180.400 ;
        RECT 146.800 177.800 147.600 180.400 ;
        RECT 150.000 177.800 150.800 180.400 ;
        RECT 154.800 176.600 155.600 180.400 ;
        RECT 159.600 176.600 160.400 180.400 ;
        RECT 166.000 177.800 166.800 180.400 ;
        RECT 169.200 175.400 170.000 180.400 ;
        RECT 174.400 175.000 175.200 180.400 ;
        RECT 178.800 176.600 179.600 180.400 ;
        RECT 185.200 176.600 186.000 180.400 ;
        RECT 193.200 176.600 194.000 180.400 ;
        RECT 198.000 177.800 198.800 180.400 ;
        RECT 202.800 176.600 203.600 180.400 ;
        RECT 206.000 177.800 206.800 180.400 ;
        RECT 209.200 177.800 210.000 180.400 ;
        RECT 210.800 177.800 211.600 180.400 ;
        RECT 215.000 175.800 215.800 180.400 ;
        RECT 218.800 177.800 219.600 180.400 ;
        RECT 220.400 177.800 221.200 180.400 ;
        RECT 226.800 175.800 227.600 180.400 ;
        RECT 238.000 177.800 238.800 180.400 ;
        RECT 241.200 177.800 242.000 180.400 ;
        RECT 250.800 175.800 251.600 180.400 ;
        RECT 255.600 177.800 256.400 180.400 ;
        RECT 258.800 177.800 259.600 180.400 ;
        RECT 260.400 177.800 261.200 180.400 ;
        RECT 264.600 175.800 265.400 180.400 ;
        RECT 274.800 175.800 275.600 180.400 ;
        RECT 284.400 177.800 285.200 180.400 ;
        RECT 287.600 177.800 288.400 180.400 ;
        RECT 298.800 175.800 299.600 180.400 ;
        RECT 305.200 177.800 306.000 180.400 ;
        RECT 308.400 175.800 309.200 180.400 ;
        RECT 311.600 175.800 312.400 180.400 ;
        RECT 316.400 175.800 317.200 180.400 ;
        RECT 319.600 176.600 320.400 180.400 ;
        RECT 327.600 175.800 328.400 180.400 ;
        RECT 337.200 177.800 338.000 180.400 ;
        RECT 340.400 177.800 341.200 180.400 ;
        RECT 351.600 175.800 352.400 180.400 ;
        RECT 358.000 177.800 358.800 180.400 ;
        RECT 359.600 177.800 360.400 180.400 ;
        RECT 366.000 175.800 366.800 180.400 ;
        RECT 377.200 177.800 378.000 180.400 ;
        RECT 380.400 177.800 381.200 180.400 ;
        RECT 390.000 175.800 390.800 180.400 ;
        RECT 396.400 175.400 397.200 180.400 ;
        RECT 401.600 175.000 402.400 180.400 ;
        RECT 406.000 175.800 406.800 180.400 ;
        RECT 409.200 175.800 410.000 180.400 ;
        RECT 415.600 177.800 416.400 180.400 ;
        RECT 422.000 175.800 422.800 180.400 ;
        RECT 433.200 177.800 434.000 180.400 ;
        RECT 436.400 177.800 437.200 180.400 ;
        RECT 446.000 175.800 446.800 180.400 ;
        RECT 450.800 175.800 451.600 180.400 ;
        RECT 455.600 177.800 456.400 180.400 ;
        RECT 462.000 175.800 462.800 180.400 ;
        RECT 465.200 175.400 466.000 180.400 ;
        RECT 470.400 175.000 471.200 180.400 ;
        RECT 474.800 175.400 475.600 180.400 ;
        RECT 480.000 175.000 480.800 180.400 ;
        RECT 484.400 177.800 485.200 180.400 ;
        RECT 489.200 176.600 490.000 180.400 ;
        RECT 494.000 177.800 494.800 180.400 ;
        RECT 495.600 177.800 496.400 180.400 ;
        RECT 498.800 175.800 499.600 180.400 ;
        RECT 502.000 175.800 502.800 180.400 ;
        RECT 508.400 175.800 509.200 180.400 ;
        RECT 518.000 177.800 518.800 180.400 ;
        RECT 521.200 177.800 522.000 180.400 ;
        RECT 532.400 175.800 533.200 180.400 ;
        RECT 538.800 177.800 539.600 180.400 ;
        RECT 540.400 175.800 541.200 180.400 ;
        RECT 543.600 175.800 544.400 180.400 ;
        RECT 548.400 175.800 549.200 180.400 ;
        RECT 551.600 175.800 552.400 180.400 ;
        RECT 554.800 177.800 555.600 180.400 ;
        RECT 559.600 176.600 560.400 180.400 ;
        RECT 562.800 175.800 563.600 180.400 ;
        RECT 573.600 175.000 574.400 180.400 ;
        RECT 578.800 175.400 579.600 180.400 ;
        RECT 585.200 176.600 586.000 180.400 ;
        RECT 590.000 177.800 590.800 180.400 ;
        RECT 593.200 176.000 594.000 180.400 ;
        RECT 598.800 177.800 599.600 180.400 ;
        RECT 602.000 177.800 603.000 180.400 ;
        RECT 607.600 175.800 608.400 180.400 ;
        RECT 612.400 177.800 613.200 180.400 ;
        RECT 615.600 176.600 616.400 180.400 ;
        RECT 623.600 176.600 624.400 180.400 ;
        RECT 628.400 175.400 629.200 180.400 ;
        RECT 633.600 175.000 634.400 180.400 ;
        RECT 639.600 175.800 640.400 180.400 ;
        RECT 641.200 177.800 642.000 180.400 ;
        RECT 644.400 177.800 645.200 180.400 ;
        RECT 646.000 177.800 646.800 180.400 ;
        RECT 649.200 177.800 650.000 180.400 ;
        RECT 652.400 177.800 653.200 180.400 ;
        RECT 654.000 177.800 654.800 180.400 ;
        RECT 660.400 175.800 661.200 180.400 ;
        RECT 671.600 177.800 672.400 180.400 ;
        RECT 674.800 177.800 675.600 180.400 ;
        RECT 684.400 175.800 685.200 180.400 ;
        RECT 2.800 141.600 3.600 144.200 ;
        RECT 6.000 141.600 6.800 145.400 ;
        RECT 14.000 141.600 14.800 145.400 ;
        RECT 17.200 141.600 18.000 146.200 ;
        RECT 20.400 141.600 21.200 146.200 ;
        RECT 23.600 141.600 24.400 146.200 ;
        RECT 26.800 141.600 27.600 146.200 ;
        RECT 31.600 141.600 32.400 145.400 ;
        RECT 39.600 141.600 40.400 145.400 ;
        RECT 44.000 141.600 44.800 147.000 ;
        RECT 49.200 141.600 50.000 146.600 ;
        RECT 53.600 141.600 54.400 147.000 ;
        RECT 58.800 141.600 59.600 146.600 ;
        RECT 63.600 141.600 64.400 145.400 ;
        RECT 71.600 141.600 72.400 145.400 ;
        RECT 74.800 141.600 75.600 146.200 ;
        RECT 78.000 141.600 78.800 146.200 ;
        RECT 82.800 141.600 83.600 145.400 ;
        RECT 90.800 141.600 91.600 145.400 ;
        RECT 95.600 141.600 96.400 146.000 ;
        RECT 101.200 141.600 102.000 144.200 ;
        RECT 104.400 141.600 105.400 144.200 ;
        RECT 110.000 141.600 110.800 146.200 ;
        RECT 119.600 141.600 120.400 146.600 ;
        RECT 124.800 141.600 125.600 147.000 ;
        RECT 129.200 141.600 130.000 145.400 ;
        RECT 135.600 141.600 136.400 146.200 ;
        RECT 138.800 141.600 139.600 146.200 ;
        RECT 142.000 141.600 142.800 146.600 ;
        RECT 147.200 141.600 148.000 147.000 ;
        RECT 151.600 141.600 152.400 145.400 ;
        RECT 159.600 141.600 160.400 145.400 ;
        RECT 164.400 141.600 165.200 146.200 ;
        RECT 169.800 141.600 170.800 144.200 ;
        RECT 173.200 141.600 174.000 144.200 ;
        RECT 178.800 141.600 179.600 146.000 ;
        RECT 182.000 141.600 182.800 144.200 ;
        RECT 186.800 141.600 187.600 146.600 ;
        RECT 192.000 141.600 192.800 147.000 ;
        RECT 196.400 141.600 197.200 146.600 ;
        RECT 201.600 141.600 202.400 147.000 ;
        RECT 206.000 141.600 206.800 145.400 ;
        RECT 214.000 141.600 214.800 145.400 ;
        RECT 218.800 141.600 219.600 146.000 ;
        RECT 224.400 141.600 225.200 144.200 ;
        RECT 227.600 141.600 228.600 144.200 ;
        RECT 233.200 141.600 234.000 146.200 ;
        RECT 238.000 141.600 238.800 146.600 ;
        RECT 243.200 141.600 244.000 147.000 ;
        RECT 247.600 141.600 248.400 146.600 ;
        RECT 252.800 141.600 253.600 147.000 ;
        RECT 257.200 142.200 258.200 145.600 ;
        RECT 257.400 141.600 258.200 142.200 ;
        RECT 263.400 141.600 264.400 145.600 ;
        RECT 274.800 141.600 275.600 146.200 ;
        RECT 284.400 141.600 285.200 144.200 ;
        RECT 287.600 141.600 288.400 144.200 ;
        RECT 298.800 141.600 299.600 146.200 ;
        RECT 305.200 141.600 306.000 144.200 ;
        RECT 308.400 141.600 309.200 145.400 ;
        RECT 316.400 141.600 317.200 146.200 ;
        RECT 326.000 141.600 326.800 144.200 ;
        RECT 329.200 141.600 330.000 144.200 ;
        RECT 340.400 141.600 341.200 146.200 ;
        RECT 346.800 141.600 347.600 144.200 ;
        RECT 348.400 141.600 349.200 144.200 ;
        RECT 354.800 141.600 355.600 146.200 ;
        RECT 366.000 141.600 366.800 144.200 ;
        RECT 369.200 141.600 370.000 144.200 ;
        RECT 378.800 141.600 379.600 146.200 ;
        RECT 386.800 141.600 387.600 146.200 ;
        RECT 396.400 141.600 397.200 144.200 ;
        RECT 399.600 141.600 400.400 144.200 ;
        RECT 410.800 141.600 411.600 146.200 ;
        RECT 417.200 141.600 418.000 144.200 ;
        RECT 425.200 141.600 426.000 144.200 ;
        RECT 428.400 141.600 429.200 145.400 ;
        RECT 433.200 141.600 434.000 146.200 ;
        RECT 441.200 141.600 442.000 146.200 ;
        RECT 450.800 141.600 451.600 144.200 ;
        RECT 454.000 141.600 454.800 144.200 ;
        RECT 465.200 141.600 466.000 146.200 ;
        RECT 471.600 141.600 472.400 144.200 ;
        RECT 474.800 141.600 475.600 144.200 ;
        RECT 479.600 141.600 480.400 146.200 ;
        RECT 489.200 141.600 490.000 144.200 ;
        RECT 492.400 141.600 493.200 144.200 ;
        RECT 503.600 141.600 504.400 146.200 ;
        RECT 510.000 141.600 510.800 144.200 ;
        RECT 511.600 141.600 512.400 144.200 ;
        RECT 518.000 141.600 518.800 145.400 ;
        RECT 522.800 141.600 523.600 145.400 ;
        RECT 530.800 141.600 531.600 145.400 ;
        RECT 534.000 141.600 534.800 144.200 ;
        RECT 537.200 141.600 538.000 144.200 ;
        RECT 538.800 141.600 539.600 144.200 ;
        RECT 543.600 141.600 544.400 145.400 ;
        RECT 550.000 141.600 550.800 146.200 ;
        RECT 554.800 141.600 555.600 146.200 ;
        RECT 556.400 141.600 557.200 146.200 ;
        RECT 559.600 141.600 560.400 146.200 ;
        RECT 566.000 141.600 566.800 145.400 ;
        RECT 577.200 141.600 578.000 145.400 ;
        RECT 582.000 141.600 582.800 145.400 ;
        RECT 590.000 141.600 590.800 145.400 ;
        RECT 594.800 141.600 595.600 146.600 ;
        RECT 600.000 141.600 600.800 147.000 ;
        RECT 604.400 141.600 605.200 146.200 ;
        RECT 607.600 141.600 608.400 146.200 ;
        RECT 610.800 141.600 611.600 145.400 ;
        RECT 615.600 141.600 616.400 146.200 ;
        RECT 618.800 141.600 619.600 146.200 ;
        RECT 626.800 141.600 627.600 148.200 ;
        RECT 630.000 141.600 630.800 146.200 ;
        RECT 633.200 141.600 634.000 146.200 ;
        RECT 636.400 141.600 637.200 146.200 ;
        RECT 639.600 141.600 640.400 146.200 ;
        RECT 642.800 141.600 643.600 144.200 ;
        RECT 646.000 141.600 646.800 146.600 ;
        RECT 651.200 141.600 652.000 147.000 ;
        RECT 655.600 141.600 656.400 146.600 ;
        RECT 660.800 141.600 661.600 147.000 ;
        RECT 665.200 141.600 666.000 145.400 ;
        RECT 671.600 141.600 672.400 146.000 ;
        RECT 677.200 141.600 678.000 144.200 ;
        RECT 680.400 141.600 681.400 144.200 ;
        RECT 686.000 141.600 686.800 146.200 ;
        RECT 0.400 140.400 689.200 141.600 ;
        RECT 2.800 135.800 3.600 140.400 ;
        RECT 8.200 137.800 9.200 140.400 ;
        RECT 11.600 137.800 12.400 140.400 ;
        RECT 17.200 136.000 18.000 140.400 ;
        RECT 23.600 136.600 24.400 140.400 ;
        RECT 30.000 136.600 30.800 140.400 ;
        RECT 34.800 135.800 35.600 140.400 ;
        RECT 40.200 137.800 41.200 140.400 ;
        RECT 43.600 137.800 44.400 140.400 ;
        RECT 49.200 136.000 50.000 140.400 ;
        RECT 54.000 136.600 54.800 140.400 ;
        RECT 62.000 136.600 62.800 140.400 ;
        RECT 66.400 135.000 67.200 140.400 ;
        RECT 71.600 135.400 72.400 140.400 ;
        RECT 76.400 136.600 77.200 140.400 ;
        RECT 84.400 136.600 85.200 140.400 ;
        RECT 87.600 137.800 88.400 140.400 ;
        RECT 92.000 135.000 92.800 140.400 ;
        RECT 97.200 135.400 98.000 140.400 ;
        RECT 100.400 133.800 101.200 140.400 ;
        RECT 110.000 136.600 110.800 140.400 ;
        RECT 118.000 135.800 118.800 140.400 ;
        RECT 126.000 136.600 126.800 140.400 ;
        RECT 130.800 137.800 131.600 140.400 ;
        RECT 132.400 133.800 133.200 140.400 ;
        RECT 138.800 137.800 139.600 140.400 ;
        RECT 143.600 136.600 144.400 140.400 ;
        RECT 151.600 136.600 152.400 140.400 ;
        RECT 156.400 136.600 157.200 140.400 ;
        RECT 162.800 137.800 163.600 140.400 ;
        RECT 166.000 135.800 166.800 140.400 ;
        RECT 169.200 135.800 170.000 140.400 ;
        RECT 175.600 133.800 176.400 140.400 ;
        RECT 180.400 136.600 181.200 140.400 ;
        RECT 186.800 135.800 187.600 140.400 ;
        RECT 191.600 136.600 192.400 140.400 ;
        RECT 196.400 136.600 197.200 140.400 ;
        RECT 201.200 137.800 202.000 140.400 ;
        RECT 207.600 135.800 208.400 140.400 ;
        RECT 218.800 137.800 219.600 140.400 ;
        RECT 222.000 137.800 222.800 140.400 ;
        RECT 231.600 135.800 232.400 140.400 ;
        RECT 241.200 133.800 242.000 140.400 ;
        RECT 244.400 136.200 245.200 140.400 ;
        RECT 247.600 137.800 248.400 140.400 ;
        RECT 249.200 137.800 250.000 140.400 ;
        RECT 252.400 137.800 253.200 140.400 ;
        RECT 254.000 135.800 254.800 140.400 ;
        RECT 257.200 135.800 258.000 140.400 ;
        RECT 260.400 135.800 261.200 140.400 ;
        RECT 266.800 135.800 267.600 140.400 ;
        RECT 270.000 135.800 270.800 140.400 ;
        RECT 273.200 135.800 274.000 140.400 ;
        RECT 276.400 135.800 277.200 140.400 ;
        RECT 282.800 135.800 283.600 140.400 ;
        RECT 287.600 136.600 288.400 140.400 ;
        RECT 294.000 135.800 294.800 140.400 ;
        RECT 297.200 136.600 298.000 140.400 ;
        RECT 305.200 135.800 306.000 140.400 ;
        RECT 306.800 137.800 307.600 140.400 ;
        RECT 313.200 135.800 314.000 140.400 ;
        RECT 324.400 137.800 325.200 140.400 ;
        RECT 327.600 137.800 328.400 140.400 ;
        RECT 337.200 135.800 338.000 140.400 ;
        RECT 342.000 137.800 342.800 140.400 ;
        RECT 345.200 137.800 346.000 140.400 ;
        RECT 346.800 137.800 347.600 140.400 ;
        RECT 350.000 137.800 350.800 140.400 ;
        RECT 354.800 135.800 355.600 140.400 ;
        RECT 364.400 137.800 365.200 140.400 ;
        RECT 367.600 137.800 368.400 140.400 ;
        RECT 378.800 135.800 379.600 140.400 ;
        RECT 385.200 137.800 386.000 140.400 ;
        RECT 386.800 135.800 387.600 140.400 ;
        RECT 390.000 135.800 390.800 140.400 ;
        RECT 393.200 137.800 394.000 140.400 ;
        RECT 399.600 135.800 400.400 140.400 ;
        RECT 410.800 137.800 411.600 140.400 ;
        RECT 414.000 137.800 414.800 140.400 ;
        RECT 423.600 135.800 424.400 140.400 ;
        RECT 434.800 135.800 435.600 140.400 ;
        RECT 438.000 137.800 438.800 140.400 ;
        RECT 444.400 135.800 445.200 140.400 ;
        RECT 454.000 137.800 454.800 140.400 ;
        RECT 457.200 137.800 458.000 140.400 ;
        RECT 468.400 135.800 469.200 140.400 ;
        RECT 474.800 137.800 475.600 140.400 ;
        RECT 479.600 135.800 480.400 140.400 ;
        RECT 489.200 137.800 490.000 140.400 ;
        RECT 492.400 137.800 493.200 140.400 ;
        RECT 503.600 135.800 504.400 140.400 ;
        RECT 510.000 137.800 510.800 140.400 ;
        RECT 514.800 136.600 515.600 140.400 ;
        RECT 519.600 136.000 520.400 140.400 ;
        RECT 525.200 137.800 526.000 140.400 ;
        RECT 528.400 137.800 529.400 140.400 ;
        RECT 534.000 135.800 534.800 140.400 ;
        RECT 538.800 135.800 539.600 140.400 ;
        RECT 542.000 135.800 542.800 140.400 ;
        RECT 545.200 136.600 546.000 140.400 ;
        RECT 553.200 136.600 554.000 140.400 ;
        RECT 556.400 137.800 557.200 140.400 ;
        RECT 559.600 137.800 560.400 140.400 ;
        RECT 562.800 135.800 563.600 140.400 ;
        RECT 568.200 137.800 569.200 140.400 ;
        RECT 571.600 137.800 572.400 140.400 ;
        RECT 577.200 136.000 578.000 140.400 ;
        RECT 588.400 135.800 589.200 140.400 ;
        RECT 594.800 133.800 595.600 140.400 ;
        RECT 599.600 136.600 600.400 140.400 ;
        RECT 604.400 135.400 605.200 140.400 ;
        RECT 609.600 135.000 610.400 140.400 ;
        RECT 614.000 136.600 614.800 140.400 ;
        RECT 620.400 136.600 621.200 140.400 ;
        RECT 626.800 136.000 627.600 140.400 ;
        RECT 632.400 137.800 633.200 140.400 ;
        RECT 635.600 137.800 636.600 140.400 ;
        RECT 641.200 135.800 642.000 140.400 ;
        RECT 646.000 137.800 646.800 140.400 ;
        RECT 649.200 135.400 650.000 140.400 ;
        RECT 654.400 135.000 655.200 140.400 ;
        RECT 658.800 135.800 659.600 140.400 ;
        RECT 662.000 135.800 662.800 140.400 ;
        RECT 665.200 136.600 666.000 140.400 ;
        RECT 671.600 136.000 672.400 140.400 ;
        RECT 677.200 137.800 678.000 140.400 ;
        RECT 680.400 137.800 681.400 140.400 ;
        RECT 686.000 135.800 686.800 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 8.200 101.600 9.200 104.200 ;
        RECT 11.600 101.600 12.400 104.200 ;
        RECT 17.200 101.600 18.000 106.000 ;
        RECT 20.400 101.600 21.200 106.200 ;
        RECT 23.600 101.600 24.400 106.200 ;
        RECT 28.400 101.600 29.200 106.600 ;
        RECT 33.600 101.600 34.400 107.000 ;
        RECT 38.000 101.600 38.800 106.200 ;
        RECT 41.200 101.600 42.000 106.200 ;
        RECT 44.400 101.600 45.200 106.200 ;
        RECT 47.600 101.600 48.400 106.200 ;
        RECT 50.800 101.600 51.600 106.200 ;
        RECT 56.200 101.600 57.200 104.200 ;
        RECT 59.600 101.600 60.400 104.200 ;
        RECT 65.200 101.600 66.000 106.000 ;
        RECT 70.000 101.600 70.800 106.600 ;
        RECT 75.200 101.600 76.000 107.000 ;
        RECT 78.000 101.600 78.800 104.200 ;
        RECT 82.800 101.600 83.600 106.200 ;
        RECT 88.200 101.600 89.200 104.200 ;
        RECT 91.600 101.600 92.400 104.200 ;
        RECT 97.200 101.600 98.000 106.000 ;
        RECT 102.000 101.600 102.800 105.400 ;
        RECT 110.000 101.600 110.800 105.400 ;
        RECT 119.600 101.600 120.400 106.200 ;
        RECT 122.800 101.600 123.600 106.200 ;
        RECT 124.400 101.600 125.200 106.200 ;
        RECT 130.800 101.600 131.600 105.400 ;
        RECT 136.800 101.600 137.600 107.000 ;
        RECT 142.000 101.600 142.800 106.600 ;
        RECT 146.800 101.600 147.600 105.400 ;
        RECT 153.200 101.600 154.000 106.200 ;
        RECT 158.600 101.600 159.600 104.200 ;
        RECT 162.000 101.600 162.800 104.200 ;
        RECT 167.600 101.600 168.400 106.000 ;
        RECT 170.800 101.600 171.600 104.200 ;
        RECT 175.600 101.600 176.400 105.400 ;
        RECT 182.000 101.600 182.800 105.400 ;
        RECT 188.400 101.600 189.200 106.200 ;
        RECT 193.200 101.600 194.000 105.400 ;
        RECT 199.600 101.600 200.400 105.400 ;
        RECT 202.800 101.600 203.600 104.200 ;
        RECT 206.000 101.600 206.800 104.200 ;
        RECT 209.200 101.600 210.000 105.800 ;
        RECT 212.400 101.600 213.200 104.200 ;
        RECT 217.200 101.600 218.000 106.200 ;
        RECT 220.400 101.600 221.200 104.200 ;
        RECT 222.000 101.600 222.800 104.200 ;
        RECT 225.200 101.600 226.000 104.200 ;
        RECT 227.400 101.600 228.200 106.200 ;
        RECT 231.600 101.600 232.400 104.200 ;
        RECT 234.800 101.600 235.600 105.400 ;
        RECT 241.200 101.600 242.000 105.400 ;
        RECT 246.000 101.600 246.800 106.200 ;
        RECT 252.400 101.600 253.200 105.400 ;
        RECT 257.200 101.600 258.000 106.200 ;
        RECT 266.800 101.600 267.600 104.200 ;
        RECT 273.200 101.600 274.000 106.200 ;
        RECT 284.400 101.600 285.200 104.200 ;
        RECT 287.600 101.600 288.400 104.200 ;
        RECT 297.200 101.600 298.000 106.200 ;
        RECT 303.600 101.600 304.400 106.200 ;
        RECT 306.800 101.600 307.600 106.200 ;
        RECT 310.000 101.600 310.800 106.200 ;
        RECT 314.800 101.600 315.600 104.200 ;
        RECT 318.000 101.600 318.800 105.400 ;
        RECT 322.800 101.600 323.600 106.200 ;
        RECT 327.600 101.600 328.400 104.200 ;
        RECT 334.000 101.600 334.800 106.200 ;
        RECT 345.200 101.600 346.000 104.200 ;
        RECT 348.400 101.600 349.200 104.200 ;
        RECT 358.000 101.600 358.800 106.200 ;
        RECT 362.800 101.600 363.600 104.200 ;
        RECT 369.200 101.600 370.000 106.200 ;
        RECT 380.400 101.600 381.200 104.200 ;
        RECT 383.600 101.600 384.400 104.200 ;
        RECT 393.200 101.600 394.000 106.200 ;
        RECT 399.600 101.600 400.400 104.200 ;
        RECT 404.400 101.600 405.200 105.400 ;
        RECT 407.600 101.600 408.400 106.200 ;
        RECT 415.600 101.600 416.400 105.400 ;
        RECT 423.600 101.600 424.400 104.200 ;
        RECT 430.000 101.600 430.800 106.200 ;
        RECT 441.200 101.600 442.000 104.200 ;
        RECT 444.400 101.600 445.200 104.200 ;
        RECT 454.000 101.600 454.800 106.200 ;
        RECT 458.800 101.600 459.600 106.200 ;
        RECT 462.000 101.600 462.800 106.200 ;
        RECT 466.800 101.600 467.600 105.400 ;
        RECT 471.600 101.600 472.400 106.200 ;
        RECT 476.400 101.600 477.200 106.200 ;
        RECT 481.200 101.600 482.000 104.200 ;
        RECT 487.600 101.600 488.400 106.200 ;
        RECT 498.800 101.600 499.600 104.200 ;
        RECT 502.000 101.600 502.800 104.200 ;
        RECT 511.600 101.600 512.400 106.200 ;
        RECT 516.400 101.600 517.200 106.200 ;
        RECT 519.600 101.600 520.400 106.200 ;
        RECT 526.000 101.600 526.800 105.400 ;
        RECT 529.200 101.600 530.000 106.200 ;
        RECT 532.400 101.600 533.200 106.200 ;
        RECT 535.600 101.600 536.400 106.200 ;
        RECT 538.800 101.600 539.600 106.200 ;
        RECT 542.000 101.600 542.800 106.200 ;
        RECT 546.800 101.600 547.600 105.400 ;
        RECT 550.000 101.600 550.800 106.200 ;
        RECT 556.000 101.600 556.800 107.000 ;
        RECT 561.200 101.600 562.000 106.600 ;
        RECT 566.000 101.600 566.800 106.200 ;
        RECT 569.200 101.600 570.000 106.200 ;
        RECT 575.600 101.600 576.400 106.200 ;
        RECT 582.000 101.600 582.800 104.200 ;
        RECT 586.800 101.600 587.600 105.400 ;
        RECT 591.600 101.600 592.400 105.400 ;
        RECT 599.600 101.600 600.400 106.200 ;
        RECT 602.800 101.600 603.600 104.200 ;
        RECT 606.000 101.600 606.800 106.000 ;
        RECT 611.600 101.600 612.400 104.200 ;
        RECT 614.800 101.600 615.800 104.200 ;
        RECT 620.400 101.600 621.200 106.200 ;
        RECT 625.200 101.600 626.000 105.400 ;
        RECT 633.200 101.600 634.000 105.400 ;
        RECT 638.000 101.600 638.800 106.600 ;
        RECT 643.200 101.600 644.000 107.000 ;
        RECT 646.000 101.600 646.800 106.200 ;
        RECT 649.200 101.600 650.000 106.200 ;
        RECT 652.400 101.600 653.200 106.200 ;
        RECT 655.600 101.600 656.400 106.200 ;
        RECT 658.800 101.600 659.600 106.200 ;
        RECT 662.000 101.600 662.800 106.200 ;
        RECT 665.200 101.600 666.000 106.200 ;
        RECT 668.400 101.600 669.200 106.200 ;
        RECT 671.600 101.600 672.400 106.200 ;
        RECT 674.800 101.600 675.600 105.400 ;
        RECT 681.200 101.600 682.000 106.600 ;
        RECT 686.400 101.600 687.200 107.000 ;
        RECT 0.400 100.400 689.200 101.600 ;
        RECT 4.400 96.600 5.200 100.400 ;
        RECT 8.800 95.000 9.600 100.400 ;
        RECT 14.000 95.400 14.800 100.400 ;
        RECT 20.400 96.600 21.200 100.400 ;
        RECT 26.800 96.600 27.600 100.400 ;
        RECT 31.600 96.600 32.400 100.400 ;
        RECT 38.000 96.600 38.800 100.400 ;
        RECT 44.400 96.600 45.200 100.400 ;
        RECT 52.400 96.600 53.200 100.400 ;
        RECT 57.200 95.400 58.000 100.400 ;
        RECT 62.400 95.000 63.200 100.400 ;
        RECT 65.200 95.800 66.000 100.400 ;
        RECT 68.400 95.800 69.200 100.400 ;
        RECT 73.200 96.000 74.000 100.400 ;
        RECT 78.800 97.800 79.600 100.400 ;
        RECT 82.000 97.800 83.000 100.400 ;
        RECT 87.600 95.800 88.400 100.400 ;
        RECT 90.800 97.800 91.600 100.400 ;
        RECT 95.600 95.800 96.400 100.400 ;
        RECT 98.800 95.800 99.600 100.400 ;
        RECT 100.400 93.800 101.200 100.400 ;
        RECT 110.000 96.600 110.800 100.400 ;
        RECT 119.600 95.800 120.400 100.400 ;
        RECT 122.800 95.800 123.600 100.400 ;
        RECT 125.600 95.000 126.400 100.400 ;
        RECT 130.800 95.400 131.600 100.400 ;
        RECT 135.600 96.600 136.400 100.400 ;
        RECT 143.600 96.600 144.400 100.400 ;
        RECT 146.800 97.800 147.600 100.400 ;
        RECT 150.000 97.800 150.800 100.400 ;
        RECT 153.200 95.800 154.000 100.400 ;
        RECT 158.600 97.800 159.600 100.400 ;
        RECT 162.000 97.800 162.800 100.400 ;
        RECT 167.600 96.000 168.400 100.400 ;
        RECT 170.800 95.800 171.600 100.400 ;
        RECT 175.600 97.800 176.400 100.400 ;
        RECT 182.000 95.800 182.800 100.400 ;
        RECT 193.200 97.800 194.000 100.400 ;
        RECT 196.400 97.800 197.200 100.400 ;
        RECT 206.000 95.800 206.800 100.400 ;
        RECT 210.800 95.800 211.600 100.400 ;
        RECT 217.200 96.600 218.000 100.400 ;
        RECT 222.000 97.800 222.800 100.400 ;
        RECT 227.800 96.000 228.600 100.400 ;
        RECT 233.200 96.400 234.200 100.400 ;
        RECT 239.400 99.800 240.200 100.400 ;
        RECT 239.400 96.400 240.400 99.800 ;
        RECT 246.000 96.600 246.800 100.400 ;
        RECT 254.000 97.800 254.800 100.400 ;
        RECT 260.400 95.800 261.200 100.400 ;
        RECT 271.600 97.800 272.400 100.400 ;
        RECT 274.800 97.800 275.600 100.400 ;
        RECT 284.400 95.800 285.200 100.400 ;
        RECT 290.800 95.800 291.600 100.400 ;
        RECT 294.000 95.800 294.800 100.400 ;
        RECT 297.200 96.600 298.000 100.400 ;
        RECT 302.000 95.800 302.800 100.400 ;
        RECT 306.800 97.800 307.600 100.400 ;
        RECT 313.200 95.800 314.000 100.400 ;
        RECT 324.400 97.800 325.200 100.400 ;
        RECT 327.600 97.800 328.400 100.400 ;
        RECT 337.200 95.800 338.000 100.400 ;
        RECT 342.000 97.800 342.800 100.400 ;
        RECT 348.400 95.800 349.200 100.400 ;
        RECT 358.000 97.800 358.800 100.400 ;
        RECT 361.200 97.800 362.000 100.400 ;
        RECT 372.400 95.800 373.200 100.400 ;
        RECT 378.800 97.800 379.600 100.400 ;
        RECT 382.000 96.600 382.800 100.400 ;
        RECT 386.800 95.800 387.600 100.400 ;
        RECT 393.200 96.600 394.000 100.400 ;
        RECT 398.000 95.800 398.800 100.400 ;
        RECT 407.600 97.800 408.400 100.400 ;
        RECT 414.000 95.800 414.800 100.400 ;
        RECT 425.200 97.800 426.000 100.400 ;
        RECT 428.400 97.800 429.200 100.400 ;
        RECT 438.000 95.800 438.800 100.400 ;
        RECT 442.800 95.800 443.600 100.400 ;
        RECT 450.800 96.600 451.600 100.400 ;
        RECT 457.200 96.600 458.000 100.400 ;
        RECT 462.000 96.600 462.800 100.400 ;
        RECT 466.800 97.800 467.600 100.400 ;
        RECT 473.200 95.800 474.000 100.400 ;
        RECT 484.400 97.800 485.200 100.400 ;
        RECT 487.600 97.800 488.400 100.400 ;
        RECT 497.200 95.800 498.000 100.400 ;
        RECT 503.600 96.600 504.400 100.400 ;
        RECT 508.400 95.800 509.200 100.400 ;
        RECT 516.400 95.800 517.200 100.400 ;
        RECT 518.000 97.800 518.800 100.400 ;
        RECT 522.800 96.600 523.600 100.400 ;
        RECT 530.800 96.600 531.600 100.400 ;
        RECT 535.600 97.800 536.400 100.400 ;
        RECT 540.400 96.600 541.200 100.400 ;
        RECT 546.800 96.600 547.600 100.400 ;
        RECT 551.600 97.800 552.400 100.400 ;
        RECT 556.400 96.600 557.200 100.400 ;
        RECT 562.800 96.600 563.600 100.400 ;
        RECT 567.200 95.000 568.000 100.400 ;
        RECT 572.400 95.400 573.200 100.400 ;
        RECT 582.000 97.800 582.800 100.400 ;
        RECT 585.200 96.000 586.000 100.400 ;
        RECT 590.800 97.800 591.600 100.400 ;
        RECT 594.000 97.800 595.000 100.400 ;
        RECT 599.600 95.800 600.400 100.400 ;
        RECT 604.400 95.400 605.200 100.400 ;
        RECT 609.600 95.000 610.400 100.400 ;
        RECT 615.600 96.600 616.400 100.400 ;
        RECT 620.400 96.600 621.200 100.400 ;
        RECT 628.400 96.600 629.200 100.400 ;
        RECT 633.200 95.800 634.000 100.400 ;
        RECT 636.400 95.800 637.200 100.400 ;
        RECT 639.600 96.600 640.400 100.400 ;
        RECT 646.000 96.600 646.800 100.400 ;
        RECT 652.400 96.000 653.200 100.400 ;
        RECT 658.000 97.800 658.800 100.400 ;
        RECT 661.200 97.800 662.200 100.400 ;
        RECT 666.800 95.800 667.600 100.400 ;
        RECT 671.600 95.800 672.400 100.400 ;
        RECT 677.000 97.800 678.000 100.400 ;
        RECT 680.400 97.800 681.200 100.400 ;
        RECT 686.000 96.000 686.800 100.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 8.200 61.600 9.200 64.200 ;
        RECT 11.600 61.600 12.400 64.200 ;
        RECT 17.200 61.600 18.000 66.000 ;
        RECT 22.000 61.600 22.800 65.400 ;
        RECT 30.000 61.600 30.800 65.400 ;
        RECT 34.800 61.600 35.600 66.600 ;
        RECT 40.000 61.600 40.800 67.000 ;
        RECT 46.000 61.600 46.800 65.400 ;
        RECT 50.400 61.600 51.200 67.000 ;
        RECT 55.600 61.600 56.400 66.600 ;
        RECT 60.000 61.600 60.800 67.000 ;
        RECT 65.200 61.600 66.000 66.600 ;
        RECT 70.000 61.600 70.800 66.200 ;
        RECT 75.400 61.600 76.400 64.200 ;
        RECT 78.800 61.600 79.600 64.200 ;
        RECT 84.400 61.600 85.200 66.000 ;
        RECT 87.600 61.600 88.400 64.200 ;
        RECT 90.800 61.600 91.600 66.200 ;
        RECT 97.200 61.600 98.000 66.200 ;
        RECT 102.600 61.600 103.600 64.200 ;
        RECT 106.000 61.600 106.800 64.200 ;
        RECT 111.600 61.600 112.400 66.000 ;
        RECT 122.800 61.600 123.600 65.400 ;
        RECT 127.600 61.600 128.400 65.400 ;
        RECT 132.400 61.600 133.200 64.200 ;
        RECT 137.200 61.600 138.000 65.400 ;
        RECT 142.000 61.600 142.800 68.200 ;
        RECT 150.000 61.600 150.800 65.400 ;
        RECT 156.400 61.600 157.200 65.400 ;
        RECT 162.800 61.600 163.600 65.400 ;
        RECT 169.200 61.600 170.000 65.400 ;
        RECT 175.600 61.600 176.400 66.200 ;
        RECT 178.800 61.600 179.600 66.200 ;
        RECT 180.400 61.600 181.200 66.200 ;
        RECT 185.200 61.600 186.000 66.200 ;
        RECT 191.600 61.600 192.400 64.200 ;
        RECT 194.800 61.600 195.800 65.600 ;
        RECT 201.000 62.200 202.000 65.600 ;
        RECT 201.000 61.600 201.800 62.200 ;
        RECT 204.400 61.600 205.200 66.200 ;
        RECT 207.600 61.600 208.400 66.200 ;
        RECT 210.800 61.600 211.600 66.200 ;
        RECT 214.000 61.600 214.800 66.200 ;
        RECT 217.200 61.600 218.000 66.200 ;
        RECT 218.800 61.600 219.600 66.200 ;
        RECT 222.000 61.600 222.800 66.200 ;
        RECT 225.200 61.600 226.000 66.200 ;
        RECT 228.400 61.600 229.200 66.200 ;
        RECT 234.800 61.600 235.600 66.200 ;
        RECT 239.600 61.600 240.400 66.200 ;
        RECT 249.200 61.600 250.000 64.200 ;
        RECT 252.400 61.600 253.200 64.200 ;
        RECT 263.600 61.600 264.400 66.200 ;
        RECT 270.000 61.600 270.800 64.200 ;
        RECT 276.400 61.600 277.200 66.200 ;
        RECT 279.600 61.600 280.400 66.200 ;
        RECT 282.800 61.600 283.600 66.200 ;
        RECT 286.000 61.600 286.800 66.200 ;
        RECT 289.200 61.600 290.000 66.200 ;
        RECT 294.000 61.600 294.800 66.200 ;
        RECT 297.200 61.600 298.000 65.400 ;
        RECT 305.200 61.600 306.000 66.200 ;
        RECT 314.800 61.600 315.600 64.200 ;
        RECT 318.000 61.600 318.800 64.200 ;
        RECT 329.200 61.600 330.000 66.200 ;
        RECT 335.600 61.600 336.400 64.200 ;
        RECT 340.400 61.600 341.200 66.200 ;
        RECT 350.000 61.600 350.800 64.200 ;
        RECT 353.200 61.600 354.000 64.200 ;
        RECT 364.400 61.600 365.200 66.200 ;
        RECT 370.800 61.600 371.600 64.200 ;
        RECT 372.400 61.600 373.200 66.200 ;
        RECT 375.600 61.600 376.400 66.200 ;
        RECT 378.800 61.600 379.600 66.200 ;
        RECT 382.000 61.600 382.800 66.200 ;
        RECT 385.200 61.600 386.000 66.200 ;
        RECT 386.800 61.600 387.600 64.200 ;
        RECT 391.600 61.600 392.400 65.400 ;
        RECT 399.600 61.600 400.400 66.200 ;
        RECT 401.200 61.600 402.000 66.200 ;
        RECT 410.800 61.600 411.600 64.200 ;
        RECT 417.200 61.600 418.000 66.200 ;
        RECT 428.400 61.600 429.200 64.200 ;
        RECT 431.600 61.600 432.400 64.200 ;
        RECT 441.200 61.600 442.000 66.200 ;
        RECT 449.200 61.600 450.000 66.200 ;
        RECT 454.000 61.600 454.800 65.400 ;
        RECT 457.200 61.600 458.000 66.200 ;
        RECT 460.400 61.600 461.200 66.200 ;
        RECT 463.600 61.600 464.400 66.200 ;
        RECT 468.400 61.600 469.200 66.200 ;
        RECT 478.000 61.600 478.800 64.200 ;
        RECT 481.200 61.600 482.000 64.200 ;
        RECT 492.400 61.600 493.200 66.200 ;
        RECT 498.800 61.600 499.600 64.200 ;
        RECT 502.000 61.600 502.800 64.200 ;
        RECT 503.600 61.600 504.400 64.200 ;
        RECT 508.400 61.600 509.200 65.400 ;
        RECT 516.400 61.600 517.200 65.400 ;
        RECT 519.600 61.600 520.400 66.200 ;
        RECT 522.800 61.600 523.600 66.200 ;
        RECT 526.000 61.600 526.800 66.200 ;
        RECT 529.200 61.600 530.000 66.200 ;
        RECT 532.400 61.600 533.200 66.200 ;
        RECT 535.600 61.600 536.400 66.200 ;
        RECT 541.000 61.600 542.000 64.200 ;
        RECT 544.400 61.600 545.200 64.200 ;
        RECT 550.000 61.600 550.800 66.000 ;
        RECT 558.000 61.600 558.800 68.200 ;
        RECT 561.200 61.600 562.000 65.400 ;
        RECT 569.200 61.600 570.000 65.400 ;
        RECT 580.400 61.600 581.200 65.400 ;
        RECT 588.400 61.600 589.200 68.200 ;
        RECT 591.600 61.600 592.400 66.000 ;
        RECT 597.200 61.600 598.000 64.200 ;
        RECT 600.400 61.600 601.400 64.200 ;
        RECT 606.000 61.600 606.800 66.200 ;
        RECT 614.000 61.600 614.800 68.200 ;
        RECT 617.200 61.600 618.000 65.400 ;
        RECT 626.800 61.600 627.600 68.200 ;
        RECT 630.000 61.600 630.800 66.600 ;
        RECT 635.200 61.600 636.000 67.000 ;
        RECT 639.600 61.600 640.400 65.400 ;
        RECT 646.000 61.600 646.800 66.000 ;
        RECT 651.600 61.600 652.400 64.200 ;
        RECT 654.800 61.600 655.800 64.200 ;
        RECT 660.400 61.600 661.200 66.200 ;
        RECT 666.800 61.600 667.600 65.400 ;
        RECT 671.600 61.600 672.400 64.200 ;
        RECT 673.200 61.600 674.000 66.200 ;
        RECT 676.400 61.600 677.200 66.200 ;
        RECT 679.600 61.600 680.400 66.200 ;
        RECT 682.800 61.600 683.600 66.200 ;
        RECT 686.000 61.600 686.800 66.200 ;
        RECT 0.400 60.400 689.200 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 8.200 57.800 9.200 60.400 ;
        RECT 11.600 57.800 12.400 60.400 ;
        RECT 17.200 56.000 18.000 60.400 ;
        RECT 22.000 56.600 22.800 60.400 ;
        RECT 30.000 56.600 30.800 60.400 ;
        RECT 36.400 55.800 37.200 60.400 ;
        RECT 38.000 55.800 38.800 60.400 ;
        RECT 44.000 55.000 44.800 60.400 ;
        RECT 49.200 55.400 50.000 60.400 ;
        RECT 54.000 56.600 54.800 60.400 ;
        RECT 62.000 56.600 62.800 60.400 ;
        RECT 66.800 55.800 67.600 60.400 ;
        RECT 72.200 57.800 73.200 60.400 ;
        RECT 75.600 57.800 76.400 60.400 ;
        RECT 81.200 56.000 82.000 60.400 ;
        RECT 84.400 55.800 85.200 60.400 ;
        RECT 92.400 55.800 93.200 60.400 ;
        RECT 95.600 55.400 96.400 60.400 ;
        RECT 100.800 55.000 101.600 60.400 ;
        RECT 104.800 55.000 105.600 60.400 ;
        RECT 110.000 55.400 110.800 60.400 ;
        RECT 119.600 56.600 120.400 60.400 ;
        RECT 126.000 56.600 126.800 60.400 ;
        RECT 132.400 56.600 133.200 60.400 ;
        RECT 138.800 55.400 139.600 60.400 ;
        RECT 144.000 55.000 144.800 60.400 ;
        RECT 146.800 57.800 147.600 60.400 ;
        RECT 151.200 55.000 152.000 60.400 ;
        RECT 156.400 55.400 157.200 60.400 ;
        RECT 159.600 57.800 160.400 60.400 ;
        RECT 164.400 56.600 165.200 60.400 ;
        RECT 169.200 53.800 170.000 60.400 ;
        RECT 175.600 57.800 176.400 60.400 ;
        RECT 182.000 55.800 182.800 60.400 ;
        RECT 193.200 57.800 194.000 60.400 ;
        RECT 196.400 57.800 197.200 60.400 ;
        RECT 206.000 55.800 206.800 60.400 ;
        RECT 210.800 55.800 211.600 60.400 ;
        RECT 214.000 55.800 214.800 60.400 ;
        RECT 220.400 55.800 221.200 60.400 ;
        RECT 230.000 57.800 230.800 60.400 ;
        RECT 233.200 57.800 234.000 60.400 ;
        RECT 244.400 55.800 245.200 60.400 ;
        RECT 250.800 57.800 251.600 60.400 ;
        RECT 255.600 56.600 256.400 60.400 ;
        RECT 266.800 55.800 267.600 60.400 ;
        RECT 276.400 57.800 277.200 60.400 ;
        RECT 279.600 57.800 280.400 60.400 ;
        RECT 290.800 55.800 291.600 60.400 ;
        RECT 297.200 57.800 298.000 60.400 ;
        RECT 302.000 55.800 302.800 60.400 ;
        RECT 306.800 56.600 307.600 60.400 ;
        RECT 310.000 55.800 310.800 60.400 ;
        RECT 314.800 57.800 315.600 60.400 ;
        RECT 321.200 55.800 322.000 60.400 ;
        RECT 332.400 57.800 333.200 60.400 ;
        RECT 335.600 57.800 336.400 60.400 ;
        RECT 345.200 55.800 346.000 60.400 ;
        RECT 350.000 55.800 350.800 60.400 ;
        RECT 353.200 55.800 354.000 60.400 ;
        RECT 356.400 55.800 357.200 60.400 ;
        RECT 358.000 57.800 358.800 60.400 ;
        RECT 364.400 55.800 365.200 60.400 ;
        RECT 375.600 57.800 376.400 60.400 ;
        RECT 378.800 57.800 379.600 60.400 ;
        RECT 388.400 55.800 389.200 60.400 ;
        RECT 393.200 55.800 394.000 60.400 ;
        RECT 398.000 57.800 398.800 60.400 ;
        RECT 404.400 55.800 405.200 60.400 ;
        RECT 415.600 57.800 416.400 60.400 ;
        RECT 418.800 57.800 419.600 60.400 ;
        RECT 428.400 55.800 429.200 60.400 ;
        RECT 441.200 55.800 442.000 60.400 ;
        RECT 442.800 57.800 443.600 60.400 ;
        RECT 446.000 56.200 446.800 60.400 ;
        RECT 449.200 55.800 450.000 60.400 ;
        RECT 454.000 55.800 454.800 60.400 ;
        RECT 462.000 55.800 462.800 60.400 ;
        RECT 471.600 57.800 472.400 60.400 ;
        RECT 474.800 57.800 475.600 60.400 ;
        RECT 486.000 55.800 486.800 60.400 ;
        RECT 492.400 57.800 493.200 60.400 ;
        RECT 497.200 56.600 498.000 60.400 ;
        RECT 503.600 56.600 504.400 60.400 ;
        RECT 510.000 55.800 510.800 60.400 ;
        RECT 514.800 56.600 515.600 60.400 ;
        RECT 518.000 55.800 518.800 60.400 ;
        RECT 521.200 55.800 522.000 60.400 ;
        RECT 524.400 55.800 525.200 60.400 ;
        RECT 530.800 56.600 531.600 60.400 ;
        RECT 538.800 56.600 539.600 60.400 ;
        RECT 543.200 55.000 544.000 60.400 ;
        RECT 548.400 55.400 549.200 60.400 ;
        RECT 553.200 56.600 554.000 60.400 ;
        RECT 558.000 55.800 558.800 60.400 ;
        RECT 566.000 56.600 566.800 60.400 ;
        RECT 575.600 56.400 576.600 60.400 ;
        RECT 581.800 59.800 582.600 60.400 ;
        RECT 581.800 56.400 582.800 59.800 ;
        RECT 588.400 55.800 589.200 60.400 ;
        RECT 591.200 55.000 592.000 60.400 ;
        RECT 596.400 55.400 597.200 60.400 ;
        RECT 601.200 56.000 602.000 60.400 ;
        RECT 606.800 57.800 607.600 60.400 ;
        RECT 610.000 57.800 611.000 60.400 ;
        RECT 615.600 55.800 616.400 60.400 ;
        RECT 620.400 55.400 621.200 60.400 ;
        RECT 625.600 55.000 626.400 60.400 ;
        RECT 628.400 55.800 629.200 60.400 ;
        RECT 631.600 55.800 632.400 60.400 ;
        RECT 636.400 55.400 637.200 60.400 ;
        RECT 641.600 55.000 642.400 60.400 ;
        RECT 647.600 56.600 648.400 60.400 ;
        RECT 654.000 56.600 654.800 60.400 ;
        RECT 658.400 55.000 659.200 60.400 ;
        RECT 663.600 55.400 664.400 60.400 ;
        RECT 668.400 55.400 669.200 60.400 ;
        RECT 673.600 55.000 674.400 60.400 ;
        RECT 678.000 56.600 678.800 60.400 ;
        RECT 686.000 56.600 686.800 60.400 ;
        RECT 4.400 21.600 5.200 26.200 ;
        RECT 14.000 21.600 14.800 24.200 ;
        RECT 17.200 21.600 18.000 24.200 ;
        RECT 28.400 21.600 29.200 26.200 ;
        RECT 34.800 21.600 35.600 24.200 ;
        RECT 36.400 21.600 37.200 24.200 ;
        RECT 41.200 21.600 42.000 25.400 ;
        RECT 49.200 21.600 50.000 25.400 ;
        RECT 54.000 21.600 54.800 25.400 ;
        RECT 60.400 21.600 61.200 25.400 ;
        RECT 65.200 21.600 66.000 26.200 ;
        RECT 68.400 21.600 69.200 26.200 ;
        RECT 71.600 21.600 72.400 26.200 ;
        RECT 74.800 21.600 75.600 26.200 ;
        RECT 78.000 21.600 78.800 26.200 ;
        RECT 79.600 21.600 80.400 26.200 ;
        RECT 82.800 21.600 83.600 26.200 ;
        RECT 86.000 21.600 86.800 26.200 ;
        RECT 89.200 21.600 90.000 26.200 ;
        RECT 92.400 21.600 93.200 26.200 ;
        RECT 97.200 21.600 98.000 25.400 ;
        RECT 103.600 21.600 104.400 25.400 ;
        RECT 110.000 21.600 110.800 25.400 ;
        RECT 119.600 21.600 120.400 26.200 ;
        RECT 125.000 21.600 126.000 24.200 ;
        RECT 128.400 21.600 129.200 24.200 ;
        RECT 134.000 21.600 134.800 26.000 ;
        RECT 138.800 21.600 139.600 25.400 ;
        RECT 146.800 21.600 147.600 26.200 ;
        RECT 151.600 21.600 152.400 25.400 ;
        RECT 156.400 21.600 157.200 26.200 ;
        RECT 161.800 21.600 162.800 24.200 ;
        RECT 165.200 21.600 166.000 24.200 ;
        RECT 170.800 21.600 171.600 26.000 ;
        RECT 174.000 21.600 174.800 24.200 ;
        RECT 177.200 21.600 178.000 24.200 ;
        RECT 180.400 21.600 181.200 24.200 ;
        RECT 182.000 21.600 182.800 24.200 ;
        RECT 185.200 21.600 186.000 24.200 ;
        RECT 188.400 22.200 189.400 25.600 ;
        RECT 188.600 21.600 189.400 22.200 ;
        RECT 194.600 21.600 195.600 25.600 ;
        RECT 198.000 21.600 198.800 24.200 ;
        RECT 204.400 21.600 205.200 26.200 ;
        RECT 215.600 21.600 216.400 24.200 ;
        RECT 218.800 21.600 219.600 24.200 ;
        RECT 228.400 21.600 229.200 26.200 ;
        RECT 236.400 21.600 237.200 26.200 ;
        RECT 246.000 21.600 246.800 24.200 ;
        RECT 249.200 21.600 250.000 24.200 ;
        RECT 260.400 21.600 261.200 26.200 ;
        RECT 266.800 21.600 267.600 24.200 ;
        RECT 274.800 21.600 275.600 25.400 ;
        RECT 282.800 21.600 283.600 26.200 ;
        RECT 284.400 21.600 285.200 26.200 ;
        RECT 289.200 21.600 290.000 26.200 ;
        RECT 292.400 21.600 293.200 26.200 ;
        RECT 295.600 21.600 296.400 26.200 ;
        RECT 298.800 21.600 299.600 26.200 ;
        RECT 302.000 21.600 302.800 26.200 ;
        RECT 305.200 21.600 306.000 25.400 ;
        RECT 311.600 21.600 312.400 24.200 ;
        RECT 313.200 21.600 314.000 24.200 ;
        RECT 319.600 21.600 320.400 26.200 ;
        RECT 330.800 21.600 331.600 24.200 ;
        RECT 334.000 21.600 334.800 24.200 ;
        RECT 343.600 21.600 344.400 26.200 ;
        RECT 348.400 21.600 349.200 26.200 ;
        RECT 351.600 21.600 352.400 26.200 ;
        RECT 354.800 21.600 355.600 26.200 ;
        RECT 358.000 21.600 358.800 26.200 ;
        RECT 361.200 21.600 362.000 26.200 ;
        RECT 362.800 21.600 363.600 24.200 ;
        RECT 367.600 21.600 368.400 25.400 ;
        RECT 375.600 21.600 376.400 26.200 ;
        RECT 385.200 21.600 386.000 24.200 ;
        RECT 388.400 21.600 389.200 24.200 ;
        RECT 399.600 21.600 400.400 26.200 ;
        RECT 406.000 21.600 406.800 24.200 ;
        RECT 407.600 21.600 408.400 24.200 ;
        RECT 414.000 21.600 414.800 25.400 ;
        RECT 425.200 21.600 426.000 25.400 ;
        RECT 430.000 21.600 430.800 24.200 ;
        RECT 434.800 21.600 435.600 26.200 ;
        RECT 444.400 21.600 445.200 24.200 ;
        RECT 447.600 21.600 448.400 24.200 ;
        RECT 458.800 21.600 459.600 26.200 ;
        RECT 465.200 21.600 466.000 24.200 ;
        RECT 468.400 21.600 469.200 25.400 ;
        RECT 476.400 21.600 477.200 25.400 ;
        RECT 482.800 21.600 483.600 25.400 ;
        RECT 489.200 21.600 490.000 25.400 ;
        RECT 494.000 21.600 494.800 24.200 ;
        RECT 495.600 21.600 496.400 24.200 ;
        RECT 502.000 21.600 502.800 26.200 ;
        RECT 513.200 21.600 514.000 24.200 ;
        RECT 516.400 21.600 517.200 24.200 ;
        RECT 526.000 21.600 526.800 26.200 ;
        RECT 534.000 21.600 534.800 25.400 ;
        RECT 538.800 21.600 539.600 25.400 ;
        RECT 546.800 21.600 547.600 25.400 ;
        RECT 551.600 21.600 552.400 25.400 ;
        RECT 559.600 21.600 560.400 26.200 ;
        RECT 562.400 21.600 563.200 27.000 ;
        RECT 567.600 21.600 568.400 26.600 ;
        RECT 577.200 21.600 578.000 26.000 ;
        RECT 582.800 21.600 583.600 24.200 ;
        RECT 586.000 21.600 587.000 24.200 ;
        RECT 591.600 21.600 592.400 26.200 ;
        RECT 596.400 21.600 597.200 24.200 ;
        RECT 599.600 21.600 600.400 26.000 ;
        RECT 605.200 21.600 606.000 24.200 ;
        RECT 608.400 21.600 609.400 24.200 ;
        RECT 614.000 21.600 614.800 26.200 ;
        RECT 618.800 21.600 619.600 25.400 ;
        RECT 626.800 21.600 627.600 25.400 ;
        RECT 631.200 21.600 632.000 27.000 ;
        RECT 636.400 21.600 637.200 26.600 ;
        RECT 641.200 21.600 642.000 26.600 ;
        RECT 646.400 21.600 647.200 27.000 ;
        RECT 650.800 21.600 651.600 25.400 ;
        RECT 658.800 21.600 659.600 25.400 ;
        RECT 663.600 21.600 664.400 25.400 ;
        RECT 671.600 21.600 672.400 25.400 ;
        RECT 676.400 21.600 677.400 25.600 ;
        RECT 682.600 22.200 683.600 25.600 ;
        RECT 682.600 21.600 683.400 22.200 ;
        RECT 0.400 20.400 689.200 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 17.200 17.800 18.000 20.400 ;
        RECT 20.400 17.800 21.200 20.400 ;
        RECT 31.600 15.800 32.400 20.400 ;
        RECT 38.000 17.800 38.800 20.400 ;
        RECT 41.200 15.800 42.000 20.400 ;
        RECT 44.400 17.800 45.200 20.400 ;
        RECT 47.600 17.800 48.400 20.400 ;
        RECT 54.000 15.800 54.800 20.400 ;
        RECT 65.200 17.800 66.000 20.400 ;
        RECT 68.400 17.800 69.200 20.400 ;
        RECT 78.000 15.800 78.800 20.400 ;
        RECT 82.800 17.800 83.600 20.400 ;
        RECT 89.200 15.800 90.000 20.400 ;
        RECT 100.400 17.800 101.200 20.400 ;
        RECT 103.600 17.800 104.400 20.400 ;
        RECT 113.200 15.800 114.000 20.400 ;
        RECT 124.400 15.800 125.200 20.400 ;
        RECT 129.800 17.800 130.800 20.400 ;
        RECT 133.200 17.800 134.000 20.400 ;
        RECT 138.800 16.000 139.600 20.400 ;
        RECT 142.000 17.800 142.800 20.400 ;
        RECT 145.200 17.800 146.000 20.400 ;
        RECT 148.600 19.800 149.400 20.400 ;
        RECT 148.400 16.400 149.400 19.800 ;
        RECT 154.600 16.400 155.600 20.400 ;
        RECT 159.600 17.800 160.400 20.400 ;
        RECT 161.200 17.800 162.000 20.400 ;
        RECT 164.400 17.800 165.200 20.400 ;
        RECT 166.000 17.800 166.800 20.400 ;
        RECT 172.400 15.800 173.200 20.400 ;
        RECT 183.600 17.800 184.400 20.400 ;
        RECT 186.800 17.800 187.600 20.400 ;
        RECT 196.400 15.800 197.200 20.400 ;
        RECT 204.400 15.800 205.200 20.400 ;
        RECT 214.000 17.800 214.800 20.400 ;
        RECT 217.200 17.800 218.000 20.400 ;
        RECT 228.400 15.800 229.200 20.400 ;
        RECT 234.800 17.800 235.600 20.400 ;
        RECT 236.400 17.800 237.200 20.400 ;
        RECT 241.200 15.800 242.000 20.400 ;
        RECT 247.600 16.600 248.400 20.400 ;
        RECT 250.800 15.800 251.600 20.400 ;
        RECT 257.200 15.800 258.000 20.400 ;
        RECT 260.400 17.800 261.200 20.400 ;
        RECT 270.000 15.800 270.800 20.400 ;
        RECT 273.200 17.800 274.000 20.400 ;
        RECT 278.000 16.600 278.800 20.400 ;
        RECT 282.800 17.800 283.600 20.400 ;
        RECT 289.200 15.800 290.000 20.400 ;
        RECT 300.400 17.800 301.200 20.400 ;
        RECT 303.600 17.800 304.400 20.400 ;
        RECT 313.200 15.800 314.000 20.400 ;
        RECT 319.600 15.800 320.400 20.400 ;
        RECT 322.800 15.800 323.600 20.400 ;
        RECT 326.000 15.800 326.800 20.400 ;
        RECT 329.200 15.800 330.000 20.400 ;
        RECT 332.400 15.800 333.200 20.400 ;
        RECT 335.600 17.800 336.400 20.400 ;
        RECT 342.000 15.800 342.800 20.400 ;
        RECT 353.200 17.800 354.000 20.400 ;
        RECT 356.400 17.800 357.200 20.400 ;
        RECT 366.000 15.800 366.800 20.400 ;
        RECT 372.400 15.800 373.200 20.400 ;
        RECT 377.200 15.800 378.000 20.400 ;
        RECT 383.600 15.800 384.400 20.400 ;
        RECT 393.200 17.800 394.000 20.400 ;
        RECT 396.400 17.800 397.200 20.400 ;
        RECT 407.600 15.800 408.400 20.400 ;
        RECT 414.000 17.800 414.800 20.400 ;
        RECT 417.200 15.800 418.000 20.400 ;
        RECT 428.400 15.800 429.200 20.400 ;
        RECT 438.000 17.800 438.800 20.400 ;
        RECT 441.200 17.800 442.000 20.400 ;
        RECT 452.400 15.800 453.200 20.400 ;
        RECT 458.800 17.800 459.600 20.400 ;
        RECT 462.000 17.800 462.800 20.400 ;
        RECT 463.600 17.800 464.400 20.400 ;
        RECT 466.800 17.800 467.600 20.400 ;
        RECT 473.200 15.800 474.000 20.400 ;
        RECT 484.400 17.800 485.200 20.400 ;
        RECT 487.600 17.800 488.400 20.400 ;
        RECT 497.200 15.800 498.000 20.400 ;
        RECT 502.000 17.800 502.800 20.400 ;
        RECT 508.400 15.800 509.200 20.400 ;
        RECT 518.000 17.800 518.800 20.400 ;
        RECT 521.200 17.800 522.000 20.400 ;
        RECT 532.400 15.800 533.200 20.400 ;
        RECT 538.800 17.800 539.600 20.400 ;
        RECT 542.000 17.800 542.800 20.400 ;
        RECT 546.800 15.800 547.600 20.400 ;
        RECT 556.400 17.800 557.200 20.400 ;
        RECT 559.600 17.800 560.400 20.400 ;
        RECT 570.800 15.800 571.600 20.400 ;
        RECT 577.200 17.800 578.000 20.400 ;
        RECT 585.200 15.800 586.000 20.400 ;
        RECT 590.000 16.000 590.800 20.400 ;
        RECT 595.600 17.800 596.400 20.400 ;
        RECT 598.800 17.800 599.800 20.400 ;
        RECT 604.400 15.800 605.200 20.400 ;
        RECT 609.200 16.600 610.000 20.400 ;
        RECT 617.200 16.600 618.000 20.400 ;
        RECT 622.000 16.600 622.800 20.400 ;
        RECT 630.000 16.600 630.800 20.400 ;
        RECT 634.800 17.800 635.600 20.400 ;
        RECT 639.600 16.600 640.400 20.400 ;
        RECT 644.400 16.000 645.200 20.400 ;
        RECT 650.000 17.800 650.800 20.400 ;
        RECT 653.200 17.800 654.200 20.400 ;
        RECT 658.800 15.800 659.600 20.400 ;
        RECT 663.600 16.000 664.400 20.400 ;
        RECT 669.200 17.800 670.000 20.400 ;
        RECT 672.400 17.800 673.400 20.400 ;
        RECT 678.000 15.800 678.800 20.400 ;
        RECT 684.400 16.600 685.200 20.400 ;
      LAYER via1 ;
        RECT 263.800 500.600 264.600 501.400 ;
        RECT 265.200 500.600 266.000 501.400 ;
        RECT 266.600 500.600 267.400 501.400 ;
        RECT 572.600 500.600 573.400 501.400 ;
        RECT 574.000 500.600 574.800 501.400 ;
        RECT 575.400 500.600 576.200 501.400 ;
        RECT 263.800 460.600 264.600 461.400 ;
        RECT 265.200 460.600 266.000 461.400 ;
        RECT 266.600 460.600 267.400 461.400 ;
        RECT 572.600 460.600 573.400 461.400 ;
        RECT 574.000 460.600 574.800 461.400 ;
        RECT 575.400 460.600 576.200 461.400 ;
        RECT 263.800 420.600 264.600 421.400 ;
        RECT 265.200 420.600 266.000 421.400 ;
        RECT 266.600 420.600 267.400 421.400 ;
        RECT 572.600 420.600 573.400 421.400 ;
        RECT 574.000 420.600 574.800 421.400 ;
        RECT 575.400 420.600 576.200 421.400 ;
        RECT 263.800 380.600 264.600 381.400 ;
        RECT 265.200 380.600 266.000 381.400 ;
        RECT 266.600 380.600 267.400 381.400 ;
        RECT 572.600 380.600 573.400 381.400 ;
        RECT 574.000 380.600 574.800 381.400 ;
        RECT 575.400 380.600 576.200 381.400 ;
        RECT 263.800 340.600 264.600 341.400 ;
        RECT 265.200 340.600 266.000 341.400 ;
        RECT 266.600 340.600 267.400 341.400 ;
        RECT 572.600 340.600 573.400 341.400 ;
        RECT 574.000 340.600 574.800 341.400 ;
        RECT 575.400 340.600 576.200 341.400 ;
        RECT 354.800 303.600 355.600 304.400 ;
        RECT 263.800 300.600 264.600 301.400 ;
        RECT 265.200 300.600 266.000 301.400 ;
        RECT 266.600 300.600 267.400 301.400 ;
        RECT 572.600 300.600 573.400 301.400 ;
        RECT 574.000 300.600 574.800 301.400 ;
        RECT 575.400 300.600 576.200 301.400 ;
        RECT 329.200 267.600 330.000 268.400 ;
        RECT 329.200 263.600 330.000 264.400 ;
        RECT 263.800 260.600 264.600 261.400 ;
        RECT 265.200 260.600 266.000 261.400 ;
        RECT 266.600 260.600 267.400 261.400 ;
        RECT 572.600 260.600 573.400 261.400 ;
        RECT 574.000 260.600 574.800 261.400 ;
        RECT 575.400 260.600 576.200 261.400 ;
        RECT 358.000 257.600 358.800 258.400 ;
        RECT 380.400 259.600 381.200 260.400 ;
        RECT 393.200 259.600 394.000 260.400 ;
        RECT 281.200 227.600 282.000 228.400 ;
        RECT 263.800 220.600 264.600 221.400 ;
        RECT 265.200 220.600 266.000 221.400 ;
        RECT 266.600 220.600 267.400 221.400 ;
        RECT 572.600 220.600 573.400 221.400 ;
        RECT 574.000 220.600 574.800 221.400 ;
        RECT 575.400 220.600 576.200 221.400 ;
        RECT 281.200 219.600 282.000 220.400 ;
        RECT 319.600 217.600 320.400 218.400 ;
        RECT 263.800 180.600 264.600 181.400 ;
        RECT 265.200 180.600 266.000 181.400 ;
        RECT 266.600 180.600 267.400 181.400 ;
        RECT 572.600 180.600 573.400 181.400 ;
        RECT 574.000 180.600 574.800 181.400 ;
        RECT 575.400 180.600 576.200 181.400 ;
        RECT 263.800 140.600 264.600 141.400 ;
        RECT 265.200 140.600 266.000 141.400 ;
        RECT 266.600 140.600 267.400 141.400 ;
        RECT 572.600 140.600 573.400 141.400 ;
        RECT 574.000 140.600 574.800 141.400 ;
        RECT 575.400 140.600 576.200 141.400 ;
        RECT 263.800 100.600 264.600 101.400 ;
        RECT 265.200 100.600 266.000 101.400 ;
        RECT 266.600 100.600 267.400 101.400 ;
        RECT 572.600 100.600 573.400 101.400 ;
        RECT 574.000 100.600 574.800 101.400 ;
        RECT 575.400 100.600 576.200 101.400 ;
        RECT 263.800 60.600 264.600 61.400 ;
        RECT 265.200 60.600 266.000 61.400 ;
        RECT 266.600 60.600 267.400 61.400 ;
        RECT 572.600 60.600 573.400 61.400 ;
        RECT 574.000 60.600 574.800 61.400 ;
        RECT 575.400 60.600 576.200 61.400 ;
        RECT 263.800 20.600 264.600 21.400 ;
        RECT 265.200 20.600 266.000 21.400 ;
        RECT 266.600 20.600 267.400 21.400 ;
        RECT 572.600 20.600 573.400 21.400 ;
        RECT 574.000 20.600 574.800 21.400 ;
        RECT 575.400 20.600 576.200 21.400 ;
      LAYER metal2 ;
        RECT 263.200 500.600 268.000 501.400 ;
        RECT 572.000 500.600 576.800 501.400 ;
        RECT 263.200 460.600 268.000 461.400 ;
        RECT 572.000 460.600 576.800 461.400 ;
        RECT 263.200 420.600 268.000 421.400 ;
        RECT 572.000 420.600 576.800 421.400 ;
        RECT 263.200 380.600 268.000 381.400 ;
        RECT 572.000 380.600 576.800 381.400 ;
        RECT 263.200 340.600 268.000 341.400 ;
        RECT 572.000 340.600 576.800 341.400 ;
        RECT 351.600 311.600 352.400 312.400 ;
        RECT 351.700 304.400 352.300 311.600 ;
        RECT 351.600 303.600 352.400 304.400 ;
        RECT 354.800 303.600 355.600 304.400 ;
        RECT 263.200 300.600 268.000 301.400 ;
        RECT 572.000 300.600 576.800 301.400 ;
        RECT 380.400 271.600 381.200 272.400 ;
        RECT 329.200 267.600 330.000 268.400 ;
        RECT 329.300 264.400 329.900 267.600 ;
        RECT 329.200 263.600 330.000 264.400 ;
        RECT 263.200 260.600 268.000 261.400 ;
        RECT 380.500 260.400 381.100 271.600 ;
        RECT 572.000 260.600 576.800 261.400 ;
        RECT 380.400 259.600 381.200 260.400 ;
        RECT 393.200 259.600 394.000 260.400 ;
        RECT 358.000 257.600 358.800 258.400 ;
        RECT 358.100 252.400 358.700 257.600 ;
        RECT 393.300 256.400 393.900 259.600 ;
        RECT 393.200 255.600 394.000 256.400 ;
        RECT 358.000 251.600 358.800 252.400 ;
        RECT 281.200 227.600 282.000 228.400 ;
        RECT 263.200 220.600 268.000 221.400 ;
        RECT 281.300 220.400 281.900 227.600 ;
        RECT 343.600 223.600 344.400 224.400 ;
        RECT 281.200 219.600 282.000 220.400 ;
        RECT 319.600 217.600 320.400 218.400 ;
        RECT 319.700 214.400 320.300 217.600 ;
        RECT 343.700 214.400 344.300 223.600 ;
        RECT 572.000 220.600 576.800 221.400 ;
        RECT 319.600 213.600 320.400 214.400 ;
        RECT 343.600 213.600 344.400 214.400 ;
        RECT 263.200 180.600 268.000 181.400 ;
        RECT 572.000 180.600 576.800 181.400 ;
        RECT 263.200 140.600 268.000 141.400 ;
        RECT 572.000 140.600 576.800 141.400 ;
        RECT 263.200 100.600 268.000 101.400 ;
        RECT 572.000 100.600 576.800 101.400 ;
        RECT 263.200 60.600 268.000 61.400 ;
        RECT 572.000 60.600 576.800 61.400 ;
        RECT 263.200 20.600 268.000 21.400 ;
        RECT 572.000 20.600 576.800 21.400 ;
      LAYER via2 ;
        RECT 263.800 500.600 264.600 501.400 ;
        RECT 265.200 500.600 266.000 501.400 ;
        RECT 266.600 500.600 267.400 501.400 ;
        RECT 572.600 500.600 573.400 501.400 ;
        RECT 574.000 500.600 574.800 501.400 ;
        RECT 575.400 500.600 576.200 501.400 ;
        RECT 263.800 460.600 264.600 461.400 ;
        RECT 265.200 460.600 266.000 461.400 ;
        RECT 266.600 460.600 267.400 461.400 ;
        RECT 572.600 460.600 573.400 461.400 ;
        RECT 574.000 460.600 574.800 461.400 ;
        RECT 575.400 460.600 576.200 461.400 ;
        RECT 263.800 420.600 264.600 421.400 ;
        RECT 265.200 420.600 266.000 421.400 ;
        RECT 266.600 420.600 267.400 421.400 ;
        RECT 572.600 420.600 573.400 421.400 ;
        RECT 574.000 420.600 574.800 421.400 ;
        RECT 575.400 420.600 576.200 421.400 ;
        RECT 263.800 380.600 264.600 381.400 ;
        RECT 265.200 380.600 266.000 381.400 ;
        RECT 266.600 380.600 267.400 381.400 ;
        RECT 572.600 380.600 573.400 381.400 ;
        RECT 574.000 380.600 574.800 381.400 ;
        RECT 575.400 380.600 576.200 381.400 ;
        RECT 263.800 340.600 264.600 341.400 ;
        RECT 265.200 340.600 266.000 341.400 ;
        RECT 266.600 340.600 267.400 341.400 ;
        RECT 572.600 340.600 573.400 341.400 ;
        RECT 574.000 340.600 574.800 341.400 ;
        RECT 575.400 340.600 576.200 341.400 ;
        RECT 263.800 300.600 264.600 301.400 ;
        RECT 265.200 300.600 266.000 301.400 ;
        RECT 266.600 300.600 267.400 301.400 ;
        RECT 572.600 300.600 573.400 301.400 ;
        RECT 574.000 300.600 574.800 301.400 ;
        RECT 575.400 300.600 576.200 301.400 ;
        RECT 263.800 260.600 264.600 261.400 ;
        RECT 265.200 260.600 266.000 261.400 ;
        RECT 266.600 260.600 267.400 261.400 ;
        RECT 572.600 260.600 573.400 261.400 ;
        RECT 574.000 260.600 574.800 261.400 ;
        RECT 575.400 260.600 576.200 261.400 ;
        RECT 263.800 220.600 264.600 221.400 ;
        RECT 265.200 220.600 266.000 221.400 ;
        RECT 266.600 220.600 267.400 221.400 ;
        RECT 572.600 220.600 573.400 221.400 ;
        RECT 574.000 220.600 574.800 221.400 ;
        RECT 575.400 220.600 576.200 221.400 ;
        RECT 263.800 180.600 264.600 181.400 ;
        RECT 265.200 180.600 266.000 181.400 ;
        RECT 266.600 180.600 267.400 181.400 ;
        RECT 572.600 180.600 573.400 181.400 ;
        RECT 574.000 180.600 574.800 181.400 ;
        RECT 575.400 180.600 576.200 181.400 ;
        RECT 263.800 140.600 264.600 141.400 ;
        RECT 265.200 140.600 266.000 141.400 ;
        RECT 266.600 140.600 267.400 141.400 ;
        RECT 572.600 140.600 573.400 141.400 ;
        RECT 574.000 140.600 574.800 141.400 ;
        RECT 575.400 140.600 576.200 141.400 ;
        RECT 263.800 100.600 264.600 101.400 ;
        RECT 265.200 100.600 266.000 101.400 ;
        RECT 266.600 100.600 267.400 101.400 ;
        RECT 572.600 100.600 573.400 101.400 ;
        RECT 574.000 100.600 574.800 101.400 ;
        RECT 575.400 100.600 576.200 101.400 ;
        RECT 263.800 60.600 264.600 61.400 ;
        RECT 265.200 60.600 266.000 61.400 ;
        RECT 266.600 60.600 267.400 61.400 ;
        RECT 572.600 60.600 573.400 61.400 ;
        RECT 574.000 60.600 574.800 61.400 ;
        RECT 575.400 60.600 576.200 61.400 ;
        RECT 263.800 20.600 264.600 21.400 ;
        RECT 265.200 20.600 266.000 21.400 ;
        RECT 266.600 20.600 267.400 21.400 ;
        RECT 572.600 20.600 573.400 21.400 ;
        RECT 574.000 20.600 574.800 21.400 ;
        RECT 575.400 20.600 576.200 21.400 ;
      LAYER metal3 ;
        RECT 263.200 500.400 268.000 501.600 ;
        RECT 572.000 500.400 576.800 501.600 ;
        RECT 263.200 460.400 268.000 461.600 ;
        RECT 572.000 460.400 576.800 461.600 ;
        RECT 263.200 420.400 268.000 421.600 ;
        RECT 572.000 420.400 576.800 421.600 ;
        RECT 263.200 380.400 268.000 381.600 ;
        RECT 572.000 380.400 576.800 381.600 ;
        RECT 263.200 340.400 268.000 341.600 ;
        RECT 572.000 340.400 576.800 341.600 ;
        RECT 351.600 304.300 352.400 304.400 ;
        RECT 354.800 304.300 355.600 304.400 ;
        RECT 351.600 303.700 355.600 304.300 ;
        RECT 351.600 303.600 352.400 303.700 ;
        RECT 354.800 303.600 355.600 303.700 ;
        RECT 263.200 300.400 268.000 301.600 ;
        RECT 572.000 300.400 576.800 301.600 ;
        RECT 263.200 260.400 268.000 261.600 ;
        RECT 572.000 260.400 576.800 261.600 ;
        RECT 263.200 220.400 268.000 221.600 ;
        RECT 572.000 220.400 576.800 221.600 ;
        RECT 263.200 180.400 268.000 181.600 ;
        RECT 572.000 180.400 576.800 181.600 ;
        RECT 263.200 140.400 268.000 141.600 ;
        RECT 572.000 140.400 576.800 141.600 ;
        RECT 263.200 100.400 268.000 101.600 ;
        RECT 572.000 100.400 576.800 101.600 ;
        RECT 263.200 60.400 268.000 61.600 ;
        RECT 572.000 60.400 576.800 61.600 ;
        RECT 263.200 20.400 268.000 21.600 ;
        RECT 572.000 20.400 576.800 21.600 ;
      LAYER via3 ;
        RECT 263.600 500.600 264.400 501.400 ;
        RECT 265.200 500.600 266.000 501.400 ;
        RECT 266.800 500.600 267.600 501.400 ;
        RECT 572.400 500.600 573.200 501.400 ;
        RECT 574.000 500.600 574.800 501.400 ;
        RECT 575.600 500.600 576.400 501.400 ;
        RECT 263.600 460.600 264.400 461.400 ;
        RECT 265.200 460.600 266.000 461.400 ;
        RECT 266.800 460.600 267.600 461.400 ;
        RECT 572.400 460.600 573.200 461.400 ;
        RECT 574.000 460.600 574.800 461.400 ;
        RECT 575.600 460.600 576.400 461.400 ;
        RECT 263.600 420.600 264.400 421.400 ;
        RECT 265.200 420.600 266.000 421.400 ;
        RECT 266.800 420.600 267.600 421.400 ;
        RECT 572.400 420.600 573.200 421.400 ;
        RECT 574.000 420.600 574.800 421.400 ;
        RECT 575.600 420.600 576.400 421.400 ;
        RECT 263.600 380.600 264.400 381.400 ;
        RECT 265.200 380.600 266.000 381.400 ;
        RECT 266.800 380.600 267.600 381.400 ;
        RECT 572.400 380.600 573.200 381.400 ;
        RECT 574.000 380.600 574.800 381.400 ;
        RECT 575.600 380.600 576.400 381.400 ;
        RECT 263.600 340.600 264.400 341.400 ;
        RECT 265.200 340.600 266.000 341.400 ;
        RECT 266.800 340.600 267.600 341.400 ;
        RECT 572.400 340.600 573.200 341.400 ;
        RECT 574.000 340.600 574.800 341.400 ;
        RECT 575.600 340.600 576.400 341.400 ;
        RECT 263.600 300.600 264.400 301.400 ;
        RECT 265.200 300.600 266.000 301.400 ;
        RECT 266.800 300.600 267.600 301.400 ;
        RECT 572.400 300.600 573.200 301.400 ;
        RECT 574.000 300.600 574.800 301.400 ;
        RECT 575.600 300.600 576.400 301.400 ;
        RECT 263.600 260.600 264.400 261.400 ;
        RECT 265.200 260.600 266.000 261.400 ;
        RECT 266.800 260.600 267.600 261.400 ;
        RECT 572.400 260.600 573.200 261.400 ;
        RECT 574.000 260.600 574.800 261.400 ;
        RECT 575.600 260.600 576.400 261.400 ;
        RECT 263.600 220.600 264.400 221.400 ;
        RECT 265.200 220.600 266.000 221.400 ;
        RECT 266.800 220.600 267.600 221.400 ;
        RECT 572.400 220.600 573.200 221.400 ;
        RECT 574.000 220.600 574.800 221.400 ;
        RECT 575.600 220.600 576.400 221.400 ;
        RECT 263.600 180.600 264.400 181.400 ;
        RECT 265.200 180.600 266.000 181.400 ;
        RECT 266.800 180.600 267.600 181.400 ;
        RECT 572.400 180.600 573.200 181.400 ;
        RECT 574.000 180.600 574.800 181.400 ;
        RECT 575.600 180.600 576.400 181.400 ;
        RECT 263.600 140.600 264.400 141.400 ;
        RECT 265.200 140.600 266.000 141.400 ;
        RECT 266.800 140.600 267.600 141.400 ;
        RECT 572.400 140.600 573.200 141.400 ;
        RECT 574.000 140.600 574.800 141.400 ;
        RECT 575.600 140.600 576.400 141.400 ;
        RECT 263.600 100.600 264.400 101.400 ;
        RECT 265.200 100.600 266.000 101.400 ;
        RECT 266.800 100.600 267.600 101.400 ;
        RECT 572.400 100.600 573.200 101.400 ;
        RECT 574.000 100.600 574.800 101.400 ;
        RECT 575.600 100.600 576.400 101.400 ;
        RECT 263.600 60.600 264.400 61.400 ;
        RECT 265.200 60.600 266.000 61.400 ;
        RECT 266.800 60.600 267.600 61.400 ;
        RECT 572.400 60.600 573.200 61.400 ;
        RECT 574.000 60.600 574.800 61.400 ;
        RECT 575.600 60.600 576.400 61.400 ;
        RECT 263.600 20.600 264.400 21.400 ;
        RECT 265.200 20.600 266.000 21.400 ;
        RECT 266.800 20.600 267.600 21.400 ;
        RECT 572.400 20.600 573.200 21.400 ;
        RECT 574.000 20.600 574.800 21.400 ;
        RECT 575.600 20.600 576.400 21.400 ;
      LAYER metal4 ;
        RECT 263.200 -4.000 268.000 504.000 ;
        RECT 572.000 -4.000 576.800 504.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 207.400 332.400 208.200 333.200 ;
        RECT 493.800 332.400 494.600 333.200 ;
        RECT 207.400 331.600 208.400 332.400 ;
        RECT 493.800 331.600 494.800 332.400 ;
        RECT 186.600 270.300 187.600 270.400 ;
        RECT 188.400 270.300 189.200 270.400 ;
        RECT 186.600 269.700 189.200 270.300 ;
        RECT 186.600 269.600 187.600 269.700 ;
        RECT 188.400 269.600 189.200 269.700 ;
        RECT 186.600 268.800 187.400 269.600 ;
        RECT 510.000 189.600 511.000 190.400 ;
        RECT 510.200 188.800 511.000 189.600 ;
        RECT 404.600 172.400 405.400 173.200 ;
        RECT 404.400 171.600 405.400 172.400 ;
        RECT 215.400 52.400 216.200 53.200 ;
        RECT 215.400 51.600 216.400 52.400 ;
      LAYER via1 ;
        RECT 207.600 331.600 208.400 332.400 ;
        RECT 494.000 331.600 494.800 332.400 ;
        RECT 215.600 51.600 216.400 52.400 ;
      LAYER metal2 ;
        RECT 207.600 331.600 208.400 332.400 ;
        RECT 494.000 331.600 494.800 332.400 ;
        RECT 207.700 306.400 208.300 331.600 ;
        RECT 494.100 318.400 494.700 331.600 ;
        RECT 494.000 317.600 494.800 318.400 ;
        RECT 188.400 305.600 189.200 306.400 ;
        RECT 207.600 305.600 208.400 306.400 ;
        RECT 188.500 270.400 189.100 305.600 ;
        RECT 188.400 269.600 189.200 270.400 ;
        RECT 188.500 226.400 189.100 269.600 ;
        RECT 188.400 225.600 189.200 226.400 ;
        RECT 510.000 197.600 510.800 198.400 ;
        RECT 510.100 190.400 510.700 197.600 ;
        RECT 510.000 189.600 510.800 190.400 ;
        RECT 404.400 171.600 405.200 172.400 ;
        RECT 404.500 166.400 405.100 171.600 ;
        RECT 510.100 166.400 510.700 189.600 ;
        RECT 404.400 165.600 405.200 166.400 ;
        RECT 510.000 165.600 510.800 166.400 ;
        RECT 209.200 139.600 210.000 140.400 ;
        RECT 209.300 52.400 209.900 139.600 ;
        RECT 209.200 51.600 210.000 52.400 ;
        RECT 215.600 51.600 216.400 52.400 ;
        RECT 215.600 1.600 216.400 2.400 ;
        RECT 215.700 -2.300 216.300 1.600 ;
      LAYER metal3 ;
        RECT 494.000 317.600 494.800 318.400 ;
        RECT 188.400 306.300 189.200 306.400 ;
        RECT 207.600 306.300 208.400 306.400 ;
        RECT 188.400 305.700 208.400 306.300 ;
        RECT 188.400 305.600 189.200 305.700 ;
        RECT 207.600 305.600 208.400 305.700 ;
        RECT 188.400 226.300 189.200 226.400 ;
        RECT 193.200 226.300 194.000 226.400 ;
        RECT 188.400 225.700 194.000 226.300 ;
        RECT 188.400 225.600 189.200 225.700 ;
        RECT 193.200 225.600 194.000 225.700 ;
        RECT 494.000 198.300 494.800 198.400 ;
        RECT 510.000 198.300 510.800 198.400 ;
        RECT 494.000 197.700 510.800 198.300 ;
        RECT 494.000 197.600 494.800 197.700 ;
        RECT 510.000 197.600 510.800 197.700 ;
        RECT 193.200 166.300 194.000 166.400 ;
        RECT 404.400 166.300 405.200 166.400 ;
        RECT 510.000 166.300 510.800 166.400 ;
        RECT 193.200 165.700 510.800 166.300 ;
        RECT 193.200 165.600 194.000 165.700 ;
        RECT 404.400 165.600 405.200 165.700 ;
        RECT 510.000 165.600 510.800 165.700 ;
        RECT 193.200 140.300 194.000 140.400 ;
        RECT 209.200 140.300 210.000 140.400 ;
        RECT 193.200 139.700 210.000 140.300 ;
        RECT 193.200 139.600 194.000 139.700 ;
        RECT 209.200 139.600 210.000 139.700 ;
        RECT 209.200 52.300 210.000 52.400 ;
        RECT 215.600 52.300 216.400 52.400 ;
        RECT 209.200 51.700 216.400 52.300 ;
        RECT 209.200 51.600 210.000 51.700 ;
        RECT 215.600 51.600 216.400 51.700 ;
        RECT 215.600 1.600 216.400 2.400 ;
      LAYER metal4 ;
        RECT 193.000 139.400 194.200 226.600 ;
        RECT 493.800 197.400 495.000 318.600 ;
        RECT 215.400 1.400 216.600 52.600 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 257.200 386.800 258.000 388.400 ;
        RECT 492.400 386.800 493.200 388.400 ;
        RECT 402.800 373.600 403.600 375.200 ;
        RECT 236.400 306.800 237.200 308.400 ;
        RECT 289.200 306.800 290.000 308.400 ;
        RECT 383.600 266.800 384.400 268.400 ;
        RECT 260.400 134.300 261.200 135.200 ;
        RECT 265.200 134.300 266.000 134.400 ;
        RECT 260.400 133.700 266.000 134.300 ;
        RECT 260.400 133.600 261.200 133.700 ;
        RECT 265.200 133.600 266.000 133.700 ;
        RECT 463.600 66.800 464.400 68.400 ;
        RECT 356.400 53.600 357.200 55.200 ;
        RECT 329.200 13.600 330.000 15.200 ;
      LAYER via1 ;
        RECT 257.200 387.600 258.000 388.400 ;
        RECT 492.400 387.600 493.200 388.400 ;
        RECT 236.400 307.600 237.200 308.400 ;
        RECT 289.200 307.600 290.000 308.400 ;
        RECT 383.600 267.600 384.400 268.400 ;
        RECT 463.600 67.600 464.400 68.400 ;
      LAYER metal2 ;
        RECT 257.200 387.600 258.000 388.400 ;
        RECT 492.400 387.600 493.200 388.400 ;
        RECT 257.300 382.400 257.900 387.600 ;
        RECT 257.200 381.600 258.000 382.400 ;
        RECT 492.500 378.400 493.100 387.600 ;
        RECT 402.800 377.600 403.600 378.400 ;
        RECT 492.400 377.600 493.200 378.400 ;
        RECT 402.900 374.400 403.500 377.600 ;
        RECT 402.800 373.600 403.600 374.400 ;
        RECT 236.400 307.600 237.200 308.400 ;
        RECT 289.200 307.600 290.000 308.400 ;
        RECT 383.600 267.600 384.400 268.400 ;
        RECT 265.200 133.600 266.000 134.400 ;
        RECT 265.300 104.400 265.900 133.600 ;
        RECT 265.200 103.600 266.000 104.400 ;
        RECT 303.600 103.600 304.400 104.400 ;
        RECT 303.700 54.400 304.300 103.600 ;
        RECT 388.400 67.600 389.200 68.400 ;
        RECT 463.600 67.600 464.400 68.400 ;
        RECT 388.500 54.400 389.100 67.600 ;
        RECT 303.600 53.600 304.400 54.400 ;
        RECT 356.400 53.600 357.200 54.400 ;
        RECT 388.400 53.600 389.200 54.400 ;
        RECT 322.800 13.600 323.600 14.400 ;
        RECT 329.200 13.600 330.000 14.400 ;
        RECT 322.900 -2.300 323.500 13.600 ;
      LAYER metal3 ;
        RECT 257.200 381.600 258.000 382.400 ;
        RECT 402.800 378.300 403.600 378.400 ;
        RECT 492.400 378.300 493.200 378.400 ;
        RECT 402.800 377.700 493.200 378.300 ;
        RECT 402.800 377.600 403.600 377.700 ;
        RECT 492.400 377.600 493.200 377.700 ;
        RECT 343.600 374.300 344.400 374.400 ;
        RECT 402.800 374.300 403.600 374.400 ;
        RECT 343.600 373.700 403.600 374.300 ;
        RECT 343.600 373.600 344.400 373.700 ;
        RECT 402.800 373.600 403.600 373.700 ;
        RECT 236.400 308.300 237.200 308.400 ;
        RECT 257.200 308.300 258.000 308.400 ;
        RECT 276.400 308.300 277.200 308.400 ;
        RECT 289.200 308.300 290.000 308.400 ;
        RECT 343.600 308.300 344.400 308.400 ;
        RECT 236.400 307.700 344.400 308.300 ;
        RECT 236.400 307.600 237.200 307.700 ;
        RECT 257.200 307.600 258.000 307.700 ;
        RECT 276.400 307.600 277.200 307.700 ;
        RECT 289.200 307.600 290.000 307.700 ;
        RECT 343.600 307.600 344.400 307.700 ;
        RECT 343.600 268.300 344.400 268.400 ;
        RECT 383.600 268.300 384.400 268.400 ;
        RECT 343.600 267.700 384.400 268.300 ;
        RECT 343.600 267.600 344.400 267.700 ;
        RECT 383.600 267.600 384.400 267.700 ;
        RECT 265.200 134.300 266.000 134.400 ;
        RECT 276.400 134.300 277.200 134.400 ;
        RECT 265.200 133.700 277.200 134.300 ;
        RECT 265.200 133.600 266.000 133.700 ;
        RECT 276.400 133.600 277.200 133.700 ;
        RECT 265.200 104.300 266.000 104.400 ;
        RECT 303.600 104.300 304.400 104.400 ;
        RECT 265.200 103.700 304.400 104.300 ;
        RECT 265.200 103.600 266.000 103.700 ;
        RECT 303.600 103.600 304.400 103.700 ;
        RECT 388.400 68.300 389.200 68.400 ;
        RECT 463.600 68.300 464.400 68.400 ;
        RECT 388.400 67.700 464.400 68.300 ;
        RECT 388.400 67.600 389.200 67.700 ;
        RECT 463.600 67.600 464.400 67.700 ;
        RECT 303.600 54.300 304.400 54.400 ;
        RECT 327.600 54.300 328.400 54.400 ;
        RECT 356.400 54.300 357.200 54.400 ;
        RECT 388.400 54.300 389.200 54.400 ;
        RECT 303.600 53.700 389.200 54.300 ;
        RECT 303.600 53.600 304.400 53.700 ;
        RECT 327.600 53.600 328.400 53.700 ;
        RECT 356.400 53.600 357.200 53.700 ;
        RECT 388.400 53.600 389.200 53.700 ;
        RECT 322.800 14.300 323.600 14.400 ;
        RECT 327.600 14.300 328.400 14.400 ;
        RECT 329.200 14.300 330.000 14.400 ;
        RECT 322.800 13.700 330.000 14.300 ;
        RECT 322.800 13.600 323.600 13.700 ;
        RECT 327.600 13.600 328.400 13.700 ;
        RECT 329.200 13.600 330.000 13.700 ;
      LAYER metal4 ;
        RECT 257.000 307.400 258.200 382.600 ;
        RECT 276.200 133.400 277.400 308.600 ;
        RECT 343.400 267.400 344.600 374.600 ;
        RECT 327.400 13.400 328.600 54.600 ;
    END
  END rst
  PIN ext_data_in[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 215.600 2.000 217.200 ;
      LAYER metal2 ;
        RECT 1.200 215.600 2.000 216.400 ;
        RECT 1.300 210.400 1.900 215.600 ;
        RECT 1.200 209.600 2.000 210.400 ;
      LAYER metal3 ;
        RECT 1.200 210.300 2.000 210.400 ;
        RECT -1.900 209.700 2.000 210.300 ;
        RECT 1.200 209.600 2.000 209.700 ;
    END
  END ext_data_in[0]
  PIN ext_data_in[1]
    PORT
      LAYER metal1 ;
        RECT 36.400 24.800 37.200 26.400 ;
      LAYER via1 ;
        RECT 36.400 25.600 37.200 26.400 ;
      LAYER metal2 ;
        RECT 36.400 25.600 37.200 26.400 ;
        RECT 36.500 -2.300 37.100 25.600 ;
    END
  END ext_data_in[1]
  PIN ext_data_in[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 184.800 2.000 186.400 ;
      LAYER via1 ;
        RECT 1.200 185.600 2.000 186.400 ;
      LAYER metal2 ;
        RECT 1.200 189.600 2.000 190.400 ;
        RECT 1.300 186.400 1.900 189.600 ;
        RECT 1.200 185.600 2.000 186.400 ;
      LAYER metal3 ;
        RECT 1.200 190.300 2.000 190.400 ;
        RECT -1.900 189.700 2.000 190.300 ;
        RECT 1.200 189.600 2.000 189.700 ;
    END
  END ext_data_in[2]
  PIN ext_data_in[3]
    PORT
      LAYER metal1 ;
        RECT 44.400 15.600 45.200 17.200 ;
      LAYER metal2 ;
        RECT 44.400 16.300 45.200 16.400 ;
        RECT 42.900 15.700 45.200 16.300 ;
        RECT 42.900 -1.700 43.500 15.700 ;
        RECT 44.400 15.600 45.200 15.700 ;
        RECT 42.900 -2.300 45.100 -1.700 ;
    END
  END ext_data_in[3]
  PIN ext_data_in[4]
    PORT
      LAYER metal1 ;
        RECT 542.000 15.600 542.800 17.200 ;
      LAYER metal2 ;
        RECT 542.000 15.600 542.800 16.400 ;
        RECT 542.100 -1.700 542.700 15.600 ;
        RECT 540.500 -2.300 542.700 -1.700 ;
    END
  END ext_data_in[4]
  PIN ext_data_in[5]
    PORT
      LAYER metal1 ;
        RECT 502.000 15.600 502.800 17.200 ;
      LAYER metal2 ;
        RECT 502.000 15.600 502.800 16.400 ;
        RECT 502.100 -2.300 502.700 15.600 ;
    END
  END ext_data_in[5]
  PIN ext_data_in[6]
    PORT
      LAYER metal1 ;
        RECT 463.600 15.600 464.400 17.200 ;
      LAYER metal2 ;
        RECT 463.600 15.600 464.400 16.400 ;
        RECT 463.700 -2.300 464.300 15.600 ;
    END
  END ext_data_in[6]
  PIN ext_data_in[7]
    PORT
      LAYER metal1 ;
        RECT 494.000 24.800 494.800 26.400 ;
      LAYER via1 ;
        RECT 494.000 25.600 494.800 26.400 ;
      LAYER metal2 ;
        RECT 494.000 25.600 494.800 26.400 ;
        RECT 494.100 14.400 494.700 25.600 ;
        RECT 494.000 13.600 494.800 14.400 ;
        RECT 492.400 1.600 493.200 2.400 ;
        RECT 492.500 -2.300 493.100 1.600 ;
      LAYER metal3 ;
        RECT 494.000 13.600 494.800 14.400 ;
        RECT 492.400 2.300 493.200 2.400 ;
        RECT 494.000 2.300 494.800 2.400 ;
        RECT 492.400 1.700 494.800 2.300 ;
        RECT 492.400 1.600 493.200 1.700 ;
        RECT 494.000 1.600 494.800 1.700 ;
      LAYER metal4 ;
        RECT 493.800 1.400 495.000 14.600 ;
    END
  END ext_data_in[7]
  PIN ext_data_in[8]
    PORT
      LAYER metal1 ;
        RECT 81.200 495.600 82.000 497.200 ;
      LAYER metal2 ;
        RECT 81.300 496.400 81.900 504.300 ;
        RECT 81.200 495.600 82.000 496.400 ;
    END
  END ext_data_in[8]
  PIN ext_data_in[9]
    PORT
      LAYER metal1 ;
        RECT 1.200 295.600 2.000 297.200 ;
      LAYER metal2 ;
        RECT 1.200 295.600 2.000 296.400 ;
        RECT 1.300 290.400 1.900 295.600 ;
        RECT 1.200 289.600 2.000 290.400 ;
      LAYER metal3 ;
        RECT 1.200 290.300 2.000 290.400 ;
        RECT -1.900 289.700 2.000 290.300 ;
        RECT 1.200 289.600 2.000 289.700 ;
    END
  END ext_data_in[9]
  PIN ext_data_in[10]
    PORT
      LAYER metal1 ;
        RECT 156.400 495.600 157.200 497.200 ;
      LAYER metal2 ;
        RECT 156.500 496.400 157.100 504.300 ;
        RECT 156.400 495.600 157.200 496.400 ;
    END
  END ext_data_in[10]
  PIN ext_data_in[11]
    PORT
      LAYER metal1 ;
        RECT 44.400 495.600 45.200 497.200 ;
      LAYER metal2 ;
        RECT 42.900 503.700 45.100 504.300 ;
        RECT 44.500 496.400 45.100 503.700 ;
        RECT 44.400 495.600 45.200 496.400 ;
    END
  END ext_data_in[11]
  PIN ext_data_in[12]
    PORT
      LAYER metal1 ;
        RECT 489.200 455.600 490.000 457.200 ;
      LAYER metal2 ;
        RECT 484.500 500.400 485.100 504.300 ;
        RECT 484.400 499.600 485.200 500.400 ;
        RECT 489.200 461.600 490.000 462.400 ;
        RECT 489.300 456.400 489.900 461.600 ;
        RECT 489.200 455.600 490.000 456.400 ;
      LAYER metal3 ;
        RECT 484.400 499.600 485.200 500.400 ;
        RECT 484.400 462.300 485.200 462.400 ;
        RECT 489.200 462.300 490.000 462.400 ;
        RECT 484.400 461.700 490.000 462.300 ;
        RECT 484.400 461.600 485.200 461.700 ;
        RECT 489.200 461.600 490.000 461.700 ;
      LAYER metal4 ;
        RECT 484.200 461.400 485.400 500.600 ;
    END
  END ext_data_in[12]
  PIN ext_data_in[13]
    PORT
      LAYER metal1 ;
        RECT 484.400 495.600 485.200 497.200 ;
      LAYER metal2 ;
        RECT 487.700 498.400 488.300 504.300 ;
        RECT 484.400 497.600 485.200 498.400 ;
        RECT 487.600 497.600 488.400 498.400 ;
        RECT 484.500 496.400 485.100 497.600 ;
        RECT 484.400 495.600 485.200 496.400 ;
      LAYER metal3 ;
        RECT 484.400 498.300 485.200 498.400 ;
        RECT 487.600 498.300 488.400 498.400 ;
        RECT 484.400 497.700 488.400 498.300 ;
        RECT 484.400 497.600 485.200 497.700 ;
        RECT 487.600 497.600 488.400 497.700 ;
    END
  END ext_data_in[13]
  PIN ext_data_in[14]
    PORT
      LAYER metal1 ;
        RECT 540.400 455.600 541.200 457.200 ;
      LAYER metal2 ;
        RECT 538.900 503.700 541.100 504.300 ;
        RECT 540.500 456.400 541.100 503.700 ;
        RECT 540.400 455.600 541.200 456.400 ;
    END
  END ext_data_in[14]
  PIN ext_data_in[15]
    PORT
      LAYER metal1 ;
        RECT 479.600 495.600 480.400 497.200 ;
      LAYER metal2 ;
        RECT 479.700 496.400 480.300 504.300 ;
        RECT 479.600 495.600 480.400 496.400 ;
    END
  END ext_data_in[15]
  PIN ext_data_out[0]
    PORT
      LAYER metal1 ;
        RECT 318.000 12.400 318.800 19.800 ;
        RECT 318.000 10.200 318.600 12.400 ;
        RECT 318.000 2.200 318.800 10.200 ;
      LAYER via1 ;
        RECT 318.000 3.600 318.800 4.400 ;
      LAYER metal2 ;
        RECT 318.000 3.600 318.800 4.400 ;
        RECT 318.100 -1.700 318.700 3.600 ;
        RECT 318.100 -2.300 320.300 -1.700 ;
    END
  END ext_data_out[0]
  PIN ext_data_out[1]
    PORT
      LAYER metal1 ;
        RECT 242.800 12.400 243.600 19.800 ;
        RECT 243.000 10.200 243.600 12.400 ;
        RECT 242.800 2.200 243.600 10.200 ;
      LAYER via1 ;
        RECT 242.800 3.600 243.600 4.400 ;
      LAYER metal2 ;
        RECT 242.800 3.600 243.600 4.400 ;
        RECT 242.900 -1.700 243.500 3.600 ;
        RECT 241.300 -2.300 243.500 -1.700 ;
    END
  END ext_data_out[1]
  PIN ext_data_out[2]
    PORT
      LAYER metal1 ;
        RECT 255.600 12.400 256.400 19.800 ;
        RECT 255.600 10.200 256.200 12.400 ;
        RECT 255.600 2.200 256.400 10.200 ;
      LAYER via1 ;
        RECT 255.600 3.600 256.400 4.400 ;
      LAYER metal2 ;
        RECT 255.600 3.600 256.400 4.400 ;
        RECT 255.700 -1.700 256.300 3.600 ;
        RECT 255.700 -2.300 257.900 -1.700 ;
    END
  END ext_data_out[2]
  PIN ext_data_out[3]
    PORT
      LAYER metal1 ;
        RECT 268.400 12.400 269.200 19.800 ;
        RECT 268.400 10.200 269.000 12.400 ;
        RECT 268.400 2.200 269.200 10.200 ;
      LAYER via1 ;
        RECT 268.400 3.600 269.200 4.400 ;
      LAYER metal2 ;
        RECT 268.400 3.600 269.200 4.400 ;
        RECT 268.500 -1.700 269.100 3.600 ;
        RECT 268.500 -2.300 270.700 -1.700 ;
    END
  END ext_data_out[3]
  PIN ext_data_out[4]
    PORT
      LAYER metal1 ;
        RECT 378.800 12.400 379.600 19.800 ;
        RECT 379.000 10.200 379.600 12.400 ;
        RECT 378.800 2.200 379.600 10.200 ;
      LAYER via1 ;
        RECT 378.800 3.600 379.600 4.400 ;
      LAYER metal2 ;
        RECT 378.800 3.600 379.600 4.400 ;
        RECT 378.900 -1.700 379.500 3.600 ;
        RECT 377.300 -2.300 379.500 -1.700 ;
    END
  END ext_data_out[4]
  PIN ext_data_out[5]
    PORT
      LAYER metal1 ;
        RECT 415.600 12.400 416.400 19.800 ;
        RECT 415.600 10.200 416.200 12.400 ;
        RECT 415.600 2.200 416.400 10.200 ;
      LAYER via1 ;
        RECT 415.600 3.600 416.400 4.400 ;
      LAYER metal2 ;
        RECT 412.400 3.600 413.200 4.400 ;
        RECT 415.600 3.600 416.400 4.400 ;
        RECT 412.500 -1.700 413.100 3.600 ;
        RECT 412.500 -2.300 421.100 -1.700 ;
      LAYER metal3 ;
        RECT 412.400 4.300 413.200 4.400 ;
        RECT 415.600 4.300 416.400 4.400 ;
        RECT 412.400 3.700 416.400 4.300 ;
        RECT 412.400 3.600 413.200 3.700 ;
        RECT 415.600 3.600 416.400 3.700 ;
    END
  END ext_data_out[5]
  PIN ext_data_out[6]
    PORT
      LAYER metal1 ;
        RECT 374.000 12.400 374.800 19.800 ;
        RECT 374.200 10.200 374.800 12.400 ;
        RECT 374.000 2.200 374.800 10.200 ;
      LAYER via1 ;
        RECT 374.000 3.600 374.800 4.400 ;
      LAYER metal2 ;
        RECT 374.000 3.600 374.800 4.400 ;
        RECT 374.100 -1.700 374.700 3.600 ;
        RECT 372.500 -2.300 374.700 -1.700 ;
    END
  END ext_data_out[6]
  PIN ext_data_out[7]
    PORT
      LAYER metal1 ;
        RECT 330.800 12.400 331.600 19.800 ;
        RECT 330.800 10.200 331.400 12.400 ;
        RECT 330.800 2.200 331.600 10.200 ;
      LAYER via1 ;
        RECT 330.800 3.600 331.600 4.400 ;
      LAYER metal2 ;
        RECT 330.800 3.600 331.600 4.400 ;
        RECT 330.900 -1.700 331.500 3.600 ;
        RECT 330.900 -2.300 333.100 -1.700 ;
    END
  END ext_data_out[7]
  PIN ext_data_out[8]
    PORT
      LAYER metal1 ;
        RECT 297.200 492.400 298.000 499.800 ;
        RECT 297.400 490.200 298.000 492.400 ;
        RECT 297.200 482.200 298.000 490.200 ;
      LAYER via1 ;
        RECT 297.200 497.600 298.000 498.400 ;
      LAYER metal2 ;
        RECT 295.700 503.700 297.900 504.300 ;
        RECT 297.300 498.400 297.900 503.700 ;
        RECT 297.200 497.600 298.000 498.400 ;
    END
  END ext_data_out[8]
  PIN ext_data_out[9]
    PORT
      LAYER metal1 ;
        RECT 225.200 372.400 226.000 379.800 ;
        RECT 225.400 370.200 226.000 372.400 ;
        RECT 225.200 362.200 226.000 370.200 ;
      LAYER via1 ;
        RECT 225.200 377.600 226.000 378.400 ;
      LAYER metal2 ;
        RECT 223.700 500.400 224.300 504.300 ;
        RECT 223.600 499.600 224.400 500.400 ;
        RECT 225.200 381.600 226.000 382.400 ;
        RECT 225.300 378.400 225.900 381.600 ;
        RECT 225.200 377.600 226.000 378.400 ;
      LAYER metal3 ;
        RECT 223.600 500.300 224.400 500.400 ;
        RECT 225.200 500.300 226.000 500.400 ;
        RECT 223.600 499.700 226.000 500.300 ;
        RECT 223.600 499.600 224.400 499.700 ;
        RECT 225.200 499.600 226.000 499.700 ;
        RECT 225.200 381.600 226.000 382.400 ;
      LAYER metal4 ;
        RECT 225.000 381.400 226.200 500.600 ;
    END
  END ext_data_out[9]
  PIN ext_data_out[10]
    PORT
      LAYER metal1 ;
        RECT 6.000 252.400 6.800 259.800 ;
        RECT 6.000 250.200 6.600 252.400 ;
        RECT 6.000 242.200 6.800 250.200 ;
      LAYER via1 ;
        RECT 6.000 253.600 6.800 254.400 ;
      LAYER metal2 ;
        RECT 6.000 253.600 6.800 254.400 ;
      LAYER metal3 ;
        RECT 6.000 254.300 6.800 254.400 ;
        RECT -1.900 253.700 6.800 254.300 ;
        RECT 6.000 253.600 6.800 253.700 ;
    END
  END ext_data_out[10]
  PIN ext_data_out[11]
    PORT
      LAYER metal1 ;
        RECT 1.200 252.400 2.000 259.800 ;
        RECT 1.200 250.200 1.800 252.400 ;
        RECT 1.200 242.200 2.000 250.200 ;
      LAYER via1 ;
        RECT 1.200 247.600 2.000 248.400 ;
      LAYER metal2 ;
        RECT 1.200 249.600 2.000 250.400 ;
        RECT 1.300 248.400 1.900 249.600 ;
        RECT 1.200 247.600 2.000 248.400 ;
      LAYER metal3 ;
        RECT 1.200 250.300 2.000 250.400 ;
        RECT -1.900 249.700 2.000 250.300 ;
        RECT 1.200 249.600 2.000 249.700 ;
    END
  END ext_data_out[11]
  PIN ext_data_out[12]
    PORT
      LAYER metal1 ;
        RECT 428.400 492.400 429.200 499.800 ;
        RECT 428.600 490.200 429.200 492.400 ;
        RECT 428.400 482.200 429.200 490.200 ;
      LAYER via1 ;
        RECT 428.400 497.600 429.200 498.400 ;
      LAYER metal2 ;
        RECT 426.900 503.700 429.100 504.300 ;
        RECT 428.500 498.400 429.100 503.700 ;
        RECT 428.400 497.600 429.200 498.400 ;
    END
  END ext_data_out[12]
  PIN ext_data_out[13]
    PORT
      LAYER metal1 ;
        RECT 380.400 492.400 381.200 499.800 ;
        RECT 380.400 490.200 381.000 492.400 ;
        RECT 380.400 482.200 381.200 490.200 ;
      LAYER via1 ;
        RECT 380.400 497.600 381.200 498.400 ;
      LAYER metal2 ;
        RECT 380.500 503.700 382.700 504.300 ;
        RECT 380.500 498.400 381.100 503.700 ;
        RECT 380.400 497.600 381.200 498.400 ;
    END
  END ext_data_out[13]
  PIN ext_data_out[14]
    PORT
      LAYER metal1 ;
        RECT 550.000 231.800 550.800 239.800 ;
        RECT 550.000 229.600 550.600 231.800 ;
        RECT 550.000 222.200 550.800 229.600 ;
      LAYER via1 ;
        RECT 550.000 237.600 550.800 238.400 ;
      LAYER metal2 ;
        RECT 551.700 500.400 552.300 504.300 ;
        RECT 551.600 499.600 552.400 500.400 ;
        RECT 553.200 461.600 554.000 462.400 ;
        RECT 553.300 362.400 553.900 461.600 ;
        RECT 553.200 361.600 554.000 362.400 ;
        RECT 550.000 261.600 550.800 262.400 ;
        RECT 550.100 238.400 550.700 261.600 ;
        RECT 550.000 237.600 550.800 238.400 ;
      LAYER metal3 ;
        RECT 551.600 499.600 552.400 500.400 ;
        RECT 551.600 462.300 552.400 462.400 ;
        RECT 553.200 462.300 554.000 462.400 ;
        RECT 551.600 461.700 554.000 462.300 ;
        RECT 551.600 461.600 552.400 461.700 ;
        RECT 553.200 461.600 554.000 461.700 ;
        RECT 553.200 362.300 554.000 362.400 ;
        RECT 554.800 362.300 555.600 362.400 ;
        RECT 553.200 361.700 555.600 362.300 ;
        RECT 553.200 361.600 554.000 361.700 ;
        RECT 554.800 361.600 555.600 361.700 ;
        RECT 550.000 262.300 550.800 262.400 ;
        RECT 554.800 262.300 555.600 262.400 ;
        RECT 550.000 261.700 555.600 262.300 ;
        RECT 550.000 261.600 550.800 261.700 ;
        RECT 554.800 261.600 555.600 261.700 ;
      LAYER metal4 ;
        RECT 551.400 461.400 552.600 500.600 ;
        RECT 554.600 261.400 555.800 362.600 ;
    END
  END ext_data_out[14]
  PIN ext_data_out[15]
    PORT
      LAYER metal1 ;
        RECT 489.200 496.300 490.000 499.800 ;
        RECT 490.800 496.300 491.600 496.400 ;
        RECT 489.200 495.700 491.600 496.300 ;
        RECT 489.200 492.400 490.000 495.700 ;
        RECT 490.800 495.600 491.600 495.700 ;
        RECT 489.400 490.200 490.000 492.400 ;
        RECT 489.200 482.200 490.000 490.200 ;
      LAYER metal2 ;
        RECT 490.900 496.400 491.500 504.300 ;
        RECT 490.800 495.600 491.600 496.400 ;
    END
  END ext_data_out[15]
  PIN pe_busy[0]
    PORT
      LAYER metal1 ;
        RECT 39.600 12.400 40.400 19.800 ;
        RECT 39.600 10.200 40.200 12.400 ;
        RECT 39.600 2.200 40.400 10.200 ;
      LAYER via1 ;
        RECT 39.600 3.600 40.400 4.400 ;
      LAYER metal2 ;
        RECT 39.600 3.600 40.400 4.400 ;
        RECT 39.700 -1.700 40.300 3.600 ;
        RECT 39.700 -2.300 41.900 -1.700 ;
    END
  END pe_busy[0]
  PIN pe_busy[1]
    PORT
      LAYER metal1 ;
        RECT 586.800 12.400 587.600 19.800 ;
        RECT 587.000 10.200 587.600 12.400 ;
        RECT 586.800 2.200 587.600 10.200 ;
      LAYER via1 ;
        RECT 586.800 3.600 587.600 4.400 ;
      LAYER metal2 ;
        RECT 586.800 3.600 587.600 4.400 ;
        RECT 586.900 -1.700 587.500 3.600 ;
        RECT 585.300 -2.300 587.500 -1.700 ;
    END
  END pe_busy[1]
  PIN pe_busy[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 391.800 2.000 399.800 ;
        RECT 1.200 389.600 1.800 391.800 ;
        RECT 1.200 382.200 2.000 389.600 ;
      LAYER via1 ;
        RECT 1.200 387.600 2.000 388.400 ;
      LAYER metal2 ;
        RECT 1.200 389.600 2.000 390.400 ;
        RECT 1.300 388.400 1.900 389.600 ;
        RECT 1.200 387.600 2.000 388.400 ;
      LAYER metal3 ;
        RECT 1.200 390.300 2.000 390.400 ;
        RECT -1.900 389.700 2.000 390.300 ;
        RECT 1.200 389.600 2.000 389.700 ;
    END
  END pe_busy[2]
  PIN pe_busy[3]
    PORT
      LAYER metal1 ;
        RECT 681.200 471.800 682.000 479.800 ;
        RECT 681.400 469.600 682.000 471.800 ;
        RECT 681.200 468.300 682.000 469.600 ;
        RECT 687.600 468.300 688.400 468.400 ;
        RECT 681.200 467.700 688.400 468.300 ;
        RECT 681.200 462.200 682.000 467.700 ;
        RECT 687.600 467.600 688.400 467.700 ;
      LAYER metal2 ;
        RECT 687.600 469.600 688.400 470.400 ;
        RECT 687.700 468.400 688.300 469.600 ;
        RECT 687.600 467.600 688.400 468.400 ;
      LAYER metal3 ;
        RECT 687.600 470.300 688.400 470.400 ;
        RECT 687.600 469.700 691.500 470.300 ;
        RECT 687.600 469.600 688.400 469.700 ;
    END
  END pe_busy[3]
  OBS
      LAYER metal1 ;
        RECT 1.200 493.800 2.000 499.800 ;
        RECT 7.600 496.600 8.400 499.800 ;
        RECT 9.200 497.000 10.000 499.800 ;
        RECT 10.800 497.000 11.600 499.800 ;
        RECT 12.400 497.000 13.200 499.800 ;
        RECT 15.600 497.000 16.400 499.800 ;
        RECT 18.800 497.000 19.600 499.800 ;
        RECT 20.400 497.000 21.200 499.800 ;
        RECT 22.000 497.000 22.800 499.800 ;
        RECT 23.600 497.000 24.400 499.800 ;
        RECT 5.800 495.800 8.400 496.600 ;
        RECT 25.200 496.600 26.000 499.800 ;
        RECT 11.800 495.800 16.400 496.400 ;
        RECT 5.800 495.200 6.600 495.800 ;
        RECT 3.600 494.400 6.600 495.200 ;
        RECT 1.200 493.000 10.000 493.800 ;
        RECT 11.800 493.400 12.600 495.800 ;
        RECT 15.600 495.600 16.400 495.800 ;
        RECT 17.200 495.600 18.800 496.400 ;
        RECT 21.800 495.600 22.800 496.400 ;
        RECT 25.200 495.800 27.600 496.600 ;
        RECT 14.000 493.600 14.800 495.200 ;
        RECT 15.600 494.800 16.400 495.000 ;
        RECT 15.600 494.200 20.000 494.800 ;
        RECT 19.200 494.000 20.000 494.200 ;
        RECT 1.200 487.400 2.000 493.000 ;
        RECT 10.600 492.600 12.600 493.400 ;
        RECT 16.400 492.600 19.600 493.400 ;
        RECT 22.000 492.800 22.800 495.600 ;
        RECT 26.800 495.200 27.600 495.800 ;
        RECT 26.800 494.600 28.600 495.200 ;
        RECT 27.800 493.400 28.600 494.600 ;
        RECT 31.600 494.600 32.400 499.800 ;
        RECT 33.200 496.000 34.000 499.800 ;
        RECT 33.200 495.200 34.200 496.000 ;
        RECT 36.400 495.800 37.200 499.800 ;
        RECT 38.000 496.000 38.800 499.800 ;
        RECT 41.200 496.000 42.000 499.800 ;
        RECT 38.000 495.800 42.000 496.000 ;
        RECT 31.600 494.000 32.800 494.600 ;
        RECT 27.800 492.600 31.600 493.400 ;
        RECT 2.600 492.000 3.400 492.200 ;
        RECT 7.600 492.000 8.400 492.400 ;
        RECT 14.000 492.000 14.800 492.400 ;
        RECT 25.200 492.000 26.000 492.600 ;
        RECT 32.200 492.000 32.800 494.000 ;
        RECT 2.600 491.400 26.000 492.000 ;
        RECT 32.000 491.400 32.800 492.000 ;
        RECT 32.000 489.600 32.600 491.400 ;
        RECT 33.400 490.800 34.200 495.200 ;
        RECT 36.600 494.400 37.200 495.800 ;
        RECT 38.200 495.400 41.800 495.800 ;
        RECT 40.400 494.400 41.200 494.800 ;
        RECT 34.800 494.300 35.600 494.400 ;
        RECT 36.400 494.300 39.000 494.400 ;
        RECT 34.800 493.700 39.000 494.300 ;
        RECT 40.400 494.300 42.000 494.400 ;
        RECT 42.800 494.300 43.600 499.800 ;
        RECT 40.400 493.800 43.600 494.300 ;
        RECT 34.800 493.600 35.600 493.700 ;
        RECT 36.400 493.600 39.000 493.700 ;
        RECT 41.200 493.700 43.600 493.800 ;
        RECT 41.200 493.600 42.000 493.700 ;
        RECT 10.800 489.400 11.600 489.600 ;
        RECT 6.200 489.000 11.600 489.400 ;
        RECT 5.400 488.800 11.600 489.000 ;
        RECT 12.600 489.000 21.200 489.600 ;
        RECT 2.800 488.000 4.400 488.800 ;
        RECT 5.400 488.200 6.800 488.800 ;
        RECT 12.600 488.200 13.200 489.000 ;
        RECT 20.400 488.800 21.200 489.000 ;
        RECT 23.600 489.000 32.600 489.600 ;
        RECT 23.600 488.800 24.400 489.000 ;
        RECT 3.800 487.600 4.400 488.000 ;
        RECT 7.400 487.600 13.200 488.200 ;
        RECT 13.800 487.600 16.400 488.400 ;
        RECT 1.200 486.800 3.200 487.400 ;
        RECT 3.800 486.800 8.000 487.600 ;
        RECT 2.600 486.200 3.200 486.800 ;
        RECT 2.600 485.600 3.600 486.200 ;
        RECT 2.800 482.200 3.600 485.600 ;
        RECT 6.000 482.200 6.800 486.800 ;
        RECT 9.200 482.200 10.000 485.000 ;
        RECT 10.800 482.200 11.600 485.000 ;
        RECT 12.400 482.200 13.200 487.000 ;
        RECT 15.600 482.200 16.400 487.000 ;
        RECT 18.800 482.200 19.600 488.400 ;
        RECT 26.800 487.600 29.400 488.400 ;
        RECT 22.000 486.800 26.200 487.600 ;
        RECT 20.400 482.200 21.200 485.000 ;
        RECT 22.000 482.200 22.800 485.000 ;
        RECT 23.600 482.200 24.400 485.000 ;
        RECT 26.800 482.200 27.600 487.600 ;
        RECT 32.000 487.400 32.600 489.000 ;
        RECT 30.000 486.800 32.600 487.400 ;
        RECT 33.200 490.000 34.200 490.800 ;
        RECT 36.400 490.200 37.200 490.400 ;
        RECT 38.400 490.200 39.000 493.600 ;
        RECT 39.600 492.300 40.400 493.200 ;
        RECT 41.200 492.300 42.000 492.400 ;
        RECT 39.600 491.700 42.000 492.300 ;
        RECT 39.600 491.600 40.400 491.700 ;
        RECT 41.200 491.600 42.000 491.700 ;
        RECT 30.000 482.200 30.800 486.800 ;
        RECT 33.200 482.200 34.000 490.000 ;
        RECT 36.400 489.600 37.800 490.200 ;
        RECT 38.400 489.600 39.400 490.200 ;
        RECT 37.200 488.400 37.800 489.600 ;
        RECT 37.200 487.600 38.000 488.400 ;
        RECT 38.600 482.200 39.400 489.600 ;
        RECT 42.800 482.200 43.600 493.700 ;
        RECT 46.000 493.800 46.800 499.800 ;
        RECT 52.400 496.600 53.200 499.800 ;
        RECT 54.000 497.000 54.800 499.800 ;
        RECT 55.600 497.000 56.400 499.800 ;
        RECT 57.200 497.000 58.000 499.800 ;
        RECT 60.400 497.000 61.200 499.800 ;
        RECT 63.600 497.000 64.400 499.800 ;
        RECT 65.200 497.000 66.000 499.800 ;
        RECT 66.800 497.000 67.600 499.800 ;
        RECT 68.400 497.000 69.200 499.800 ;
        RECT 50.600 495.800 53.200 496.600 ;
        RECT 70.000 496.600 70.800 499.800 ;
        RECT 56.600 495.800 61.200 496.400 ;
        RECT 50.600 495.200 51.400 495.800 ;
        RECT 48.400 494.400 51.400 495.200 ;
        RECT 46.000 493.000 54.800 493.800 ;
        RECT 56.600 493.400 57.400 495.800 ;
        RECT 60.400 495.600 61.200 495.800 ;
        RECT 62.000 495.600 63.600 496.400 ;
        RECT 66.600 495.600 67.600 496.400 ;
        RECT 70.000 495.800 72.400 496.600 ;
        RECT 58.800 493.600 59.600 495.200 ;
        RECT 60.400 494.800 61.200 495.000 ;
        RECT 60.400 494.200 64.800 494.800 ;
        RECT 64.000 494.000 64.800 494.200 ;
        RECT 46.000 487.400 46.800 493.000 ;
        RECT 55.400 492.600 57.400 493.400 ;
        RECT 61.200 492.600 64.400 493.400 ;
        RECT 66.800 492.800 67.600 495.600 ;
        RECT 71.600 495.200 72.400 495.800 ;
        RECT 71.600 494.600 73.400 495.200 ;
        RECT 72.600 493.400 73.400 494.600 ;
        RECT 76.400 494.600 77.200 499.800 ;
        RECT 78.000 496.000 78.800 499.800 ;
        RECT 78.000 495.200 79.000 496.000 ;
        RECT 76.400 494.000 77.600 494.600 ;
        RECT 72.600 492.600 76.400 493.400 ;
        RECT 47.400 492.000 48.200 492.200 ;
        RECT 49.200 492.000 50.000 492.400 ;
        RECT 52.400 492.000 53.200 492.400 ;
        RECT 70.000 492.000 70.800 492.600 ;
        RECT 77.000 492.000 77.600 494.000 ;
        RECT 47.400 491.400 70.800 492.000 ;
        RECT 76.800 491.400 77.600 492.000 ;
        RECT 76.800 489.600 77.400 491.400 ;
        RECT 78.200 490.800 79.000 495.200 ;
        RECT 55.600 489.400 56.400 489.600 ;
        RECT 51.000 489.000 56.400 489.400 ;
        RECT 50.200 488.800 56.400 489.000 ;
        RECT 57.400 489.000 66.000 489.600 ;
        RECT 47.600 488.000 49.200 488.800 ;
        RECT 50.200 488.200 51.600 488.800 ;
        RECT 57.400 488.200 58.000 489.000 ;
        RECT 65.200 488.800 66.000 489.000 ;
        RECT 68.400 489.000 77.400 489.600 ;
        RECT 68.400 488.800 69.200 489.000 ;
        RECT 48.600 487.600 49.200 488.000 ;
        RECT 52.200 487.600 58.000 488.200 ;
        RECT 58.600 487.600 61.200 488.400 ;
        RECT 46.000 486.800 48.000 487.400 ;
        RECT 48.600 486.800 52.800 487.600 ;
        RECT 47.400 486.200 48.000 486.800 ;
        RECT 47.400 485.600 48.400 486.200 ;
        RECT 47.600 482.200 48.400 485.600 ;
        RECT 50.800 482.200 51.600 486.800 ;
        RECT 54.000 482.200 54.800 485.000 ;
        RECT 55.600 482.200 56.400 485.000 ;
        RECT 57.200 482.200 58.000 487.000 ;
        RECT 60.400 482.200 61.200 487.000 ;
        RECT 63.600 482.200 64.400 488.400 ;
        RECT 71.600 487.600 74.200 488.400 ;
        RECT 66.800 486.800 71.000 487.600 ;
        RECT 65.200 482.200 66.000 485.000 ;
        RECT 66.800 482.200 67.600 485.000 ;
        RECT 68.400 482.200 69.200 485.000 ;
        RECT 71.600 482.200 72.400 487.600 ;
        RECT 76.800 487.400 77.400 489.000 ;
        RECT 74.800 486.800 77.400 487.400 ;
        RECT 78.000 490.000 79.000 490.800 ;
        RECT 82.800 494.300 83.600 499.800 ;
        RECT 84.400 496.000 85.200 499.800 ;
        RECT 87.600 496.000 88.400 499.800 ;
        RECT 84.400 495.800 88.400 496.000 ;
        RECT 89.200 495.800 90.000 499.800 ;
        RECT 90.800 495.800 91.600 499.800 ;
        RECT 92.400 496.000 93.200 499.800 ;
        RECT 95.600 496.000 96.400 499.800 ;
        RECT 92.400 495.800 96.400 496.000 ;
        RECT 84.600 495.400 88.200 495.800 ;
        RECT 85.200 494.400 86.000 494.800 ;
        RECT 89.200 494.400 89.800 495.800 ;
        RECT 91.000 494.400 91.600 495.800 ;
        RECT 92.600 495.400 96.200 495.800 ;
        RECT 98.800 495.200 99.600 499.800 ;
        RECT 102.000 495.200 102.800 499.800 ;
        RECT 105.200 495.200 106.000 499.800 ;
        RECT 108.400 495.200 109.200 499.800 ;
        RECT 94.800 494.400 95.600 494.800 ;
        RECT 97.200 494.400 99.600 495.200 ;
        RECT 100.600 494.400 102.800 495.200 ;
        RECT 103.800 494.400 106.000 495.200 ;
        RECT 107.400 494.400 109.200 495.200 ;
        RECT 116.400 495.000 117.200 499.800 ;
        RECT 120.800 498.400 121.600 499.800 ;
        RECT 119.600 497.800 121.600 498.400 ;
        RECT 125.200 497.800 126.000 499.800 ;
        RECT 129.400 498.400 130.600 499.800 ;
        RECT 129.200 497.800 130.600 498.400 ;
        RECT 119.600 497.000 120.400 497.800 ;
        RECT 125.200 497.200 125.800 497.800 ;
        RECT 121.200 496.400 122.000 497.200 ;
        RECT 123.000 496.600 125.800 497.200 ;
        RECT 129.200 497.000 130.000 497.800 ;
        RECT 123.000 496.400 123.800 496.600 ;
        RECT 84.400 494.300 86.000 494.400 ;
        RECT 82.800 493.800 86.000 494.300 ;
        RECT 82.800 493.700 85.200 493.800 ;
        RECT 74.800 482.200 75.600 486.800 ;
        RECT 78.000 482.200 78.800 490.000 ;
        RECT 82.800 482.200 83.600 493.700 ;
        RECT 84.400 493.600 85.200 493.700 ;
        RECT 87.400 493.600 90.000 494.400 ;
        RECT 90.800 493.600 93.400 494.400 ;
        RECT 94.800 493.800 96.400 494.400 ;
        RECT 95.600 493.600 96.400 493.800 ;
        RECT 86.000 491.600 86.800 493.200 ;
        RECT 87.400 490.200 88.000 493.600 ;
        RECT 92.800 492.300 93.400 493.600 ;
        RECT 89.300 491.700 93.400 492.300 ;
        RECT 89.300 490.400 89.900 491.700 ;
        RECT 89.200 490.200 90.000 490.400 ;
        RECT 87.000 489.600 88.000 490.200 ;
        RECT 88.600 489.600 90.000 490.200 ;
        RECT 90.800 490.200 91.600 490.400 ;
        RECT 92.800 490.200 93.400 491.700 ;
        RECT 94.000 491.600 94.800 493.200 ;
        RECT 97.200 491.600 98.000 494.400 ;
        RECT 100.600 493.800 101.400 494.400 ;
        RECT 103.800 493.800 104.600 494.400 ;
        RECT 107.400 493.800 108.200 494.400 ;
        RECT 110.000 493.800 110.800 494.400 ;
        RECT 98.800 493.000 101.400 493.800 ;
        RECT 102.200 493.000 104.600 493.800 ;
        RECT 105.600 493.000 108.200 493.800 ;
        RECT 109.000 493.000 110.800 493.800 ;
        RECT 117.200 494.200 118.800 494.400 ;
        RECT 121.400 494.200 122.000 496.400 ;
        RECT 131.000 495.400 131.800 495.600 ;
        RECT 134.000 495.400 134.800 499.800 ;
        RECT 131.000 494.800 134.800 495.400 ;
        RECT 137.200 495.200 138.000 499.800 ;
        RECT 140.400 495.200 141.200 499.800 ;
        RECT 143.600 495.200 144.400 499.800 ;
        RECT 146.800 495.200 147.600 499.800 ;
        RECT 150.000 496.000 150.800 499.800 ;
        RECT 153.200 496.000 154.000 499.800 ;
        RECT 150.000 495.800 154.000 496.000 ;
        RECT 154.800 495.800 155.600 499.800 ;
        RECT 150.200 495.400 153.800 495.800 ;
        RECT 127.000 494.200 127.800 494.400 ;
        RECT 117.200 493.600 128.200 494.200 ;
        RECT 120.200 493.400 121.000 493.600 ;
        RECT 100.600 491.600 101.400 493.000 ;
        RECT 103.800 491.600 104.600 493.000 ;
        RECT 107.400 491.600 108.200 493.000 ;
        RECT 118.600 492.400 119.400 492.600 ;
        RECT 127.600 492.400 128.200 493.600 ;
        RECT 129.200 492.800 130.000 493.000 ;
        RECT 118.600 492.300 123.600 492.400 ;
        RECT 124.400 492.300 125.200 492.400 ;
        RECT 118.600 491.800 125.200 492.300 ;
        RECT 122.800 491.700 125.200 491.800 ;
        RECT 122.800 491.600 123.600 491.700 ;
        RECT 124.400 491.600 125.200 491.700 ;
        RECT 127.600 491.600 128.400 492.400 ;
        RECT 129.200 492.200 133.000 492.800 ;
        RECT 132.200 492.000 133.000 492.200 ;
        RECT 97.200 490.800 99.600 491.600 ;
        RECT 100.600 490.800 102.800 491.600 ;
        RECT 103.800 490.800 106.000 491.600 ;
        RECT 107.400 490.800 109.200 491.600 ;
        RECT 90.800 489.600 92.200 490.200 ;
        RECT 92.800 489.600 93.800 490.200 ;
        RECT 87.000 482.200 87.800 489.600 ;
        RECT 88.600 488.400 89.200 489.600 ;
        RECT 88.400 487.600 89.200 488.400 ;
        RECT 91.600 488.400 92.200 489.600 ;
        RECT 91.600 487.600 92.400 488.400 ;
        RECT 93.000 482.200 93.800 489.600 ;
        RECT 98.800 482.200 99.600 490.800 ;
        RECT 102.000 482.200 102.800 490.800 ;
        RECT 105.200 482.200 106.000 490.800 ;
        RECT 108.400 482.200 109.200 490.800 ;
        RECT 116.400 491.000 122.000 491.200 ;
        RECT 116.400 490.800 122.200 491.000 ;
        RECT 116.400 490.600 126.200 490.800 ;
        RECT 116.400 482.200 117.200 490.600 ;
        RECT 121.400 490.200 126.200 490.600 ;
        RECT 119.600 489.000 125.000 489.600 ;
        RECT 119.600 488.800 120.400 489.000 ;
        RECT 124.200 488.800 125.000 489.000 ;
        RECT 125.600 489.000 126.200 490.200 ;
        RECT 127.600 490.400 128.200 491.600 ;
        RECT 130.600 491.400 131.400 491.600 ;
        RECT 134.000 491.400 134.800 494.800 ;
        RECT 130.600 490.800 134.800 491.400 ;
        RECT 135.600 494.400 138.000 495.200 ;
        RECT 139.000 494.400 141.200 495.200 ;
        RECT 142.200 494.400 144.400 495.200 ;
        RECT 145.800 494.400 147.600 495.200 ;
        RECT 150.800 494.400 151.600 494.800 ;
        RECT 154.800 494.400 155.400 495.800 ;
        RECT 135.600 491.600 136.400 494.400 ;
        RECT 139.000 493.800 139.800 494.400 ;
        RECT 142.200 493.800 143.000 494.400 ;
        RECT 145.800 493.800 146.600 494.400 ;
        RECT 148.400 493.800 149.200 494.400 ;
        RECT 137.200 493.000 139.800 493.800 ;
        RECT 140.600 493.000 143.000 493.800 ;
        RECT 144.000 493.000 146.600 493.800 ;
        RECT 147.400 493.000 149.200 493.800 ;
        RECT 150.000 493.800 151.600 494.400 ;
        RECT 150.000 493.600 150.800 493.800 ;
        RECT 153.000 493.600 155.600 494.400 ;
        RECT 158.000 494.300 158.800 499.800 ;
        RECT 159.600 496.000 160.400 499.800 ;
        RECT 162.800 496.000 163.600 499.800 ;
        RECT 159.600 495.800 163.600 496.000 ;
        RECT 164.400 495.800 165.200 499.800 ;
        RECT 167.600 496.000 168.400 499.800 ;
        RECT 159.800 495.400 163.400 495.800 ;
        RECT 160.400 494.400 161.200 494.800 ;
        RECT 164.400 494.400 165.000 495.800 ;
        RECT 167.400 495.200 168.400 496.000 ;
        RECT 159.600 494.300 161.200 494.400 ;
        RECT 158.000 493.800 161.200 494.300 ;
        RECT 158.000 493.700 160.400 493.800 ;
        RECT 139.000 491.600 139.800 493.000 ;
        RECT 142.200 491.600 143.000 493.000 ;
        RECT 145.800 491.600 146.600 493.000 ;
        RECT 151.600 491.600 152.400 493.200 ;
        RECT 153.000 492.300 153.600 493.600 ;
        RECT 156.400 492.300 157.200 492.400 ;
        RECT 153.000 491.700 157.200 492.300 ;
        RECT 135.600 490.800 138.000 491.600 ;
        RECT 139.000 490.800 141.200 491.600 ;
        RECT 142.200 490.800 144.400 491.600 ;
        RECT 145.800 490.800 147.600 491.600 ;
        RECT 127.600 489.800 130.000 490.400 ;
        RECT 127.000 489.000 127.800 489.200 ;
        RECT 125.600 488.400 127.800 489.000 ;
        RECT 129.400 488.800 130.000 489.800 ;
        RECT 129.400 488.000 130.800 488.800 ;
        RECT 123.000 487.400 123.800 487.600 ;
        RECT 125.800 487.400 126.600 487.600 ;
        RECT 119.600 486.200 120.400 487.000 ;
        RECT 123.000 486.800 126.600 487.400 ;
        RECT 125.200 486.200 125.800 486.800 ;
        RECT 129.200 486.200 130.000 487.000 ;
        RECT 119.600 485.600 121.600 486.200 ;
        RECT 120.800 482.200 121.600 485.600 ;
        RECT 125.200 482.200 126.000 486.200 ;
        RECT 129.400 482.200 130.600 486.200 ;
        RECT 134.000 482.200 134.800 490.800 ;
        RECT 137.200 482.200 138.000 490.800 ;
        RECT 140.400 482.200 141.200 490.800 ;
        RECT 143.600 482.200 144.400 490.800 ;
        RECT 146.800 482.200 147.600 490.800 ;
        RECT 153.000 490.200 153.600 491.700 ;
        RECT 156.400 491.600 157.200 491.700 ;
        RECT 154.800 490.200 155.600 490.400 ;
        RECT 152.600 489.600 153.600 490.200 ;
        RECT 154.200 489.600 155.600 490.200 ;
        RECT 152.600 482.200 153.400 489.600 ;
        RECT 154.200 488.400 154.800 489.600 ;
        RECT 154.000 487.600 154.800 488.400 ;
        RECT 158.000 482.200 158.800 493.700 ;
        RECT 159.600 493.600 160.400 493.700 ;
        RECT 162.600 493.600 165.200 494.400 ;
        RECT 161.200 491.600 162.000 493.200 ;
        RECT 162.600 492.300 163.200 493.600 ;
        RECT 166.000 492.300 166.800 492.400 ;
        RECT 162.600 491.700 166.800 492.300 ;
        RECT 162.600 490.200 163.200 491.700 ;
        RECT 166.000 491.600 166.800 491.700 ;
        RECT 167.400 490.800 168.200 495.200 ;
        RECT 169.200 494.600 170.000 499.800 ;
        RECT 175.600 496.600 176.400 499.800 ;
        RECT 177.200 497.000 178.000 499.800 ;
        RECT 178.800 497.000 179.600 499.800 ;
        RECT 180.400 497.000 181.200 499.800 ;
        RECT 182.000 497.000 182.800 499.800 ;
        RECT 185.200 497.000 186.000 499.800 ;
        RECT 188.400 497.000 189.200 499.800 ;
        RECT 190.000 497.000 190.800 499.800 ;
        RECT 191.600 497.000 192.400 499.800 ;
        RECT 174.000 495.800 176.400 496.600 ;
        RECT 193.200 496.600 194.000 499.800 ;
        RECT 174.000 495.200 174.800 495.800 ;
        RECT 168.800 494.000 170.000 494.600 ;
        RECT 173.000 494.600 174.800 495.200 ;
        RECT 178.800 495.600 179.800 496.400 ;
        RECT 182.800 495.600 184.400 496.400 ;
        RECT 185.200 495.800 189.800 496.400 ;
        RECT 193.200 495.800 195.800 496.600 ;
        RECT 185.200 495.600 186.000 495.800 ;
        RECT 168.800 492.000 169.400 494.000 ;
        RECT 173.000 493.400 173.800 494.600 ;
        RECT 170.000 492.600 173.800 493.400 ;
        RECT 178.800 492.800 179.600 495.600 ;
        RECT 185.200 494.800 186.000 495.000 ;
        RECT 181.600 494.200 186.000 494.800 ;
        RECT 181.600 494.000 182.400 494.200 ;
        RECT 186.800 493.600 187.600 495.200 ;
        RECT 189.000 493.400 189.800 495.800 ;
        RECT 195.000 495.200 195.800 495.800 ;
        RECT 195.000 494.400 198.000 495.200 ;
        RECT 199.600 493.800 200.400 499.800 ;
        RECT 201.200 495.600 202.000 497.200 ;
        RECT 182.000 492.600 185.200 493.400 ;
        RECT 189.000 492.600 191.000 493.400 ;
        RECT 191.600 493.000 200.400 493.800 ;
        RECT 175.600 492.000 176.400 492.600 ;
        RECT 193.200 492.000 194.000 492.400 ;
        RECT 198.000 492.200 198.800 492.400 ;
        RECT 198.000 492.000 199.000 492.200 ;
        RECT 168.800 491.400 169.600 492.000 ;
        RECT 175.600 491.400 199.000 492.000 ;
        RECT 164.400 490.200 165.200 490.400 ;
        RECT 162.200 489.600 163.200 490.200 ;
        RECT 163.800 489.600 165.200 490.200 ;
        RECT 167.400 490.000 168.400 490.800 ;
        RECT 162.200 482.200 163.000 489.600 ;
        RECT 163.800 488.400 164.400 489.600 ;
        RECT 163.600 487.600 164.400 488.400 ;
        RECT 167.600 482.200 168.400 490.000 ;
        RECT 169.000 489.600 169.600 491.400 ;
        RECT 169.000 489.000 178.000 489.600 ;
        RECT 169.000 487.400 169.600 489.000 ;
        RECT 177.200 488.800 178.000 489.000 ;
        RECT 180.400 489.000 189.000 489.600 ;
        RECT 180.400 488.800 181.200 489.000 ;
        RECT 172.200 487.600 174.800 488.400 ;
        RECT 169.000 486.800 171.600 487.400 ;
        RECT 170.800 482.200 171.600 486.800 ;
        RECT 174.000 482.200 174.800 487.600 ;
        RECT 175.400 486.800 179.600 487.600 ;
        RECT 177.200 482.200 178.000 485.000 ;
        RECT 178.800 482.200 179.600 485.000 ;
        RECT 180.400 482.200 181.200 485.000 ;
        RECT 182.000 482.200 182.800 488.400 ;
        RECT 185.200 487.600 187.800 488.400 ;
        RECT 188.400 488.200 189.000 489.000 ;
        RECT 190.000 489.400 190.800 489.600 ;
        RECT 190.000 489.000 195.400 489.400 ;
        RECT 190.000 488.800 196.200 489.000 ;
        RECT 194.800 488.200 196.200 488.800 ;
        RECT 188.400 487.600 194.200 488.200 ;
        RECT 197.200 488.000 198.800 488.800 ;
        RECT 197.200 487.600 197.800 488.000 ;
        RECT 185.200 482.200 186.000 487.000 ;
        RECT 188.400 482.200 189.200 487.000 ;
        RECT 193.600 486.800 197.800 487.600 ;
        RECT 199.600 487.400 200.400 493.000 ;
        RECT 198.400 486.800 200.400 487.400 ;
        RECT 202.800 494.300 203.600 499.800 ;
        RECT 206.000 496.000 206.800 499.800 ;
        RECT 205.800 495.200 206.800 496.000 ;
        RECT 204.400 494.300 205.200 494.400 ;
        RECT 202.800 493.700 205.200 494.300 ;
        RECT 190.000 482.200 190.800 485.000 ;
        RECT 191.600 482.200 192.400 485.000 ;
        RECT 194.800 482.200 195.600 486.800 ;
        RECT 198.400 486.200 199.000 486.800 ;
        RECT 198.000 485.600 199.000 486.200 ;
        RECT 198.000 482.200 198.800 485.600 ;
        RECT 202.800 482.200 203.600 493.700 ;
        RECT 204.400 493.600 205.200 493.700 ;
        RECT 205.800 490.800 206.600 495.200 ;
        RECT 207.600 494.600 208.400 499.800 ;
        RECT 214.000 496.600 214.800 499.800 ;
        RECT 215.600 497.000 216.400 499.800 ;
        RECT 217.200 497.000 218.000 499.800 ;
        RECT 218.800 497.000 219.600 499.800 ;
        RECT 220.400 497.000 221.200 499.800 ;
        RECT 223.600 497.000 224.400 499.800 ;
        RECT 226.800 497.000 227.600 499.800 ;
        RECT 228.400 497.000 229.200 499.800 ;
        RECT 230.000 497.000 230.800 499.800 ;
        RECT 212.400 495.800 214.800 496.600 ;
        RECT 231.600 496.600 232.400 499.800 ;
        RECT 212.400 495.200 213.200 495.800 ;
        RECT 207.200 494.000 208.400 494.600 ;
        RECT 211.400 494.600 213.200 495.200 ;
        RECT 217.200 495.600 218.200 496.400 ;
        RECT 221.200 495.600 222.800 496.400 ;
        RECT 223.600 495.800 228.200 496.400 ;
        RECT 231.600 495.800 234.200 496.600 ;
        RECT 223.600 495.600 224.400 495.800 ;
        RECT 207.200 492.000 207.800 494.000 ;
        RECT 211.400 493.400 212.200 494.600 ;
        RECT 208.400 492.600 212.200 493.400 ;
        RECT 217.200 492.800 218.000 495.600 ;
        RECT 223.600 494.800 224.400 495.000 ;
        RECT 220.000 494.200 224.400 494.800 ;
        RECT 220.000 494.000 220.800 494.200 ;
        RECT 225.200 493.600 226.000 495.200 ;
        RECT 227.400 493.400 228.200 495.800 ;
        RECT 233.400 495.200 234.200 495.800 ;
        RECT 233.400 494.400 236.400 495.200 ;
        RECT 238.000 493.800 238.800 499.800 ;
        RECT 241.200 495.200 242.000 499.800 ;
        RECT 244.400 495.200 245.200 499.800 ;
        RECT 247.600 495.200 248.400 499.800 ;
        RECT 250.800 495.200 251.600 499.800 ;
        RECT 220.400 492.600 223.600 493.400 ;
        RECT 227.400 492.600 229.400 493.400 ;
        RECT 230.000 493.000 238.800 493.800 ;
        RECT 214.000 492.000 214.800 492.600 ;
        RECT 231.600 492.000 232.400 492.400 ;
        RECT 236.400 492.200 237.200 492.400 ;
        RECT 236.400 492.000 237.400 492.200 ;
        RECT 207.200 491.400 208.000 492.000 ;
        RECT 214.000 491.400 237.400 492.000 ;
        RECT 205.800 490.000 206.800 490.800 ;
        RECT 206.000 482.200 206.800 490.000 ;
        RECT 207.400 489.600 208.000 491.400 ;
        RECT 207.400 489.000 216.400 489.600 ;
        RECT 207.400 487.400 208.000 489.000 ;
        RECT 215.600 488.800 216.400 489.000 ;
        RECT 218.800 489.000 227.400 489.600 ;
        RECT 218.800 488.800 219.600 489.000 ;
        RECT 210.600 487.600 213.200 488.400 ;
        RECT 207.400 486.800 210.000 487.400 ;
        RECT 209.200 482.200 210.000 486.800 ;
        RECT 212.400 482.200 213.200 487.600 ;
        RECT 213.800 486.800 218.000 487.600 ;
        RECT 215.600 482.200 216.400 485.000 ;
        RECT 217.200 482.200 218.000 485.000 ;
        RECT 218.800 482.200 219.600 485.000 ;
        RECT 220.400 482.200 221.200 488.400 ;
        RECT 223.600 487.600 226.200 488.400 ;
        RECT 226.800 488.200 227.400 489.000 ;
        RECT 228.400 489.400 229.200 489.600 ;
        RECT 228.400 489.000 233.800 489.400 ;
        RECT 228.400 488.800 234.600 489.000 ;
        RECT 233.200 488.200 234.600 488.800 ;
        RECT 226.800 487.600 232.600 488.200 ;
        RECT 235.600 488.000 237.200 488.800 ;
        RECT 235.600 487.600 236.200 488.000 ;
        RECT 223.600 482.200 224.400 487.000 ;
        RECT 226.800 482.200 227.600 487.000 ;
        RECT 232.000 486.800 236.200 487.600 ;
        RECT 238.000 487.400 238.800 493.000 ;
        RECT 239.600 494.400 242.000 495.200 ;
        RECT 243.000 494.400 245.200 495.200 ;
        RECT 246.200 494.400 248.400 495.200 ;
        RECT 249.800 494.400 251.600 495.200 ;
        RECT 239.600 491.600 240.400 494.400 ;
        RECT 243.000 493.800 243.800 494.400 ;
        RECT 246.200 493.800 247.000 494.400 ;
        RECT 249.800 493.800 250.600 494.400 ;
        RECT 252.400 493.800 253.200 494.400 ;
        RECT 241.200 493.000 243.800 493.800 ;
        RECT 244.600 493.000 247.000 493.800 ;
        RECT 248.000 493.000 250.600 493.800 ;
        RECT 251.400 493.000 253.200 493.800 ;
        RECT 258.800 493.800 259.600 499.800 ;
        RECT 265.200 496.600 266.000 499.800 ;
        RECT 266.800 497.000 267.600 499.800 ;
        RECT 268.400 497.000 269.200 499.800 ;
        RECT 270.000 497.000 270.800 499.800 ;
        RECT 273.200 497.000 274.000 499.800 ;
        RECT 276.400 497.000 277.200 499.800 ;
        RECT 278.000 497.000 278.800 499.800 ;
        RECT 279.600 497.000 280.400 499.800 ;
        RECT 281.200 497.000 282.000 499.800 ;
        RECT 263.400 495.800 266.000 496.600 ;
        RECT 282.800 496.600 283.600 499.800 ;
        RECT 269.400 495.800 274.000 496.400 ;
        RECT 263.400 495.200 264.200 495.800 ;
        RECT 261.200 494.400 264.200 495.200 ;
        RECT 258.800 493.000 267.600 493.800 ;
        RECT 269.400 493.400 270.200 495.800 ;
        RECT 273.200 495.600 274.000 495.800 ;
        RECT 274.800 495.600 276.400 496.400 ;
        RECT 279.400 495.600 280.400 496.400 ;
        RECT 282.800 495.800 285.200 496.600 ;
        RECT 271.600 493.600 272.400 495.200 ;
        RECT 273.200 494.800 274.000 495.000 ;
        RECT 273.200 494.200 277.600 494.800 ;
        RECT 276.800 494.000 277.600 494.200 ;
        RECT 243.000 491.600 243.800 493.000 ;
        RECT 246.200 491.600 247.000 493.000 ;
        RECT 249.800 491.600 250.600 493.000 ;
        RECT 239.600 490.800 242.000 491.600 ;
        RECT 243.000 490.800 245.200 491.600 ;
        RECT 246.200 490.800 248.400 491.600 ;
        RECT 249.800 490.800 251.600 491.600 ;
        RECT 236.800 486.800 238.800 487.400 ;
        RECT 228.400 482.200 229.200 485.000 ;
        RECT 230.000 482.200 230.800 485.000 ;
        RECT 233.200 482.200 234.000 486.800 ;
        RECT 236.800 486.200 237.400 486.800 ;
        RECT 236.400 485.600 237.400 486.200 ;
        RECT 236.400 482.200 237.200 485.600 ;
        RECT 241.200 482.200 242.000 490.800 ;
        RECT 244.400 482.200 245.200 490.800 ;
        RECT 247.600 482.200 248.400 490.800 ;
        RECT 250.800 482.200 251.600 490.800 ;
        RECT 258.800 487.400 259.600 493.000 ;
        RECT 268.200 492.600 270.200 493.400 ;
        RECT 274.000 492.600 277.200 493.400 ;
        RECT 279.600 492.800 280.400 495.600 ;
        RECT 284.400 495.200 285.200 495.800 ;
        RECT 284.400 494.600 286.200 495.200 ;
        RECT 285.400 493.400 286.200 494.600 ;
        RECT 289.200 494.600 290.000 499.800 ;
        RECT 290.800 496.000 291.600 499.800 ;
        RECT 290.800 495.200 291.800 496.000 ;
        RECT 289.200 494.000 290.400 494.600 ;
        RECT 285.400 492.600 289.200 493.400 ;
        RECT 260.200 492.000 261.000 492.200 ;
        RECT 262.000 492.000 262.800 492.400 ;
        RECT 265.200 492.000 266.000 492.400 ;
        RECT 282.800 492.000 283.600 492.600 ;
        RECT 289.800 492.000 290.400 494.000 ;
        RECT 260.200 491.400 283.600 492.000 ;
        RECT 289.600 491.400 290.400 492.000 ;
        RECT 291.000 492.300 291.800 495.200 ;
        RECT 294.000 495.200 294.800 499.800 ;
        RECT 294.000 494.600 296.200 495.200 ;
        RECT 294.000 492.300 294.800 493.200 ;
        RECT 291.000 491.700 294.800 492.300 ;
        RECT 289.600 489.600 290.200 491.400 ;
        RECT 291.000 490.800 291.800 491.700 ;
        RECT 294.000 491.600 294.800 491.700 ;
        RECT 295.600 491.600 296.200 494.600 ;
        RECT 298.800 493.800 299.600 499.800 ;
        RECT 305.200 496.600 306.000 499.800 ;
        RECT 306.800 497.000 307.600 499.800 ;
        RECT 308.400 497.000 309.200 499.800 ;
        RECT 310.000 497.000 310.800 499.800 ;
        RECT 313.200 497.000 314.000 499.800 ;
        RECT 316.400 497.000 317.200 499.800 ;
        RECT 318.000 497.000 318.800 499.800 ;
        RECT 319.600 497.000 320.400 499.800 ;
        RECT 321.200 497.000 322.000 499.800 ;
        RECT 303.400 495.800 306.000 496.600 ;
        RECT 322.800 496.600 323.600 499.800 ;
        RECT 309.400 495.800 314.000 496.400 ;
        RECT 303.400 495.200 304.200 495.800 ;
        RECT 301.200 494.400 304.200 495.200 ;
        RECT 298.800 493.000 307.600 493.800 ;
        RECT 309.400 493.400 310.200 495.800 ;
        RECT 313.200 495.600 314.000 495.800 ;
        RECT 314.800 495.600 316.400 496.400 ;
        RECT 319.400 495.600 320.400 496.400 ;
        RECT 322.800 495.800 325.200 496.600 ;
        RECT 311.600 493.600 312.400 495.200 ;
        RECT 313.200 494.800 314.000 495.000 ;
        RECT 313.200 494.200 317.600 494.800 ;
        RECT 316.800 494.000 317.600 494.200 ;
        RECT 268.400 489.400 269.200 489.600 ;
        RECT 263.800 489.000 269.200 489.400 ;
        RECT 263.000 488.800 269.200 489.000 ;
        RECT 270.200 489.000 278.800 489.600 ;
        RECT 260.400 488.000 262.000 488.800 ;
        RECT 263.000 488.200 264.400 488.800 ;
        RECT 270.200 488.200 270.800 489.000 ;
        RECT 278.000 488.800 278.800 489.000 ;
        RECT 281.200 489.000 290.200 489.600 ;
        RECT 281.200 488.800 282.000 489.000 ;
        RECT 261.400 487.600 262.000 488.000 ;
        RECT 265.000 487.600 270.800 488.200 ;
        RECT 271.400 487.600 274.000 488.400 ;
        RECT 258.800 486.800 260.800 487.400 ;
        RECT 261.400 486.800 265.600 487.600 ;
        RECT 260.200 486.200 260.800 486.800 ;
        RECT 260.200 485.600 261.200 486.200 ;
        RECT 260.400 482.200 261.200 485.600 ;
        RECT 263.600 482.200 264.400 486.800 ;
        RECT 266.800 482.200 267.600 485.000 ;
        RECT 268.400 482.200 269.200 485.000 ;
        RECT 270.000 482.200 270.800 487.000 ;
        RECT 273.200 482.200 274.000 487.000 ;
        RECT 276.400 482.200 277.200 488.400 ;
        RECT 284.400 487.600 287.000 488.400 ;
        RECT 279.600 486.800 283.800 487.600 ;
        RECT 278.000 482.200 278.800 485.000 ;
        RECT 279.600 482.200 280.400 485.000 ;
        RECT 281.200 482.200 282.000 485.000 ;
        RECT 284.400 482.200 285.200 487.600 ;
        RECT 289.600 487.400 290.200 489.000 ;
        RECT 287.600 486.800 290.200 487.400 ;
        RECT 290.800 490.000 291.800 490.800 ;
        RECT 295.600 490.800 296.800 491.600 ;
        RECT 295.600 490.200 296.200 490.800 ;
        RECT 287.600 482.200 288.400 486.800 ;
        RECT 290.800 482.200 291.600 490.000 ;
        RECT 294.000 489.600 296.200 490.200 ;
        RECT 294.000 482.200 294.800 489.600 ;
        RECT 298.800 487.400 299.600 493.000 ;
        RECT 308.200 492.600 310.200 493.400 ;
        RECT 314.000 492.600 317.200 493.400 ;
        RECT 319.600 492.800 320.400 495.600 ;
        RECT 324.400 495.200 325.200 495.800 ;
        RECT 324.400 494.600 326.200 495.200 ;
        RECT 325.400 493.400 326.200 494.600 ;
        RECT 329.200 494.600 330.000 499.800 ;
        RECT 330.800 496.000 331.600 499.800 ;
        RECT 330.800 495.200 331.800 496.000 ;
        RECT 334.000 495.800 334.800 499.800 ;
        RECT 338.400 496.200 340.000 499.800 ;
        RECT 334.000 495.200 336.200 495.800 ;
        RECT 337.200 495.400 338.800 495.600 ;
        RECT 329.200 494.000 330.400 494.600 ;
        RECT 325.400 492.600 329.200 493.400 ;
        RECT 300.200 492.000 301.000 492.200 ;
        RECT 302.000 492.000 302.800 492.400 ;
        RECT 305.200 492.000 306.000 492.400 ;
        RECT 322.800 492.000 323.600 492.600 ;
        RECT 329.800 492.000 330.400 494.000 ;
        RECT 300.200 491.400 323.600 492.000 ;
        RECT 329.600 491.400 330.400 492.000 ;
        RECT 329.600 489.600 330.200 491.400 ;
        RECT 331.000 490.800 331.800 495.200 ;
        RECT 335.400 495.000 336.200 495.200 ;
        RECT 336.800 494.800 338.800 495.400 ;
        RECT 336.800 494.400 337.400 494.800 ;
        RECT 334.000 493.800 337.400 494.400 ;
        RECT 334.000 493.600 335.600 493.800 ;
        RECT 338.000 493.400 338.800 494.200 ;
        RECT 338.000 492.800 338.600 493.400 ;
        RECT 336.000 492.200 338.600 492.800 ;
        RECT 339.400 492.800 340.000 496.200 ;
        RECT 343.600 495.800 344.400 499.800 ;
        RECT 346.800 496.000 347.600 499.800 ;
        RECT 340.600 494.800 341.400 495.600 ;
        RECT 342.000 495.200 344.400 495.800 ;
        RECT 346.600 495.200 347.600 496.000 ;
        RECT 342.000 495.000 342.800 495.200 ;
        RECT 340.800 494.400 341.400 494.800 ;
        RECT 340.800 493.600 341.600 494.400 ;
        RECT 342.800 494.300 344.400 494.400 ;
        RECT 346.600 494.300 347.400 495.200 ;
        RECT 348.400 494.600 349.200 499.800 ;
        RECT 354.800 496.600 355.600 499.800 ;
        RECT 356.400 497.000 357.200 499.800 ;
        RECT 358.000 497.000 358.800 499.800 ;
        RECT 359.600 497.000 360.400 499.800 ;
        RECT 361.200 497.000 362.000 499.800 ;
        RECT 364.400 497.000 365.200 499.800 ;
        RECT 367.600 497.000 368.400 499.800 ;
        RECT 369.200 497.000 370.000 499.800 ;
        RECT 370.800 497.000 371.600 499.800 ;
        RECT 353.200 495.800 355.600 496.600 ;
        RECT 372.400 496.600 373.200 499.800 ;
        RECT 353.200 495.200 354.000 495.800 ;
        RECT 342.800 493.700 347.400 494.300 ;
        RECT 342.800 493.600 344.400 493.700 ;
        RECT 339.400 492.400 340.400 492.800 ;
        RECT 339.400 492.300 341.200 492.400 ;
        RECT 345.200 492.300 346.000 492.400 ;
        RECT 339.400 492.200 346.000 492.300 ;
        RECT 336.000 492.000 336.800 492.200 ;
        RECT 339.800 491.700 346.000 492.200 ;
        RECT 339.800 491.600 341.200 491.700 ;
        RECT 345.200 491.600 346.000 491.700 ;
        RECT 338.200 491.400 339.000 491.600 ;
        RECT 308.400 489.400 309.200 489.600 ;
        RECT 303.800 489.000 309.200 489.400 ;
        RECT 303.000 488.800 309.200 489.000 ;
        RECT 310.200 489.000 318.800 489.600 ;
        RECT 300.400 488.000 302.000 488.800 ;
        RECT 303.000 488.200 304.400 488.800 ;
        RECT 310.200 488.200 310.800 489.000 ;
        RECT 318.000 488.800 318.800 489.000 ;
        RECT 321.200 489.000 330.200 489.600 ;
        RECT 321.200 488.800 322.000 489.000 ;
        RECT 301.400 487.600 302.000 488.000 ;
        RECT 305.000 487.600 310.800 488.200 ;
        RECT 311.400 487.600 314.000 488.400 ;
        RECT 298.800 486.800 300.800 487.400 ;
        RECT 301.400 486.800 305.600 487.600 ;
        RECT 300.200 486.200 300.800 486.800 ;
        RECT 300.200 485.600 301.200 486.200 ;
        RECT 300.400 482.200 301.200 485.600 ;
        RECT 303.600 482.200 304.400 486.800 ;
        RECT 306.800 482.200 307.600 485.000 ;
        RECT 308.400 482.200 309.200 485.000 ;
        RECT 310.000 482.200 310.800 487.000 ;
        RECT 313.200 482.200 314.000 487.000 ;
        RECT 316.400 482.200 317.200 488.400 ;
        RECT 324.400 487.600 327.000 488.400 ;
        RECT 319.600 486.800 323.800 487.600 ;
        RECT 318.000 482.200 318.800 485.000 ;
        RECT 319.600 482.200 320.400 485.000 ;
        RECT 321.200 482.200 322.000 485.000 ;
        RECT 324.400 482.200 325.200 487.600 ;
        RECT 329.600 487.400 330.200 489.000 ;
        RECT 327.600 486.800 330.200 487.400 ;
        RECT 330.800 490.000 331.800 490.800 ;
        RECT 335.600 490.800 339.000 491.400 ;
        RECT 335.600 490.200 336.200 490.800 ;
        RECT 339.800 490.200 340.400 491.600 ;
        RECT 346.600 490.800 347.400 493.700 ;
        RECT 348.000 494.000 349.200 494.600 ;
        RECT 352.200 494.600 354.000 495.200 ;
        RECT 358.000 495.600 359.000 496.400 ;
        RECT 362.000 495.600 363.600 496.400 ;
        RECT 364.400 495.800 369.000 496.400 ;
        RECT 372.400 495.800 375.000 496.600 ;
        RECT 364.400 495.600 365.200 495.800 ;
        RECT 348.000 492.000 348.600 494.000 ;
        RECT 352.200 493.400 353.000 494.600 ;
        RECT 349.200 492.600 353.000 493.400 ;
        RECT 358.000 492.800 358.800 495.600 ;
        RECT 364.400 494.800 365.200 495.000 ;
        RECT 360.800 494.200 365.200 494.800 ;
        RECT 360.800 494.000 361.600 494.200 ;
        RECT 366.000 493.600 366.800 495.200 ;
        RECT 368.200 493.400 369.000 495.800 ;
        RECT 374.200 495.200 375.000 495.800 ;
        RECT 374.200 494.400 377.200 495.200 ;
        RECT 378.800 493.800 379.600 499.800 ;
        RECT 383.600 495.200 384.400 499.800 ;
        RECT 386.800 496.000 387.600 499.800 ;
        RECT 361.200 492.600 364.400 493.400 ;
        RECT 368.200 492.600 370.200 493.400 ;
        RECT 370.800 493.000 379.600 493.800 ;
        RECT 354.800 492.000 355.600 492.600 ;
        RECT 372.400 492.000 373.200 492.400 ;
        RECT 377.400 492.000 378.200 492.200 ;
        RECT 348.000 491.400 348.800 492.000 ;
        RECT 354.800 491.400 378.200 492.000 ;
        RECT 327.600 482.200 328.400 486.800 ;
        RECT 330.800 482.200 331.600 490.000 ;
        RECT 334.000 489.600 336.200 490.200 ;
        RECT 334.000 482.200 334.800 489.600 ;
        RECT 335.400 489.400 336.200 489.600 ;
        RECT 338.400 489.600 340.400 490.200 ;
        RECT 342.000 489.600 344.400 490.200 ;
        RECT 346.600 490.000 347.600 490.800 ;
        RECT 338.400 482.200 340.000 489.600 ;
        RECT 342.000 489.400 342.800 489.600 ;
        RECT 343.600 482.200 344.400 489.600 ;
        RECT 346.800 482.200 347.600 490.000 ;
        RECT 348.200 489.600 348.800 491.400 ;
        RECT 348.200 489.000 357.200 489.600 ;
        RECT 348.200 487.400 348.800 489.000 ;
        RECT 356.400 488.800 357.200 489.000 ;
        RECT 359.600 489.000 368.200 489.600 ;
        RECT 359.600 488.800 360.400 489.000 ;
        RECT 351.400 487.600 354.000 488.400 ;
        RECT 348.200 486.800 350.800 487.400 ;
        RECT 350.000 482.200 350.800 486.800 ;
        RECT 353.200 482.200 354.000 487.600 ;
        RECT 354.600 486.800 358.800 487.600 ;
        RECT 356.400 482.200 357.200 485.000 ;
        RECT 358.000 482.200 358.800 485.000 ;
        RECT 359.600 482.200 360.400 485.000 ;
        RECT 361.200 482.200 362.000 488.400 ;
        RECT 364.400 487.600 367.000 488.400 ;
        RECT 367.600 488.200 368.200 489.000 ;
        RECT 369.200 489.400 370.000 489.600 ;
        RECT 369.200 489.000 374.600 489.400 ;
        RECT 369.200 488.800 375.400 489.000 ;
        RECT 374.000 488.200 375.400 488.800 ;
        RECT 367.600 487.600 373.400 488.200 ;
        RECT 376.400 488.000 378.000 488.800 ;
        RECT 376.400 487.600 377.000 488.000 ;
        RECT 364.400 482.200 365.200 487.000 ;
        RECT 367.600 482.200 368.400 487.000 ;
        RECT 372.800 486.800 377.000 487.600 ;
        RECT 378.800 487.400 379.600 493.000 ;
        RECT 382.200 494.600 384.400 495.200 ;
        RECT 386.600 495.200 387.600 496.000 ;
        RECT 382.200 491.600 382.800 494.600 ;
        RECT 383.600 492.300 384.400 493.200 ;
        RECT 386.600 492.300 387.400 495.200 ;
        RECT 388.400 494.600 389.200 499.800 ;
        RECT 394.800 496.600 395.600 499.800 ;
        RECT 396.400 497.000 397.200 499.800 ;
        RECT 398.000 497.000 398.800 499.800 ;
        RECT 399.600 497.000 400.400 499.800 ;
        RECT 401.200 497.000 402.000 499.800 ;
        RECT 404.400 497.000 405.200 499.800 ;
        RECT 407.600 497.000 408.400 499.800 ;
        RECT 409.200 497.000 410.000 499.800 ;
        RECT 410.800 497.000 411.600 499.800 ;
        RECT 393.200 495.800 395.600 496.600 ;
        RECT 412.400 496.600 413.200 499.800 ;
        RECT 393.200 495.200 394.000 495.800 ;
        RECT 383.600 491.700 387.400 492.300 ;
        RECT 383.600 491.600 384.400 491.700 ;
        RECT 381.600 490.800 382.800 491.600 ;
        RECT 382.200 490.200 382.800 490.800 ;
        RECT 386.600 490.800 387.400 491.700 ;
        RECT 388.000 494.000 389.200 494.600 ;
        RECT 392.200 494.600 394.000 495.200 ;
        RECT 398.000 495.600 399.000 496.400 ;
        RECT 402.000 495.600 403.600 496.400 ;
        RECT 404.400 495.800 409.000 496.400 ;
        RECT 412.400 495.800 415.000 496.600 ;
        RECT 404.400 495.600 405.200 495.800 ;
        RECT 388.000 492.000 388.600 494.000 ;
        RECT 392.200 493.400 393.000 494.600 ;
        RECT 389.200 492.600 393.000 493.400 ;
        RECT 398.000 492.800 398.800 495.600 ;
        RECT 404.400 494.800 405.200 495.000 ;
        RECT 400.800 494.200 405.200 494.800 ;
        RECT 400.800 494.000 401.600 494.200 ;
        RECT 406.000 493.600 406.800 495.200 ;
        RECT 408.200 493.400 409.000 495.800 ;
        RECT 414.200 495.200 415.000 495.800 ;
        RECT 414.200 494.400 417.200 495.200 ;
        RECT 418.800 493.800 419.600 499.800 ;
        RECT 425.200 495.200 426.000 499.800 ;
        RECT 430.000 495.600 430.800 497.200 ;
        RECT 425.200 494.600 427.400 495.200 ;
        RECT 401.200 492.600 404.400 493.400 ;
        RECT 408.200 492.600 410.200 493.400 ;
        RECT 410.800 493.000 419.600 493.800 ;
        RECT 394.800 492.000 395.600 492.600 ;
        RECT 406.000 492.000 406.800 492.400 ;
        RECT 412.400 492.000 413.200 492.400 ;
        RECT 417.400 492.000 418.200 492.200 ;
        RECT 388.000 491.400 388.800 492.000 ;
        RECT 394.800 491.400 418.200 492.000 ;
        RECT 382.200 489.600 384.400 490.200 ;
        RECT 386.600 490.000 387.600 490.800 ;
        RECT 377.600 486.800 379.600 487.400 ;
        RECT 369.200 482.200 370.000 485.000 ;
        RECT 370.800 482.200 371.600 485.000 ;
        RECT 374.000 482.200 374.800 486.800 ;
        RECT 377.600 486.200 378.200 486.800 ;
        RECT 377.200 485.600 378.200 486.200 ;
        RECT 377.200 482.200 378.000 485.600 ;
        RECT 383.600 482.200 384.400 489.600 ;
        RECT 386.800 482.200 387.600 490.000 ;
        RECT 388.200 489.600 388.800 491.400 ;
        RECT 388.200 489.000 397.200 489.600 ;
        RECT 388.200 487.400 388.800 489.000 ;
        RECT 396.400 488.800 397.200 489.000 ;
        RECT 399.600 489.000 408.200 489.600 ;
        RECT 399.600 488.800 400.400 489.000 ;
        RECT 391.400 487.600 394.000 488.400 ;
        RECT 388.200 486.800 390.800 487.400 ;
        RECT 390.000 482.200 390.800 486.800 ;
        RECT 393.200 482.200 394.000 487.600 ;
        RECT 394.600 486.800 398.800 487.600 ;
        RECT 396.400 482.200 397.200 485.000 ;
        RECT 398.000 482.200 398.800 485.000 ;
        RECT 399.600 482.200 400.400 485.000 ;
        RECT 401.200 482.200 402.000 488.400 ;
        RECT 404.400 487.600 407.000 488.400 ;
        RECT 407.600 488.200 408.200 489.000 ;
        RECT 409.200 489.400 410.000 489.600 ;
        RECT 409.200 489.000 414.600 489.400 ;
        RECT 409.200 488.800 415.400 489.000 ;
        RECT 414.000 488.200 415.400 488.800 ;
        RECT 407.600 487.600 413.400 488.200 ;
        RECT 416.400 488.000 418.000 488.800 ;
        RECT 416.400 487.600 417.000 488.000 ;
        RECT 404.400 482.200 405.200 487.000 ;
        RECT 407.600 482.200 408.400 487.000 ;
        RECT 412.800 486.800 417.000 487.600 ;
        RECT 418.800 487.400 419.600 493.000 ;
        RECT 422.000 492.300 422.800 492.400 ;
        RECT 425.200 492.300 426.000 493.200 ;
        RECT 422.000 491.700 426.000 492.300 ;
        RECT 422.000 491.600 422.800 491.700 ;
        RECT 425.200 491.600 426.000 491.700 ;
        RECT 426.800 491.600 427.400 494.600 ;
        RECT 431.600 492.300 432.400 499.800 ;
        RECT 433.200 496.000 434.000 499.800 ;
        RECT 436.400 496.000 437.200 499.800 ;
        RECT 433.200 495.800 437.200 496.000 ;
        RECT 438.000 495.800 438.800 499.800 ;
        RECT 442.200 496.400 443.000 499.800 ;
        RECT 441.200 495.800 443.000 496.400 ;
        RECT 446.000 496.000 446.800 499.800 ;
        RECT 433.400 495.400 437.000 495.800 ;
        RECT 434.000 494.400 434.800 494.800 ;
        RECT 438.000 494.400 438.600 495.800 ;
        RECT 433.200 493.800 434.800 494.400 ;
        RECT 433.200 493.600 434.000 493.800 ;
        RECT 436.200 493.600 438.800 494.400 ;
        RECT 439.600 493.600 440.400 495.200 ;
        RECT 434.800 492.300 435.600 493.200 ;
        RECT 431.600 491.700 435.600 492.300 ;
        RECT 426.800 490.800 428.000 491.600 ;
        RECT 426.800 490.200 427.400 490.800 ;
        RECT 417.600 486.800 419.600 487.400 ;
        RECT 425.200 489.600 427.400 490.200 ;
        RECT 409.200 482.200 410.000 485.000 ;
        RECT 410.800 482.200 411.600 485.000 ;
        RECT 414.000 482.200 414.800 486.800 ;
        RECT 417.600 486.200 418.200 486.800 ;
        RECT 417.200 485.600 418.200 486.200 ;
        RECT 417.200 482.200 418.000 485.600 ;
        RECT 425.200 482.200 426.000 489.600 ;
        RECT 431.600 482.200 432.400 491.700 ;
        RECT 434.800 491.600 435.600 491.700 ;
        RECT 436.200 492.400 436.800 493.600 ;
        RECT 436.200 491.600 437.200 492.400 ;
        RECT 436.200 490.200 436.800 491.600 ;
        RECT 438.000 490.300 438.800 490.400 ;
        RECT 441.200 490.300 442.000 495.800 ;
        RECT 445.800 495.200 446.800 496.000 ;
        RECT 445.800 490.800 446.600 495.200 ;
        RECT 447.600 494.600 448.400 499.800 ;
        RECT 454.000 496.600 454.800 499.800 ;
        RECT 455.600 497.000 456.400 499.800 ;
        RECT 457.200 497.000 458.000 499.800 ;
        RECT 458.800 497.000 459.600 499.800 ;
        RECT 460.400 497.000 461.200 499.800 ;
        RECT 463.600 497.000 464.400 499.800 ;
        RECT 466.800 497.000 467.600 499.800 ;
        RECT 468.400 497.000 469.200 499.800 ;
        RECT 470.000 497.000 470.800 499.800 ;
        RECT 452.400 495.800 454.800 496.600 ;
        RECT 471.600 496.600 472.400 499.800 ;
        RECT 452.400 495.200 453.200 495.800 ;
        RECT 447.200 494.000 448.400 494.600 ;
        RECT 451.400 494.600 453.200 495.200 ;
        RECT 457.200 495.600 458.200 496.400 ;
        RECT 461.200 495.600 462.800 496.400 ;
        RECT 463.600 495.800 468.200 496.400 ;
        RECT 471.600 495.800 474.200 496.600 ;
        RECT 463.600 495.600 464.400 495.800 ;
        RECT 447.200 492.000 447.800 494.000 ;
        RECT 451.400 493.400 452.200 494.600 ;
        RECT 448.400 492.600 452.200 493.400 ;
        RECT 457.200 492.800 458.000 495.600 ;
        RECT 463.600 494.800 464.400 495.000 ;
        RECT 460.000 494.200 464.400 494.800 ;
        RECT 460.000 494.000 460.800 494.200 ;
        RECT 465.200 493.600 466.000 495.200 ;
        RECT 467.400 493.400 468.200 495.800 ;
        RECT 473.400 495.200 474.200 495.800 ;
        RECT 473.400 494.400 476.400 495.200 ;
        RECT 478.000 493.800 478.800 499.800 ;
        RECT 460.400 492.600 463.600 493.400 ;
        RECT 467.400 492.600 469.400 493.400 ;
        RECT 470.000 493.000 478.800 493.800 ;
        RECT 454.000 492.000 454.800 492.600 ;
        RECT 471.600 492.000 472.400 492.400 ;
        RECT 476.600 492.000 477.400 492.200 ;
        RECT 447.200 491.400 448.000 492.000 ;
        RECT 454.000 491.400 477.400 492.000 ;
        RECT 438.000 490.200 442.000 490.300 ;
        RECT 435.800 489.600 436.800 490.200 ;
        RECT 437.400 489.700 442.000 490.200 ;
        RECT 437.400 489.600 438.800 489.700 ;
        RECT 435.800 482.200 436.600 489.600 ;
        RECT 437.400 488.400 438.000 489.600 ;
        RECT 437.200 487.600 438.000 488.400 ;
        RECT 441.200 482.200 442.000 489.700 ;
        RECT 442.800 490.300 443.600 490.400 ;
        RECT 445.800 490.300 446.800 490.800 ;
        RECT 442.800 489.700 446.800 490.300 ;
        RECT 442.800 488.800 443.600 489.700 ;
        RECT 446.000 482.200 446.800 489.700 ;
        RECT 447.400 489.600 448.000 491.400 ;
        RECT 447.400 489.000 456.400 489.600 ;
        RECT 447.400 487.400 448.000 489.000 ;
        RECT 455.600 488.800 456.400 489.000 ;
        RECT 458.800 489.000 467.400 489.600 ;
        RECT 458.800 488.800 459.600 489.000 ;
        RECT 450.600 487.600 453.200 488.400 ;
        RECT 447.400 486.800 450.000 487.400 ;
        RECT 449.200 482.200 450.000 486.800 ;
        RECT 452.400 482.200 453.200 487.600 ;
        RECT 453.800 486.800 458.000 487.600 ;
        RECT 455.600 482.200 456.400 485.000 ;
        RECT 457.200 482.200 458.000 485.000 ;
        RECT 458.800 482.200 459.600 485.000 ;
        RECT 460.400 482.200 461.200 488.400 ;
        RECT 463.600 487.600 466.200 488.400 ;
        RECT 466.800 488.200 467.400 489.000 ;
        RECT 468.400 489.400 469.200 489.600 ;
        RECT 468.400 489.000 473.800 489.400 ;
        RECT 468.400 488.800 474.600 489.000 ;
        RECT 473.200 488.200 474.600 488.800 ;
        RECT 466.800 487.600 472.600 488.200 ;
        RECT 475.600 488.000 477.200 488.800 ;
        RECT 475.600 487.600 476.200 488.000 ;
        RECT 463.600 482.200 464.400 487.000 ;
        RECT 466.800 482.200 467.600 487.000 ;
        RECT 472.000 486.800 476.200 487.600 ;
        RECT 478.000 487.400 478.800 493.000 ;
        RECT 476.800 486.800 478.800 487.400 ;
        RECT 468.400 482.200 469.200 485.000 ;
        RECT 470.000 482.200 470.800 485.000 ;
        RECT 473.200 482.200 474.000 486.800 ;
        RECT 476.800 486.200 477.400 486.800 ;
        RECT 476.400 485.600 477.400 486.200 ;
        RECT 476.400 482.200 477.200 485.600 ;
        RECT 481.200 482.200 482.000 499.800 ;
        RECT 482.800 482.200 483.600 499.800 ;
        RECT 486.000 495.200 486.800 499.800 ;
        RECT 492.400 496.000 493.200 499.800 ;
        RECT 492.200 495.200 493.200 496.000 ;
        RECT 486.000 494.600 488.200 495.200 ;
        RECT 486.000 491.600 486.800 493.200 ;
        RECT 487.600 491.600 488.200 494.600 ;
        RECT 487.600 490.800 488.800 491.600 ;
        RECT 492.200 490.800 493.000 495.200 ;
        RECT 494.000 494.600 494.800 499.800 ;
        RECT 500.400 496.600 501.200 499.800 ;
        RECT 502.000 497.000 502.800 499.800 ;
        RECT 503.600 497.000 504.400 499.800 ;
        RECT 505.200 497.000 506.000 499.800 ;
        RECT 506.800 497.000 507.600 499.800 ;
        RECT 510.000 497.000 510.800 499.800 ;
        RECT 513.200 497.000 514.000 499.800 ;
        RECT 514.800 497.000 515.600 499.800 ;
        RECT 516.400 497.000 517.200 499.800 ;
        RECT 498.800 495.800 501.200 496.600 ;
        RECT 518.000 496.600 518.800 499.800 ;
        RECT 498.800 495.200 499.600 495.800 ;
        RECT 493.600 494.000 494.800 494.600 ;
        RECT 497.800 494.600 499.600 495.200 ;
        RECT 503.600 495.600 504.600 496.400 ;
        RECT 507.600 495.600 509.200 496.400 ;
        RECT 510.000 495.800 514.600 496.400 ;
        RECT 518.000 495.800 520.600 496.600 ;
        RECT 510.000 495.600 510.800 495.800 ;
        RECT 493.600 492.000 494.200 494.000 ;
        RECT 497.800 493.400 498.600 494.600 ;
        RECT 494.800 492.600 498.600 493.400 ;
        RECT 503.600 492.800 504.400 495.600 ;
        RECT 510.000 494.800 510.800 495.000 ;
        RECT 506.400 494.200 510.800 494.800 ;
        RECT 506.400 494.000 507.200 494.200 ;
        RECT 511.600 493.600 512.400 495.200 ;
        RECT 513.800 493.400 514.600 495.800 ;
        RECT 519.800 495.200 520.600 495.800 ;
        RECT 519.800 494.400 522.800 495.200 ;
        RECT 524.400 493.800 525.200 499.800 ;
        RECT 526.000 495.600 526.800 497.200 ;
        RECT 506.800 492.600 510.000 493.400 ;
        RECT 513.800 492.600 515.800 493.400 ;
        RECT 516.400 493.000 525.200 493.800 ;
        RECT 500.400 492.000 501.200 492.600 ;
        RECT 518.000 492.000 518.800 492.400 ;
        RECT 522.800 492.200 523.600 492.400 ;
        RECT 522.800 492.000 523.800 492.200 ;
        RECT 493.600 491.400 494.400 492.000 ;
        RECT 500.400 491.400 523.800 492.000 ;
        RECT 487.600 490.200 488.200 490.800 ;
        RECT 486.000 489.600 488.200 490.200 ;
        RECT 492.200 490.000 493.200 490.800 ;
        RECT 486.000 482.200 486.800 489.600 ;
        RECT 492.400 482.200 493.200 490.000 ;
        RECT 493.800 489.600 494.400 491.400 ;
        RECT 493.800 489.000 502.800 489.600 ;
        RECT 493.800 487.400 494.400 489.000 ;
        RECT 502.000 488.800 502.800 489.000 ;
        RECT 505.200 489.000 513.800 489.600 ;
        RECT 505.200 488.800 506.000 489.000 ;
        RECT 497.000 487.600 499.600 488.400 ;
        RECT 493.800 486.800 496.400 487.400 ;
        RECT 495.600 482.200 496.400 486.800 ;
        RECT 498.800 482.200 499.600 487.600 ;
        RECT 500.200 486.800 504.400 487.600 ;
        RECT 502.000 482.200 502.800 485.000 ;
        RECT 503.600 482.200 504.400 485.000 ;
        RECT 505.200 482.200 506.000 485.000 ;
        RECT 506.800 482.200 507.600 488.400 ;
        RECT 510.000 487.600 512.600 488.400 ;
        RECT 513.200 488.200 513.800 489.000 ;
        RECT 514.800 489.400 515.600 489.600 ;
        RECT 514.800 489.000 520.200 489.400 ;
        RECT 514.800 488.800 521.000 489.000 ;
        RECT 519.600 488.200 521.000 488.800 ;
        RECT 513.200 487.600 519.000 488.200 ;
        RECT 522.000 488.000 523.600 488.800 ;
        RECT 522.000 487.600 522.600 488.000 ;
        RECT 510.000 482.200 510.800 487.000 ;
        RECT 513.200 482.200 514.000 487.000 ;
        RECT 518.400 486.800 522.600 487.600 ;
        RECT 524.400 487.400 525.200 493.000 ;
        RECT 523.200 486.800 525.200 487.400 ;
        RECT 527.600 492.300 528.400 499.800 ;
        RECT 529.200 496.000 530.000 499.800 ;
        RECT 532.400 496.000 533.200 499.800 ;
        RECT 529.200 495.800 533.200 496.000 ;
        RECT 534.000 495.800 534.800 499.800 ;
        RECT 536.200 496.400 537.000 499.800 ;
        RECT 536.200 495.800 538.000 496.400 ;
        RECT 540.400 495.800 541.200 499.800 ;
        RECT 542.000 496.000 542.800 499.800 ;
        RECT 545.200 496.000 546.000 499.800 ;
        RECT 542.000 495.800 546.000 496.000 ;
        RECT 529.400 495.400 533.000 495.800 ;
        RECT 530.000 494.400 530.800 494.800 ;
        RECT 534.000 494.400 534.600 495.800 ;
        RECT 529.200 493.800 530.800 494.400 ;
        RECT 529.200 493.600 530.000 493.800 ;
        RECT 532.200 493.600 534.800 494.400 ;
        RECT 530.800 492.300 531.600 493.200 ;
        RECT 527.600 491.700 531.600 492.300 ;
        RECT 514.800 482.200 515.600 485.000 ;
        RECT 516.400 482.200 517.200 485.000 ;
        RECT 519.600 482.200 520.400 486.800 ;
        RECT 523.200 486.200 523.800 486.800 ;
        RECT 522.800 485.600 523.800 486.200 ;
        RECT 522.800 482.200 523.600 485.600 ;
        RECT 527.600 482.200 528.400 491.700 ;
        RECT 530.800 491.600 531.600 491.700 ;
        RECT 532.200 490.200 532.800 493.600 ;
        RECT 537.200 492.300 538.000 495.800 ;
        RECT 538.800 493.600 539.600 495.200 ;
        RECT 540.600 494.400 541.200 495.800 ;
        RECT 542.200 495.400 545.800 495.800 ;
        RECT 544.400 494.400 545.200 494.800 ;
        RECT 540.400 493.600 543.000 494.400 ;
        RECT 544.400 493.800 546.000 494.400 ;
        RECT 545.200 493.600 546.000 493.800 ;
        RECT 542.400 492.400 543.000 493.600 ;
        RECT 534.100 491.700 538.000 492.300 ;
        RECT 534.100 490.400 534.700 491.700 ;
        RECT 534.000 490.200 534.800 490.400 ;
        RECT 531.800 489.600 532.800 490.200 ;
        RECT 533.400 489.600 534.800 490.200 ;
        RECT 531.800 482.200 532.600 489.600 ;
        RECT 533.400 488.400 534.000 489.600 ;
        RECT 535.600 488.800 536.400 490.400 ;
        RECT 533.200 487.600 534.000 488.400 ;
        RECT 537.200 482.200 538.000 491.700 ;
        RECT 542.000 491.600 543.000 492.400 ;
        RECT 543.600 492.300 544.400 493.200 ;
        RECT 546.800 492.300 547.600 499.800 ;
        RECT 548.400 496.300 549.200 497.200 ;
        RECT 551.600 496.300 552.400 499.800 ;
        RECT 548.400 495.700 552.400 496.300 ;
        RECT 548.400 495.600 549.200 495.700 ;
        RECT 543.600 491.700 547.600 492.300 ;
        RECT 543.600 491.600 544.400 491.700 ;
        RECT 538.800 490.300 539.600 490.400 ;
        RECT 540.400 490.300 541.200 490.400 ;
        RECT 538.800 490.200 541.200 490.300 ;
        RECT 542.400 490.200 543.000 491.600 ;
        RECT 538.800 489.700 541.800 490.200 ;
        RECT 538.800 489.600 539.600 489.700 ;
        RECT 540.400 489.600 541.800 489.700 ;
        RECT 542.400 489.600 543.400 490.200 ;
        RECT 541.200 488.400 541.800 489.600 ;
        RECT 541.200 487.600 542.000 488.400 ;
        RECT 542.600 482.200 543.400 489.600 ;
        RECT 546.800 482.200 547.600 491.700 ;
        RECT 551.400 495.200 552.400 495.700 ;
        RECT 551.400 490.800 552.200 495.200 ;
        RECT 553.200 494.600 554.000 499.800 ;
        RECT 559.600 496.600 560.400 499.800 ;
        RECT 561.200 497.000 562.000 499.800 ;
        RECT 562.800 497.000 563.600 499.800 ;
        RECT 564.400 497.000 565.200 499.800 ;
        RECT 566.000 497.000 566.800 499.800 ;
        RECT 569.200 497.000 570.000 499.800 ;
        RECT 572.400 497.000 573.200 499.800 ;
        RECT 574.000 497.000 574.800 499.800 ;
        RECT 575.600 497.000 576.400 499.800 ;
        RECT 558.000 495.800 560.400 496.600 ;
        RECT 577.200 496.600 578.000 499.800 ;
        RECT 558.000 495.200 558.800 495.800 ;
        RECT 552.800 494.000 554.000 494.600 ;
        RECT 557.000 494.600 558.800 495.200 ;
        RECT 562.800 495.600 563.800 496.400 ;
        RECT 566.800 495.600 568.400 496.400 ;
        RECT 569.200 495.800 573.800 496.400 ;
        RECT 577.200 495.800 579.800 496.600 ;
        RECT 569.200 495.600 570.000 495.800 ;
        RECT 552.800 492.000 553.400 494.000 ;
        RECT 557.000 493.400 557.800 494.600 ;
        RECT 554.000 492.600 557.800 493.400 ;
        RECT 562.800 492.800 563.600 495.600 ;
        RECT 569.200 494.800 570.000 495.000 ;
        RECT 565.600 494.200 570.000 494.800 ;
        RECT 565.600 494.000 566.400 494.200 ;
        RECT 570.800 493.600 571.600 495.200 ;
        RECT 573.000 493.400 573.800 495.800 ;
        RECT 579.000 495.200 579.800 495.800 ;
        RECT 579.000 494.400 582.000 495.200 ;
        RECT 583.600 493.800 584.400 499.800 ;
        RECT 566.000 492.600 569.200 493.400 ;
        RECT 573.000 492.600 575.000 493.400 ;
        RECT 575.600 493.000 584.400 493.800 ;
        RECT 559.600 492.000 560.400 492.600 ;
        RECT 577.200 492.000 578.000 492.400 ;
        RECT 582.200 492.000 583.000 492.200 ;
        RECT 552.800 491.400 553.600 492.000 ;
        RECT 559.600 491.400 583.000 492.000 ;
        RECT 551.400 490.000 552.400 490.800 ;
        RECT 551.600 482.200 552.400 490.000 ;
        RECT 553.000 489.600 553.600 491.400 ;
        RECT 553.000 489.000 562.000 489.600 ;
        RECT 553.000 487.400 553.600 489.000 ;
        RECT 561.200 488.800 562.000 489.000 ;
        RECT 564.400 489.000 573.000 489.600 ;
        RECT 564.400 488.800 565.200 489.000 ;
        RECT 556.200 487.600 558.800 488.400 ;
        RECT 553.000 486.800 555.600 487.400 ;
        RECT 554.800 482.200 555.600 486.800 ;
        RECT 558.000 482.200 558.800 487.600 ;
        RECT 559.400 486.800 563.600 487.600 ;
        RECT 561.200 482.200 562.000 485.000 ;
        RECT 562.800 482.200 563.600 485.000 ;
        RECT 564.400 482.200 565.200 485.000 ;
        RECT 566.000 482.200 566.800 488.400 ;
        RECT 569.200 487.600 571.800 488.400 ;
        RECT 572.400 488.200 573.000 489.000 ;
        RECT 574.000 489.400 574.800 489.600 ;
        RECT 574.000 489.000 579.400 489.400 ;
        RECT 574.000 488.800 580.200 489.000 ;
        RECT 578.800 488.200 580.200 488.800 ;
        RECT 572.400 487.600 578.200 488.200 ;
        RECT 581.200 488.000 582.800 488.800 ;
        RECT 581.200 487.600 581.800 488.000 ;
        RECT 569.200 482.200 570.000 487.000 ;
        RECT 572.400 482.200 573.200 487.000 ;
        RECT 577.600 486.800 581.800 487.600 ;
        RECT 583.600 487.400 584.400 493.000 ;
        RECT 582.400 486.800 584.400 487.400 ;
        RECT 590.000 493.800 590.800 499.800 ;
        RECT 596.400 496.600 597.200 499.800 ;
        RECT 598.000 497.000 598.800 499.800 ;
        RECT 599.600 497.000 600.400 499.800 ;
        RECT 601.200 497.000 602.000 499.800 ;
        RECT 604.400 497.000 605.200 499.800 ;
        RECT 607.600 497.000 608.400 499.800 ;
        RECT 609.200 497.000 610.000 499.800 ;
        RECT 610.800 497.000 611.600 499.800 ;
        RECT 612.400 497.000 613.200 499.800 ;
        RECT 594.600 495.800 597.200 496.600 ;
        RECT 614.000 496.600 614.800 499.800 ;
        RECT 600.600 495.800 605.200 496.400 ;
        RECT 594.600 495.200 595.400 495.800 ;
        RECT 592.400 494.400 595.400 495.200 ;
        RECT 590.000 493.000 598.800 493.800 ;
        RECT 600.600 493.400 601.400 495.800 ;
        RECT 604.400 495.600 605.200 495.800 ;
        RECT 606.000 495.600 607.600 496.400 ;
        RECT 610.600 495.600 611.600 496.400 ;
        RECT 614.000 495.800 616.400 496.600 ;
        RECT 602.800 493.600 603.600 495.200 ;
        RECT 604.400 494.800 605.200 495.000 ;
        RECT 604.400 494.200 608.800 494.800 ;
        RECT 608.000 494.000 608.800 494.200 ;
        RECT 590.000 487.400 590.800 493.000 ;
        RECT 599.400 492.600 601.400 493.400 ;
        RECT 605.200 492.600 608.400 493.400 ;
        RECT 610.800 492.800 611.600 495.600 ;
        RECT 615.600 495.200 616.400 495.800 ;
        RECT 615.600 494.600 617.400 495.200 ;
        RECT 616.600 493.400 617.400 494.600 ;
        RECT 620.400 494.600 621.200 499.800 ;
        RECT 622.000 496.000 622.800 499.800 ;
        RECT 622.000 495.200 623.000 496.000 ;
        RECT 625.200 495.800 626.000 499.800 ;
        RECT 629.600 498.400 631.200 499.800 ;
        RECT 629.600 497.600 632.400 498.400 ;
        RECT 629.600 496.200 631.200 497.600 ;
        RECT 625.200 495.200 627.800 495.800 ;
        RECT 620.400 494.000 621.600 494.600 ;
        RECT 616.600 492.600 620.400 493.400 ;
        RECT 591.400 492.000 592.200 492.200 ;
        RECT 594.800 492.000 595.600 492.400 ;
        RECT 596.400 492.000 597.200 492.400 ;
        RECT 614.000 492.000 614.800 492.600 ;
        RECT 621.000 492.000 621.600 494.000 ;
        RECT 591.400 491.400 614.800 492.000 ;
        RECT 620.800 491.400 621.600 492.000 ;
        RECT 620.800 489.600 621.400 491.400 ;
        RECT 622.200 490.800 623.000 495.200 ;
        RECT 627.000 495.000 627.800 495.200 ;
        RECT 628.400 494.800 630.000 495.600 ;
        RECT 625.200 494.200 626.800 494.400 ;
        RECT 630.600 494.200 631.200 496.200 ;
        RECT 634.800 495.800 635.600 499.800 ;
        RECT 631.800 494.800 632.600 495.600 ;
        RECT 633.200 495.200 635.600 495.800 ;
        RECT 638.000 495.200 638.800 499.800 ;
        RECT 641.200 495.200 642.000 499.800 ;
        RECT 644.400 495.200 645.200 499.800 ;
        RECT 647.600 495.200 648.400 499.800 ;
        RECT 652.400 496.000 653.200 499.800 ;
        RECT 652.200 495.200 653.200 496.000 ;
        RECT 633.200 495.000 634.000 495.200 ;
        RECT 625.200 494.000 627.400 494.200 ;
        RECT 625.200 493.600 629.600 494.000 ;
        RECT 626.800 493.400 629.600 493.600 ;
        RECT 628.800 493.200 629.600 493.400 ;
        RECT 630.200 493.600 631.200 494.200 ;
        RECT 632.000 494.400 632.600 494.800 ;
        RECT 638.000 494.400 639.800 495.200 ;
        RECT 641.200 494.400 643.400 495.200 ;
        RECT 644.400 494.400 646.600 495.200 ;
        RECT 647.600 494.400 650.000 495.200 ;
        RECT 632.000 493.600 632.800 494.400 ;
        RECT 634.000 493.600 635.600 494.400 ;
        RECT 636.400 493.800 637.200 494.400 ;
        RECT 639.000 493.800 639.800 494.400 ;
        RECT 642.600 493.800 643.400 494.400 ;
        RECT 645.800 493.800 646.600 494.400 ;
        RECT 630.200 492.400 630.800 493.600 ;
        RECT 636.400 493.000 638.200 493.800 ;
        RECT 639.000 493.000 641.600 493.800 ;
        RECT 642.600 493.000 645.000 493.800 ;
        RECT 645.800 493.000 648.400 493.800 ;
        RECT 627.400 492.200 628.200 492.400 ;
        RECT 627.400 491.600 629.000 492.200 ;
        RECT 630.000 491.600 630.800 492.400 ;
        RECT 639.000 491.600 639.800 493.000 ;
        RECT 642.600 491.600 643.400 493.000 ;
        RECT 645.800 491.600 646.600 493.000 ;
        RECT 649.200 491.600 650.000 494.400 ;
        RECT 628.200 491.400 629.000 491.600 ;
        RECT 599.600 489.400 600.400 489.600 ;
        RECT 595.000 489.000 600.400 489.400 ;
        RECT 594.200 488.800 600.400 489.000 ;
        RECT 601.400 489.000 610.000 489.600 ;
        RECT 591.600 488.000 593.200 488.800 ;
        RECT 594.200 488.200 595.600 488.800 ;
        RECT 601.400 488.200 602.000 489.000 ;
        RECT 609.200 488.800 610.000 489.000 ;
        RECT 612.400 489.000 621.400 489.600 ;
        RECT 612.400 488.800 613.200 489.000 ;
        RECT 592.600 487.600 593.200 488.000 ;
        RECT 596.200 487.600 602.000 488.200 ;
        RECT 602.600 487.600 605.200 488.400 ;
        RECT 590.000 486.800 592.000 487.400 ;
        RECT 592.600 486.800 596.800 487.600 ;
        RECT 574.000 482.200 574.800 485.000 ;
        RECT 575.600 482.200 576.400 485.000 ;
        RECT 578.800 482.200 579.600 486.800 ;
        RECT 582.400 486.200 583.000 486.800 ;
        RECT 582.000 485.600 583.000 486.200 ;
        RECT 591.400 486.200 592.000 486.800 ;
        RECT 591.400 485.600 592.400 486.200 ;
        RECT 582.000 482.200 582.800 485.600 ;
        RECT 591.600 482.200 592.400 485.600 ;
        RECT 594.800 482.200 595.600 486.800 ;
        RECT 598.000 482.200 598.800 485.000 ;
        RECT 599.600 482.200 600.400 485.000 ;
        RECT 601.200 482.200 602.000 487.000 ;
        RECT 604.400 482.200 605.200 487.000 ;
        RECT 607.600 482.200 608.400 488.400 ;
        RECT 615.600 487.600 618.200 488.400 ;
        RECT 610.800 486.800 615.000 487.600 ;
        RECT 609.200 482.200 610.000 485.000 ;
        RECT 610.800 482.200 611.600 485.000 ;
        RECT 612.400 482.200 613.200 485.000 ;
        RECT 615.600 482.200 616.400 487.600 ;
        RECT 620.800 487.400 621.400 489.000 ;
        RECT 618.800 486.800 621.400 487.400 ;
        RECT 622.000 490.000 623.000 490.800 ;
        RECT 630.200 490.200 630.800 491.600 ;
        RECT 638.000 490.800 639.800 491.600 ;
        RECT 641.200 490.800 643.400 491.600 ;
        RECT 644.400 490.800 646.600 491.600 ;
        RECT 647.600 490.800 650.000 491.600 ;
        RECT 652.200 490.800 653.000 495.200 ;
        RECT 654.000 494.600 654.800 499.800 ;
        RECT 660.400 496.600 661.200 499.800 ;
        RECT 662.000 497.000 662.800 499.800 ;
        RECT 663.600 497.000 664.400 499.800 ;
        RECT 665.200 497.000 666.000 499.800 ;
        RECT 666.800 497.000 667.600 499.800 ;
        RECT 670.000 497.000 670.800 499.800 ;
        RECT 673.200 497.000 674.000 499.800 ;
        RECT 674.800 497.000 675.600 499.800 ;
        RECT 676.400 497.000 677.200 499.800 ;
        RECT 658.800 495.800 661.200 496.600 ;
        RECT 678.000 496.600 678.800 499.800 ;
        RECT 658.800 495.200 659.600 495.800 ;
        RECT 653.600 494.000 654.800 494.600 ;
        RECT 657.800 494.600 659.600 495.200 ;
        RECT 663.600 495.600 664.600 496.400 ;
        RECT 667.600 495.600 669.200 496.400 ;
        RECT 670.000 495.800 674.600 496.400 ;
        RECT 678.000 495.800 680.600 496.600 ;
        RECT 670.000 495.600 670.800 495.800 ;
        RECT 653.600 492.000 654.200 494.000 ;
        RECT 657.800 493.400 658.600 494.600 ;
        RECT 654.800 492.600 658.600 493.400 ;
        RECT 663.600 492.800 664.400 495.600 ;
        RECT 670.000 494.800 670.800 495.000 ;
        RECT 666.400 494.200 670.800 494.800 ;
        RECT 666.400 494.000 667.200 494.200 ;
        RECT 671.600 493.600 672.400 495.200 ;
        RECT 673.800 493.400 674.600 495.800 ;
        RECT 679.800 495.200 680.600 495.800 ;
        RECT 679.800 494.400 682.800 495.200 ;
        RECT 684.400 493.800 685.200 499.800 ;
        RECT 666.800 492.600 670.000 493.400 ;
        RECT 673.800 492.600 675.800 493.400 ;
        RECT 676.400 493.000 685.200 493.800 ;
        RECT 660.400 492.000 661.200 492.600 ;
        RECT 678.000 492.000 678.800 492.400 ;
        RECT 683.000 492.000 683.800 492.200 ;
        RECT 653.600 491.400 654.400 492.000 ;
        RECT 660.400 491.400 683.800 492.000 ;
        RECT 618.800 482.200 619.600 486.800 ;
        RECT 622.000 482.200 622.800 490.000 ;
        RECT 625.200 489.600 627.800 490.200 ;
        RECT 625.200 482.200 626.000 489.600 ;
        RECT 627.000 489.400 627.800 489.600 ;
        RECT 629.600 482.200 631.200 490.200 ;
        RECT 633.200 489.600 635.600 490.200 ;
        RECT 633.200 489.400 634.000 489.600 ;
        RECT 634.800 482.200 635.600 489.600 ;
        RECT 638.000 482.200 638.800 490.800 ;
        RECT 641.200 482.200 642.000 490.800 ;
        RECT 644.400 482.200 645.200 490.800 ;
        RECT 647.600 482.200 648.400 490.800 ;
        RECT 652.200 490.000 653.200 490.800 ;
        RECT 652.400 482.200 653.200 490.000 ;
        RECT 653.800 489.600 654.400 491.400 ;
        RECT 653.800 489.000 662.800 489.600 ;
        RECT 653.800 487.400 654.400 489.000 ;
        RECT 662.000 488.800 662.800 489.000 ;
        RECT 665.200 489.000 673.800 489.600 ;
        RECT 665.200 488.800 666.000 489.000 ;
        RECT 657.000 487.600 659.600 488.400 ;
        RECT 653.800 486.800 656.400 487.400 ;
        RECT 655.600 482.200 656.400 486.800 ;
        RECT 658.800 482.200 659.600 487.600 ;
        RECT 660.200 486.800 664.400 487.600 ;
        RECT 662.000 482.200 662.800 485.000 ;
        RECT 663.600 482.200 664.400 485.000 ;
        RECT 665.200 482.200 666.000 485.000 ;
        RECT 666.800 482.200 667.600 488.400 ;
        RECT 670.000 487.600 672.600 488.400 ;
        RECT 673.200 488.200 673.800 489.000 ;
        RECT 674.800 489.400 675.600 489.600 ;
        RECT 674.800 489.000 680.200 489.400 ;
        RECT 674.800 488.800 681.000 489.000 ;
        RECT 679.600 488.200 681.000 488.800 ;
        RECT 673.200 487.600 679.000 488.200 ;
        RECT 682.000 488.000 683.600 488.800 ;
        RECT 682.000 487.600 682.600 488.000 ;
        RECT 670.000 482.200 670.800 487.000 ;
        RECT 673.200 482.200 674.000 487.000 ;
        RECT 678.400 486.800 682.600 487.600 ;
        RECT 684.400 487.400 685.200 493.000 ;
        RECT 683.200 486.800 685.200 487.400 ;
        RECT 674.800 482.200 675.600 485.000 ;
        RECT 676.400 482.200 677.200 485.000 ;
        RECT 679.600 482.200 680.400 486.800 ;
        RECT 683.200 486.200 683.800 486.800 ;
        RECT 682.800 485.600 683.800 486.200 ;
        RECT 682.800 482.200 683.600 485.600 ;
        RECT 2.800 472.000 3.600 479.800 ;
        RECT 6.000 475.200 6.800 479.800 ;
        RECT 2.600 471.200 3.600 472.000 ;
        RECT 4.200 474.600 6.800 475.200 ;
        RECT 4.200 473.000 4.800 474.600 ;
        RECT 9.200 474.400 10.000 479.800 ;
        RECT 12.400 477.000 13.200 479.800 ;
        RECT 14.000 477.000 14.800 479.800 ;
        RECT 15.600 477.000 16.400 479.800 ;
        RECT 10.600 474.400 14.800 475.200 ;
        RECT 7.400 473.600 10.000 474.400 ;
        RECT 17.200 473.600 18.000 479.800 ;
        RECT 20.400 475.000 21.200 479.800 ;
        RECT 23.600 475.000 24.400 479.800 ;
        RECT 25.200 477.000 26.000 479.800 ;
        RECT 26.800 477.000 27.600 479.800 ;
        RECT 30.000 475.200 30.800 479.800 ;
        RECT 33.200 476.400 34.000 479.800 ;
        RECT 38.600 478.400 39.400 479.800 ;
        RECT 38.600 477.600 40.400 478.400 ;
        RECT 33.200 475.800 34.200 476.400 ;
        RECT 33.600 475.200 34.200 475.800 ;
        RECT 28.800 474.400 33.000 475.200 ;
        RECT 33.600 474.600 35.600 475.200 ;
        RECT 20.400 473.600 23.000 474.400 ;
        RECT 23.600 473.800 29.400 474.400 ;
        RECT 32.400 474.000 33.000 474.400 ;
        RECT 12.400 473.000 13.200 473.200 ;
        RECT 4.200 472.400 13.200 473.000 ;
        RECT 15.600 473.000 16.400 473.200 ;
        RECT 23.600 473.000 24.200 473.800 ;
        RECT 30.000 473.200 31.400 473.800 ;
        RECT 32.400 473.200 34.000 474.000 ;
        RECT 15.600 472.400 24.200 473.000 ;
        RECT 25.200 473.000 31.400 473.200 ;
        RECT 25.200 472.600 30.600 473.000 ;
        RECT 25.200 472.400 26.000 472.600 ;
        RECT 2.600 466.800 3.400 471.200 ;
        RECT 4.200 470.600 4.800 472.400 ;
        RECT 4.000 470.000 4.800 470.600 ;
        RECT 10.800 470.000 34.200 470.600 ;
        RECT 4.000 468.000 4.600 470.000 ;
        RECT 10.800 469.400 11.600 470.000 ;
        RECT 28.400 469.600 29.200 470.000 ;
        RECT 33.400 469.800 34.200 470.000 ;
        RECT 5.200 468.600 9.000 469.400 ;
        RECT 4.000 467.400 5.200 468.000 ;
        RECT 2.600 466.000 3.600 466.800 ;
        RECT 2.800 462.200 3.600 466.000 ;
        RECT 4.400 462.200 5.200 467.400 ;
        RECT 8.200 467.400 9.000 468.600 ;
        RECT 8.200 466.800 10.000 467.400 ;
        RECT 9.200 466.200 10.000 466.800 ;
        RECT 14.000 466.400 14.800 469.200 ;
        RECT 17.200 468.600 20.400 469.400 ;
        RECT 24.200 468.600 26.200 469.400 ;
        RECT 34.800 469.000 35.600 474.600 ;
        RECT 37.200 473.600 38.000 474.400 ;
        RECT 37.200 472.400 37.800 473.600 ;
        RECT 38.600 472.400 39.400 477.600 ;
        RECT 36.400 471.800 37.800 472.400 ;
        RECT 38.400 471.800 39.400 472.400 ;
        RECT 36.400 471.600 37.200 471.800 ;
        RECT 16.800 467.800 17.600 468.000 ;
        RECT 16.800 467.200 21.200 467.800 ;
        RECT 20.400 467.000 21.200 467.200 ;
        RECT 22.000 466.800 22.800 468.400 ;
        RECT 9.200 465.400 11.600 466.200 ;
        RECT 14.000 465.600 15.000 466.400 ;
        RECT 18.000 465.600 19.600 466.400 ;
        RECT 20.400 466.200 21.200 466.400 ;
        RECT 24.200 466.200 25.000 468.600 ;
        RECT 26.800 468.200 35.600 469.000 ;
        RECT 38.400 468.400 39.000 471.800 ;
        RECT 42.800 471.600 43.600 473.200 ;
        RECT 39.600 468.800 40.400 470.400 ;
        RECT 30.200 466.800 33.200 467.600 ;
        RECT 30.200 466.200 31.000 466.800 ;
        RECT 20.400 465.600 25.000 466.200 ;
        RECT 10.800 462.200 11.600 465.400 ;
        RECT 28.400 465.400 31.000 466.200 ;
        RECT 12.400 462.200 13.200 465.000 ;
        RECT 14.000 462.200 14.800 465.000 ;
        RECT 15.600 462.200 16.400 465.000 ;
        RECT 17.200 462.200 18.000 465.000 ;
        RECT 20.400 462.200 21.200 465.000 ;
        RECT 23.600 462.200 24.400 465.000 ;
        RECT 25.200 462.200 26.000 465.000 ;
        RECT 26.800 462.200 27.600 465.000 ;
        RECT 28.400 462.200 29.200 465.400 ;
        RECT 34.800 462.200 35.600 468.200 ;
        RECT 36.400 467.600 39.000 468.400 ;
        RECT 41.200 468.200 42.000 468.400 ;
        RECT 40.400 467.600 42.000 468.200 ;
        RECT 36.600 466.200 37.200 467.600 ;
        RECT 40.400 467.200 41.200 467.600 ;
        RECT 38.200 466.200 41.800 466.600 ;
        RECT 44.400 466.200 45.200 479.800 ;
        RECT 47.600 471.400 48.400 479.800 ;
        RECT 52.000 476.400 52.800 479.800 ;
        RECT 50.800 475.800 52.800 476.400 ;
        RECT 56.400 475.800 57.200 479.800 ;
        RECT 60.600 475.800 61.800 479.800 ;
        RECT 50.800 475.000 51.600 475.800 ;
        RECT 56.400 475.200 57.000 475.800 ;
        RECT 54.200 474.600 57.800 475.200 ;
        RECT 60.400 475.000 61.200 475.800 ;
        RECT 54.200 474.400 55.000 474.600 ;
        RECT 57.000 474.400 57.800 474.600 ;
        RECT 61.400 474.000 62.800 474.400 ;
        RECT 60.600 473.600 62.800 474.000 ;
        RECT 50.800 473.000 51.600 473.200 ;
        RECT 55.400 473.000 56.200 473.200 ;
        RECT 50.800 472.400 56.200 473.000 ;
        RECT 56.800 473.000 59.000 473.600 ;
        RECT 56.800 471.800 57.400 473.000 ;
        RECT 58.200 472.800 59.000 473.000 ;
        RECT 60.600 473.200 62.000 473.600 ;
        RECT 60.600 472.200 61.200 473.200 ;
        RECT 52.600 471.400 57.400 471.800 ;
        RECT 47.600 471.200 57.400 471.400 ;
        RECT 58.800 471.600 61.200 472.200 ;
        RECT 47.600 471.000 53.400 471.200 ;
        RECT 47.600 470.800 53.200 471.000 ;
        RECT 54.000 470.200 54.800 470.400 ;
        RECT 49.800 469.600 54.800 470.200 ;
        RECT 49.800 469.400 50.600 469.600 ;
        RECT 52.400 469.400 53.200 469.600 ;
        RECT 51.400 468.400 52.200 468.600 ;
        RECT 58.800 468.400 59.400 471.600 ;
        RECT 65.200 471.200 66.000 479.800 ;
        RECT 70.600 474.400 71.400 479.800 ;
        RECT 74.800 475.000 75.600 479.000 ;
        RECT 70.600 473.600 72.400 474.400 ;
        RECT 70.600 472.800 71.400 473.600 ;
        RECT 69.800 472.200 71.400 472.800 ;
        RECT 61.800 470.600 66.000 471.200 ;
        RECT 61.800 470.400 62.600 470.600 ;
        RECT 63.400 469.800 64.200 470.000 ;
        RECT 60.400 469.200 64.200 469.800 ;
        RECT 60.400 469.000 61.200 469.200 ;
        RECT 46.000 466.800 46.800 468.400 ;
        RECT 48.400 467.800 59.400 468.400 ;
        RECT 48.400 467.600 50.000 467.800 ;
        RECT 36.400 462.200 37.200 466.200 ;
        RECT 38.000 466.000 42.000 466.200 ;
        RECT 38.000 462.200 38.800 466.000 ;
        RECT 41.200 462.200 42.000 466.000 ;
        RECT 43.400 465.600 45.200 466.200 ;
        RECT 43.400 464.400 44.200 465.600 ;
        RECT 42.800 463.600 44.200 464.400 ;
        RECT 43.400 462.200 44.200 463.600 ;
        RECT 47.600 462.200 48.400 467.000 ;
        RECT 52.600 465.600 53.200 467.800 ;
        RECT 55.600 467.600 56.400 467.800 ;
        RECT 58.200 467.600 59.000 467.800 ;
        RECT 65.200 467.200 66.000 470.600 ;
        RECT 68.400 469.600 69.200 471.200 ;
        RECT 69.800 468.400 70.400 472.200 ;
        RECT 75.000 471.600 75.600 475.000 ;
        RECT 79.000 472.400 79.800 479.800 ;
        RECT 80.400 473.600 81.200 474.400 ;
        RECT 80.600 472.400 81.200 473.600 ;
        RECT 83.600 473.600 84.400 474.400 ;
        RECT 83.600 472.400 84.200 473.600 ;
        RECT 85.000 472.400 85.800 479.800 ;
        RECT 79.000 471.800 80.000 472.400 ;
        RECT 80.600 471.800 82.000 472.400 ;
        RECT 71.800 471.000 75.600 471.600 ;
        RECT 71.800 469.000 72.400 471.000 ;
        RECT 68.400 467.600 70.400 468.400 ;
        RECT 71.000 468.200 72.400 469.000 ;
        RECT 73.200 468.800 74.000 470.400 ;
        RECT 74.800 468.800 75.600 470.400 ;
        RECT 78.000 468.800 78.800 470.400 ;
        RECT 79.400 468.400 80.000 471.800 ;
        RECT 81.200 471.600 82.000 471.800 ;
        RECT 82.800 471.800 84.200 472.400 ;
        RECT 84.800 471.800 85.800 472.400 ;
        RECT 82.800 471.600 83.600 471.800 ;
        RECT 81.300 470.300 81.900 471.600 ;
        RECT 84.800 470.300 85.400 471.800 ;
        RECT 89.200 471.600 90.000 474.400 ;
        RECT 81.300 469.700 85.400 470.300 ;
        RECT 84.800 468.400 85.400 469.700 ;
        RECT 86.000 468.800 86.800 470.400 ;
        RECT 62.200 466.600 66.000 467.200 ;
        RECT 62.200 466.400 63.000 466.600 ;
        RECT 50.800 464.200 51.600 465.000 ;
        RECT 52.400 464.800 53.200 465.600 ;
        RECT 54.200 465.400 55.000 465.600 ;
        RECT 54.200 464.800 57.000 465.400 ;
        RECT 56.400 464.200 57.000 464.800 ;
        RECT 60.400 464.200 61.200 465.000 ;
        RECT 50.800 463.600 52.800 464.200 ;
        RECT 52.000 462.200 52.800 463.600 ;
        RECT 56.400 462.200 57.200 464.200 ;
        RECT 60.400 463.600 61.800 464.200 ;
        RECT 60.600 462.200 61.800 463.600 ;
        RECT 65.200 462.200 66.000 466.600 ;
        RECT 69.800 467.000 70.400 467.600 ;
        RECT 71.400 467.800 72.400 468.200 ;
        RECT 76.400 468.200 77.200 468.400 ;
        RECT 71.400 467.200 75.600 467.800 ;
        RECT 76.400 467.600 78.000 468.200 ;
        RECT 79.400 467.600 82.000 468.400 ;
        RECT 82.800 467.600 85.400 468.400 ;
        RECT 87.600 468.200 88.400 468.400 ;
        RECT 86.800 467.600 88.400 468.200 ;
        RECT 77.200 467.200 78.000 467.600 ;
        RECT 69.800 466.600 70.600 467.000 ;
        RECT 69.800 466.000 71.400 466.600 ;
        RECT 70.600 463.000 71.400 466.000 ;
        RECT 75.000 465.000 75.600 467.200 ;
        RECT 76.600 466.200 80.200 466.600 ;
        RECT 81.200 466.200 81.800 467.600 ;
        RECT 83.000 466.200 83.600 467.600 ;
        RECT 86.800 467.200 87.600 467.600 ;
        RECT 84.600 466.200 88.200 466.600 ;
        RECT 90.800 466.200 91.600 479.800 ;
        RECT 94.000 471.400 94.800 479.800 ;
        RECT 98.400 476.400 99.200 479.800 ;
        RECT 97.200 475.800 99.200 476.400 ;
        RECT 102.800 475.800 103.600 479.800 ;
        RECT 107.000 475.800 108.200 479.800 ;
        RECT 97.200 475.000 98.000 475.800 ;
        RECT 102.800 475.200 103.400 475.800 ;
        RECT 100.600 474.600 104.200 475.200 ;
        RECT 106.800 475.000 107.600 475.800 ;
        RECT 100.600 474.400 101.400 474.600 ;
        RECT 103.400 474.400 104.200 474.600 ;
        RECT 97.200 473.000 98.000 473.200 ;
        RECT 101.800 473.000 102.600 473.200 ;
        RECT 97.200 472.400 102.600 473.000 ;
        RECT 103.200 473.000 105.400 473.600 ;
        RECT 103.200 471.800 103.800 473.000 ;
        RECT 104.600 472.800 105.400 473.000 ;
        RECT 107.000 473.200 108.400 474.000 ;
        RECT 107.000 472.200 107.600 473.200 ;
        RECT 99.000 471.400 103.800 471.800 ;
        RECT 94.000 471.200 103.800 471.400 ;
        RECT 105.200 471.600 107.600 472.200 ;
        RECT 94.000 471.000 99.800 471.200 ;
        RECT 94.000 470.800 99.600 471.000 ;
        RECT 105.200 470.400 105.800 471.600 ;
        RECT 111.600 471.200 112.400 479.800 ;
        RECT 120.600 472.400 121.400 479.800 ;
        RECT 122.000 473.600 122.800 474.400 ;
        RECT 122.200 472.400 122.800 473.600 ;
        RECT 125.200 473.600 126.000 474.400 ;
        RECT 125.200 472.400 125.800 473.600 ;
        RECT 126.600 472.400 127.400 479.800 ;
        RECT 120.600 471.800 121.600 472.400 ;
        RECT 122.200 471.800 123.600 472.400 ;
        RECT 108.200 470.600 112.400 471.200 ;
        RECT 108.200 470.400 109.000 470.600 ;
        RECT 100.400 470.200 101.200 470.400 ;
        RECT 96.200 469.600 101.200 470.200 ;
        RECT 105.200 469.600 106.000 470.400 ;
        RECT 109.800 469.800 110.600 470.000 ;
        RECT 96.200 469.400 97.000 469.600 ;
        RECT 98.800 469.400 99.600 469.600 ;
        RECT 97.800 468.400 98.600 468.600 ;
        RECT 105.200 468.400 105.800 469.600 ;
        RECT 106.800 469.200 110.600 469.800 ;
        RECT 106.800 469.000 107.600 469.200 ;
        RECT 92.400 466.800 93.200 468.400 ;
        RECT 94.800 467.800 105.800 468.400 ;
        RECT 94.800 467.600 96.400 467.800 ;
        RECT 74.800 463.000 75.600 465.000 ;
        RECT 76.400 466.000 80.400 466.200 ;
        RECT 76.400 462.200 77.200 466.000 ;
        RECT 79.600 462.200 80.400 466.000 ;
        RECT 81.200 462.200 82.000 466.200 ;
        RECT 82.800 462.200 83.600 466.200 ;
        RECT 84.400 466.000 88.400 466.200 ;
        RECT 84.400 462.200 85.200 466.000 ;
        RECT 87.600 462.200 88.400 466.000 ;
        RECT 89.800 465.600 91.600 466.200 ;
        RECT 89.800 464.400 90.600 465.600 ;
        RECT 89.800 463.600 91.600 464.400 ;
        RECT 89.800 462.200 90.600 463.600 ;
        RECT 94.000 462.200 94.800 467.000 ;
        RECT 99.000 465.600 99.600 467.800 ;
        RECT 104.600 467.600 105.400 467.800 ;
        RECT 111.600 467.200 112.400 470.600 ;
        RECT 119.600 468.800 120.400 470.400 ;
        RECT 121.000 470.300 121.600 471.800 ;
        RECT 122.800 471.600 123.600 471.800 ;
        RECT 124.400 471.800 125.800 472.400 ;
        RECT 126.400 471.800 127.400 472.400 ;
        RECT 130.800 475.000 131.600 479.000 ;
        RECT 124.400 471.600 125.200 471.800 ;
        RECT 124.500 470.300 125.100 471.600 ;
        RECT 121.000 469.700 125.100 470.300 ;
        RECT 121.000 468.400 121.600 469.700 ;
        RECT 126.400 468.400 127.000 471.800 ;
        RECT 130.800 471.600 131.400 475.000 ;
        RECT 135.000 472.800 135.800 479.800 ;
        RECT 135.000 472.200 136.600 472.800 ;
        RECT 130.800 471.000 134.600 471.600 ;
        RECT 127.600 468.800 128.400 470.400 ;
        RECT 130.800 468.800 131.600 470.400 ;
        RECT 132.400 468.800 133.200 470.400 ;
        RECT 134.000 469.000 134.600 471.000 ;
        RECT 118.000 468.200 118.800 468.400 ;
        RECT 118.000 467.600 119.600 468.200 ;
        RECT 121.000 467.600 123.600 468.400 ;
        RECT 124.400 467.600 127.000 468.400 ;
        RECT 129.200 468.200 130.000 468.400 ;
        RECT 128.400 467.600 130.000 468.200 ;
        RECT 134.000 468.200 135.400 469.000 ;
        RECT 136.000 468.400 136.600 472.200 ;
        RECT 140.400 471.200 141.200 479.800 ;
        RECT 144.600 475.800 145.800 479.800 ;
        RECT 149.200 475.800 150.000 479.800 ;
        RECT 153.600 476.400 154.400 479.800 ;
        RECT 153.600 475.800 155.600 476.400 ;
        RECT 145.200 475.000 146.000 475.800 ;
        RECT 149.400 475.200 150.000 475.800 ;
        RECT 148.600 474.600 152.200 475.200 ;
        RECT 154.800 475.000 155.600 475.800 ;
        RECT 148.600 474.400 149.400 474.600 ;
        RECT 151.400 474.400 152.200 474.600 ;
        RECT 144.400 473.200 145.800 474.000 ;
        RECT 145.200 472.200 145.800 473.200 ;
        RECT 147.400 473.000 149.600 473.600 ;
        RECT 147.400 472.800 148.200 473.000 ;
        RECT 145.200 471.600 147.600 472.200 ;
        RECT 137.200 469.600 138.000 471.200 ;
        RECT 140.400 470.600 144.600 471.200 ;
        RECT 134.000 467.800 135.000 468.200 ;
        RECT 118.800 467.200 119.600 467.600 ;
        RECT 108.600 466.600 112.400 467.200 ;
        RECT 108.600 466.400 109.400 466.600 ;
        RECT 97.200 464.200 98.000 465.000 ;
        RECT 98.800 464.800 99.600 465.600 ;
        RECT 100.600 465.400 101.400 465.600 ;
        RECT 100.600 464.800 103.400 465.400 ;
        RECT 102.800 464.200 103.400 464.800 ;
        RECT 106.800 464.200 107.600 465.000 ;
        RECT 97.200 463.600 99.200 464.200 ;
        RECT 98.400 462.200 99.200 463.600 ;
        RECT 102.800 462.200 103.600 464.200 ;
        RECT 106.800 463.600 108.200 464.200 ;
        RECT 107.000 462.200 108.200 463.600 ;
        RECT 111.600 462.200 112.400 466.600 ;
        RECT 118.200 466.200 121.800 466.600 ;
        RECT 122.800 466.200 123.400 467.600 ;
        RECT 124.600 466.200 125.200 467.600 ;
        RECT 128.400 467.200 129.200 467.600 ;
        RECT 130.800 467.200 135.000 467.800 ;
        RECT 136.000 467.600 138.000 468.400 ;
        RECT 126.200 466.200 129.800 466.600 ;
        RECT 118.000 466.000 122.000 466.200 ;
        RECT 118.000 462.200 118.800 466.000 ;
        RECT 121.200 462.200 122.000 466.000 ;
        RECT 122.800 462.200 123.600 466.200 ;
        RECT 124.400 462.200 125.200 466.200 ;
        RECT 126.000 466.000 130.000 466.200 ;
        RECT 126.000 462.200 126.800 466.000 ;
        RECT 129.200 462.200 130.000 466.000 ;
        RECT 130.800 465.000 131.400 467.200 ;
        RECT 136.000 467.000 136.600 467.600 ;
        RECT 135.800 466.600 136.600 467.000 ;
        RECT 135.000 466.000 136.600 466.600 ;
        RECT 140.400 467.200 141.200 470.600 ;
        RECT 143.800 470.400 144.600 470.600 ;
        RECT 142.200 469.800 143.000 470.000 ;
        RECT 142.200 469.200 146.000 469.800 ;
        RECT 145.200 469.000 146.000 469.200 ;
        RECT 147.000 468.400 147.600 471.600 ;
        RECT 149.000 471.800 149.600 473.000 ;
        RECT 150.200 473.000 151.000 473.200 ;
        RECT 154.800 473.000 155.600 473.200 ;
        RECT 150.200 472.400 155.600 473.000 ;
        RECT 149.000 471.400 153.800 471.800 ;
        RECT 158.000 471.400 158.800 479.800 ;
        RECT 149.000 471.200 158.800 471.400 ;
        RECT 153.000 471.000 158.800 471.200 ;
        RECT 153.200 470.800 158.800 471.000 ;
        RECT 151.600 470.200 152.400 470.400 ;
        RECT 151.600 469.600 156.600 470.200 ;
        RECT 153.200 469.400 154.000 469.600 ;
        RECT 155.800 469.400 156.600 469.600 ;
        RECT 154.200 468.400 155.000 468.600 ;
        RECT 147.000 467.800 158.000 468.400 ;
        RECT 147.400 467.600 148.200 467.800 ;
        RECT 140.400 466.600 144.200 467.200 ;
        RECT 130.800 463.000 131.600 465.000 ;
        RECT 135.000 464.400 135.800 466.000 ;
        RECT 134.000 463.600 135.800 464.400 ;
        RECT 135.000 463.000 135.800 463.600 ;
        RECT 140.400 462.200 141.200 466.600 ;
        RECT 143.400 466.400 144.200 466.600 ;
        RECT 153.200 465.600 153.800 467.800 ;
        RECT 156.400 467.600 158.000 467.800 ;
        RECT 151.400 465.400 152.200 465.600 ;
        RECT 145.200 464.200 146.000 465.000 ;
        RECT 149.400 464.800 152.200 465.400 ;
        RECT 153.200 464.800 154.000 465.600 ;
        RECT 149.400 464.200 150.000 464.800 ;
        RECT 154.800 464.200 155.600 465.000 ;
        RECT 144.600 463.600 146.000 464.200 ;
        RECT 144.600 462.200 145.800 463.600 ;
        RECT 149.200 462.200 150.000 464.200 ;
        RECT 153.600 463.600 155.600 464.200 ;
        RECT 153.600 462.200 154.400 463.600 ;
        RECT 158.000 462.200 158.800 467.000 ;
        RECT 159.600 466.800 160.400 468.400 ;
        RECT 161.200 466.200 162.000 479.800 ;
        RECT 164.400 474.300 165.200 474.400 ;
        RECT 162.800 473.700 165.200 474.300 ;
        RECT 162.800 471.600 163.600 473.700 ;
        RECT 164.400 473.600 165.200 473.700 ;
        RECT 162.800 470.300 163.600 470.400 ;
        RECT 166.000 470.300 166.800 479.800 ;
        RECT 167.600 471.600 168.400 473.200 ;
        RECT 169.800 472.600 170.600 479.800 ;
        RECT 176.600 472.600 177.400 479.800 ;
        RECT 169.800 471.800 171.600 472.600 ;
        RECT 175.600 471.800 177.400 472.600 ;
        RECT 167.700 470.400 168.300 471.600 ;
        RECT 162.800 469.700 166.800 470.300 ;
        RECT 162.800 469.600 163.600 469.700 ;
        RECT 164.400 466.800 165.200 468.400 ;
        RECT 166.000 466.200 166.800 469.700 ;
        RECT 167.600 470.300 168.400 470.400 ;
        RECT 169.200 470.300 170.000 471.200 ;
        RECT 167.600 469.700 170.000 470.300 ;
        RECT 167.600 469.600 168.400 469.700 ;
        RECT 169.200 469.600 170.000 469.700 ;
        RECT 170.800 468.400 171.400 471.800 ;
        RECT 175.800 468.400 176.400 471.800 ;
        RECT 177.200 469.600 178.000 471.200 ;
        RECT 170.800 467.600 171.600 468.400 ;
        RECT 175.600 467.600 176.400 468.400 ;
        RECT 161.200 465.600 163.000 466.200 ;
        RECT 166.000 465.600 167.800 466.200 ;
        RECT 162.200 464.400 163.000 465.600 ;
        RECT 162.200 463.600 163.600 464.400 ;
        RECT 162.200 462.200 163.000 463.600 ;
        RECT 167.000 462.200 167.800 465.600 ;
        RECT 170.800 464.400 171.400 467.600 ;
        RECT 172.400 464.800 173.200 466.400 ;
        RECT 174.000 464.800 174.800 466.400 ;
        RECT 175.800 464.400 176.400 467.600 ;
        RECT 170.800 462.200 171.600 464.400 ;
        RECT 175.600 462.200 176.400 464.400 ;
        RECT 178.800 462.200 179.600 479.800 ;
        RECT 180.400 472.300 181.200 472.400 ;
        RECT 182.000 472.300 182.800 479.800 ;
        RECT 180.400 471.700 182.800 472.300 ;
        RECT 186.800 472.000 187.600 479.800 ;
        RECT 190.000 475.200 190.800 479.800 ;
        RECT 180.400 471.600 181.200 471.700 ;
        RECT 182.000 468.300 182.800 471.700 ;
        RECT 186.600 471.200 187.600 472.000 ;
        RECT 188.200 474.600 190.800 475.200 ;
        RECT 188.200 473.000 188.800 474.600 ;
        RECT 193.200 474.400 194.000 479.800 ;
        RECT 196.400 477.000 197.200 479.800 ;
        RECT 198.000 477.000 198.800 479.800 ;
        RECT 199.600 477.000 200.400 479.800 ;
        RECT 194.600 474.400 198.800 475.200 ;
        RECT 191.400 473.600 194.000 474.400 ;
        RECT 201.200 473.600 202.000 479.800 ;
        RECT 204.400 475.000 205.200 479.800 ;
        RECT 207.600 475.000 208.400 479.800 ;
        RECT 209.200 477.000 210.000 479.800 ;
        RECT 210.800 477.000 211.600 479.800 ;
        RECT 214.000 475.200 214.800 479.800 ;
        RECT 217.200 476.400 218.000 479.800 ;
        RECT 217.200 475.800 218.200 476.400 ;
        RECT 217.600 475.200 218.200 475.800 ;
        RECT 212.800 474.400 217.000 475.200 ;
        RECT 217.600 474.600 219.600 475.200 ;
        RECT 204.400 473.600 207.000 474.400 ;
        RECT 207.600 473.800 213.400 474.400 ;
        RECT 216.400 474.000 217.000 474.400 ;
        RECT 196.400 473.000 197.200 473.200 ;
        RECT 188.200 472.400 197.200 473.000 ;
        RECT 199.600 473.000 200.400 473.200 ;
        RECT 207.600 473.000 208.200 473.800 ;
        RECT 214.000 473.200 215.400 473.800 ;
        RECT 216.400 473.200 218.000 474.000 ;
        RECT 199.600 472.400 208.200 473.000 ;
        RECT 209.200 473.000 215.400 473.200 ;
        RECT 209.200 472.600 214.600 473.000 ;
        RECT 209.200 472.400 210.000 472.600 ;
        RECT 185.200 468.300 186.000 468.400 ;
        RECT 182.000 467.700 186.000 468.300 ;
        RECT 180.400 464.800 181.200 466.400 ;
        RECT 182.000 462.200 182.800 467.700 ;
        RECT 185.200 467.600 186.000 467.700 ;
        RECT 186.600 466.800 187.400 471.200 ;
        RECT 188.200 470.600 188.800 472.400 ;
        RECT 188.000 470.000 188.800 470.600 ;
        RECT 194.800 470.000 218.200 470.600 ;
        RECT 188.000 468.000 188.600 470.000 ;
        RECT 194.800 469.400 195.600 470.000 ;
        RECT 212.400 469.600 213.200 470.000 ;
        RECT 215.600 469.600 216.400 470.000 ;
        RECT 217.400 469.800 218.200 470.000 ;
        RECT 189.200 468.600 193.000 469.400 ;
        RECT 188.000 467.400 189.200 468.000 ;
        RECT 183.600 466.300 184.400 466.400 ;
        RECT 186.600 466.300 187.600 466.800 ;
        RECT 183.600 465.700 187.600 466.300 ;
        RECT 183.600 464.800 184.400 465.700 ;
        RECT 186.800 462.200 187.600 465.700 ;
        RECT 188.400 462.200 189.200 467.400 ;
        RECT 192.200 467.400 193.000 468.600 ;
        RECT 192.200 466.800 194.000 467.400 ;
        RECT 193.200 466.200 194.000 466.800 ;
        RECT 198.000 466.400 198.800 469.200 ;
        RECT 201.200 468.600 204.400 469.400 ;
        RECT 208.200 468.600 210.200 469.400 ;
        RECT 218.800 469.000 219.600 474.600 ;
        RECT 220.400 472.400 221.200 479.800 ;
        RECT 221.800 472.400 222.600 472.600 ;
        RECT 220.400 471.800 222.600 472.400 ;
        RECT 224.800 472.400 226.400 479.800 ;
        RECT 228.400 472.400 229.200 472.600 ;
        RECT 230.000 472.400 230.800 479.800 ;
        RECT 224.800 471.800 226.800 472.400 ;
        RECT 228.400 471.800 230.800 472.400 ;
        RECT 233.200 472.000 234.000 479.800 ;
        RECT 236.400 475.200 237.200 479.800 ;
        RECT 222.000 471.200 222.600 471.800 ;
        RECT 222.000 470.600 225.400 471.200 ;
        RECT 224.600 470.400 225.400 470.600 ;
        RECT 226.200 470.400 226.800 471.800 ;
        RECT 233.000 471.200 234.000 472.000 ;
        RECT 234.600 474.600 237.200 475.200 ;
        RECT 234.600 473.000 235.200 474.600 ;
        RECT 239.600 474.400 240.400 479.800 ;
        RECT 242.800 477.000 243.600 479.800 ;
        RECT 244.400 477.000 245.200 479.800 ;
        RECT 246.000 477.000 246.800 479.800 ;
        RECT 241.000 474.400 245.200 475.200 ;
        RECT 237.800 473.600 240.400 474.400 ;
        RECT 247.600 473.600 248.400 479.800 ;
        RECT 250.800 475.000 251.600 479.800 ;
        RECT 254.000 475.000 254.800 479.800 ;
        RECT 255.600 477.000 256.400 479.800 ;
        RECT 257.200 477.000 258.000 479.800 ;
        RECT 260.400 475.200 261.200 479.800 ;
        RECT 263.600 476.400 264.400 479.800 ;
        RECT 274.200 478.400 275.000 479.800 ;
        RECT 273.200 477.600 275.000 478.400 ;
        RECT 263.600 475.800 264.600 476.400 ;
        RECT 264.000 475.200 264.600 475.800 ;
        RECT 259.200 474.400 263.400 475.200 ;
        RECT 264.000 474.600 266.000 475.200 ;
        RECT 250.800 473.600 253.400 474.400 ;
        RECT 254.000 473.800 259.800 474.400 ;
        RECT 262.800 474.000 263.400 474.400 ;
        RECT 242.800 473.000 243.600 473.200 ;
        RECT 234.600 472.400 243.600 473.000 ;
        RECT 246.000 473.000 246.800 473.200 ;
        RECT 254.000 473.000 254.600 473.800 ;
        RECT 260.400 473.200 261.800 473.800 ;
        RECT 262.800 473.200 264.400 474.000 ;
        RECT 246.000 472.400 254.600 473.000 ;
        RECT 255.600 473.000 261.800 473.200 ;
        RECT 255.600 472.600 261.000 473.000 ;
        RECT 255.600 472.400 256.400 472.600 ;
        RECT 226.200 470.300 227.600 470.400 ;
        RECT 231.600 470.300 232.400 470.400 ;
        RECT 222.400 469.800 223.200 470.000 ;
        RECT 226.200 469.800 232.400 470.300 ;
        RECT 222.400 469.200 225.000 469.800 ;
        RECT 200.800 467.800 201.600 468.000 ;
        RECT 200.800 467.200 205.200 467.800 ;
        RECT 204.400 467.000 205.200 467.200 ;
        RECT 206.000 466.800 206.800 468.400 ;
        RECT 193.200 465.400 195.600 466.200 ;
        RECT 198.000 465.600 199.000 466.400 ;
        RECT 202.000 465.600 203.600 466.400 ;
        RECT 204.400 466.200 205.200 466.400 ;
        RECT 208.200 466.200 209.000 468.600 ;
        RECT 210.800 468.200 219.600 469.000 ;
        RECT 224.400 468.600 225.000 469.200 ;
        RECT 225.800 469.700 232.400 469.800 ;
        RECT 225.800 469.600 227.600 469.700 ;
        RECT 231.600 469.600 232.400 469.700 ;
        RECT 225.800 469.200 226.800 469.600 ;
        RECT 214.200 466.800 217.200 467.600 ;
        RECT 214.200 466.200 215.000 466.800 ;
        RECT 204.400 465.600 209.000 466.200 ;
        RECT 194.800 462.200 195.600 465.400 ;
        RECT 212.400 465.400 215.000 466.200 ;
        RECT 196.400 462.200 197.200 465.000 ;
        RECT 198.000 462.200 198.800 465.000 ;
        RECT 199.600 462.200 200.400 465.000 ;
        RECT 201.200 462.200 202.000 465.000 ;
        RECT 204.400 462.200 205.200 465.000 ;
        RECT 207.600 462.200 208.400 465.000 ;
        RECT 209.200 462.200 210.000 465.000 ;
        RECT 210.800 462.200 211.600 465.000 ;
        RECT 212.400 462.200 213.200 465.400 ;
        RECT 218.800 462.200 219.600 468.200 ;
        RECT 220.400 468.200 222.000 468.400 ;
        RECT 220.400 467.600 223.800 468.200 ;
        RECT 224.400 467.800 225.200 468.600 ;
        RECT 223.200 467.200 223.800 467.600 ;
        RECT 221.800 466.800 222.600 467.000 ;
        RECT 220.400 466.200 222.600 466.800 ;
        RECT 223.200 466.600 225.200 467.200 ;
        RECT 223.600 466.400 225.200 466.600 ;
        RECT 220.400 462.200 221.200 466.200 ;
        RECT 225.800 465.800 226.400 469.200 ;
        RECT 227.200 467.600 228.000 468.400 ;
        RECT 229.200 468.300 230.800 468.400 ;
        RECT 233.000 468.300 233.800 471.200 ;
        RECT 234.600 470.600 235.200 472.400 ;
        RECT 229.200 467.700 233.800 468.300 ;
        RECT 229.200 467.600 230.800 467.700 ;
        RECT 227.200 467.200 227.800 467.600 ;
        RECT 227.000 466.400 227.800 467.200 ;
        RECT 228.400 466.800 229.200 467.000 ;
        RECT 233.000 466.800 233.800 467.700 ;
        RECT 234.400 470.000 235.200 470.600 ;
        RECT 241.200 470.000 264.600 470.600 ;
        RECT 234.400 468.000 235.000 470.000 ;
        RECT 241.200 469.400 242.000 470.000 ;
        RECT 258.800 469.600 259.600 470.000 ;
        RECT 260.400 469.600 261.200 470.000 ;
        RECT 263.800 469.800 264.600 470.000 ;
        RECT 235.600 468.600 239.400 469.400 ;
        RECT 234.400 467.400 235.600 468.000 ;
        RECT 228.400 466.200 230.800 466.800 ;
        RECT 224.800 462.200 226.400 465.800 ;
        RECT 230.000 462.200 230.800 466.200 ;
        RECT 233.000 466.000 234.000 466.800 ;
        RECT 233.200 462.200 234.000 466.000 ;
        RECT 234.800 462.200 235.600 467.400 ;
        RECT 238.600 467.400 239.400 468.600 ;
        RECT 238.600 466.800 240.400 467.400 ;
        RECT 239.600 466.200 240.400 466.800 ;
        RECT 244.400 466.400 245.200 469.200 ;
        RECT 247.600 468.600 250.800 469.400 ;
        RECT 254.600 468.600 256.600 469.400 ;
        RECT 265.200 469.000 266.000 474.600 ;
        RECT 274.200 472.400 275.000 477.600 ;
        RECT 275.600 473.600 276.400 474.400 ;
        RECT 275.800 472.400 276.400 473.600 ;
        RECT 274.200 471.800 275.200 472.400 ;
        RECT 275.800 471.800 277.200 472.400 ;
        RECT 247.200 467.800 248.000 468.000 ;
        RECT 247.200 467.200 251.600 467.800 ;
        RECT 250.800 467.000 251.600 467.200 ;
        RECT 252.400 466.800 253.200 468.400 ;
        RECT 239.600 465.400 242.000 466.200 ;
        RECT 244.400 465.600 245.400 466.400 ;
        RECT 248.400 465.600 250.000 466.400 ;
        RECT 250.800 466.200 251.600 466.400 ;
        RECT 254.600 466.200 255.400 468.600 ;
        RECT 257.200 468.200 266.000 469.000 ;
        RECT 273.200 468.800 274.000 470.400 ;
        RECT 274.600 468.400 275.200 471.800 ;
        RECT 276.400 471.600 277.200 471.800 ;
        RECT 276.400 470.300 277.200 470.400 ;
        RECT 278.000 470.300 278.800 479.800 ;
        RECT 282.800 471.200 283.600 479.800 ;
        RECT 286.000 471.200 286.800 479.800 ;
        RECT 289.200 471.200 290.000 479.800 ;
        RECT 292.400 471.200 293.200 479.800 ;
        RECT 298.200 474.300 299.000 479.800 ;
        RECT 302.600 478.400 303.400 479.800 ;
        RECT 302.600 477.600 304.400 478.400 ;
        RECT 301.200 474.300 302.000 474.400 ;
        RECT 298.200 473.700 302.000 474.300 ;
        RECT 298.200 472.600 299.000 473.700 ;
        RECT 297.200 471.800 299.000 472.600 ;
        RECT 301.200 473.600 302.000 473.700 ;
        RECT 301.200 472.400 301.800 473.600 ;
        RECT 302.600 472.400 303.400 477.600 ;
        RECT 309.400 472.600 310.200 479.800 ;
        RECT 314.200 472.600 315.000 479.800 ;
        RECT 300.400 471.800 301.800 472.400 ;
        RECT 302.400 471.800 303.400 472.400 ;
        RECT 308.400 471.800 310.200 472.600 ;
        RECT 313.200 471.800 315.000 472.600 ;
        RECT 282.800 470.400 284.600 471.200 ;
        RECT 286.000 470.400 288.200 471.200 ;
        RECT 289.200 470.400 291.400 471.200 ;
        RECT 292.400 470.400 294.800 471.200 ;
        RECT 276.400 469.700 278.800 470.300 ;
        RECT 276.400 469.600 277.200 469.700 ;
        RECT 260.600 466.800 263.600 467.600 ;
        RECT 260.600 466.200 261.400 466.800 ;
        RECT 250.800 465.600 255.400 466.200 ;
        RECT 241.200 462.200 242.000 465.400 ;
        RECT 258.800 465.400 261.400 466.200 ;
        RECT 242.800 462.200 243.600 465.000 ;
        RECT 244.400 462.200 245.200 465.000 ;
        RECT 246.000 462.200 246.800 465.000 ;
        RECT 247.600 462.200 248.400 465.000 ;
        RECT 250.800 462.200 251.600 465.000 ;
        RECT 254.000 462.200 254.800 465.000 ;
        RECT 255.600 462.200 256.400 465.000 ;
        RECT 257.200 462.200 258.000 465.000 ;
        RECT 258.800 462.200 259.600 465.400 ;
        RECT 265.200 462.200 266.000 468.200 ;
        RECT 271.600 468.200 272.400 468.400 ;
        RECT 271.600 467.600 273.200 468.200 ;
        RECT 274.600 467.600 277.200 468.400 ;
        RECT 272.400 467.200 273.200 467.600 ;
        RECT 271.800 466.200 275.400 466.600 ;
        RECT 276.400 466.200 277.000 467.600 ;
        RECT 271.600 466.000 275.600 466.200 ;
        RECT 271.600 462.200 272.400 466.000 ;
        RECT 274.800 462.200 275.600 466.000 ;
        RECT 276.400 462.200 277.200 466.200 ;
        RECT 278.000 462.200 278.800 469.700 ;
        RECT 283.800 469.000 284.600 470.400 ;
        RECT 287.400 469.000 288.200 470.400 ;
        RECT 290.600 469.000 291.400 470.400 ;
        RECT 281.200 468.200 283.000 469.000 ;
        RECT 283.800 468.200 286.400 469.000 ;
        RECT 287.400 468.200 289.800 469.000 ;
        RECT 290.600 468.200 293.200 469.000 ;
        RECT 281.200 467.600 282.000 468.200 ;
        RECT 283.800 467.600 284.600 468.200 ;
        RECT 287.400 467.600 288.200 468.200 ;
        RECT 290.600 467.600 291.400 468.200 ;
        RECT 294.000 467.600 294.800 470.400 ;
        RECT 297.400 468.400 298.000 471.800 ;
        RECT 300.400 471.600 301.200 471.800 ;
        RECT 298.800 469.600 299.600 471.200 ;
        RECT 302.400 468.400 303.000 471.800 ;
        RECT 303.600 470.300 304.400 470.400 ;
        RECT 308.600 470.300 309.200 471.800 ;
        RECT 303.600 469.700 309.200 470.300 ;
        RECT 303.600 468.800 304.400 469.700 ;
        RECT 308.600 468.400 309.200 469.700 ;
        RECT 310.000 469.600 310.800 471.200 ;
        RECT 311.600 470.300 312.400 470.400 ;
        RECT 313.400 470.300 314.000 471.800 ;
        RECT 316.400 471.600 317.200 473.200 ;
        RECT 311.600 469.700 314.000 470.300 ;
        RECT 311.600 469.600 312.400 469.700 ;
        RECT 313.400 468.400 314.000 469.700 ;
        RECT 314.800 470.300 315.600 471.200 ;
        RECT 316.400 470.300 317.200 470.400 ;
        RECT 314.800 469.700 317.200 470.300 ;
        RECT 314.800 469.600 315.600 469.700 ;
        RECT 316.400 469.600 317.200 469.700 ;
        RECT 297.200 467.600 298.000 468.400 ;
        RECT 300.400 467.600 303.000 468.400 ;
        RECT 305.200 468.200 306.000 468.400 ;
        RECT 304.400 467.600 306.000 468.200 ;
        RECT 308.400 467.600 309.200 468.400 ;
        RECT 313.200 467.600 314.000 468.400 ;
        RECT 282.800 466.800 284.600 467.600 ;
        RECT 286.000 466.800 288.200 467.600 ;
        RECT 289.200 466.800 291.400 467.600 ;
        RECT 292.400 466.800 294.800 467.600 ;
        RECT 279.600 464.800 280.400 466.400 ;
        RECT 282.800 462.200 283.600 466.800 ;
        RECT 286.000 462.200 286.800 466.800 ;
        RECT 289.200 462.200 290.000 466.800 ;
        RECT 292.400 462.200 293.200 466.800 ;
        RECT 295.600 464.800 296.400 466.400 ;
        RECT 297.400 464.200 298.000 467.600 ;
        RECT 300.600 466.200 301.200 467.600 ;
        RECT 304.400 467.200 305.200 467.600 ;
        RECT 302.200 466.200 305.800 466.600 ;
        RECT 297.200 462.200 298.000 464.200 ;
        RECT 300.400 462.200 301.200 466.200 ;
        RECT 302.000 466.000 306.000 466.200 ;
        RECT 302.000 462.200 302.800 466.000 ;
        RECT 305.200 462.200 306.000 466.000 ;
        RECT 306.800 464.800 307.600 466.400 ;
        RECT 308.600 464.200 309.200 467.600 ;
        RECT 310.000 466.300 310.800 466.400 ;
        RECT 311.600 466.300 312.400 466.400 ;
        RECT 310.000 465.700 312.400 466.300 ;
        RECT 310.000 465.600 310.800 465.700 ;
        RECT 311.600 464.800 312.400 465.700 ;
        RECT 313.400 464.200 314.000 467.600 ;
        RECT 314.800 466.300 315.600 466.400 ;
        RECT 318.000 466.300 318.800 479.800 ;
        RECT 319.600 472.300 320.400 472.400 ;
        RECT 321.200 472.300 322.000 479.800 ;
        RECT 319.600 471.700 322.000 472.300 ;
        RECT 322.800 472.400 323.600 479.800 ;
        RECT 326.000 472.400 326.800 479.800 ;
        RECT 322.800 471.800 326.800 472.400 ;
        RECT 319.600 471.600 320.400 471.700 ;
        RECT 321.400 470.400 322.000 471.700 ;
        RECT 325.200 470.400 326.000 470.800 ;
        RECT 321.200 469.800 323.600 470.400 ;
        RECT 325.200 469.800 326.800 470.400 ;
        RECT 321.200 469.600 322.000 469.800 ;
        RECT 319.600 466.800 320.400 468.400 ;
        RECT 314.800 465.700 318.800 466.300 ;
        RECT 314.800 465.600 315.600 465.700 ;
        RECT 317.000 465.600 318.800 465.700 ;
        RECT 321.200 465.600 322.000 466.400 ;
        RECT 323.000 466.200 323.600 469.800 ;
        RECT 326.000 469.600 326.800 469.800 ;
        RECT 324.400 467.600 325.200 469.200 ;
        RECT 327.600 466.800 328.400 468.400 ;
        RECT 308.400 462.200 309.200 464.200 ;
        RECT 313.200 462.200 314.000 464.200 ;
        RECT 317.000 462.200 317.800 465.600 ;
        RECT 321.400 464.800 322.200 465.600 ;
        RECT 322.800 462.200 323.600 466.200 ;
        RECT 329.200 466.200 330.000 479.800 ;
        RECT 330.800 471.600 331.600 473.200 ;
        RECT 332.400 466.800 333.200 468.400 ;
        RECT 334.000 466.200 334.800 479.800 ;
        RECT 335.600 471.600 336.400 473.200 ;
        RECT 339.800 472.400 340.600 479.800 ;
        RECT 341.200 473.600 342.000 474.400 ;
        RECT 341.400 472.400 342.000 473.600 ;
        RECT 339.800 471.800 340.800 472.400 ;
        RECT 341.400 472.300 342.800 472.400 ;
        RECT 345.200 472.300 346.000 479.800 ;
        RECT 341.400 471.800 346.000 472.300 ;
        RECT 338.800 468.800 339.600 470.400 ;
        RECT 340.200 470.300 340.800 471.800 ;
        RECT 342.000 471.700 346.000 471.800 ;
        RECT 342.000 471.600 342.800 471.700 ;
        RECT 343.600 470.300 344.400 470.400 ;
        RECT 340.200 469.700 344.400 470.300 ;
        RECT 340.200 468.400 340.800 469.700 ;
        RECT 343.600 469.600 344.400 469.700 ;
        RECT 335.600 468.300 336.400 468.400 ;
        RECT 337.200 468.300 338.000 468.400 ;
        RECT 335.600 468.200 338.000 468.300 ;
        RECT 335.600 467.700 338.800 468.200 ;
        RECT 335.600 467.600 336.400 467.700 ;
        RECT 337.200 467.600 338.800 467.700 ;
        RECT 340.200 467.600 342.800 468.400 ;
        RECT 338.000 467.200 338.800 467.600 ;
        RECT 337.400 466.200 341.000 466.600 ;
        RECT 342.000 466.200 342.600 467.600 ;
        RECT 343.600 466.800 344.400 468.400 ;
        RECT 345.200 466.200 346.000 471.700 ;
        RECT 346.800 471.600 347.600 473.200 ;
        RECT 346.800 468.300 347.600 468.400 ;
        RECT 348.400 468.300 349.200 468.400 ;
        RECT 346.800 467.700 349.200 468.300 ;
        RECT 346.800 467.600 347.600 467.700 ;
        RECT 348.400 466.800 349.200 467.700 ;
        RECT 329.200 465.600 331.000 466.200 ;
        RECT 334.000 465.600 335.800 466.200 ;
        RECT 330.200 464.400 331.000 465.600 ;
        RECT 335.000 464.400 335.800 465.600 ;
        RECT 337.200 466.000 341.200 466.200 ;
        RECT 330.200 463.600 331.600 464.400 ;
        RECT 335.000 463.600 336.400 464.400 ;
        RECT 330.200 462.200 331.000 463.600 ;
        RECT 335.000 462.200 335.800 463.600 ;
        RECT 337.200 462.200 338.000 466.000 ;
        RECT 340.400 462.200 341.200 466.000 ;
        RECT 342.000 462.200 342.800 466.200 ;
        RECT 345.200 465.600 347.000 466.200 ;
        RECT 346.200 462.200 347.000 465.600 ;
        RECT 350.000 462.200 350.800 479.800 ;
        RECT 353.200 471.600 354.000 473.200 ;
        RECT 354.800 466.200 355.600 479.800 ;
        RECT 356.400 468.300 357.200 468.400 ;
        RECT 358.000 468.300 358.800 479.800 ;
        RECT 356.400 467.700 358.800 468.300 ;
        RECT 356.400 466.800 357.200 467.700 ;
        RECT 353.800 465.600 355.600 466.200 ;
        RECT 353.800 464.400 354.600 465.600 ;
        RECT 353.800 463.600 355.600 464.400 ;
        RECT 353.800 462.200 354.600 463.600 ;
        RECT 358.000 462.200 358.800 467.700 ;
        RECT 359.600 468.300 360.400 468.400 ;
        RECT 361.200 468.300 362.000 468.400 ;
        RECT 359.600 467.700 362.000 468.300 ;
        RECT 359.600 466.800 360.400 467.700 ;
        RECT 361.200 466.800 362.000 467.700 ;
        RECT 362.800 466.200 363.600 479.800 ;
        RECT 366.800 473.600 367.600 474.400 ;
        RECT 364.400 471.600 365.200 473.200 ;
        RECT 366.800 472.400 367.400 473.600 ;
        RECT 368.200 472.400 369.000 479.800 ;
        RECT 366.000 471.800 367.400 472.400 ;
        RECT 368.000 471.800 369.000 472.400 ;
        RECT 372.400 472.300 373.200 472.400 ;
        RECT 374.000 472.300 374.800 479.800 ;
        RECT 378.800 476.400 379.600 479.800 ;
        RECT 378.600 475.800 379.600 476.400 ;
        RECT 378.600 475.200 379.200 475.800 ;
        RECT 382.000 475.200 382.800 479.800 ;
        RECT 385.200 477.000 386.000 479.800 ;
        RECT 386.800 477.000 387.600 479.800 ;
        RECT 377.200 474.600 379.200 475.200 ;
        RECT 366.000 471.600 366.800 471.800 ;
        RECT 364.500 470.300 365.100 471.600 ;
        RECT 368.000 470.300 368.600 471.800 ;
        RECT 372.400 471.700 374.800 472.300 ;
        RECT 372.400 471.600 373.200 471.700 ;
        RECT 364.500 469.700 368.600 470.300 ;
        RECT 368.000 468.400 368.600 469.700 ;
        RECT 369.200 468.800 370.000 470.400 ;
        RECT 366.000 467.600 368.600 468.400 ;
        RECT 370.800 468.300 371.600 468.400 ;
        RECT 372.400 468.300 373.200 468.400 ;
        RECT 370.800 468.200 373.200 468.300 ;
        RECT 370.000 467.700 373.200 468.200 ;
        RECT 370.000 467.600 371.600 467.700 ;
        RECT 366.200 466.200 366.800 467.600 ;
        RECT 370.000 467.200 370.800 467.600 ;
        RECT 372.400 466.800 373.200 467.700 ;
        RECT 367.800 466.200 371.400 466.600 ;
        RECT 374.000 466.200 374.800 471.700 ;
        RECT 375.600 471.600 376.400 473.200 ;
        RECT 377.200 469.000 378.000 474.600 ;
        RECT 379.800 474.400 384.000 475.200 ;
        RECT 388.400 475.000 389.200 479.800 ;
        RECT 391.600 475.000 392.400 479.800 ;
        RECT 379.800 474.000 380.400 474.400 ;
        RECT 378.800 473.200 380.400 474.000 ;
        RECT 383.400 473.800 389.200 474.400 ;
        RECT 381.400 473.200 382.800 473.800 ;
        RECT 381.400 473.000 387.600 473.200 ;
        RECT 382.200 472.600 387.600 473.000 ;
        RECT 386.800 472.400 387.600 472.600 ;
        RECT 388.600 473.000 389.200 473.800 ;
        RECT 389.800 473.600 392.400 474.400 ;
        RECT 394.800 473.600 395.600 479.800 ;
        RECT 396.400 477.000 397.200 479.800 ;
        RECT 398.000 477.000 398.800 479.800 ;
        RECT 399.600 477.000 400.400 479.800 ;
        RECT 398.000 474.400 402.200 475.200 ;
        RECT 402.800 474.400 403.600 479.800 ;
        RECT 406.000 475.200 406.800 479.800 ;
        RECT 406.000 474.600 408.600 475.200 ;
        RECT 402.800 473.600 405.400 474.400 ;
        RECT 396.400 473.000 397.200 473.200 ;
        RECT 388.600 472.400 397.200 473.000 ;
        RECT 399.600 473.000 400.400 473.200 ;
        RECT 408.000 473.000 408.600 474.600 ;
        RECT 399.600 472.400 408.600 473.000 ;
        RECT 408.000 470.600 408.600 472.400 ;
        RECT 409.200 472.000 410.000 479.800 ;
        RECT 409.200 471.200 410.200 472.000 ;
        RECT 378.600 470.000 402.000 470.600 ;
        RECT 408.000 470.000 408.800 470.600 ;
        RECT 378.600 469.800 379.400 470.000 ;
        RECT 383.600 469.600 384.400 470.000 ;
        RECT 401.200 469.400 402.000 470.000 ;
        RECT 377.200 468.200 386.000 469.000 ;
        RECT 386.600 468.600 388.600 469.400 ;
        RECT 392.400 468.600 395.600 469.400 ;
        RECT 362.800 465.600 364.600 466.200 ;
        RECT 363.800 464.400 364.600 465.600 ;
        RECT 363.800 463.600 365.200 464.400 ;
        RECT 363.800 462.200 364.600 463.600 ;
        RECT 366.000 462.200 366.800 466.200 ;
        RECT 367.600 466.000 371.600 466.200 ;
        RECT 367.600 462.200 368.400 466.000 ;
        RECT 370.800 462.200 371.600 466.000 ;
        RECT 374.000 465.600 375.800 466.200 ;
        RECT 375.000 462.200 375.800 465.600 ;
        RECT 377.200 462.200 378.000 468.200 ;
        RECT 379.600 466.800 382.600 467.600 ;
        RECT 381.800 466.200 382.600 466.800 ;
        RECT 387.800 466.200 388.600 468.600 ;
        RECT 390.000 466.800 390.800 468.400 ;
        RECT 395.200 467.800 396.000 468.000 ;
        RECT 391.600 467.200 396.000 467.800 ;
        RECT 391.600 467.000 392.400 467.200 ;
        RECT 398.000 466.400 398.800 469.200 ;
        RECT 403.800 468.600 407.600 469.400 ;
        RECT 403.800 467.400 404.600 468.600 ;
        RECT 408.200 468.000 408.800 470.000 ;
        RECT 391.600 466.200 392.400 466.400 ;
        RECT 381.800 465.400 384.400 466.200 ;
        RECT 387.800 465.600 392.400 466.200 ;
        RECT 393.200 465.600 394.800 466.400 ;
        RECT 397.800 465.600 398.800 466.400 ;
        RECT 402.800 466.800 404.600 467.400 ;
        RECT 407.600 467.400 408.800 468.000 ;
        RECT 402.800 466.200 403.600 466.800 ;
        RECT 383.600 462.200 384.400 465.400 ;
        RECT 401.200 465.400 403.600 466.200 ;
        RECT 385.200 462.200 386.000 465.000 ;
        RECT 386.800 462.200 387.600 465.000 ;
        RECT 388.400 462.200 389.200 465.000 ;
        RECT 391.600 462.200 392.400 465.000 ;
        RECT 394.800 462.200 395.600 465.000 ;
        RECT 396.400 462.200 397.200 465.000 ;
        RECT 398.000 462.200 398.800 465.000 ;
        RECT 399.600 462.200 400.400 465.000 ;
        RECT 401.200 462.200 402.000 465.400 ;
        RECT 407.600 462.200 408.400 467.400 ;
        RECT 409.400 466.800 410.200 471.200 ;
        RECT 409.200 466.300 410.200 466.800 ;
        RECT 414.000 470.300 414.800 479.800 ;
        RECT 421.200 473.600 422.000 474.400 ;
        RECT 421.200 472.400 421.800 473.600 ;
        RECT 422.600 472.400 423.400 479.800 ;
        RECT 420.400 471.800 421.800 472.400 ;
        RECT 422.400 471.800 423.400 472.400 ;
        RECT 420.400 471.600 421.200 471.800 ;
        RECT 420.400 470.300 421.200 470.400 ;
        RECT 414.000 469.700 421.200 470.300 ;
        RECT 412.400 466.300 413.200 466.400 ;
        RECT 409.200 465.700 413.200 466.300 ;
        RECT 409.200 462.200 410.000 465.700 ;
        RECT 412.400 464.800 413.200 465.700 ;
        RECT 414.000 462.200 414.800 469.700 ;
        RECT 420.400 469.600 421.200 469.700 ;
        RECT 422.400 468.400 423.000 471.800 ;
        RECT 426.800 471.600 427.600 473.200 ;
        RECT 423.600 468.800 424.400 470.400 ;
        RECT 415.600 468.300 416.400 468.400 ;
        RECT 420.400 468.300 423.000 468.400 ;
        RECT 415.600 467.700 423.000 468.300 ;
        RECT 425.200 468.300 426.000 468.400 ;
        RECT 426.800 468.300 427.600 468.400 ;
        RECT 425.200 468.200 427.600 468.300 ;
        RECT 415.600 467.600 416.400 467.700 ;
        RECT 420.400 467.600 423.000 467.700 ;
        RECT 424.400 467.700 427.600 468.200 ;
        RECT 424.400 467.600 426.000 467.700 ;
        RECT 426.800 467.600 427.600 467.700 ;
        RECT 420.600 466.200 421.200 467.600 ;
        RECT 424.400 467.200 425.200 467.600 ;
        RECT 422.200 466.200 425.800 466.600 ;
        RECT 428.400 466.200 429.200 479.800 ;
        RECT 432.400 473.600 433.200 474.400 ;
        RECT 432.400 472.400 433.000 473.600 ;
        RECT 433.800 472.400 434.600 479.800 ;
        RECT 430.000 472.300 430.800 472.400 ;
        RECT 431.600 472.300 433.000 472.400 ;
        RECT 430.000 471.800 433.000 472.300 ;
        RECT 433.600 471.800 434.600 472.400 ;
        RECT 440.600 472.400 441.400 479.800 ;
        RECT 442.000 473.600 443.600 474.400 ;
        RECT 442.200 472.400 442.800 473.600 ;
        RECT 440.600 471.800 441.600 472.400 ;
        RECT 442.200 471.800 443.600 472.400 ;
        RECT 446.000 472.000 446.800 479.800 ;
        RECT 449.200 475.200 450.000 479.800 ;
        RECT 430.000 471.700 432.400 471.800 ;
        RECT 430.000 471.600 430.800 471.700 ;
        RECT 431.600 471.600 432.400 471.700 ;
        RECT 433.600 468.400 434.200 471.800 ;
        RECT 434.800 470.300 435.600 470.400 ;
        RECT 439.600 470.300 440.400 470.400 ;
        RECT 434.800 469.700 440.400 470.300 ;
        RECT 434.800 468.800 435.600 469.700 ;
        RECT 439.600 468.800 440.400 469.700 ;
        RECT 441.000 468.400 441.600 471.800 ;
        RECT 442.800 471.600 443.600 471.800 ;
        RECT 445.800 471.200 446.800 472.000 ;
        RECT 447.400 474.600 450.000 475.200 ;
        RECT 447.400 473.000 448.000 474.600 ;
        RECT 452.400 474.400 453.200 479.800 ;
        RECT 455.600 477.000 456.400 479.800 ;
        RECT 457.200 477.000 458.000 479.800 ;
        RECT 458.800 477.000 459.600 479.800 ;
        RECT 453.800 474.400 458.000 475.200 ;
        RECT 450.600 473.600 453.200 474.400 ;
        RECT 460.400 473.600 461.200 479.800 ;
        RECT 463.600 475.000 464.400 479.800 ;
        RECT 466.800 475.000 467.600 479.800 ;
        RECT 468.400 477.000 469.200 479.800 ;
        RECT 470.000 477.000 470.800 479.800 ;
        RECT 473.200 475.200 474.000 479.800 ;
        RECT 476.400 476.400 477.200 479.800 ;
        RECT 481.200 476.400 482.000 479.800 ;
        RECT 476.400 475.800 477.400 476.400 ;
        RECT 476.800 475.200 477.400 475.800 ;
        RECT 481.000 475.800 482.000 476.400 ;
        RECT 481.000 475.200 481.600 475.800 ;
        RECT 484.400 475.200 485.200 479.800 ;
        RECT 487.600 477.000 488.400 479.800 ;
        RECT 489.200 477.000 490.000 479.800 ;
        RECT 472.000 474.400 476.200 475.200 ;
        RECT 476.800 474.600 478.800 475.200 ;
        RECT 463.600 473.600 466.200 474.400 ;
        RECT 466.800 473.800 472.600 474.400 ;
        RECT 475.600 474.000 476.200 474.400 ;
        RECT 455.600 473.000 456.400 473.200 ;
        RECT 447.400 472.400 456.400 473.000 ;
        RECT 458.800 473.000 459.600 473.200 ;
        RECT 466.800 473.000 467.400 473.800 ;
        RECT 473.200 473.200 474.600 473.800 ;
        RECT 475.600 473.200 477.200 474.000 ;
        RECT 458.800 472.400 467.400 473.000 ;
        RECT 468.400 473.000 474.600 473.200 ;
        RECT 468.400 472.600 473.800 473.000 ;
        RECT 468.400 472.400 469.200 472.600 ;
        RECT 430.000 466.800 430.800 468.400 ;
        RECT 431.600 467.600 434.200 468.400 ;
        RECT 436.400 468.300 437.200 468.400 ;
        RECT 438.000 468.300 438.800 468.400 ;
        RECT 436.400 468.200 438.800 468.300 ;
        RECT 435.600 467.700 439.600 468.200 ;
        RECT 435.600 467.600 437.200 467.700 ;
        RECT 438.000 467.600 439.600 467.700 ;
        RECT 441.000 467.600 443.600 468.400 ;
        RECT 431.800 466.200 432.400 467.600 ;
        RECT 435.600 467.200 436.400 467.600 ;
        RECT 438.800 467.200 439.600 467.600 ;
        RECT 433.400 466.200 437.000 466.600 ;
        RECT 438.200 466.200 441.800 466.600 ;
        RECT 442.800 466.200 443.400 467.600 ;
        RECT 445.800 466.800 446.600 471.200 ;
        RECT 447.400 470.600 448.000 472.400 ;
        RECT 447.200 470.000 448.000 470.600 ;
        RECT 454.000 470.000 477.400 470.600 ;
        RECT 447.200 468.000 447.800 470.000 ;
        RECT 454.000 469.400 454.800 470.000 ;
        RECT 471.600 469.600 472.400 470.000 ;
        RECT 474.800 469.600 475.600 470.000 ;
        RECT 476.600 469.800 477.400 470.000 ;
        RECT 448.400 468.600 452.200 469.400 ;
        RECT 447.200 467.400 448.400 468.000 ;
        RECT 420.400 462.200 421.200 466.200 ;
        RECT 422.000 466.000 426.000 466.200 ;
        RECT 422.000 462.200 422.800 466.000 ;
        RECT 425.200 462.200 426.000 466.000 ;
        RECT 427.400 465.600 429.200 466.200 ;
        RECT 427.400 462.200 428.200 465.600 ;
        RECT 431.600 462.200 432.400 466.200 ;
        RECT 433.200 466.000 437.200 466.200 ;
        RECT 433.200 462.200 434.000 466.000 ;
        RECT 436.400 462.200 437.200 466.000 ;
        RECT 438.000 466.000 442.000 466.200 ;
        RECT 438.000 462.200 438.800 466.000 ;
        RECT 441.200 462.200 442.000 466.000 ;
        RECT 442.800 462.200 443.600 466.200 ;
        RECT 445.800 466.000 446.800 466.800 ;
        RECT 446.000 462.200 446.800 466.000 ;
        RECT 447.600 462.200 448.400 467.400 ;
        RECT 451.400 467.400 452.200 468.600 ;
        RECT 451.400 466.800 453.200 467.400 ;
        RECT 452.400 466.200 453.200 466.800 ;
        RECT 457.200 466.400 458.000 469.200 ;
        RECT 460.400 468.600 463.600 469.400 ;
        RECT 467.400 468.600 469.400 469.400 ;
        RECT 478.000 469.000 478.800 474.600 ;
        RECT 460.000 467.800 460.800 468.000 ;
        RECT 460.000 467.200 464.400 467.800 ;
        RECT 463.600 467.000 464.400 467.200 ;
        RECT 465.200 466.800 466.000 468.400 ;
        RECT 452.400 465.400 454.800 466.200 ;
        RECT 457.200 465.600 458.200 466.400 ;
        RECT 461.200 465.600 462.800 466.400 ;
        RECT 463.600 466.200 464.400 466.400 ;
        RECT 467.400 466.200 468.200 468.600 ;
        RECT 470.000 468.200 478.800 469.000 ;
        RECT 473.400 466.800 476.400 467.600 ;
        RECT 473.400 466.200 474.200 466.800 ;
        RECT 463.600 465.600 468.200 466.200 ;
        RECT 454.000 462.200 454.800 465.400 ;
        RECT 471.600 465.400 474.200 466.200 ;
        RECT 455.600 462.200 456.400 465.000 ;
        RECT 457.200 462.200 458.000 465.000 ;
        RECT 458.800 462.200 459.600 465.000 ;
        RECT 460.400 462.200 461.200 465.000 ;
        RECT 463.600 462.200 464.400 465.000 ;
        RECT 466.800 462.200 467.600 465.000 ;
        RECT 468.400 462.200 469.200 465.000 ;
        RECT 470.000 462.200 470.800 465.000 ;
        RECT 471.600 462.200 472.400 465.400 ;
        RECT 478.000 462.200 478.800 468.200 ;
        RECT 479.600 474.600 481.600 475.200 ;
        RECT 479.600 469.000 480.400 474.600 ;
        RECT 482.200 474.400 486.400 475.200 ;
        RECT 490.800 475.000 491.600 479.800 ;
        RECT 494.000 475.000 494.800 479.800 ;
        RECT 482.200 474.000 482.800 474.400 ;
        RECT 481.200 473.200 482.800 474.000 ;
        RECT 485.800 473.800 491.600 474.400 ;
        RECT 483.800 473.200 485.200 473.800 ;
        RECT 483.800 473.000 490.000 473.200 ;
        RECT 484.600 472.600 490.000 473.000 ;
        RECT 489.200 472.400 490.000 472.600 ;
        RECT 491.000 473.000 491.600 473.800 ;
        RECT 492.200 473.600 494.800 474.400 ;
        RECT 497.200 473.600 498.000 479.800 ;
        RECT 498.800 477.000 499.600 479.800 ;
        RECT 500.400 477.000 501.200 479.800 ;
        RECT 502.000 477.000 502.800 479.800 ;
        RECT 500.400 474.400 504.600 475.200 ;
        RECT 505.200 474.400 506.000 479.800 ;
        RECT 508.400 475.200 509.200 479.800 ;
        RECT 508.400 474.600 511.000 475.200 ;
        RECT 505.200 473.600 507.800 474.400 ;
        RECT 498.800 473.000 499.600 473.200 ;
        RECT 491.000 472.400 499.600 473.000 ;
        RECT 502.000 473.000 502.800 473.200 ;
        RECT 510.400 473.000 511.000 474.600 ;
        RECT 502.000 472.400 511.000 473.000 ;
        RECT 510.400 470.600 511.000 472.400 ;
        RECT 511.600 474.300 512.400 479.800 ;
        RECT 515.600 474.300 516.400 474.400 ;
        RECT 511.600 473.700 516.400 474.300 ;
        RECT 511.600 472.000 512.400 473.700 ;
        RECT 515.600 473.600 516.400 473.700 ;
        RECT 515.600 472.400 516.200 473.600 ;
        RECT 517.000 472.400 517.800 479.800 ;
        RECT 511.600 471.200 512.600 472.000 ;
        RECT 514.800 471.800 516.200 472.400 ;
        RECT 516.800 471.800 517.800 472.400 ;
        RECT 523.800 472.400 524.600 479.800 ;
        RECT 525.200 473.600 526.000 474.400 ;
        RECT 525.400 472.400 526.000 473.600 ;
        RECT 523.800 471.800 524.800 472.400 ;
        RECT 525.400 471.800 526.800 472.400 ;
        RECT 514.800 471.600 515.600 471.800 ;
        RECT 481.000 470.000 504.400 470.600 ;
        RECT 510.400 470.000 511.200 470.600 ;
        RECT 481.000 469.800 481.800 470.000 ;
        RECT 484.400 469.600 485.200 470.000 ;
        RECT 486.000 469.600 486.800 470.000 ;
        RECT 503.600 469.400 504.400 470.000 ;
        RECT 479.600 468.200 488.400 469.000 ;
        RECT 489.000 468.600 491.000 469.400 ;
        RECT 494.800 468.600 498.000 469.400 ;
        RECT 479.600 462.200 480.400 468.200 ;
        RECT 482.000 466.800 485.000 467.600 ;
        RECT 484.200 466.200 485.000 466.800 ;
        RECT 490.200 466.200 491.000 468.600 ;
        RECT 492.400 466.800 493.200 468.400 ;
        RECT 497.600 467.800 498.400 468.000 ;
        RECT 494.000 467.200 498.400 467.800 ;
        RECT 494.000 467.000 494.800 467.200 ;
        RECT 500.400 466.400 501.200 469.200 ;
        RECT 506.200 468.600 510.000 469.400 ;
        RECT 506.200 467.400 507.000 468.600 ;
        RECT 510.600 468.000 511.200 470.000 ;
        RECT 494.000 466.200 494.800 466.400 ;
        RECT 484.200 465.400 486.800 466.200 ;
        RECT 490.200 465.600 494.800 466.200 ;
        RECT 495.600 465.600 497.200 466.400 ;
        RECT 500.200 465.600 501.200 466.400 ;
        RECT 505.200 466.800 507.000 467.400 ;
        RECT 510.000 467.400 511.200 468.000 ;
        RECT 505.200 466.200 506.000 466.800 ;
        RECT 486.000 462.200 486.800 465.400 ;
        RECT 503.600 465.400 506.000 466.200 ;
        RECT 487.600 462.200 488.400 465.000 ;
        RECT 489.200 462.200 490.000 465.000 ;
        RECT 490.800 462.200 491.600 465.000 ;
        RECT 494.000 462.200 494.800 465.000 ;
        RECT 497.200 462.200 498.000 465.000 ;
        RECT 498.800 462.200 499.600 465.000 ;
        RECT 500.400 462.200 501.200 465.000 ;
        RECT 502.000 462.200 502.800 465.000 ;
        RECT 503.600 462.200 504.400 465.400 ;
        RECT 510.000 462.200 510.800 467.400 ;
        RECT 511.800 466.800 512.600 471.200 ;
        RECT 516.800 468.400 517.400 471.800 ;
        RECT 518.000 470.300 518.800 470.400 ;
        RECT 522.800 470.300 523.600 470.400 ;
        RECT 518.000 469.700 523.600 470.300 ;
        RECT 518.000 468.800 518.800 469.700 ;
        RECT 522.800 468.800 523.600 469.700 ;
        RECT 524.200 468.400 524.800 471.800 ;
        RECT 526.000 471.600 526.800 471.800 ;
        RECT 514.800 467.600 517.400 468.400 ;
        RECT 519.600 468.300 520.400 468.400 ;
        RECT 521.200 468.300 522.000 468.400 ;
        RECT 519.600 468.200 522.000 468.300 ;
        RECT 518.800 467.700 522.800 468.200 ;
        RECT 518.800 467.600 520.400 467.700 ;
        RECT 521.200 467.600 522.800 467.700 ;
        RECT 524.200 467.600 526.800 468.400 ;
        RECT 511.600 466.000 512.600 466.800 ;
        RECT 515.000 466.200 515.600 467.600 ;
        RECT 518.800 467.200 519.600 467.600 ;
        RECT 522.000 467.200 522.800 467.600 ;
        RECT 516.600 466.200 520.200 466.600 ;
        RECT 521.400 466.200 525.000 466.600 ;
        RECT 526.000 466.200 526.600 467.600 ;
        RECT 527.600 466.800 528.400 468.400 ;
        RECT 529.200 466.200 530.000 479.800 ;
        RECT 534.000 474.300 534.800 479.800 ;
        RECT 537.200 475.200 538.000 479.800 ;
        RECT 530.800 473.700 534.800 474.300 ;
        RECT 530.800 471.600 531.600 473.700 ;
        RECT 534.000 472.000 534.800 473.700 ;
        RECT 533.800 471.200 534.800 472.000 ;
        RECT 535.400 474.600 538.000 475.200 ;
        RECT 535.400 473.000 536.000 474.600 ;
        RECT 540.400 474.400 541.200 479.800 ;
        RECT 543.600 477.000 544.400 479.800 ;
        RECT 545.200 477.000 546.000 479.800 ;
        RECT 546.800 477.000 547.600 479.800 ;
        RECT 541.800 474.400 546.000 475.200 ;
        RECT 538.600 473.600 541.200 474.400 ;
        RECT 548.400 473.600 549.200 479.800 ;
        RECT 551.600 475.000 552.400 479.800 ;
        RECT 554.800 475.000 555.600 479.800 ;
        RECT 556.400 477.000 557.200 479.800 ;
        RECT 558.000 477.000 558.800 479.800 ;
        RECT 561.200 475.200 562.000 479.800 ;
        RECT 564.400 476.400 565.200 479.800 ;
        RECT 564.400 475.800 565.400 476.400 ;
        RECT 564.800 475.200 565.400 475.800 ;
        RECT 560.000 474.400 564.200 475.200 ;
        RECT 564.800 474.600 566.800 475.200 ;
        RECT 551.600 473.600 554.200 474.400 ;
        RECT 554.800 473.800 560.600 474.400 ;
        RECT 563.600 474.000 564.200 474.400 ;
        RECT 543.600 473.000 544.400 473.200 ;
        RECT 535.400 472.400 544.400 473.000 ;
        RECT 546.800 473.000 547.600 473.200 ;
        RECT 554.800 473.000 555.400 473.800 ;
        RECT 561.200 473.200 562.600 473.800 ;
        RECT 563.600 473.200 565.200 474.000 ;
        RECT 546.800 472.400 555.400 473.000 ;
        RECT 556.400 473.000 562.600 473.200 ;
        RECT 556.400 472.600 561.800 473.000 ;
        RECT 556.400 472.400 557.200 472.600 ;
        RECT 533.800 466.800 534.600 471.200 ;
        RECT 535.400 470.600 536.000 472.400 ;
        RECT 535.200 470.000 536.000 470.600 ;
        RECT 542.000 470.000 565.400 470.600 ;
        RECT 535.200 468.000 535.800 470.000 ;
        RECT 542.000 469.400 542.800 470.000 ;
        RECT 559.600 469.600 560.400 470.000 ;
        RECT 562.800 469.600 563.600 470.000 ;
        RECT 564.600 469.800 565.400 470.000 ;
        RECT 536.400 468.600 540.200 469.400 ;
        RECT 535.200 467.400 536.400 468.000 ;
        RECT 511.600 462.200 512.400 466.000 ;
        RECT 514.800 462.200 515.600 466.200 ;
        RECT 516.400 466.000 520.400 466.200 ;
        RECT 516.400 462.200 517.200 466.000 ;
        RECT 519.600 462.200 520.400 466.000 ;
        RECT 521.200 466.000 525.200 466.200 ;
        RECT 521.200 462.200 522.000 466.000 ;
        RECT 524.400 462.200 525.200 466.000 ;
        RECT 526.000 462.200 526.800 466.200 ;
        RECT 529.200 465.600 531.000 466.200 ;
        RECT 533.800 466.000 534.800 466.800 ;
        RECT 530.200 462.200 531.000 465.600 ;
        RECT 534.000 462.200 534.800 466.000 ;
        RECT 535.600 462.200 536.400 467.400 ;
        RECT 539.400 467.400 540.200 468.600 ;
        RECT 539.400 466.800 541.200 467.400 ;
        RECT 540.400 466.200 541.200 466.800 ;
        RECT 545.200 466.400 546.000 469.200 ;
        RECT 548.400 468.600 551.600 469.400 ;
        RECT 555.400 468.600 557.400 469.400 ;
        RECT 566.000 469.000 566.800 474.600 ;
        RECT 567.600 471.200 568.400 479.800 ;
        RECT 571.800 472.400 572.600 479.800 ;
        RECT 581.400 472.400 582.200 479.800 ;
        RECT 582.800 473.600 583.600 474.400 ;
        RECT 583.000 472.400 583.600 473.600 ;
        RECT 571.800 471.800 573.200 472.400 ;
        RECT 581.400 471.800 582.400 472.400 ;
        RECT 583.000 471.800 584.400 472.400 ;
        RECT 567.600 470.800 571.600 471.200 ;
        RECT 567.600 470.600 571.800 470.800 ;
        RECT 571.000 470.000 571.800 470.600 ;
        RECT 572.600 470.400 573.200 471.800 ;
        RECT 548.000 467.800 548.800 468.000 ;
        RECT 548.000 467.200 552.400 467.800 ;
        RECT 551.600 467.000 552.400 467.200 ;
        RECT 553.200 466.800 554.000 468.400 ;
        RECT 540.400 465.400 542.800 466.200 ;
        RECT 545.200 465.600 546.200 466.400 ;
        RECT 549.200 465.600 550.800 466.400 ;
        RECT 551.600 466.200 552.400 466.400 ;
        RECT 555.400 466.200 556.200 468.600 ;
        RECT 558.000 468.200 566.800 469.000 ;
        RECT 569.600 468.400 570.400 469.200 ;
        RECT 561.400 466.800 564.400 467.600 ;
        RECT 561.400 466.200 562.200 466.800 ;
        RECT 551.600 465.600 556.200 466.200 ;
        RECT 542.000 462.200 542.800 465.400 ;
        RECT 559.600 465.400 562.200 466.200 ;
        RECT 543.600 462.200 544.400 465.000 ;
        RECT 545.200 462.200 546.000 465.000 ;
        RECT 546.800 462.200 547.600 465.000 ;
        RECT 548.400 462.200 549.200 465.000 ;
        RECT 551.600 462.200 552.400 465.000 ;
        RECT 554.800 462.200 555.600 465.000 ;
        RECT 556.400 462.200 557.200 465.000 ;
        RECT 558.000 462.200 558.800 465.000 ;
        RECT 559.600 462.200 560.400 465.400 ;
        RECT 566.000 462.200 566.800 468.200 ;
        RECT 569.200 467.600 570.200 468.400 ;
        RECT 571.200 467.000 571.800 470.000 ;
        RECT 572.400 469.600 573.200 470.400 ;
        RECT 575.600 470.300 576.400 470.400 ;
        RECT 580.400 470.300 581.200 470.400 ;
        RECT 575.600 469.700 581.200 470.300 ;
        RECT 575.600 469.600 576.400 469.700 ;
        RECT 569.400 466.400 571.800 467.000 ;
        RECT 567.600 464.800 568.400 466.400 ;
        RECT 569.400 464.200 570.000 466.400 ;
        RECT 572.600 466.300 573.200 469.600 ;
        RECT 580.400 468.800 581.200 469.700 ;
        RECT 581.800 470.300 582.400 471.800 ;
        RECT 583.600 471.600 584.400 471.800 ;
        RECT 585.200 470.300 586.000 470.400 ;
        RECT 581.800 469.700 586.000 470.300 ;
        RECT 581.800 468.400 582.400 469.700 ;
        RECT 585.200 469.600 586.000 469.700 ;
        RECT 577.200 468.300 578.000 468.400 ;
        RECT 578.800 468.300 579.600 468.400 ;
        RECT 577.200 468.200 579.600 468.300 ;
        RECT 577.200 467.700 580.400 468.200 ;
        RECT 577.200 467.600 578.000 467.700 ;
        RECT 578.800 467.600 580.400 467.700 ;
        RECT 581.800 467.600 584.400 468.400 ;
        RECT 579.600 467.200 580.400 467.600 ;
        RECT 577.200 466.300 578.000 466.400 ;
        RECT 572.500 466.200 578.000 466.300 ;
        RECT 579.000 466.200 582.600 466.600 ;
        RECT 583.600 466.200 584.200 467.600 ;
        RECT 585.200 466.800 586.000 468.400 ;
        RECT 586.800 466.200 587.600 479.800 ;
        RECT 590.800 473.600 591.600 474.400 ;
        RECT 588.400 471.600 589.200 473.200 ;
        RECT 590.800 472.400 591.400 473.600 ;
        RECT 592.200 472.400 593.000 479.800 ;
        RECT 590.000 471.800 591.400 472.400 ;
        RECT 592.000 471.800 593.000 472.400 ;
        RECT 596.400 471.800 597.200 479.800 ;
        RECT 599.600 475.800 600.400 479.800 ;
        RECT 590.000 471.600 590.800 471.800 ;
        RECT 588.500 470.300 589.100 471.600 ;
        RECT 592.000 470.300 592.600 471.800 ;
        RECT 596.400 470.400 597.000 471.800 ;
        RECT 599.600 471.600 600.200 475.800 ;
        RECT 597.800 471.000 600.200 471.600 ;
        RECT 588.500 469.700 592.600 470.300 ;
        RECT 592.000 468.400 592.600 469.700 ;
        RECT 593.200 468.800 594.000 470.400 ;
        RECT 596.400 470.300 597.200 470.400 ;
        RECT 594.900 469.700 597.200 470.300 ;
        RECT 594.900 468.400 595.500 469.700 ;
        RECT 596.400 469.600 597.200 469.700 ;
        RECT 590.000 467.600 592.600 468.400 ;
        RECT 594.800 468.200 595.600 468.400 ;
        RECT 594.000 467.600 595.600 468.200 ;
        RECT 590.200 466.200 590.800 467.600 ;
        RECT 594.000 467.200 594.800 467.600 ;
        RECT 591.800 466.200 595.400 466.600 ;
        RECT 596.400 466.200 597.000 469.600 ;
        RECT 597.800 467.600 598.400 471.000 ;
        RECT 599.600 469.600 600.400 470.400 ;
        RECT 599.600 468.800 600.200 469.600 ;
        RECT 599.200 468.200 600.200 468.800 ;
        RECT 599.200 468.000 600.000 468.200 ;
        RECT 601.200 467.600 602.000 469.200 ;
        RECT 597.600 467.400 598.400 467.600 ;
        RECT 597.600 467.000 600.600 467.400 ;
        RECT 597.600 466.800 601.800 467.000 ;
        RECT 600.000 466.400 601.800 466.800 ;
        RECT 601.200 466.200 601.800 466.400 ;
        RECT 569.200 462.200 570.000 464.200 ;
        RECT 572.400 465.700 578.000 466.200 ;
        RECT 572.400 462.200 573.200 465.700 ;
        RECT 577.200 465.600 578.000 465.700 ;
        RECT 578.800 466.000 582.800 466.200 ;
        RECT 578.800 462.200 579.600 466.000 ;
        RECT 582.000 462.200 582.800 466.000 ;
        RECT 583.600 462.200 584.400 466.200 ;
        RECT 586.800 465.600 588.600 466.200 ;
        RECT 587.800 462.200 588.600 465.600 ;
        RECT 590.000 462.200 590.800 466.200 ;
        RECT 591.600 466.000 595.600 466.200 ;
        RECT 591.600 462.200 592.400 466.000 ;
        RECT 594.800 462.200 595.600 466.000 ;
        RECT 596.400 465.200 597.800 466.200 ;
        RECT 597.000 462.200 597.800 465.200 ;
        RECT 601.200 462.200 602.000 466.200 ;
        RECT 602.800 462.200 603.600 479.800 ;
        RECT 606.800 473.600 607.600 474.400 ;
        RECT 606.800 472.400 607.400 473.600 ;
        RECT 608.200 472.400 609.000 479.800 ;
        RECT 606.000 471.800 607.400 472.400 ;
        RECT 608.000 471.800 609.000 472.400 ;
        RECT 606.000 471.600 606.800 471.800 ;
        RECT 608.000 468.400 608.600 471.800 ;
        RECT 609.200 468.800 610.000 470.400 ;
        RECT 606.000 467.600 608.600 468.400 ;
        RECT 610.800 468.200 611.600 468.400 ;
        RECT 610.000 467.600 611.600 468.200 ;
        RECT 604.400 466.300 605.200 466.400 ;
        RECT 606.200 466.300 606.800 467.600 ;
        RECT 610.000 467.200 610.800 467.600 ;
        RECT 612.400 466.800 613.200 468.400 ;
        RECT 604.400 465.700 606.800 466.300 ;
        RECT 607.800 466.200 611.400 466.600 ;
        RECT 614.000 466.200 614.800 479.800 ;
        RECT 615.600 471.600 616.400 473.200 ;
        RECT 617.200 471.600 618.000 473.200 ;
        RECT 615.700 470.300 616.300 471.600 ;
        RECT 618.800 470.300 619.600 479.800 ;
        RECT 622.000 472.400 622.800 479.800 ;
        RECT 623.600 472.400 624.400 472.600 ;
        RECT 622.000 471.800 624.400 472.400 ;
        RECT 626.400 471.800 628.000 479.800 ;
        RECT 629.800 472.400 630.600 472.600 ;
        RECT 631.600 472.400 632.400 479.800 ;
        RECT 629.800 471.800 632.400 472.400 ;
        RECT 633.200 475.000 634.000 479.000 ;
        RECT 615.700 469.700 619.600 470.300 ;
        RECT 618.800 466.200 619.600 469.700 ;
        RECT 626.800 470.400 627.400 471.800 ;
        RECT 633.200 471.600 633.800 475.000 ;
        RECT 637.400 472.800 638.200 479.800 ;
        RECT 642.800 475.000 643.600 479.000 ;
        RECT 637.400 472.200 639.000 472.800 ;
        RECT 633.200 471.000 637.000 471.600 ;
        RECT 628.600 470.400 629.400 470.600 ;
        RECT 626.800 469.600 627.600 470.400 ;
        RECT 628.600 469.800 630.200 470.400 ;
        RECT 629.400 469.600 630.200 469.800 ;
        RECT 626.800 468.400 627.400 469.600 ;
        RECT 633.200 468.800 634.000 470.400 ;
        RECT 634.800 468.800 635.600 470.400 ;
        RECT 636.400 469.000 637.000 471.000 ;
        RECT 620.400 466.800 621.200 468.400 ;
        RECT 622.000 467.600 623.600 468.400 ;
        RECT 624.800 467.600 625.600 468.400 ;
        RECT 625.000 467.200 625.600 467.600 ;
        RECT 626.400 467.800 627.400 468.400 ;
        RECT 628.000 468.600 628.800 468.800 ;
        RECT 628.000 468.400 630.800 468.600 ;
        RECT 628.000 468.000 632.400 468.400 ;
        RECT 630.200 467.800 632.400 468.000 ;
        RECT 636.400 468.200 637.800 469.000 ;
        RECT 638.400 468.400 639.000 472.200 ;
        RECT 642.800 471.600 643.400 475.000 ;
        RECT 647.000 472.800 647.800 479.800 ;
        RECT 653.200 473.600 654.000 474.400 ;
        RECT 647.000 472.200 648.600 472.800 ;
        RECT 653.200 472.400 653.800 473.600 ;
        RECT 654.600 472.400 655.400 479.800 ;
        RECT 639.600 469.600 640.400 471.200 ;
        RECT 642.800 471.000 646.600 471.600 ;
        RECT 642.800 468.800 643.600 470.400 ;
        RECT 644.400 468.800 645.200 470.400 ;
        RECT 646.000 469.000 646.600 471.000 ;
        RECT 638.400 468.300 640.400 468.400 ;
        RECT 641.200 468.300 642.000 468.400 ;
        RECT 636.400 467.800 637.400 468.200 ;
        RECT 623.600 466.800 624.400 467.000 ;
        RECT 604.400 464.800 605.200 465.700 ;
        RECT 606.000 462.200 606.800 465.700 ;
        RECT 607.600 466.000 611.600 466.200 ;
        RECT 607.600 462.200 608.400 466.000 ;
        RECT 610.800 462.200 611.600 466.000 ;
        RECT 614.000 465.600 615.800 466.200 ;
        RECT 615.000 464.400 615.800 465.600 ;
        RECT 614.000 463.600 615.800 464.400 ;
        RECT 615.000 462.200 615.800 463.600 ;
        RECT 617.800 465.600 619.600 466.200 ;
        RECT 622.000 466.200 624.400 466.800 ;
        RECT 625.000 466.400 625.800 467.200 ;
        RECT 617.800 462.200 618.600 465.600 ;
        RECT 622.000 462.200 622.800 466.200 ;
        RECT 626.400 465.800 627.000 467.800 ;
        RECT 630.800 467.600 632.400 467.800 ;
        RECT 633.200 467.200 637.400 467.800 ;
        RECT 638.400 467.700 642.000 468.300 ;
        RECT 646.000 468.200 647.400 469.000 ;
        RECT 648.000 468.400 648.600 472.200 ;
        RECT 652.400 471.800 653.800 472.400 ;
        RECT 654.400 471.800 655.400 472.400 ;
        RECT 652.400 471.600 653.200 471.800 ;
        RECT 649.200 469.600 650.000 471.200 ;
        RECT 654.400 468.400 655.000 471.800 ;
        RECT 658.800 471.200 659.600 479.800 ;
        RECT 663.000 475.800 664.200 479.800 ;
        RECT 667.600 475.800 668.400 479.800 ;
        RECT 672.000 476.400 672.800 479.800 ;
        RECT 672.000 475.800 674.000 476.400 ;
        RECT 663.600 475.000 664.400 475.800 ;
        RECT 667.800 475.200 668.400 475.800 ;
        RECT 667.000 474.600 670.600 475.200 ;
        RECT 673.200 475.000 674.000 475.800 ;
        RECT 667.000 474.400 667.800 474.600 ;
        RECT 669.800 474.400 670.600 474.600 ;
        RECT 662.800 473.200 664.200 474.000 ;
        RECT 663.600 472.200 664.200 473.200 ;
        RECT 665.800 473.000 668.000 473.600 ;
        RECT 665.800 472.800 666.600 473.000 ;
        RECT 663.600 471.600 666.000 472.200 ;
        RECT 658.800 470.600 663.000 471.200 ;
        RECT 655.600 468.800 656.400 470.400 ;
        RECT 646.000 467.800 647.000 468.200 ;
        RECT 638.400 467.600 640.400 467.700 ;
        RECT 641.200 467.600 642.000 467.700 ;
        RECT 627.600 466.400 629.200 467.200 ;
        RECT 629.800 466.800 630.600 467.000 ;
        RECT 629.800 466.200 632.400 466.800 ;
        RECT 626.400 462.200 628.000 465.800 ;
        RECT 631.600 462.200 632.400 466.200 ;
        RECT 633.200 465.000 633.800 467.200 ;
        RECT 638.400 467.000 639.000 467.600 ;
        RECT 638.200 466.600 639.000 467.000 ;
        RECT 637.400 466.000 639.000 466.600 ;
        RECT 642.800 467.200 647.000 467.800 ;
        RECT 648.000 467.600 650.000 468.400 ;
        RECT 652.400 467.600 655.000 468.400 ;
        RECT 657.200 468.200 658.000 468.400 ;
        RECT 656.400 467.600 658.000 468.200 ;
        RECT 633.200 463.000 634.000 465.000 ;
        RECT 637.400 463.000 638.200 466.000 ;
        RECT 642.800 465.000 643.400 467.200 ;
        RECT 648.000 467.000 648.600 467.600 ;
        RECT 647.800 466.600 648.600 467.000 ;
        RECT 647.000 466.000 648.600 466.600 ;
        RECT 652.600 466.200 653.200 467.600 ;
        RECT 656.400 467.200 657.200 467.600 ;
        RECT 658.800 467.200 659.600 470.600 ;
        RECT 662.200 470.400 663.000 470.600 ;
        RECT 660.600 469.800 661.400 470.000 ;
        RECT 660.600 469.200 664.400 469.800 ;
        RECT 663.600 469.000 664.400 469.200 ;
        RECT 665.400 468.400 666.000 471.600 ;
        RECT 667.400 471.800 668.000 473.000 ;
        RECT 668.600 473.000 669.400 473.200 ;
        RECT 673.200 473.000 674.000 473.200 ;
        RECT 668.600 472.400 674.000 473.000 ;
        RECT 667.400 471.400 672.200 471.800 ;
        RECT 676.400 471.400 677.200 479.800 ;
        RECT 678.000 472.400 678.800 479.800 ;
        RECT 678.000 471.800 680.200 472.400 ;
        RECT 667.400 471.200 677.200 471.400 ;
        RECT 671.400 471.000 677.200 471.200 ;
        RECT 671.600 470.800 677.200 471.000 ;
        RECT 679.600 471.200 680.200 471.800 ;
        RECT 679.600 470.400 680.800 471.200 ;
        RECT 670.000 470.200 670.800 470.400 ;
        RECT 670.000 469.600 675.000 470.200 ;
        RECT 674.200 469.400 675.000 469.600 ;
        RECT 678.000 468.800 678.800 470.400 ;
        RECT 672.600 468.400 673.400 468.600 ;
        RECT 665.400 467.800 676.400 468.400 ;
        RECT 665.800 467.600 666.600 467.800 ;
        RECT 658.800 466.600 662.600 467.200 ;
        RECT 654.200 466.200 657.800 466.600 ;
        RECT 642.800 463.000 643.600 465.000 ;
        RECT 647.000 464.400 647.800 466.000 ;
        RECT 647.000 463.600 648.400 464.400 ;
        RECT 647.000 463.000 647.800 463.600 ;
        RECT 652.400 462.200 653.200 466.200 ;
        RECT 654.000 466.000 658.000 466.200 ;
        RECT 654.000 462.200 654.800 466.000 ;
        RECT 657.200 462.200 658.000 466.000 ;
        RECT 658.800 462.200 659.600 466.600 ;
        RECT 661.800 466.400 662.600 466.600 ;
        RECT 671.600 465.600 672.200 467.800 ;
        RECT 674.800 467.600 676.400 467.800 ;
        RECT 679.600 467.400 680.200 470.400 ;
        RECT 669.800 465.400 670.600 465.600 ;
        RECT 663.600 464.200 664.400 465.000 ;
        RECT 667.800 464.800 670.600 465.400 ;
        RECT 671.600 464.800 672.400 465.600 ;
        RECT 667.800 464.200 668.400 464.800 ;
        RECT 673.200 464.200 674.000 465.000 ;
        RECT 663.000 463.600 664.400 464.200 ;
        RECT 663.000 462.200 664.200 463.600 ;
        RECT 667.600 462.200 668.400 464.200 ;
        RECT 672.000 463.600 674.000 464.200 ;
        RECT 672.000 462.200 672.800 463.600 ;
        RECT 676.400 462.200 677.200 467.000 ;
        RECT 678.000 466.800 680.200 467.400 ;
        RECT 678.000 462.200 678.800 466.800 ;
        RECT 1.200 455.400 2.000 459.800 ;
        RECT 5.400 458.400 6.600 459.800 ;
        RECT 5.400 457.800 6.800 458.400 ;
        RECT 10.000 457.800 10.800 459.800 ;
        RECT 14.400 458.400 15.200 459.800 ;
        RECT 14.400 457.800 16.400 458.400 ;
        RECT 6.000 457.000 6.800 457.800 ;
        RECT 10.200 457.200 10.800 457.800 ;
        RECT 10.200 456.600 13.000 457.200 ;
        RECT 12.200 456.400 13.000 456.600 ;
        RECT 14.000 456.400 14.800 457.200 ;
        RECT 15.600 457.000 16.400 457.800 ;
        RECT 4.200 455.400 5.000 455.600 ;
        RECT 1.200 454.800 5.000 455.400 ;
        RECT 1.200 451.400 2.000 454.800 ;
        RECT 8.200 454.200 9.000 454.400 ;
        RECT 14.000 454.200 14.600 456.400 ;
        RECT 18.800 455.000 19.600 459.800 ;
        RECT 20.400 456.000 21.200 459.800 ;
        RECT 23.600 456.000 24.400 459.800 ;
        RECT 20.400 455.800 24.400 456.000 ;
        RECT 25.200 455.800 26.000 459.800 ;
        RECT 26.800 455.800 27.600 459.800 ;
        RECT 28.400 456.000 29.200 459.800 ;
        RECT 31.600 456.000 32.400 459.800 ;
        RECT 28.400 455.800 32.400 456.000 ;
        RECT 33.200 456.000 34.000 459.800 ;
        RECT 36.400 456.000 37.200 459.800 ;
        RECT 33.200 455.800 37.200 456.000 ;
        RECT 38.000 455.800 38.800 459.800 ;
        RECT 40.200 456.400 41.000 459.800 ;
        RECT 40.200 455.800 42.000 456.400 ;
        RECT 44.400 456.000 45.200 459.800 ;
        RECT 47.600 456.000 48.400 459.800 ;
        RECT 44.400 455.800 48.400 456.000 ;
        RECT 49.200 455.800 50.000 459.800 ;
        RECT 50.800 455.800 51.600 459.800 ;
        RECT 52.400 456.000 53.200 459.800 ;
        RECT 55.600 456.000 56.400 459.800 ;
        RECT 61.000 456.000 61.800 459.000 ;
        RECT 65.200 457.000 66.000 459.000 ;
        RECT 52.400 455.800 56.400 456.000 ;
        RECT 20.600 455.400 24.200 455.800 ;
        RECT 21.200 454.400 22.000 454.800 ;
        RECT 25.200 454.400 25.800 455.800 ;
        RECT 27.000 454.400 27.600 455.800 ;
        RECT 28.600 455.400 32.200 455.800 ;
        RECT 33.400 455.400 37.000 455.800 ;
        RECT 30.800 454.400 31.600 454.800 ;
        RECT 34.000 454.400 34.800 454.800 ;
        RECT 38.000 454.400 38.600 455.800 ;
        RECT 17.200 454.200 18.800 454.400 ;
        RECT 7.800 453.600 18.800 454.200 ;
        RECT 20.400 453.800 22.000 454.400 ;
        RECT 20.400 453.600 21.200 453.800 ;
        RECT 23.400 453.600 26.000 454.400 ;
        RECT 26.800 453.600 29.400 454.400 ;
        RECT 30.800 454.300 32.400 454.400 ;
        RECT 33.200 454.300 34.800 454.400 ;
        RECT 30.800 453.800 34.800 454.300 ;
        RECT 31.600 453.700 34.000 453.800 ;
        RECT 31.600 453.600 32.400 453.700 ;
        RECT 33.200 453.600 34.000 453.700 ;
        RECT 36.200 453.600 38.800 454.400 ;
        RECT 6.000 452.800 6.800 453.000 ;
        RECT 3.000 452.200 6.800 452.800 ;
        RECT 3.000 452.000 3.800 452.200 ;
        RECT 4.600 451.400 5.400 451.600 ;
        RECT 1.200 450.800 5.400 451.400 ;
        RECT 1.200 442.200 2.000 450.800 ;
        RECT 7.800 450.400 8.400 453.600 ;
        RECT 15.000 453.400 15.800 453.600 ;
        RECT 14.000 452.400 14.800 452.600 ;
        RECT 16.600 452.400 17.400 452.600 ;
        RECT 12.400 451.800 17.400 452.400 ;
        RECT 12.400 451.600 13.200 451.800 ;
        RECT 22.000 451.600 22.800 453.200 ;
        RECT 14.000 451.000 19.600 451.200 ;
        RECT 13.800 450.800 19.600 451.000 ;
        RECT 6.000 449.800 8.400 450.400 ;
        RECT 9.800 450.600 19.600 450.800 ;
        RECT 9.800 450.200 14.600 450.600 ;
        RECT 6.000 448.800 6.600 449.800 ;
        RECT 5.200 448.000 6.600 448.800 ;
        RECT 8.200 449.000 9.000 449.200 ;
        RECT 9.800 449.000 10.400 450.200 ;
        RECT 8.200 448.400 10.400 449.000 ;
        RECT 11.000 449.000 16.400 449.600 ;
        RECT 11.000 448.800 11.800 449.000 ;
        RECT 15.600 448.800 16.400 449.000 ;
        RECT 9.400 447.400 10.200 447.600 ;
        RECT 12.200 447.400 13.000 447.600 ;
        RECT 6.000 446.200 6.800 447.000 ;
        RECT 9.400 446.800 13.000 447.400 ;
        RECT 10.200 446.200 10.800 446.800 ;
        RECT 15.600 446.200 16.400 447.000 ;
        RECT 5.400 442.200 6.600 446.200 ;
        RECT 10.000 442.200 10.800 446.200 ;
        RECT 14.400 445.600 16.400 446.200 ;
        RECT 14.400 442.200 15.200 445.600 ;
        RECT 18.800 442.200 19.600 450.600 ;
        RECT 23.400 450.400 24.000 453.600 ;
        RECT 28.800 452.300 29.400 453.600 ;
        RECT 25.300 451.700 29.400 452.300 ;
        RECT 25.300 450.400 25.900 451.700 ;
        RECT 22.000 449.600 24.000 450.400 ;
        RECT 25.200 450.200 26.000 450.400 ;
        RECT 24.600 449.600 26.000 450.200 ;
        RECT 26.800 450.200 27.600 450.400 ;
        RECT 28.800 450.200 29.400 451.700 ;
        RECT 30.000 451.600 30.800 453.200 ;
        RECT 34.800 451.600 35.600 453.200 ;
        RECT 36.200 450.200 36.800 453.600 ;
        RECT 41.200 452.300 42.000 455.800 ;
        RECT 44.600 455.400 48.200 455.800 ;
        RECT 42.800 454.300 43.600 455.200 ;
        RECT 45.200 454.400 46.000 454.800 ;
        RECT 49.200 454.400 49.800 455.800 ;
        RECT 51.000 454.400 51.600 455.800 ;
        RECT 52.600 455.400 56.200 455.800 ;
        RECT 60.200 455.400 61.800 456.000 ;
        RECT 60.200 455.000 61.000 455.400 ;
        RECT 54.800 454.400 55.600 454.800 ;
        RECT 60.200 454.400 60.800 455.000 ;
        RECT 65.400 454.800 66.000 457.000 ;
        RECT 66.800 455.800 67.600 459.800 ;
        RECT 68.400 456.000 69.200 459.800 ;
        RECT 71.600 456.000 72.400 459.800 ;
        RECT 68.400 455.800 72.400 456.000 ;
        RECT 73.200 455.800 74.000 459.800 ;
        RECT 74.800 456.000 75.600 459.800 ;
        RECT 78.000 456.000 78.800 459.800 ;
        RECT 74.800 455.800 78.800 456.000 ;
        RECT 44.400 454.300 46.000 454.400 ;
        RECT 42.800 453.800 46.000 454.300 ;
        RECT 42.800 453.700 45.200 453.800 ;
        RECT 42.800 453.600 43.600 453.700 ;
        RECT 44.400 453.600 45.200 453.700 ;
        RECT 47.400 453.600 50.000 454.400 ;
        RECT 50.800 453.600 53.400 454.400 ;
        RECT 54.800 453.800 56.400 454.400 ;
        RECT 58.800 454.300 60.800 454.400 ;
        RECT 55.600 453.600 56.400 453.800 ;
        RECT 57.300 453.700 60.800 454.300 ;
        RECT 61.800 454.200 66.000 454.800 ;
        RECT 67.000 454.400 67.600 455.800 ;
        RECT 68.600 455.400 72.200 455.800 ;
        RECT 70.800 454.400 71.600 454.800 ;
        RECT 73.400 454.400 74.000 455.800 ;
        RECT 75.000 455.400 78.600 455.800 ;
        RECT 79.600 455.000 80.400 459.800 ;
        RECT 84.000 458.400 84.800 459.800 ;
        RECT 82.800 457.800 84.800 458.400 ;
        RECT 88.400 457.800 89.200 459.800 ;
        RECT 92.600 458.400 93.800 459.800 ;
        RECT 92.400 457.800 93.800 458.400 ;
        RECT 82.800 457.000 83.600 457.800 ;
        RECT 88.400 457.200 89.000 457.800 ;
        RECT 84.400 455.600 85.200 457.200 ;
        RECT 86.200 456.600 89.000 457.200 ;
        RECT 92.400 457.000 93.200 457.800 ;
        RECT 86.200 456.400 87.000 456.600 ;
        RECT 77.200 454.400 78.000 454.800 ;
        RECT 61.800 453.800 62.800 454.200 ;
        RECT 38.100 451.700 42.000 452.300 ;
        RECT 38.100 450.400 38.700 451.700 ;
        RECT 38.000 450.200 38.800 450.400 ;
        RECT 26.800 449.600 28.200 450.200 ;
        RECT 28.800 449.600 29.800 450.200 ;
        RECT 23.000 442.200 23.800 449.600 ;
        RECT 24.600 448.400 25.200 449.600 ;
        RECT 24.400 447.600 25.200 448.400 ;
        RECT 27.600 448.400 28.200 449.600 ;
        RECT 27.600 447.600 28.400 448.400 ;
        RECT 29.000 442.200 29.800 449.600 ;
        RECT 35.800 449.600 36.800 450.200 ;
        RECT 37.400 449.600 38.800 450.200 ;
        RECT 35.800 442.200 36.600 449.600 ;
        RECT 37.400 448.400 38.000 449.600 ;
        RECT 39.600 448.800 40.400 450.400 ;
        RECT 37.200 447.600 38.000 448.400 ;
        RECT 41.200 442.200 42.000 451.700 ;
        RECT 44.400 452.300 45.200 452.400 ;
        RECT 46.000 452.300 46.800 453.200 ;
        RECT 44.400 451.700 46.800 452.300 ;
        RECT 44.400 451.600 45.200 451.700 ;
        RECT 46.000 451.600 46.800 451.700 ;
        RECT 47.400 452.300 48.000 453.600 ;
        RECT 47.400 451.700 51.500 452.300 ;
        RECT 47.400 450.200 48.000 451.700 ;
        RECT 50.900 450.400 51.500 451.700 ;
        RECT 49.200 450.200 50.000 450.400 ;
        RECT 47.000 449.600 48.000 450.200 ;
        RECT 48.600 449.600 50.000 450.200 ;
        RECT 50.800 450.200 51.600 450.400 ;
        RECT 52.800 450.200 53.400 453.600 ;
        RECT 54.000 452.300 54.800 453.200 ;
        RECT 57.300 452.300 57.900 453.700 ;
        RECT 58.800 453.600 60.800 453.700 ;
        RECT 54.000 451.700 57.900 452.300 ;
        RECT 54.000 451.600 54.800 451.700 ;
        RECT 58.800 450.800 59.600 452.400 ;
        RECT 50.800 449.600 52.200 450.200 ;
        RECT 52.800 449.600 53.800 450.200 ;
        RECT 47.000 442.200 47.800 449.600 ;
        RECT 48.600 448.400 49.200 449.600 ;
        RECT 48.400 447.600 49.200 448.400 ;
        RECT 51.600 448.400 52.200 449.600 ;
        RECT 51.600 447.600 52.400 448.400 ;
        RECT 53.000 442.200 53.800 449.600 ;
        RECT 60.200 449.800 60.800 453.600 ;
        RECT 61.400 453.000 62.800 453.800 ;
        RECT 66.800 453.600 69.400 454.400 ;
        RECT 70.800 453.800 72.400 454.400 ;
        RECT 71.600 453.600 72.400 453.800 ;
        RECT 73.200 453.600 75.800 454.400 ;
        RECT 77.200 453.800 78.800 454.400 ;
        RECT 78.000 453.600 78.800 453.800 ;
        RECT 80.400 454.200 82.000 454.400 ;
        RECT 84.600 454.200 85.200 455.600 ;
        RECT 94.200 455.400 95.000 455.600 ;
        RECT 97.200 455.400 98.000 459.800 ;
        RECT 98.800 456.000 99.600 459.800 ;
        RECT 102.000 456.000 102.800 459.800 ;
        RECT 98.800 455.800 102.800 456.000 ;
        RECT 103.600 455.800 104.400 459.800 ;
        RECT 105.200 455.800 106.000 459.800 ;
        RECT 106.800 456.000 107.600 459.800 ;
        RECT 110.000 456.000 110.800 459.800 ;
        RECT 106.800 455.800 110.800 456.000 ;
        RECT 99.000 455.400 102.600 455.800 ;
        RECT 94.200 454.800 98.000 455.400 ;
        RECT 90.200 454.200 91.000 454.400 ;
        RECT 80.400 453.600 91.400 454.200 ;
        RECT 62.200 451.000 62.800 453.000 ;
        RECT 63.600 451.600 64.400 453.200 ;
        RECT 65.200 451.600 66.000 453.200 ;
        RECT 62.200 450.400 66.000 451.000 ;
        RECT 68.800 450.400 69.400 453.600 ;
        RECT 70.000 451.600 70.800 453.200 ;
        RECT 73.200 452.300 74.000 452.400 ;
        RECT 75.200 452.300 75.800 453.600 ;
        RECT 83.400 453.400 84.200 453.600 ;
        RECT 73.200 451.700 75.800 452.300 ;
        RECT 73.200 451.600 74.000 451.700 ;
        RECT 60.200 449.200 61.800 449.800 ;
        RECT 61.000 442.200 61.800 449.200 ;
        RECT 65.400 447.000 66.000 450.400 ;
        RECT 66.800 450.200 67.600 450.400 ;
        RECT 66.800 449.600 68.200 450.200 ;
        RECT 68.800 449.600 70.800 450.400 ;
        RECT 73.200 450.200 74.000 450.400 ;
        RECT 75.200 450.200 75.800 451.700 ;
        RECT 76.400 451.600 77.200 453.200 ;
        RECT 81.800 452.400 82.600 452.600 ;
        RECT 84.400 452.400 85.200 452.600 ;
        RECT 81.800 451.800 86.800 452.400 ;
        RECT 86.000 451.600 86.800 451.800 ;
        RECT 79.600 451.000 85.200 451.200 ;
        RECT 79.600 450.800 85.400 451.000 ;
        RECT 79.600 450.600 89.400 450.800 ;
        RECT 73.200 449.600 74.600 450.200 ;
        RECT 75.200 449.600 76.200 450.200 ;
        RECT 67.600 448.400 68.200 449.600 ;
        RECT 67.600 447.600 68.400 448.400 ;
        RECT 65.200 443.000 66.000 447.000 ;
        RECT 69.000 442.200 69.800 449.600 ;
        RECT 74.000 448.400 74.600 449.600 ;
        RECT 74.000 447.600 74.800 448.400 ;
        RECT 75.400 442.200 76.200 449.600 ;
        RECT 79.600 442.200 80.400 450.600 ;
        RECT 84.600 450.200 89.400 450.600 ;
        RECT 82.800 449.000 88.200 449.600 ;
        RECT 82.800 448.800 83.600 449.000 ;
        RECT 87.400 448.800 88.200 449.000 ;
        RECT 88.800 449.000 89.400 450.200 ;
        RECT 90.800 450.400 91.400 453.600 ;
        RECT 92.400 452.800 93.200 453.000 ;
        RECT 92.400 452.200 96.200 452.800 ;
        RECT 95.400 452.000 96.200 452.200 ;
        RECT 93.800 451.400 94.600 451.600 ;
        RECT 97.200 451.400 98.000 454.800 ;
        RECT 99.600 454.400 100.400 454.800 ;
        RECT 103.600 454.400 104.200 455.800 ;
        RECT 105.400 454.400 106.000 455.800 ;
        RECT 107.000 455.400 110.600 455.800 ;
        RECT 116.400 455.400 117.200 459.800 ;
        RECT 120.600 458.400 121.800 459.800 ;
        RECT 120.600 457.800 122.000 458.400 ;
        RECT 125.200 457.800 126.000 459.800 ;
        RECT 129.600 458.400 130.400 459.800 ;
        RECT 129.600 457.800 131.600 458.400 ;
        RECT 121.200 457.000 122.000 457.800 ;
        RECT 125.400 457.200 126.000 457.800 ;
        RECT 125.400 456.600 128.200 457.200 ;
        RECT 127.400 456.400 128.200 456.600 ;
        RECT 129.200 456.400 130.000 457.200 ;
        RECT 130.800 457.000 131.600 457.800 ;
        RECT 119.400 455.400 120.200 455.600 ;
        RECT 116.400 454.800 120.200 455.400 ;
        RECT 109.200 454.400 110.000 454.800 ;
        RECT 98.800 453.800 100.400 454.400 ;
        RECT 98.800 453.600 99.600 453.800 ;
        RECT 101.800 453.600 104.400 454.400 ;
        RECT 105.200 453.600 107.800 454.400 ;
        RECT 109.200 453.800 110.800 454.400 ;
        RECT 110.000 453.600 110.800 453.800 ;
        RECT 100.400 451.600 101.200 453.200 ;
        RECT 101.800 452.300 102.400 453.600 ;
        RECT 107.200 452.400 107.800 453.600 ;
        RECT 101.800 451.700 105.900 452.300 ;
        RECT 93.800 450.800 98.000 451.400 ;
        RECT 90.800 449.800 93.200 450.400 ;
        RECT 90.200 449.000 91.000 449.200 ;
        RECT 88.800 448.400 91.000 449.000 ;
        RECT 92.600 448.800 93.200 449.800 ;
        RECT 92.600 448.000 94.000 448.800 ;
        RECT 86.200 447.400 87.000 447.600 ;
        RECT 89.000 447.400 89.800 447.600 ;
        RECT 82.800 446.200 83.600 447.000 ;
        RECT 86.200 446.800 89.800 447.400 ;
        RECT 88.400 446.200 89.000 446.800 ;
        RECT 92.400 446.200 93.200 447.000 ;
        RECT 82.800 445.600 84.800 446.200 ;
        RECT 84.000 442.200 84.800 445.600 ;
        RECT 88.400 442.200 89.200 446.200 ;
        RECT 92.600 442.200 93.800 446.200 ;
        RECT 97.200 442.200 98.000 450.800 ;
        RECT 101.800 450.200 102.400 451.700 ;
        RECT 105.300 450.400 105.900 451.700 ;
        RECT 106.800 451.600 107.800 452.400 ;
        RECT 108.400 451.600 109.200 453.200 ;
        RECT 103.600 450.200 104.400 450.400 ;
        RECT 101.400 449.600 102.400 450.200 ;
        RECT 103.000 449.600 104.400 450.200 ;
        RECT 105.200 450.200 106.000 450.400 ;
        RECT 107.200 450.200 107.800 451.600 ;
        RECT 116.400 451.400 117.200 454.800 ;
        RECT 123.400 454.200 124.200 454.400 ;
        RECT 126.000 454.200 126.800 454.400 ;
        RECT 129.200 454.200 129.800 456.400 ;
        RECT 134.000 455.000 134.800 459.800 ;
        RECT 132.400 454.200 134.000 454.400 ;
        RECT 123.000 453.600 134.000 454.200 ;
        RECT 121.200 452.800 122.000 453.000 ;
        RECT 118.200 452.200 122.000 452.800 ;
        RECT 118.200 452.000 119.000 452.200 ;
        RECT 119.800 451.400 120.600 451.600 ;
        RECT 116.400 450.800 120.600 451.400 ;
        RECT 105.200 449.600 106.600 450.200 ;
        RECT 107.200 449.600 108.200 450.200 ;
        RECT 101.400 442.200 102.200 449.600 ;
        RECT 103.000 448.400 103.600 449.600 ;
        RECT 102.800 447.600 103.600 448.400 ;
        RECT 106.000 448.400 106.600 449.600 ;
        RECT 106.000 447.600 106.800 448.400 ;
        RECT 107.400 442.200 108.200 449.600 ;
        RECT 116.400 442.200 117.200 450.800 ;
        RECT 123.000 450.400 123.600 453.600 ;
        RECT 130.200 453.400 131.000 453.600 ;
        RECT 131.800 452.400 132.600 452.600 ;
        RECT 127.600 451.800 132.600 452.400 ;
        RECT 127.600 451.600 128.400 451.800 ;
        RECT 129.200 451.000 134.800 451.200 ;
        RECT 129.000 450.800 134.800 451.000 ;
        RECT 121.200 449.800 123.600 450.400 ;
        RECT 125.000 450.600 134.800 450.800 ;
        RECT 125.000 450.200 129.800 450.600 ;
        RECT 121.200 448.800 121.800 449.800 ;
        RECT 120.400 448.000 121.800 448.800 ;
        RECT 123.400 449.000 124.200 449.200 ;
        RECT 125.000 449.000 125.600 450.200 ;
        RECT 123.400 448.400 125.600 449.000 ;
        RECT 126.200 449.000 131.600 449.600 ;
        RECT 126.200 448.800 127.000 449.000 ;
        RECT 130.800 448.800 131.600 449.000 ;
        RECT 124.600 447.400 125.400 447.600 ;
        RECT 127.400 447.400 128.200 447.600 ;
        RECT 121.200 446.200 122.000 447.000 ;
        RECT 124.600 446.800 128.200 447.400 ;
        RECT 125.400 446.200 126.000 446.800 ;
        RECT 130.800 446.200 131.600 447.000 ;
        RECT 120.600 442.200 121.800 446.200 ;
        RECT 125.200 442.200 126.000 446.200 ;
        RECT 129.600 445.600 131.600 446.200 ;
        RECT 129.600 442.200 130.400 445.600 ;
        RECT 134.000 442.200 134.800 450.600 ;
        RECT 135.600 442.200 136.400 459.800 ;
        RECT 137.200 455.600 138.000 457.200 ;
        RECT 138.800 457.000 139.600 459.000 ;
        RECT 138.800 454.800 139.400 457.000 ;
        RECT 143.000 456.000 143.800 459.000 ;
        RECT 148.400 456.000 149.200 459.800 ;
        RECT 151.600 456.000 152.400 459.800 ;
        RECT 143.000 455.400 144.600 456.000 ;
        RECT 148.400 455.800 152.400 456.000 ;
        RECT 153.200 455.800 154.000 459.800 ;
        RECT 154.800 457.000 155.600 459.000 ;
        RECT 148.600 455.400 152.200 455.800 ;
        RECT 143.800 455.000 144.600 455.400 ;
        RECT 138.800 454.200 143.000 454.800 ;
        RECT 142.000 453.800 143.000 454.200 ;
        RECT 144.000 454.400 144.600 455.000 ;
        RECT 149.200 454.400 150.000 454.800 ;
        RECT 153.200 454.400 153.800 455.800 ;
        RECT 154.800 454.800 155.400 457.000 ;
        RECT 159.000 456.000 159.800 459.000 ;
        RECT 166.000 457.800 166.800 459.800 ;
        RECT 159.000 455.400 160.600 456.000 ;
        RECT 164.400 455.600 165.200 457.200 ;
        RECT 159.800 455.000 160.600 455.400 ;
        RECT 138.800 451.600 139.600 453.200 ;
        RECT 140.400 451.600 141.200 453.200 ;
        RECT 142.000 453.000 143.400 453.800 ;
        RECT 144.000 453.600 146.000 454.400 ;
        RECT 148.400 453.800 150.000 454.400 ;
        RECT 148.400 453.600 149.200 453.800 ;
        RECT 151.400 453.600 154.000 454.400 ;
        RECT 154.800 454.200 159.000 454.800 ;
        RECT 158.000 453.800 159.000 454.200 ;
        RECT 160.000 454.400 160.600 455.000 ;
        RECT 166.200 454.400 166.800 457.800 ;
        RECT 169.200 456.000 170.000 459.800 ;
        RECT 172.400 456.000 173.200 459.800 ;
        RECT 169.200 455.800 173.200 456.000 ;
        RECT 174.000 455.800 174.800 459.800 ;
        RECT 169.400 455.400 173.000 455.800 ;
        RECT 170.000 454.400 170.800 454.800 ;
        RECT 174.000 454.400 174.600 455.800 ;
        RECT 175.600 455.000 176.400 459.800 ;
        RECT 180.000 458.400 180.800 459.800 ;
        RECT 178.800 457.800 180.800 458.400 ;
        RECT 184.400 457.800 185.200 459.800 ;
        RECT 188.600 458.400 189.800 459.800 ;
        RECT 188.400 457.800 189.800 458.400 ;
        RECT 178.800 457.000 179.600 457.800 ;
        RECT 184.400 457.200 185.000 457.800 ;
        RECT 180.400 456.400 181.200 457.200 ;
        RECT 182.200 456.600 185.000 457.200 ;
        RECT 188.400 457.000 189.200 457.800 ;
        RECT 182.200 456.400 183.000 456.600 ;
        RECT 160.000 454.300 162.000 454.400 ;
        RECT 164.400 454.300 165.200 454.400 ;
        RECT 142.000 451.000 142.600 453.000 ;
        RECT 138.800 450.400 142.600 451.000 ;
        RECT 138.800 447.000 139.400 450.400 ;
        RECT 144.000 449.800 144.600 453.600 ;
        RECT 145.200 452.300 146.000 452.400 ;
        RECT 146.800 452.300 147.600 452.400 ;
        RECT 145.200 451.700 147.600 452.300 ;
        RECT 145.200 450.800 146.000 451.700 ;
        RECT 146.800 451.600 147.600 451.700 ;
        RECT 150.000 451.600 150.800 453.200 ;
        RECT 151.400 450.200 152.000 453.600 ;
        RECT 154.800 451.600 155.600 453.200 ;
        RECT 156.400 451.600 157.200 453.200 ;
        RECT 158.000 453.000 159.400 453.800 ;
        RECT 160.000 453.700 165.200 454.300 ;
        RECT 160.000 453.600 162.000 453.700 ;
        RECT 164.400 453.600 165.200 453.700 ;
        RECT 166.000 453.600 166.800 454.400 ;
        RECT 169.200 453.800 170.800 454.400 ;
        RECT 169.200 453.600 170.000 453.800 ;
        RECT 172.200 453.600 174.800 454.400 ;
        RECT 176.400 454.200 178.000 454.400 ;
        RECT 180.600 454.200 181.200 456.400 ;
        RECT 190.200 455.400 191.000 455.600 ;
        RECT 193.200 455.400 194.000 459.800 ;
        RECT 196.400 457.800 197.200 459.800 ;
        RECT 194.800 455.600 195.600 457.200 ;
        RECT 190.200 454.800 194.000 455.400 ;
        RECT 182.000 454.200 182.800 454.400 ;
        RECT 186.200 454.200 187.000 454.400 ;
        RECT 176.400 453.600 187.400 454.200 ;
        RECT 158.000 451.000 158.600 453.000 ;
        RECT 154.800 450.400 158.600 451.000 ;
        RECT 153.200 450.200 154.000 450.400 ;
        RECT 143.000 449.200 144.600 449.800 ;
        RECT 151.000 449.600 152.000 450.200 ;
        RECT 152.600 449.600 154.000 450.200 ;
        RECT 138.800 443.000 139.600 447.000 ;
        RECT 143.000 442.200 143.800 449.200 ;
        RECT 151.000 442.200 151.800 449.600 ;
        RECT 152.600 448.400 153.200 449.600 ;
        RECT 152.400 447.600 153.200 448.400 ;
        RECT 154.800 447.000 155.400 450.400 ;
        RECT 160.000 449.800 160.600 453.600 ;
        RECT 161.200 450.800 162.000 452.400 ;
        RECT 162.800 452.300 163.600 452.400 ;
        RECT 166.200 452.300 166.800 453.600 ;
        RECT 162.800 451.700 166.800 452.300 ;
        RECT 162.800 451.600 163.600 451.700 ;
        RECT 166.200 450.200 166.800 451.700 ;
        RECT 167.600 450.800 168.400 452.400 ;
        RECT 170.800 451.600 171.600 453.200 ;
        RECT 172.200 452.300 172.800 453.600 ;
        RECT 179.400 453.400 180.200 453.600 ;
        RECT 177.800 452.400 178.600 452.600 ;
        RECT 180.400 452.400 181.200 452.600 ;
        RECT 174.000 452.300 174.800 452.400 ;
        RECT 172.200 451.700 174.800 452.300 ;
        RECT 177.800 451.800 182.800 452.400 ;
        RECT 172.200 450.200 172.800 451.700 ;
        RECT 174.000 451.600 174.800 451.700 ;
        RECT 182.000 451.600 182.800 451.800 ;
        RECT 175.600 451.000 181.200 451.200 ;
        RECT 175.600 450.800 181.400 451.000 ;
        RECT 175.600 450.600 185.400 450.800 ;
        RECT 174.000 450.200 174.800 450.400 ;
        RECT 159.000 449.200 160.600 449.800 ;
        RECT 166.000 449.400 167.800 450.200 ;
        RECT 154.800 443.000 155.600 447.000 ;
        RECT 159.000 442.200 159.800 449.200 ;
        RECT 167.000 442.200 167.800 449.400 ;
        RECT 171.800 449.600 172.800 450.200 ;
        RECT 173.400 449.600 174.800 450.200 ;
        RECT 171.800 442.200 172.600 449.600 ;
        RECT 173.400 448.400 174.000 449.600 ;
        RECT 173.200 447.600 174.000 448.400 ;
        RECT 175.600 442.200 176.400 450.600 ;
        RECT 180.600 450.200 185.400 450.600 ;
        RECT 178.800 449.000 184.200 449.600 ;
        RECT 178.800 448.800 179.600 449.000 ;
        RECT 183.400 448.800 184.200 449.000 ;
        RECT 184.800 449.000 185.400 450.200 ;
        RECT 186.800 450.400 187.400 453.600 ;
        RECT 188.400 452.800 189.200 453.000 ;
        RECT 188.400 452.200 192.200 452.800 ;
        RECT 191.400 452.000 192.200 452.200 ;
        RECT 189.800 451.400 190.600 451.600 ;
        RECT 193.200 451.400 194.000 454.800 ;
        RECT 196.600 454.400 197.200 457.800 ;
        RECT 199.600 455.800 200.400 459.800 ;
        RECT 204.000 458.400 205.600 459.800 ;
        RECT 204.000 457.600 206.800 458.400 ;
        RECT 204.000 456.200 205.600 457.600 ;
        RECT 199.600 455.200 202.000 455.800 ;
        RECT 201.200 455.000 202.000 455.200 ;
        RECT 202.600 454.800 203.400 455.600 ;
        RECT 202.600 454.400 203.200 454.800 ;
        RECT 196.400 453.600 197.200 454.400 ;
        RECT 199.600 453.600 201.200 454.400 ;
        RECT 202.400 453.600 203.200 454.400 ;
        RECT 196.600 452.400 197.200 453.600 ;
        RECT 204.000 452.800 204.600 456.200 ;
        RECT 209.200 455.800 210.000 459.800 ;
        RECT 205.200 455.400 206.800 455.600 ;
        RECT 205.200 454.800 207.200 455.400 ;
        RECT 207.800 455.200 210.000 455.800 ;
        RECT 207.800 455.000 208.600 455.200 ;
        RECT 206.600 454.400 207.200 454.800 ;
        RECT 205.200 453.400 206.000 454.200 ;
        RECT 206.600 453.800 210.000 454.400 ;
        RECT 212.000 454.200 212.800 459.800 ;
        RECT 217.200 456.000 218.000 459.800 ;
        RECT 220.400 456.000 221.200 459.800 ;
        RECT 217.200 455.800 221.200 456.000 ;
        RECT 222.000 456.300 222.800 459.800 ;
        RECT 223.600 456.300 224.400 457.200 ;
        RECT 217.400 455.400 221.000 455.800 ;
        RECT 222.000 455.700 224.400 456.300 ;
        RECT 218.000 454.400 218.800 454.800 ;
        RECT 222.000 454.400 222.600 455.700 ;
        RECT 223.600 455.600 224.400 455.700 ;
        RECT 208.400 453.600 210.000 453.800 ;
        RECT 211.000 453.800 212.800 454.200 ;
        RECT 217.200 453.800 218.800 454.400 ;
        RECT 211.000 453.600 212.600 453.800 ;
        RECT 217.200 453.600 218.000 453.800 ;
        RECT 220.200 453.600 222.800 454.400 ;
        RECT 203.600 452.400 204.600 452.800 ;
        RECT 196.400 451.600 197.200 452.400 ;
        RECT 189.800 450.800 194.000 451.400 ;
        RECT 186.800 449.800 189.200 450.400 ;
        RECT 186.200 449.000 187.000 449.200 ;
        RECT 184.800 448.400 187.000 449.000 ;
        RECT 188.600 448.800 189.200 449.800 ;
        RECT 188.600 448.400 190.000 448.800 ;
        RECT 188.600 448.000 190.800 448.400 ;
        RECT 189.400 447.600 190.800 448.000 ;
        RECT 182.200 447.400 183.000 447.600 ;
        RECT 185.000 447.400 185.800 447.600 ;
        RECT 178.800 446.200 179.600 447.000 ;
        RECT 182.200 446.800 185.800 447.400 ;
        RECT 184.400 446.200 185.000 446.800 ;
        RECT 188.400 446.200 189.200 447.000 ;
        RECT 178.800 445.600 180.800 446.200 ;
        RECT 180.000 442.200 180.800 445.600 ;
        RECT 184.400 442.200 185.200 446.200 ;
        RECT 188.600 442.200 189.800 446.200 ;
        RECT 193.200 442.200 194.000 450.800 ;
        RECT 196.600 450.200 197.200 451.600 ;
        RECT 198.000 450.800 198.800 452.400 ;
        RECT 202.800 452.200 204.600 452.400 ;
        RECT 205.400 452.800 206.000 453.400 ;
        RECT 205.400 452.200 208.000 452.800 ;
        RECT 202.800 451.600 204.200 452.200 ;
        RECT 207.200 452.000 208.000 452.200 ;
        RECT 203.600 450.200 204.200 451.600 ;
        RECT 205.000 451.400 205.800 451.600 ;
        RECT 205.000 450.800 208.400 451.400 ;
        RECT 207.800 450.200 208.400 450.800 ;
        RECT 211.000 450.400 211.600 453.600 ;
        RECT 213.200 451.600 214.800 452.400 ;
        RECT 217.300 452.300 217.900 453.600 ;
        RECT 215.600 451.700 217.900 452.300 ;
        RECT 196.400 449.400 198.200 450.200 ;
        RECT 197.400 442.200 198.200 449.400 ;
        RECT 199.600 449.600 202.000 450.200 ;
        RECT 203.600 449.600 205.600 450.200 ;
        RECT 199.600 442.200 200.400 449.600 ;
        RECT 201.200 449.400 202.000 449.600 ;
        RECT 204.000 442.200 205.600 449.600 ;
        RECT 207.800 449.600 210.000 450.200 ;
        RECT 210.800 449.600 211.600 450.400 ;
        RECT 215.600 449.600 216.400 451.700 ;
        RECT 218.800 451.600 219.600 453.200 ;
        RECT 220.200 450.200 220.800 453.600 ;
        RECT 222.000 450.200 222.800 450.400 ;
        RECT 219.800 449.600 220.800 450.200 ;
        RECT 221.400 449.600 222.800 450.200 ;
        RECT 207.800 449.400 208.600 449.600 ;
        RECT 209.200 442.200 210.000 449.600 ;
        RECT 211.000 447.000 211.600 449.600 ;
        RECT 212.400 448.300 213.200 449.200 ;
        RECT 214.000 448.300 214.800 448.400 ;
        RECT 212.400 447.700 214.800 448.300 ;
        RECT 212.400 447.600 213.200 447.700 ;
        RECT 214.000 447.600 214.800 447.700 ;
        RECT 211.000 446.400 214.600 447.000 ;
        RECT 211.000 446.200 211.600 446.400 ;
        RECT 210.800 442.200 211.600 446.200 ;
        RECT 214.000 446.200 214.600 446.400 ;
        RECT 214.000 442.200 214.800 446.200 ;
        RECT 219.800 442.200 220.600 449.600 ;
        RECT 221.400 448.400 222.000 449.600 ;
        RECT 221.200 447.600 222.000 448.400 ;
        RECT 225.200 442.200 226.000 459.800 ;
        RECT 228.400 456.000 229.200 459.800 ;
        RECT 228.200 455.200 229.200 456.000 ;
        RECT 228.200 450.800 229.000 455.200 ;
        RECT 230.000 454.600 230.800 459.800 ;
        RECT 236.400 456.600 237.200 459.800 ;
        RECT 238.000 457.000 238.800 459.800 ;
        RECT 239.600 457.000 240.400 459.800 ;
        RECT 241.200 457.000 242.000 459.800 ;
        RECT 242.800 457.000 243.600 459.800 ;
        RECT 246.000 457.000 246.800 459.800 ;
        RECT 249.200 457.000 250.000 459.800 ;
        RECT 250.800 457.000 251.600 459.800 ;
        RECT 252.400 457.000 253.200 459.800 ;
        RECT 234.800 455.800 237.200 456.600 ;
        RECT 254.000 456.600 254.800 459.800 ;
        RECT 234.800 455.200 235.600 455.800 ;
        RECT 229.600 454.000 230.800 454.600 ;
        RECT 233.800 454.600 235.600 455.200 ;
        RECT 239.600 455.600 240.600 456.400 ;
        RECT 243.600 455.600 245.200 456.400 ;
        RECT 246.000 455.800 250.600 456.400 ;
        RECT 254.000 455.800 256.600 456.600 ;
        RECT 246.000 455.600 246.800 455.800 ;
        RECT 229.600 452.000 230.200 454.000 ;
        RECT 233.800 453.400 234.600 454.600 ;
        RECT 230.800 452.600 234.600 453.400 ;
        RECT 239.600 452.800 240.400 455.600 ;
        RECT 246.000 454.800 246.800 455.000 ;
        RECT 242.400 454.200 246.800 454.800 ;
        RECT 242.400 454.000 243.200 454.200 ;
        RECT 247.600 453.600 248.400 455.200 ;
        RECT 249.800 453.400 250.600 455.800 ;
        RECT 255.800 455.200 256.600 455.800 ;
        RECT 255.800 454.400 258.800 455.200 ;
        RECT 260.400 453.800 261.200 459.800 ;
        RECT 242.800 452.600 246.000 453.400 ;
        RECT 249.800 452.600 251.800 453.400 ;
        RECT 252.400 453.000 261.200 453.800 ;
        RECT 236.400 452.000 237.200 452.600 ;
        RECT 254.000 452.000 254.800 452.400 ;
        RECT 257.200 452.000 258.000 452.400 ;
        RECT 259.000 452.000 259.800 452.200 ;
        RECT 229.600 451.400 230.400 452.000 ;
        RECT 236.400 451.400 259.800 452.000 ;
        RECT 228.200 450.000 229.200 450.800 ;
        RECT 226.800 448.300 227.600 448.400 ;
        RECT 228.400 448.300 229.200 450.000 ;
        RECT 226.800 447.700 229.200 448.300 ;
        RECT 226.800 447.600 227.600 447.700 ;
        RECT 228.400 442.200 229.200 447.700 ;
        RECT 229.800 449.600 230.400 451.400 ;
        RECT 229.800 449.000 238.800 449.600 ;
        RECT 229.800 447.400 230.400 449.000 ;
        RECT 238.000 448.800 238.800 449.000 ;
        RECT 241.200 449.000 249.800 449.600 ;
        RECT 241.200 448.800 242.000 449.000 ;
        RECT 233.000 447.600 235.600 448.400 ;
        RECT 229.800 446.800 232.400 447.400 ;
        RECT 231.600 442.200 232.400 446.800 ;
        RECT 234.800 442.200 235.600 447.600 ;
        RECT 236.200 446.800 240.400 447.600 ;
        RECT 238.000 442.200 238.800 445.000 ;
        RECT 239.600 442.200 240.400 445.000 ;
        RECT 241.200 442.200 242.000 445.000 ;
        RECT 242.800 442.200 243.600 448.400 ;
        RECT 246.000 447.600 248.600 448.400 ;
        RECT 249.200 448.200 249.800 449.000 ;
        RECT 250.800 449.400 251.600 449.600 ;
        RECT 250.800 449.000 256.200 449.400 ;
        RECT 250.800 448.800 257.000 449.000 ;
        RECT 255.600 448.200 257.000 448.800 ;
        RECT 249.200 447.600 255.000 448.200 ;
        RECT 258.000 448.000 259.600 448.800 ;
        RECT 258.000 447.600 258.600 448.000 ;
        RECT 246.000 442.200 246.800 447.000 ;
        RECT 249.200 442.200 250.000 447.000 ;
        RECT 254.400 446.800 258.600 447.600 ;
        RECT 260.400 447.400 261.200 453.000 ;
        RECT 259.200 446.800 261.200 447.400 ;
        RECT 266.800 453.800 267.600 459.800 ;
        RECT 273.200 456.600 274.000 459.800 ;
        RECT 274.800 457.000 275.600 459.800 ;
        RECT 276.400 457.000 277.200 459.800 ;
        RECT 278.000 457.000 278.800 459.800 ;
        RECT 281.200 457.000 282.000 459.800 ;
        RECT 284.400 457.000 285.200 459.800 ;
        RECT 286.000 457.000 286.800 459.800 ;
        RECT 287.600 457.000 288.400 459.800 ;
        RECT 289.200 457.000 290.000 459.800 ;
        RECT 271.400 455.800 274.000 456.600 ;
        RECT 290.800 456.600 291.600 459.800 ;
        RECT 277.400 455.800 282.000 456.400 ;
        RECT 271.400 455.200 272.200 455.800 ;
        RECT 269.200 454.400 272.200 455.200 ;
        RECT 266.800 453.000 275.600 453.800 ;
        RECT 277.400 453.400 278.200 455.800 ;
        RECT 281.200 455.600 282.000 455.800 ;
        RECT 282.800 455.600 284.400 456.400 ;
        RECT 287.400 455.600 288.400 456.400 ;
        RECT 290.800 455.800 293.200 456.600 ;
        RECT 279.600 453.600 280.400 455.200 ;
        RECT 281.200 454.800 282.000 455.000 ;
        RECT 281.200 454.200 285.600 454.800 ;
        RECT 284.800 454.000 285.600 454.200 ;
        RECT 266.800 447.400 267.600 453.000 ;
        RECT 276.200 452.600 278.200 453.400 ;
        RECT 282.000 452.600 285.200 453.400 ;
        RECT 287.600 452.800 288.400 455.600 ;
        RECT 292.400 455.200 293.200 455.800 ;
        RECT 292.400 454.600 294.200 455.200 ;
        RECT 293.400 453.400 294.200 454.600 ;
        RECT 297.200 454.600 298.000 459.800 ;
        RECT 298.800 456.300 299.600 459.800 ;
        RECT 300.400 456.300 301.200 456.400 ;
        RECT 298.800 455.700 301.200 456.300 ;
        RECT 302.000 455.800 302.800 459.800 ;
        RECT 303.600 456.000 304.400 459.800 ;
        RECT 306.800 456.000 307.600 459.800 ;
        RECT 308.600 456.400 309.400 457.200 ;
        RECT 303.600 455.800 307.600 456.000 ;
        RECT 298.800 455.200 299.800 455.700 ;
        RECT 300.400 455.600 301.200 455.700 ;
        RECT 297.200 454.000 298.400 454.600 ;
        RECT 293.400 452.600 297.200 453.400 ;
        RECT 268.200 452.000 269.000 452.200 ;
        RECT 273.200 452.000 274.000 452.400 ;
        RECT 290.800 452.000 291.600 452.600 ;
        RECT 297.800 452.000 298.400 454.000 ;
        RECT 268.200 451.400 291.600 452.000 ;
        RECT 297.600 451.400 298.400 452.000 ;
        RECT 297.600 449.600 298.200 451.400 ;
        RECT 299.000 450.800 299.800 455.200 ;
        RECT 302.200 454.400 302.800 455.800 ;
        RECT 303.800 455.400 307.400 455.800 ;
        RECT 308.400 455.600 309.200 456.400 ;
        RECT 310.000 455.800 310.800 459.800 ;
        RECT 306.000 454.400 306.800 454.800 ;
        RECT 300.400 454.300 301.200 454.400 ;
        RECT 302.000 454.300 304.600 454.400 ;
        RECT 300.400 453.700 304.600 454.300 ;
        RECT 306.000 454.300 307.600 454.400 ;
        RECT 308.400 454.300 309.200 454.400 ;
        RECT 306.000 453.800 309.200 454.300 ;
        RECT 300.400 453.600 301.200 453.700 ;
        RECT 302.000 453.600 304.600 453.700 ;
        RECT 306.800 453.700 309.200 453.800 ;
        RECT 306.800 453.600 307.600 453.700 ;
        RECT 308.400 453.600 309.200 453.700 ;
        RECT 276.400 449.400 277.200 449.600 ;
        RECT 271.800 449.000 277.200 449.400 ;
        RECT 271.000 448.800 277.200 449.000 ;
        RECT 278.200 449.000 286.800 449.600 ;
        RECT 268.400 448.000 270.000 448.800 ;
        RECT 271.000 448.200 272.400 448.800 ;
        RECT 278.200 448.200 278.800 449.000 ;
        RECT 286.000 448.800 286.800 449.000 ;
        RECT 289.200 449.000 298.200 449.600 ;
        RECT 289.200 448.800 290.000 449.000 ;
        RECT 269.400 447.600 270.000 448.000 ;
        RECT 273.000 447.600 278.800 448.200 ;
        RECT 279.400 447.600 282.000 448.400 ;
        RECT 266.800 446.800 268.800 447.400 ;
        RECT 269.400 446.800 273.600 447.600 ;
        RECT 250.800 442.200 251.600 445.000 ;
        RECT 252.400 442.200 253.200 445.000 ;
        RECT 255.600 442.200 256.400 446.800 ;
        RECT 259.200 446.200 259.800 446.800 ;
        RECT 258.800 445.600 259.800 446.200 ;
        RECT 268.200 446.200 268.800 446.800 ;
        RECT 268.200 445.600 269.200 446.200 ;
        RECT 258.800 442.200 259.600 445.600 ;
        RECT 268.400 442.200 269.200 445.600 ;
        RECT 271.600 442.200 272.400 446.800 ;
        RECT 274.800 442.200 275.600 445.000 ;
        RECT 276.400 442.200 277.200 445.000 ;
        RECT 278.000 442.200 278.800 447.000 ;
        RECT 281.200 442.200 282.000 447.000 ;
        RECT 284.400 442.200 285.200 448.400 ;
        RECT 292.400 447.600 295.000 448.400 ;
        RECT 287.600 446.800 291.800 447.600 ;
        RECT 286.000 442.200 286.800 445.000 ;
        RECT 287.600 442.200 288.400 445.000 ;
        RECT 289.200 442.200 290.000 445.000 ;
        RECT 292.400 442.200 293.200 447.600 ;
        RECT 297.600 447.400 298.200 449.000 ;
        RECT 295.600 446.800 298.200 447.400 ;
        RECT 298.800 450.000 299.800 450.800 ;
        RECT 300.400 450.300 301.200 450.400 ;
        RECT 302.000 450.300 302.800 450.400 ;
        RECT 300.400 450.200 302.800 450.300 ;
        RECT 304.000 450.200 304.600 453.600 ;
        RECT 305.200 452.300 306.000 453.200 ;
        RECT 308.400 452.300 309.200 452.400 ;
        RECT 305.200 452.200 309.200 452.300 ;
        RECT 310.200 452.200 310.800 455.800 ;
        RECT 316.400 457.600 317.200 459.800 ;
        RECT 316.400 454.400 317.000 457.600 ;
        RECT 318.000 455.600 318.800 457.200 ;
        RECT 320.800 454.400 321.600 459.800 ;
        RECT 326.000 455.800 326.800 459.800 ;
        RECT 327.600 456.000 328.400 459.800 ;
        RECT 330.800 456.000 331.600 459.800 ;
        RECT 327.600 455.800 331.600 456.000 ;
        RECT 332.400 455.800 333.200 459.800 ;
        RECT 334.000 456.000 334.800 459.800 ;
        RECT 337.200 456.000 338.000 459.800 ;
        RECT 340.400 457.600 341.200 459.800 ;
        RECT 334.000 455.800 338.000 456.000 ;
        RECT 326.200 454.400 326.800 455.800 ;
        RECT 327.800 455.400 331.400 455.800 ;
        RECT 330.000 454.400 330.800 454.800 ;
        RECT 332.600 454.400 333.200 455.800 ;
        RECT 334.200 455.400 337.800 455.800 ;
        RECT 338.800 455.600 339.600 457.200 ;
        RECT 336.400 454.400 337.200 454.800 ;
        RECT 340.600 454.400 341.200 457.600 ;
        RECT 343.600 456.000 344.400 459.800 ;
        RECT 346.800 459.200 350.800 459.800 ;
        RECT 346.800 456.000 347.600 459.200 ;
        RECT 343.600 455.800 347.600 456.000 ;
        RECT 348.400 455.800 349.200 458.600 ;
        RECT 350.000 455.800 350.800 459.200 ;
        RECT 351.600 456.000 352.400 459.800 ;
        RECT 354.800 459.200 358.800 459.800 ;
        RECT 354.800 456.000 355.600 459.200 ;
        RECT 351.600 455.800 355.600 456.000 ;
        RECT 343.800 455.400 347.400 455.800 ;
        RECT 344.400 454.400 345.200 454.800 ;
        RECT 348.600 454.400 349.200 455.800 ;
        RECT 351.800 455.400 355.400 455.800 ;
        RECT 356.400 455.600 357.200 458.600 ;
        RECT 358.000 455.800 358.800 459.200 ;
        RECT 352.400 454.400 353.200 454.800 ;
        RECT 356.600 454.400 357.200 455.600 ;
        RECT 311.600 452.800 312.400 454.400 ;
        RECT 314.800 454.300 315.600 454.400 ;
        RECT 313.300 453.700 315.600 454.300 ;
        RECT 313.300 452.400 313.900 453.700 ;
        RECT 314.800 453.600 315.600 453.700 ;
        RECT 316.400 453.600 317.200 454.400 ;
        RECT 319.600 453.800 321.600 454.400 ;
        RECT 319.600 453.600 321.400 453.800 ;
        RECT 326.000 453.600 328.600 454.400 ;
        RECT 330.000 453.800 331.600 454.400 ;
        RECT 330.800 453.600 331.600 453.800 ;
        RECT 332.400 453.600 335.000 454.400 ;
        RECT 336.400 454.300 338.000 454.400 ;
        RECT 338.800 454.300 339.600 454.400 ;
        RECT 336.400 453.800 339.600 454.300 ;
        RECT 337.200 453.700 339.600 453.800 ;
        RECT 337.200 453.600 338.000 453.700 ;
        RECT 338.800 453.600 339.600 453.700 ;
        RECT 340.400 453.600 341.200 454.400 ;
        RECT 343.600 453.800 345.200 454.400 ;
        RECT 346.800 453.800 349.200 454.400 ;
        RECT 350.000 454.300 350.800 454.400 ;
        RECT 351.600 454.300 353.200 454.400 ;
        RECT 350.000 453.800 353.200 454.300 ;
        RECT 354.800 453.800 357.200 454.400 ;
        RECT 358.000 454.300 358.800 454.400 ;
        RECT 359.600 454.300 360.400 459.800 ;
        RECT 361.200 455.600 362.000 457.200 ;
        RECT 343.600 453.600 344.400 453.800 ;
        RECT 346.800 453.600 347.600 453.800 ;
        RECT 350.000 453.700 352.400 453.800 ;
        RECT 313.200 452.200 314.000 452.400 ;
        RECT 305.200 451.700 310.800 452.200 ;
        RECT 305.200 451.600 306.000 451.700 ;
        RECT 308.400 451.600 310.800 451.700 ;
        RECT 312.400 451.600 314.000 452.200 ;
        RECT 308.600 450.200 309.200 451.600 ;
        RECT 312.400 451.200 313.200 451.600 ;
        RECT 314.800 450.800 315.600 452.400 ;
        RECT 316.400 450.200 317.000 453.600 ;
        RECT 319.800 450.400 320.400 453.600 ;
        RECT 328.000 452.400 328.600 453.600 ;
        RECT 322.000 451.600 323.600 452.400 ;
        RECT 327.600 451.600 328.600 452.400 ;
        RECT 329.200 451.600 330.000 453.200 ;
        RECT 295.600 442.200 296.400 446.800 ;
        RECT 298.800 442.200 299.600 450.000 ;
        RECT 300.400 449.700 303.400 450.200 ;
        RECT 300.400 449.600 301.200 449.700 ;
        RECT 302.000 449.600 303.400 449.700 ;
        RECT 304.000 449.600 305.000 450.200 ;
        RECT 302.800 448.400 303.400 449.600 ;
        RECT 302.800 447.600 303.600 448.400 ;
        RECT 304.200 442.200 305.000 449.600 ;
        RECT 308.400 442.200 309.200 450.200 ;
        RECT 310.000 449.600 314.000 450.200 ;
        RECT 310.000 442.200 310.800 449.600 ;
        RECT 313.200 442.200 314.000 449.600 ;
        RECT 315.400 449.400 317.200 450.200 ;
        RECT 319.600 449.600 320.400 450.400 ;
        RECT 322.800 450.300 323.600 450.400 ;
        RECT 324.400 450.300 325.200 451.200 ;
        RECT 322.800 449.700 325.200 450.300 ;
        RECT 322.800 449.600 323.600 449.700 ;
        RECT 324.400 449.600 325.200 449.700 ;
        RECT 326.000 450.200 326.800 450.400 ;
        RECT 328.000 450.200 328.600 451.600 ;
        RECT 332.400 450.200 333.200 450.400 ;
        RECT 334.400 450.200 335.000 453.600 ;
        RECT 335.600 451.600 336.400 453.200 ;
        RECT 340.600 450.200 341.200 453.600 ;
        RECT 342.000 450.800 342.800 452.400 ;
        RECT 345.200 451.600 346.000 453.200 ;
        RECT 346.800 450.200 347.400 453.600 ;
        RECT 348.400 451.600 349.200 453.200 ;
        RECT 350.000 452.800 350.800 453.700 ;
        RECT 351.600 453.600 352.400 453.700 ;
        RECT 354.800 453.600 355.600 453.800 ;
        RECT 358.000 453.700 360.400 454.300 ;
        RECT 364.000 454.200 364.800 459.800 ;
        RECT 370.400 454.200 371.200 459.800 ;
        RECT 377.200 457.600 378.000 459.800 ;
        RECT 375.600 455.600 376.400 457.200 ;
        RECT 377.400 454.400 378.000 457.600 ;
        RECT 384.000 454.400 384.800 459.800 ;
        RECT 351.600 452.300 352.400 452.400 ;
        RECT 353.200 452.300 354.000 453.200 ;
        RECT 351.600 451.700 354.000 452.300 ;
        RECT 351.600 451.600 352.400 451.700 ;
        RECT 353.200 451.600 354.000 451.700 ;
        RECT 354.800 450.200 355.400 453.600 ;
        RECT 356.400 451.600 357.200 453.200 ;
        RECT 358.000 452.800 358.800 453.700 ;
        RECT 326.000 449.600 327.400 450.200 ;
        RECT 328.000 449.600 329.000 450.200 ;
        RECT 332.400 449.600 333.800 450.200 ;
        RECT 334.400 449.600 335.400 450.200 ;
        RECT 315.400 442.200 316.200 449.400 ;
        RECT 319.800 447.000 320.400 449.600 ;
        RECT 321.200 447.600 322.000 449.200 ;
        RECT 326.800 448.400 327.400 449.600 ;
        RECT 326.800 447.600 327.600 448.400 ;
        RECT 319.800 446.400 323.400 447.000 ;
        RECT 319.800 446.200 320.400 446.400 ;
        RECT 319.600 442.200 320.400 446.200 ;
        RECT 322.800 446.200 323.400 446.400 ;
        RECT 322.800 442.200 323.600 446.200 ;
        RECT 328.200 442.200 329.000 449.600 ;
        RECT 333.200 448.400 333.800 449.600 ;
        RECT 333.200 447.600 334.000 448.400 ;
        RECT 334.600 442.200 335.400 449.600 ;
        RECT 340.400 449.400 342.200 450.200 ;
        RECT 341.400 442.200 342.200 449.400 ;
        RECT 346.200 442.200 348.200 450.200 ;
        RECT 354.200 442.200 356.200 450.200 ;
        RECT 359.600 442.200 360.400 453.700 ;
        RECT 363.000 453.800 364.800 454.200 ;
        RECT 369.400 453.800 371.200 454.200 ;
        RECT 363.000 453.600 364.600 453.800 ;
        RECT 369.400 453.600 371.000 453.800 ;
        RECT 377.200 453.600 378.000 454.400 ;
        RECT 382.000 454.300 382.800 454.400 ;
        RECT 383.600 454.300 384.800 454.400 ;
        RECT 382.000 454.200 384.800 454.300 ;
        RECT 390.400 454.200 391.200 459.800 ;
        RECT 394.800 456.000 395.600 459.800 ;
        RECT 394.600 455.200 395.600 456.000 ;
        RECT 382.000 453.700 385.800 454.200 ;
        RECT 390.400 453.800 392.200 454.200 ;
        RECT 382.000 453.600 382.800 453.700 ;
        RECT 384.200 453.600 385.800 453.700 ;
        RECT 390.600 453.600 392.200 453.800 ;
        RECT 363.000 450.400 363.600 453.600 ;
        RECT 365.200 451.600 366.800 452.400 ;
        RECT 362.800 449.600 363.600 450.400 ;
        RECT 367.600 449.600 368.400 451.200 ;
        RECT 369.400 450.400 370.000 453.600 ;
        RECT 371.600 451.600 373.200 452.400 ;
        RECT 369.200 449.600 370.000 450.400 ;
        RECT 374.000 449.600 374.800 451.200 ;
        RECT 377.400 450.200 378.000 453.600 ;
        RECT 378.800 450.800 379.600 452.400 ;
        RECT 382.000 451.600 383.600 452.400 ;
        RECT 363.000 447.000 363.600 449.600 ;
        RECT 364.400 447.600 365.200 449.200 ;
        RECT 369.400 447.000 370.000 449.600 ;
        RECT 377.200 449.400 379.000 450.200 ;
        RECT 380.400 449.600 381.200 451.200 ;
        RECT 385.200 450.400 385.800 453.600 ;
        RECT 388.400 451.600 390.000 452.400 ;
        RECT 385.200 449.600 386.000 450.400 ;
        RECT 386.800 449.600 387.600 451.200 ;
        RECT 391.600 450.400 392.200 453.600 ;
        RECT 394.600 450.800 395.400 455.200 ;
        RECT 396.400 454.600 397.200 459.800 ;
        RECT 402.800 456.600 403.600 459.800 ;
        RECT 404.400 457.000 405.200 459.800 ;
        RECT 406.000 457.000 406.800 459.800 ;
        RECT 407.600 457.000 408.400 459.800 ;
        RECT 409.200 457.000 410.000 459.800 ;
        RECT 412.400 457.000 413.200 459.800 ;
        RECT 415.600 457.000 416.400 459.800 ;
        RECT 417.200 457.000 418.000 459.800 ;
        RECT 418.800 457.000 419.600 459.800 ;
        RECT 401.200 455.800 403.600 456.600 ;
        RECT 420.400 456.600 421.200 459.800 ;
        RECT 401.200 455.200 402.000 455.800 ;
        RECT 396.000 454.000 397.200 454.600 ;
        RECT 400.200 454.600 402.000 455.200 ;
        RECT 406.000 455.600 407.000 456.400 ;
        RECT 410.000 455.600 411.600 456.400 ;
        RECT 412.400 455.800 417.000 456.400 ;
        RECT 420.400 455.800 423.000 456.600 ;
        RECT 412.400 455.600 413.200 455.800 ;
        RECT 396.000 452.000 396.600 454.000 ;
        RECT 400.200 453.400 401.000 454.600 ;
        RECT 397.200 452.600 401.000 453.400 ;
        RECT 406.000 452.800 406.800 455.600 ;
        RECT 412.400 454.800 413.200 455.000 ;
        RECT 408.800 454.200 413.200 454.800 ;
        RECT 408.800 454.000 409.600 454.200 ;
        RECT 414.000 453.600 414.800 455.200 ;
        RECT 416.200 453.400 417.000 455.800 ;
        RECT 422.200 455.200 423.000 455.800 ;
        RECT 422.200 454.400 425.200 455.200 ;
        RECT 426.800 453.800 427.600 459.800 ;
        RECT 435.800 458.400 436.600 459.800 ;
        RECT 435.800 457.600 437.200 458.400 ;
        RECT 435.800 456.400 436.600 457.600 ;
        RECT 434.800 455.800 436.600 456.400 ;
        RECT 409.200 452.600 412.400 453.400 ;
        RECT 416.200 452.600 418.200 453.400 ;
        RECT 418.800 453.000 427.600 453.800 ;
        RECT 431.600 454.300 432.400 454.400 ;
        RECT 433.200 454.300 434.000 455.200 ;
        RECT 431.600 453.700 434.000 454.300 ;
        RECT 431.600 453.600 432.400 453.700 ;
        RECT 433.200 453.600 434.000 453.700 ;
        RECT 402.800 452.000 403.600 452.600 ;
        RECT 420.400 452.000 421.200 452.400 ;
        RECT 423.600 452.000 424.400 452.400 ;
        RECT 425.400 452.000 426.200 452.200 ;
        RECT 396.000 451.400 396.800 452.000 ;
        RECT 402.800 451.400 426.200 452.000 ;
        RECT 391.600 449.600 392.400 450.400 ;
        RECT 394.600 450.000 395.600 450.800 ;
        RECT 370.800 447.600 371.600 449.200 ;
        RECT 363.000 446.400 366.600 447.000 ;
        RECT 362.800 442.200 363.600 446.400 ;
        RECT 366.000 446.200 366.600 446.400 ;
        RECT 369.400 446.400 373.000 447.000 ;
        RECT 369.400 446.200 370.000 446.400 ;
        RECT 366.000 442.200 366.800 446.200 ;
        RECT 369.200 442.200 370.000 446.200 ;
        RECT 372.400 442.200 373.200 446.400 ;
        RECT 378.200 444.400 379.000 449.400 ;
        RECT 383.600 447.600 384.400 449.200 ;
        RECT 385.200 447.000 385.800 449.600 ;
        RECT 390.000 447.600 390.800 449.200 ;
        RECT 391.600 447.000 392.200 449.600 ;
        RECT 382.200 446.400 385.800 447.000 ;
        RECT 388.600 446.400 392.200 447.000 ;
        RECT 382.200 446.200 382.800 446.400 ;
        RECT 378.200 443.600 379.600 444.400 ;
        RECT 378.200 442.200 379.000 443.600 ;
        RECT 382.000 442.200 382.800 446.200 ;
        RECT 385.200 446.200 385.800 446.400 ;
        RECT 385.200 442.200 386.000 446.200 ;
        RECT 388.400 442.200 389.200 446.400 ;
        RECT 391.600 446.200 392.200 446.400 ;
        RECT 391.600 442.200 392.400 446.200 ;
        RECT 394.800 442.200 395.600 450.000 ;
        RECT 396.200 449.600 396.800 451.400 ;
        RECT 396.200 449.000 405.200 449.600 ;
        RECT 396.200 447.400 396.800 449.000 ;
        RECT 404.400 448.800 405.200 449.000 ;
        RECT 407.600 449.000 416.200 449.600 ;
        RECT 407.600 448.800 408.400 449.000 ;
        RECT 399.400 447.600 402.000 448.400 ;
        RECT 396.200 446.800 398.800 447.400 ;
        RECT 398.000 442.200 398.800 446.800 ;
        RECT 401.200 442.200 402.000 447.600 ;
        RECT 402.600 446.800 406.800 447.600 ;
        RECT 404.400 442.200 405.200 445.000 ;
        RECT 406.000 442.200 406.800 445.000 ;
        RECT 407.600 442.200 408.400 445.000 ;
        RECT 409.200 442.200 410.000 448.400 ;
        RECT 412.400 447.600 415.000 448.400 ;
        RECT 415.600 448.200 416.200 449.000 ;
        RECT 417.200 449.400 418.000 449.600 ;
        RECT 417.200 449.000 422.600 449.400 ;
        RECT 417.200 448.800 423.400 449.000 ;
        RECT 422.000 448.200 423.400 448.800 ;
        RECT 415.600 447.600 421.400 448.200 ;
        RECT 424.400 448.000 426.000 448.800 ;
        RECT 424.400 447.600 425.000 448.000 ;
        RECT 412.400 442.200 413.200 447.000 ;
        RECT 415.600 442.200 416.400 447.000 ;
        RECT 420.800 446.800 425.000 447.600 ;
        RECT 426.800 447.400 427.600 453.000 ;
        RECT 425.600 446.800 427.600 447.400 ;
        RECT 417.200 442.200 418.000 445.000 ;
        RECT 418.800 442.200 419.600 445.000 ;
        RECT 422.000 442.200 422.800 446.800 ;
        RECT 425.600 446.200 426.200 446.800 ;
        RECT 425.200 445.600 426.200 446.200 ;
        RECT 425.200 442.200 426.000 445.600 ;
        RECT 434.800 442.200 435.600 455.800 ;
        RECT 438.000 453.800 438.800 459.800 ;
        RECT 444.400 456.600 445.200 459.800 ;
        RECT 446.000 457.000 446.800 459.800 ;
        RECT 447.600 457.000 448.400 459.800 ;
        RECT 449.200 457.000 450.000 459.800 ;
        RECT 452.400 457.000 453.200 459.800 ;
        RECT 455.600 457.000 456.400 459.800 ;
        RECT 457.200 457.000 458.000 459.800 ;
        RECT 458.800 457.000 459.600 459.800 ;
        RECT 460.400 457.000 461.200 459.800 ;
        RECT 442.600 455.800 445.200 456.600 ;
        RECT 462.000 456.600 462.800 459.800 ;
        RECT 448.600 455.800 453.200 456.400 ;
        RECT 442.600 455.200 443.400 455.800 ;
        RECT 440.400 454.400 443.400 455.200 ;
        RECT 438.000 453.000 446.800 453.800 ;
        RECT 448.600 453.400 449.400 455.800 ;
        RECT 452.400 455.600 453.200 455.800 ;
        RECT 454.000 455.600 455.600 456.400 ;
        RECT 458.600 455.600 459.600 456.400 ;
        RECT 462.000 455.800 464.400 456.600 ;
        RECT 450.800 453.600 451.600 455.200 ;
        RECT 452.400 454.800 453.200 455.000 ;
        RECT 452.400 454.200 456.800 454.800 ;
        RECT 456.000 454.000 456.800 454.200 ;
        RECT 436.400 448.800 437.200 450.400 ;
        RECT 438.000 447.400 438.800 453.000 ;
        RECT 447.400 452.600 449.400 453.400 ;
        RECT 453.200 452.600 456.400 453.400 ;
        RECT 458.800 452.800 459.600 455.600 ;
        RECT 463.600 455.200 464.400 455.800 ;
        RECT 463.600 454.600 465.400 455.200 ;
        RECT 464.600 453.400 465.400 454.600 ;
        RECT 468.400 454.600 469.200 459.800 ;
        RECT 470.000 456.000 470.800 459.800 ;
        RECT 475.800 458.400 476.600 459.800 ;
        RECT 475.800 457.600 477.200 458.400 ;
        RECT 475.800 456.400 476.600 457.600 ;
        RECT 470.000 455.200 471.000 456.000 ;
        RECT 474.800 455.800 476.600 456.400 ;
        RECT 468.400 454.000 469.600 454.600 ;
        RECT 464.600 452.600 468.400 453.400 ;
        RECT 439.400 452.000 440.200 452.200 ;
        RECT 444.400 452.000 445.200 452.400 ;
        RECT 450.800 452.000 451.600 452.400 ;
        RECT 462.000 452.000 462.800 452.600 ;
        RECT 469.000 452.000 469.600 454.000 ;
        RECT 439.400 451.400 462.800 452.000 ;
        RECT 468.800 451.400 469.600 452.000 ;
        RECT 468.800 449.600 469.400 451.400 ;
        RECT 470.200 450.800 471.000 455.200 ;
        RECT 473.200 453.600 474.000 455.200 ;
        RECT 447.600 449.400 448.400 449.600 ;
        RECT 443.000 449.000 448.400 449.400 ;
        RECT 442.200 448.800 448.400 449.000 ;
        RECT 449.400 449.000 458.000 449.600 ;
        RECT 439.600 448.000 441.200 448.800 ;
        RECT 442.200 448.200 443.600 448.800 ;
        RECT 449.400 448.200 450.000 449.000 ;
        RECT 457.200 448.800 458.000 449.000 ;
        RECT 460.400 449.000 469.400 449.600 ;
        RECT 460.400 448.800 461.200 449.000 ;
        RECT 440.600 447.600 441.200 448.000 ;
        RECT 444.200 447.600 450.000 448.200 ;
        RECT 450.600 447.600 453.200 448.400 ;
        RECT 438.000 446.800 440.000 447.400 ;
        RECT 440.600 446.800 444.800 447.600 ;
        RECT 439.400 446.200 440.000 446.800 ;
        RECT 439.400 445.600 440.400 446.200 ;
        RECT 439.600 442.200 440.400 445.600 ;
        RECT 442.800 442.200 443.600 446.800 ;
        RECT 446.000 442.200 446.800 445.000 ;
        RECT 447.600 442.200 448.400 445.000 ;
        RECT 449.200 442.200 450.000 447.000 ;
        RECT 452.400 442.200 453.200 447.000 ;
        RECT 455.600 442.200 456.400 448.400 ;
        RECT 463.600 447.600 466.200 448.400 ;
        RECT 458.800 446.800 463.000 447.600 ;
        RECT 457.200 442.200 458.000 445.000 ;
        RECT 458.800 442.200 459.600 445.000 ;
        RECT 460.400 442.200 461.200 445.000 ;
        RECT 463.600 442.200 464.400 447.600 ;
        RECT 468.800 447.400 469.400 449.000 ;
        RECT 466.800 446.800 469.400 447.400 ;
        RECT 470.000 450.000 471.000 450.800 ;
        RECT 466.800 442.200 467.600 446.800 ;
        RECT 470.000 442.200 470.800 450.000 ;
        RECT 474.800 442.200 475.600 455.800 ;
        RECT 476.400 448.800 477.200 450.400 ;
        RECT 478.000 442.200 478.800 459.800 ;
        RECT 479.600 455.600 480.400 457.200 ;
        RECT 481.200 456.000 482.000 459.800 ;
        RECT 484.400 456.000 485.200 459.800 ;
        RECT 481.200 455.800 485.200 456.000 ;
        RECT 486.000 455.800 486.800 459.800 ;
        RECT 481.400 455.400 485.000 455.800 ;
        RECT 482.000 454.400 482.800 454.800 ;
        RECT 486.000 454.400 486.600 455.800 ;
        RECT 481.200 453.800 482.800 454.400 ;
        RECT 481.200 453.600 482.000 453.800 ;
        RECT 484.200 453.600 486.800 454.400 ;
        RECT 479.600 452.300 480.400 452.400 ;
        RECT 482.800 452.300 483.600 453.200 ;
        RECT 479.600 451.700 483.600 452.300 ;
        RECT 479.600 451.600 480.400 451.700 ;
        RECT 482.800 451.600 483.600 451.700 ;
        RECT 484.200 452.400 484.800 453.600 ;
        RECT 484.200 451.600 485.200 452.400 ;
        RECT 484.200 450.200 484.800 451.600 ;
        RECT 486.000 450.200 486.800 450.400 ;
        RECT 483.800 449.600 484.800 450.200 ;
        RECT 485.400 449.600 486.800 450.200 ;
        RECT 483.800 442.200 484.600 449.600 ;
        RECT 485.400 448.400 486.000 449.600 ;
        RECT 485.200 447.600 486.000 448.400 ;
        RECT 487.600 448.300 488.400 459.800 ;
        RECT 492.400 456.400 493.200 459.800 ;
        RECT 492.200 455.800 493.200 456.400 ;
        RECT 492.200 454.400 492.800 455.800 ;
        RECT 495.600 455.200 496.400 459.800 ;
        RECT 493.800 454.600 496.400 455.200 ;
        RECT 492.200 453.600 493.200 454.400 ;
        RECT 492.200 450.200 492.800 453.600 ;
        RECT 493.800 453.000 494.400 454.600 ;
        RECT 497.200 453.800 498.000 459.800 ;
        RECT 503.600 456.600 504.400 459.800 ;
        RECT 505.200 457.000 506.000 459.800 ;
        RECT 506.800 457.000 507.600 459.800 ;
        RECT 508.400 457.000 509.200 459.800 ;
        RECT 511.600 457.000 512.400 459.800 ;
        RECT 514.800 457.000 515.600 459.800 ;
        RECT 516.400 457.000 517.200 459.800 ;
        RECT 518.000 457.000 518.800 459.800 ;
        RECT 519.600 457.000 520.400 459.800 ;
        RECT 501.800 455.800 504.400 456.600 ;
        RECT 521.200 456.600 522.000 459.800 ;
        RECT 507.800 455.800 512.400 456.400 ;
        RECT 501.800 455.200 502.600 455.800 ;
        RECT 499.600 454.400 502.600 455.200 ;
        RECT 493.400 452.200 494.400 453.000 ;
        RECT 493.800 450.200 494.400 452.200 ;
        RECT 495.400 452.400 496.200 453.200 ;
        RECT 497.200 453.000 506.000 453.800 ;
        RECT 507.800 453.400 508.600 455.800 ;
        RECT 511.600 455.600 512.400 455.800 ;
        RECT 513.200 455.600 514.800 456.400 ;
        RECT 517.800 455.600 518.800 456.400 ;
        RECT 521.200 455.800 523.600 456.600 ;
        RECT 510.000 453.600 510.800 455.200 ;
        RECT 511.600 454.800 512.400 455.000 ;
        RECT 511.600 454.200 516.000 454.800 ;
        RECT 515.200 454.000 516.000 454.200 ;
        RECT 495.400 451.600 496.400 452.400 ;
        RECT 492.200 449.200 493.200 450.200 ;
        RECT 493.800 449.600 496.400 450.200 ;
        RECT 489.200 448.300 490.000 448.400 ;
        RECT 487.600 447.700 490.000 448.300 ;
        RECT 487.600 442.200 488.400 447.700 ;
        RECT 489.200 447.600 490.000 447.700 ;
        RECT 492.400 442.200 493.200 449.200 ;
        RECT 495.600 442.200 496.400 449.600 ;
        RECT 497.200 447.400 498.000 453.000 ;
        RECT 506.600 452.600 508.600 453.400 ;
        RECT 512.400 452.600 515.600 453.400 ;
        RECT 518.000 452.800 518.800 455.600 ;
        RECT 522.800 455.200 523.600 455.800 ;
        RECT 522.800 454.600 524.600 455.200 ;
        RECT 523.800 453.400 524.600 454.600 ;
        RECT 527.600 454.600 528.400 459.800 ;
        RECT 529.200 456.000 530.000 459.800 ;
        RECT 530.800 456.300 531.600 456.400 ;
        RECT 532.400 456.300 533.200 459.800 ;
        RECT 529.200 455.200 530.200 456.000 ;
        RECT 530.800 455.700 533.200 456.300 ;
        RECT 534.000 456.000 534.800 459.800 ;
        RECT 537.200 456.000 538.000 459.800 ;
        RECT 534.000 455.800 538.000 456.000 ;
        RECT 530.800 455.600 531.600 455.700 ;
        RECT 527.600 454.000 528.800 454.600 ;
        RECT 523.800 452.600 527.600 453.400 ;
        RECT 498.600 452.000 499.400 452.200 ;
        RECT 502.000 452.000 502.800 452.400 ;
        RECT 503.600 452.000 504.400 452.400 ;
        RECT 521.200 452.000 522.000 452.600 ;
        RECT 528.200 452.000 528.800 454.000 ;
        RECT 498.600 451.400 522.000 452.000 ;
        RECT 528.000 451.400 528.800 452.000 ;
        RECT 528.000 449.600 528.600 451.400 ;
        RECT 529.400 450.800 530.200 455.200 ;
        RECT 532.600 454.400 533.200 455.700 ;
        RECT 534.200 455.400 537.800 455.800 ;
        RECT 536.400 454.400 537.200 454.800 ;
        RECT 532.400 453.600 535.000 454.400 ;
        RECT 536.400 454.300 538.000 454.400 ;
        RECT 538.800 454.300 539.600 459.800 ;
        RECT 544.600 458.400 545.400 459.800 ;
        RECT 543.600 457.600 545.400 458.400 ;
        RECT 544.600 456.400 545.400 457.600 ;
        RECT 549.400 458.400 550.200 459.800 ;
        RECT 549.400 457.600 550.800 458.400 ;
        RECT 553.200 457.800 554.000 459.800 ;
        RECT 549.400 456.400 550.200 457.600 ;
        RECT 543.600 455.800 545.400 456.400 ;
        RECT 548.400 455.800 550.200 456.400 ;
        RECT 536.400 453.800 539.600 454.300 ;
        RECT 537.200 453.700 539.600 453.800 ;
        RECT 537.200 453.600 538.000 453.700 ;
        RECT 506.800 449.400 507.600 449.600 ;
        RECT 502.200 449.000 507.600 449.400 ;
        RECT 501.400 448.800 507.600 449.000 ;
        RECT 508.600 449.000 517.200 449.600 ;
        RECT 498.800 448.000 500.400 448.800 ;
        RECT 501.400 448.200 502.800 448.800 ;
        RECT 508.600 448.200 509.200 449.000 ;
        RECT 516.400 448.800 517.200 449.000 ;
        RECT 519.600 449.000 528.600 449.600 ;
        RECT 519.600 448.800 520.400 449.000 ;
        RECT 499.800 447.600 500.400 448.000 ;
        RECT 503.400 447.600 509.200 448.200 ;
        RECT 509.800 447.600 512.400 448.400 ;
        RECT 497.200 446.800 499.200 447.400 ;
        RECT 499.800 446.800 504.000 447.600 ;
        RECT 498.600 446.200 499.200 446.800 ;
        RECT 498.600 445.600 499.600 446.200 ;
        RECT 498.800 442.200 499.600 445.600 ;
        RECT 502.000 442.200 502.800 446.800 ;
        RECT 505.200 442.200 506.000 445.000 ;
        RECT 506.800 442.200 507.600 445.000 ;
        RECT 508.400 442.200 509.200 447.000 ;
        RECT 511.600 442.200 512.400 447.000 ;
        RECT 514.800 442.200 515.600 448.400 ;
        RECT 522.800 447.600 525.400 448.400 ;
        RECT 518.000 446.800 522.200 447.600 ;
        RECT 516.400 442.200 517.200 445.000 ;
        RECT 518.000 442.200 518.800 445.000 ;
        RECT 519.600 442.200 520.400 445.000 ;
        RECT 522.800 442.200 523.600 447.600 ;
        RECT 528.000 447.400 528.600 449.000 ;
        RECT 526.000 446.800 528.600 447.400 ;
        RECT 529.200 450.000 530.200 450.800 ;
        RECT 530.800 450.300 531.600 450.400 ;
        RECT 532.400 450.300 533.200 450.400 ;
        RECT 530.800 450.200 533.200 450.300 ;
        RECT 534.400 450.200 535.000 453.600 ;
        RECT 535.600 452.300 536.400 453.200 ;
        RECT 537.200 452.300 538.000 452.400 ;
        RECT 535.600 451.700 538.000 452.300 ;
        RECT 535.600 451.600 536.400 451.700 ;
        RECT 537.200 451.600 538.000 451.700 ;
        RECT 529.200 448.300 530.000 450.000 ;
        RECT 530.800 449.700 533.800 450.200 ;
        RECT 530.800 449.600 531.600 449.700 ;
        RECT 532.400 449.600 533.800 449.700 ;
        RECT 534.400 449.600 535.400 450.200 ;
        RECT 533.200 448.400 533.800 449.600 ;
        RECT 530.800 448.300 531.600 448.400 ;
        RECT 529.200 447.700 531.600 448.300 ;
        RECT 526.000 442.200 526.800 446.800 ;
        RECT 529.200 442.200 530.000 447.700 ;
        RECT 530.800 447.600 531.600 447.700 ;
        RECT 533.200 447.600 534.000 448.400 ;
        RECT 534.600 442.200 535.400 449.600 ;
        RECT 538.800 442.200 539.600 453.700 ;
        RECT 542.000 453.600 542.800 455.200 ;
        RECT 543.600 442.200 544.400 455.800 ;
        RECT 546.800 453.600 547.600 455.200 ;
        RECT 545.200 450.300 546.000 450.400 ;
        RECT 546.800 450.300 547.600 450.400 ;
        RECT 545.200 449.700 547.600 450.300 ;
        RECT 545.200 448.800 546.000 449.700 ;
        RECT 546.800 449.600 547.600 449.700 ;
        RECT 548.400 442.200 549.200 455.800 ;
        RECT 551.600 455.600 552.400 457.200 ;
        RECT 553.400 454.400 554.000 457.800 ;
        RECT 562.800 456.000 563.600 459.800 ;
        RECT 553.200 453.600 554.000 454.400 ;
        RECT 550.000 448.800 550.800 450.400 ;
        RECT 553.400 450.200 554.000 453.600 ;
        RECT 562.600 455.200 563.600 456.000 ;
        RECT 554.800 452.300 555.600 452.400 ;
        RECT 559.600 452.300 560.400 452.400 ;
        RECT 554.800 451.700 560.400 452.300 ;
        RECT 554.800 450.800 555.600 451.700 ;
        RECT 559.600 451.600 560.400 451.700 ;
        RECT 562.600 450.800 563.400 455.200 ;
        RECT 564.400 454.600 565.200 459.800 ;
        RECT 570.800 456.600 571.600 459.800 ;
        RECT 572.400 457.000 573.200 459.800 ;
        RECT 574.000 457.000 574.800 459.800 ;
        RECT 575.600 457.000 576.400 459.800 ;
        RECT 577.200 457.000 578.000 459.800 ;
        RECT 580.400 457.000 581.200 459.800 ;
        RECT 583.600 457.000 584.400 459.800 ;
        RECT 585.200 457.000 586.000 459.800 ;
        RECT 586.800 457.000 587.600 459.800 ;
        RECT 569.200 455.800 571.600 456.600 ;
        RECT 588.400 456.600 589.200 459.800 ;
        RECT 569.200 455.200 570.000 455.800 ;
        RECT 564.000 454.000 565.200 454.600 ;
        RECT 568.200 454.600 570.000 455.200 ;
        RECT 574.000 455.600 575.000 456.400 ;
        RECT 578.000 455.600 579.600 456.400 ;
        RECT 580.400 455.800 585.000 456.400 ;
        RECT 588.400 455.800 591.000 456.600 ;
        RECT 580.400 455.600 581.200 455.800 ;
        RECT 564.000 452.000 564.600 454.000 ;
        RECT 568.200 453.400 569.000 454.600 ;
        RECT 565.200 452.600 569.000 453.400 ;
        RECT 574.000 452.800 574.800 455.600 ;
        RECT 580.400 454.800 581.200 455.000 ;
        RECT 576.800 454.200 581.200 454.800 ;
        RECT 576.800 454.000 577.600 454.200 ;
        RECT 582.000 453.600 582.800 455.200 ;
        RECT 584.200 453.400 585.000 455.800 ;
        RECT 590.200 455.200 591.000 455.800 ;
        RECT 590.200 454.400 593.200 455.200 ;
        RECT 594.800 453.800 595.600 459.800 ;
        RECT 596.400 455.800 597.200 459.800 ;
        RECT 598.000 456.000 598.800 459.800 ;
        RECT 601.200 456.000 602.000 459.800 ;
        RECT 598.000 455.800 602.000 456.000 ;
        RECT 596.600 454.400 597.200 455.800 ;
        RECT 598.200 455.400 601.800 455.800 ;
        RECT 602.800 455.200 603.600 459.800 ;
        RECT 606.000 456.400 606.800 459.800 ;
        RECT 609.400 456.400 610.200 457.200 ;
        RECT 606.000 455.800 607.000 456.400 ;
        RECT 600.400 454.400 601.200 454.800 ;
        RECT 602.800 454.600 605.400 455.200 ;
        RECT 577.200 452.600 580.400 453.400 ;
        RECT 584.200 452.600 586.200 453.400 ;
        RECT 586.800 453.000 595.600 453.800 ;
        RECT 596.400 453.600 599.000 454.400 ;
        RECT 600.400 453.800 602.000 454.400 ;
        RECT 601.200 453.600 602.000 453.800 ;
        RECT 570.800 452.000 571.600 452.600 ;
        RECT 588.400 452.000 589.200 452.400 ;
        RECT 591.600 452.000 592.400 452.400 ;
        RECT 593.400 452.000 594.200 452.200 ;
        RECT 564.000 451.400 564.800 452.000 ;
        RECT 570.800 451.400 594.200 452.000 ;
        RECT 553.200 449.400 555.000 450.200 ;
        RECT 562.600 450.000 563.600 450.800 ;
        RECT 554.200 444.400 555.000 449.400 ;
        RECT 561.200 448.300 562.000 448.400 ;
        RECT 562.800 448.300 563.600 450.000 ;
        RECT 561.200 447.700 563.600 448.300 ;
        RECT 561.200 447.600 562.000 447.700 ;
        RECT 554.200 443.600 555.600 444.400 ;
        RECT 554.200 442.200 555.000 443.600 ;
        RECT 562.800 442.200 563.600 447.700 ;
        RECT 564.200 449.600 564.800 451.400 ;
        RECT 564.200 449.000 573.200 449.600 ;
        RECT 564.200 447.400 564.800 449.000 ;
        RECT 572.400 448.800 573.200 449.000 ;
        RECT 575.600 449.000 584.200 449.600 ;
        RECT 575.600 448.800 576.400 449.000 ;
        RECT 567.400 447.600 570.000 448.400 ;
        RECT 564.200 446.800 566.800 447.400 ;
        RECT 566.000 442.200 566.800 446.800 ;
        RECT 569.200 442.200 570.000 447.600 ;
        RECT 570.600 446.800 574.800 447.600 ;
        RECT 572.400 442.200 573.200 445.000 ;
        RECT 574.000 442.200 574.800 445.000 ;
        RECT 575.600 442.200 576.400 445.000 ;
        RECT 577.200 442.200 578.000 448.400 ;
        RECT 580.400 447.600 583.000 448.400 ;
        RECT 583.600 448.200 584.200 449.000 ;
        RECT 585.200 449.400 586.000 449.600 ;
        RECT 585.200 449.000 590.600 449.400 ;
        RECT 585.200 448.800 591.400 449.000 ;
        RECT 590.000 448.200 591.400 448.800 ;
        RECT 583.600 447.600 589.400 448.200 ;
        RECT 592.400 448.000 594.000 448.800 ;
        RECT 592.400 447.600 593.000 448.000 ;
        RECT 580.400 442.200 581.200 447.000 ;
        RECT 583.600 442.200 584.400 447.000 ;
        RECT 588.800 446.800 593.000 447.600 ;
        RECT 594.800 447.400 595.600 453.000 ;
        RECT 596.400 450.200 597.200 450.400 ;
        RECT 598.400 450.200 599.000 453.600 ;
        RECT 599.600 451.600 600.400 453.200 ;
        RECT 603.000 452.400 603.800 453.200 ;
        RECT 602.800 451.600 603.800 452.400 ;
        RECT 604.800 453.000 605.400 454.600 ;
        RECT 606.400 454.400 607.000 455.800 ;
        RECT 609.200 455.600 610.000 456.400 ;
        RECT 610.800 455.800 611.600 459.800 ;
        RECT 617.200 457.800 618.000 459.800 ;
        RECT 606.000 453.600 607.000 454.400 ;
        RECT 604.800 452.200 605.800 453.000 ;
        RECT 604.800 450.200 605.400 452.200 ;
        RECT 606.400 450.200 607.000 453.600 ;
        RECT 609.200 452.200 610.000 452.400 ;
        RECT 611.000 452.200 611.600 455.800 ;
        RECT 615.600 455.600 616.400 457.200 ;
        RECT 617.400 454.400 618.000 457.800 ;
        RECT 612.400 452.800 613.200 454.400 ;
        RECT 617.200 453.600 618.000 454.400 ;
        RECT 614.000 452.200 614.800 452.400 ;
        RECT 609.200 451.600 611.600 452.200 ;
        RECT 613.200 451.600 614.800 452.200 ;
        RECT 609.400 450.200 610.000 451.600 ;
        RECT 613.200 451.200 614.000 451.600 ;
        RECT 617.400 450.400 618.000 453.600 ;
        RECT 622.000 457.800 622.800 459.800 ;
        RECT 622.000 454.400 622.600 457.800 ;
        RECT 623.600 455.600 624.400 457.200 ;
        RECT 625.200 455.600 626.000 457.200 ;
        RECT 622.000 453.600 622.800 454.400 ;
        RECT 623.700 454.300 624.300 455.600 ;
        RECT 626.800 454.300 627.600 459.800 ;
        RECT 623.700 453.700 627.600 454.300 ;
        RECT 629.600 454.200 630.400 459.800 ;
        RECT 636.400 456.000 637.200 459.800 ;
        RECT 622.000 452.400 622.600 453.600 ;
        RECT 618.800 452.300 619.600 452.400 ;
        RECT 620.400 452.300 621.200 452.400 ;
        RECT 618.800 451.700 621.200 452.300 ;
        RECT 618.800 450.800 619.600 451.700 ;
        RECT 620.400 450.800 621.200 451.700 ;
        RECT 622.000 451.600 622.800 452.400 ;
        RECT 617.200 450.200 618.000 450.400 ;
        RECT 622.000 450.200 622.600 451.600 ;
        RECT 596.400 449.600 597.800 450.200 ;
        RECT 598.400 449.600 599.400 450.200 ;
        RECT 597.200 448.400 597.800 449.600 ;
        RECT 597.200 447.600 598.000 448.400 ;
        RECT 593.600 446.800 595.600 447.400 ;
        RECT 585.200 442.200 586.000 445.000 ;
        RECT 586.800 442.200 587.600 445.000 ;
        RECT 590.000 442.200 590.800 446.800 ;
        RECT 593.600 446.200 594.200 446.800 ;
        RECT 593.200 445.600 594.200 446.200 ;
        RECT 593.200 442.200 594.000 445.600 ;
        RECT 598.600 442.200 599.400 449.600 ;
        RECT 602.800 449.600 605.400 450.200 ;
        RECT 602.800 442.200 603.600 449.600 ;
        RECT 606.000 449.200 607.000 450.200 ;
        RECT 606.000 442.200 606.800 449.200 ;
        RECT 609.200 442.200 610.000 450.200 ;
        RECT 610.800 449.600 614.800 450.200 ;
        RECT 610.800 442.200 611.600 449.600 ;
        RECT 614.000 442.200 614.800 449.600 ;
        RECT 617.200 449.400 619.000 450.200 ;
        RECT 618.200 442.200 619.000 449.400 ;
        RECT 621.000 449.400 622.800 450.200 ;
        RECT 621.000 442.200 621.800 449.400 ;
        RECT 626.800 442.200 627.600 453.700 ;
        RECT 628.600 453.800 630.400 454.200 ;
        RECT 636.200 455.200 637.200 456.000 ;
        RECT 628.600 453.600 630.200 453.800 ;
        RECT 628.600 450.400 629.200 453.600 ;
        RECT 630.800 451.600 632.400 452.400 ;
        RECT 628.400 449.600 629.200 450.400 ;
        RECT 633.200 450.300 634.000 451.200 ;
        RECT 636.200 450.800 637.000 455.200 ;
        RECT 638.000 454.600 638.800 459.800 ;
        RECT 644.400 456.600 645.200 459.800 ;
        RECT 646.000 457.000 646.800 459.800 ;
        RECT 647.600 457.000 648.400 459.800 ;
        RECT 649.200 457.000 650.000 459.800 ;
        RECT 650.800 457.000 651.600 459.800 ;
        RECT 654.000 457.000 654.800 459.800 ;
        RECT 657.200 457.000 658.000 459.800 ;
        RECT 658.800 457.000 659.600 459.800 ;
        RECT 660.400 457.000 661.200 459.800 ;
        RECT 642.800 455.800 645.200 456.600 ;
        RECT 662.000 456.600 662.800 459.800 ;
        RECT 642.800 455.200 643.600 455.800 ;
        RECT 637.600 454.000 638.800 454.600 ;
        RECT 641.800 454.600 643.600 455.200 ;
        RECT 647.600 455.600 648.600 456.400 ;
        RECT 651.600 455.600 653.200 456.400 ;
        RECT 654.000 455.800 658.600 456.400 ;
        RECT 662.000 455.800 664.600 456.600 ;
        RECT 654.000 455.600 654.800 455.800 ;
        RECT 637.600 452.000 638.200 454.000 ;
        RECT 641.800 453.400 642.600 454.600 ;
        RECT 638.800 452.600 642.600 453.400 ;
        RECT 647.600 452.800 648.400 455.600 ;
        RECT 654.000 454.800 654.800 455.000 ;
        RECT 650.400 454.200 654.800 454.800 ;
        RECT 650.400 454.000 651.200 454.200 ;
        RECT 655.600 453.600 656.400 455.200 ;
        RECT 657.800 453.400 658.600 455.800 ;
        RECT 663.800 455.200 664.600 455.800 ;
        RECT 663.800 454.400 666.800 455.200 ;
        RECT 668.400 453.800 669.200 459.800 ;
        RECT 671.600 455.200 672.400 459.800 ;
        RECT 674.800 455.200 675.600 459.800 ;
        RECT 678.000 455.200 678.800 459.800 ;
        RECT 681.200 455.200 682.000 459.800 ;
        RECT 671.600 454.400 673.400 455.200 ;
        RECT 674.800 454.400 677.000 455.200 ;
        RECT 678.000 454.400 680.200 455.200 ;
        RECT 681.200 454.400 683.600 455.200 ;
        RECT 650.800 452.600 654.000 453.400 ;
        RECT 657.800 452.600 659.800 453.400 ;
        RECT 660.400 453.000 669.200 453.800 ;
        RECT 670.000 453.800 670.800 454.400 ;
        RECT 672.600 453.800 673.400 454.400 ;
        RECT 676.200 453.800 677.000 454.400 ;
        RECT 679.400 453.800 680.200 454.400 ;
        RECT 670.000 453.000 671.800 453.800 ;
        RECT 672.600 453.000 675.200 453.800 ;
        RECT 676.200 453.000 678.600 453.800 ;
        RECT 679.400 453.000 682.000 453.800 ;
        RECT 644.400 452.000 645.200 452.600 ;
        RECT 662.000 452.000 662.800 452.400 ;
        RECT 667.000 452.000 667.800 452.200 ;
        RECT 637.600 451.400 638.400 452.000 ;
        RECT 644.400 451.400 667.800 452.000 ;
        RECT 636.200 450.300 637.200 450.800 ;
        RECT 633.200 449.700 637.200 450.300 ;
        RECT 633.200 449.600 634.000 449.700 ;
        RECT 628.600 447.000 629.200 449.600 ;
        RECT 630.000 447.600 630.800 449.200 ;
        RECT 628.600 446.400 632.200 447.000 ;
        RECT 628.400 442.200 629.200 446.400 ;
        RECT 631.600 446.200 632.200 446.400 ;
        RECT 631.600 442.200 632.400 446.200 ;
        RECT 636.400 442.200 637.200 449.700 ;
        RECT 637.800 449.600 638.400 451.400 ;
        RECT 637.800 449.000 646.800 449.600 ;
        RECT 637.800 447.400 638.400 449.000 ;
        RECT 646.000 448.800 646.800 449.000 ;
        RECT 649.200 449.000 657.800 449.600 ;
        RECT 649.200 448.800 650.000 449.000 ;
        RECT 641.000 447.600 643.600 448.400 ;
        RECT 637.800 446.800 640.400 447.400 ;
        RECT 639.600 442.200 640.400 446.800 ;
        RECT 642.800 442.200 643.600 447.600 ;
        RECT 644.200 446.800 648.400 447.600 ;
        RECT 646.000 442.200 646.800 445.000 ;
        RECT 647.600 442.200 648.400 445.000 ;
        RECT 649.200 442.200 650.000 445.000 ;
        RECT 650.800 442.200 651.600 448.400 ;
        RECT 654.000 447.600 656.600 448.400 ;
        RECT 657.200 448.200 657.800 449.000 ;
        RECT 658.800 449.400 659.600 449.600 ;
        RECT 658.800 449.000 664.200 449.400 ;
        RECT 658.800 448.800 665.000 449.000 ;
        RECT 663.600 448.200 665.000 448.800 ;
        RECT 657.200 447.600 663.000 448.200 ;
        RECT 666.000 448.000 667.600 448.800 ;
        RECT 666.000 447.600 666.600 448.000 ;
        RECT 654.000 442.200 654.800 447.000 ;
        RECT 657.200 442.200 658.000 447.000 ;
        RECT 662.400 446.800 666.600 447.600 ;
        RECT 668.400 447.400 669.200 453.000 ;
        RECT 672.600 451.600 673.400 453.000 ;
        RECT 676.200 451.600 677.000 453.000 ;
        RECT 679.400 451.600 680.200 453.000 ;
        RECT 682.800 451.600 683.600 454.400 ;
        RECT 667.200 446.800 669.200 447.400 ;
        RECT 671.600 450.800 673.400 451.600 ;
        RECT 674.800 450.800 677.000 451.600 ;
        RECT 678.000 450.800 680.200 451.600 ;
        RECT 681.200 450.800 683.600 451.600 ;
        RECT 658.800 442.200 659.600 445.000 ;
        RECT 660.400 442.200 661.200 445.000 ;
        RECT 663.600 442.200 664.400 446.800 ;
        RECT 667.200 446.200 667.800 446.800 ;
        RECT 666.800 445.600 667.800 446.200 ;
        RECT 666.800 442.200 667.600 445.600 ;
        RECT 671.600 442.200 672.400 450.800 ;
        RECT 674.800 442.200 675.600 450.800 ;
        RECT 678.000 442.200 678.800 450.800 ;
        RECT 681.200 442.200 682.000 450.800 ;
        RECT 1.200 431.200 2.000 439.800 ;
        RECT 5.400 435.800 6.600 439.800 ;
        RECT 10.000 435.800 10.800 439.800 ;
        RECT 14.400 436.400 15.200 439.800 ;
        RECT 14.400 435.800 16.400 436.400 ;
        RECT 6.000 435.000 6.800 435.800 ;
        RECT 10.200 435.200 10.800 435.800 ;
        RECT 9.400 434.600 13.000 435.200 ;
        RECT 15.600 435.000 16.400 435.800 ;
        RECT 9.400 434.400 10.200 434.600 ;
        RECT 12.200 434.400 13.000 434.600 ;
        RECT 5.200 433.200 6.600 434.000 ;
        RECT 6.000 432.200 6.600 433.200 ;
        RECT 8.200 433.000 10.400 433.600 ;
        RECT 8.200 432.800 9.000 433.000 ;
        RECT 6.000 431.600 8.400 432.200 ;
        RECT 1.200 430.600 5.400 431.200 ;
        RECT 1.200 427.200 2.000 430.600 ;
        RECT 4.600 430.400 5.400 430.600 ;
        RECT 3.000 429.800 3.800 430.000 ;
        RECT 3.000 429.200 6.800 429.800 ;
        RECT 6.000 429.000 6.800 429.200 ;
        RECT 7.800 428.400 8.400 431.600 ;
        RECT 9.800 431.800 10.400 433.000 ;
        RECT 11.000 433.000 11.800 433.200 ;
        RECT 15.600 433.000 16.400 433.200 ;
        RECT 11.000 432.400 16.400 433.000 ;
        RECT 9.800 431.400 14.600 431.800 ;
        RECT 18.800 431.400 19.600 439.800 ;
        RECT 23.000 432.400 23.800 439.800 ;
        RECT 24.400 433.600 25.200 434.400 ;
        RECT 24.600 432.400 25.200 433.600 ;
        RECT 27.600 433.600 28.400 434.400 ;
        RECT 27.600 432.400 28.200 433.600 ;
        RECT 29.000 432.400 29.800 439.800 ;
        RECT 37.000 438.400 37.800 439.800 ;
        RECT 36.400 437.600 37.800 438.400 ;
        RECT 37.000 432.800 37.800 437.600 ;
        RECT 41.200 435.000 42.000 439.000 ;
        RECT 23.000 431.800 24.000 432.400 ;
        RECT 24.600 431.800 26.000 432.400 ;
        RECT 9.800 431.200 19.600 431.400 ;
        RECT 13.800 431.000 19.600 431.200 ;
        RECT 14.000 430.800 19.600 431.000 ;
        RECT 23.400 430.400 24.000 431.800 ;
        RECT 25.200 431.600 26.000 431.800 ;
        RECT 26.800 431.800 28.200 432.400 ;
        RECT 28.800 431.800 29.800 432.400 ;
        RECT 36.200 432.200 37.800 432.800 ;
        RECT 26.800 431.600 27.600 431.800 ;
        RECT 12.400 430.200 13.200 430.400 ;
        RECT 12.400 429.600 17.400 430.200 ;
        RECT 14.000 429.400 14.800 429.600 ;
        RECT 16.600 429.400 17.400 429.600 ;
        RECT 22.000 428.800 22.800 430.400 ;
        RECT 23.400 429.600 24.400 430.400 ;
        RECT 25.300 430.300 25.900 431.600 ;
        RECT 28.800 430.300 29.400 431.800 ;
        RECT 25.300 429.700 29.400 430.300 ;
        RECT 15.000 428.400 15.800 428.600 ;
        RECT 23.400 428.400 24.000 429.600 ;
        RECT 28.800 428.400 29.400 429.700 ;
        RECT 30.000 428.800 30.800 430.400 ;
        RECT 34.800 429.600 35.600 431.200 ;
        RECT 36.200 428.400 36.800 432.200 ;
        RECT 41.400 431.600 42.000 435.000 ;
        RECT 43.600 433.600 44.400 434.400 ;
        RECT 43.600 432.400 44.200 433.600 ;
        RECT 45.000 432.400 45.800 439.800 ;
        RECT 50.800 432.800 51.600 439.800 ;
        RECT 42.800 431.800 44.200 432.400 ;
        RECT 44.800 431.800 45.800 432.400 ;
        RECT 50.600 431.800 51.600 432.800 ;
        RECT 54.000 432.400 54.800 439.800 ;
        RECT 52.200 431.800 54.800 432.400 ;
        RECT 55.600 435.000 56.400 439.000 ;
        RECT 42.800 431.600 43.600 431.800 ;
        RECT 38.200 431.000 42.000 431.600 ;
        RECT 38.200 429.000 38.800 431.000 ;
        RECT 7.800 427.800 18.800 428.400 ;
        RECT 8.200 427.600 9.000 427.800 ;
        RECT 1.200 426.600 5.000 427.200 ;
        RECT 1.200 422.200 2.000 426.600 ;
        RECT 4.200 426.400 5.000 426.600 ;
        RECT 14.000 425.600 14.600 427.800 ;
        RECT 17.200 427.600 18.800 427.800 ;
        RECT 20.400 428.200 21.200 428.400 ;
        RECT 20.400 427.600 22.000 428.200 ;
        RECT 23.400 427.600 26.000 428.400 ;
        RECT 26.800 427.600 29.400 428.400 ;
        RECT 31.600 428.200 32.400 428.400 ;
        RECT 30.800 427.600 32.400 428.200 ;
        RECT 34.800 427.600 36.800 428.400 ;
        RECT 37.400 428.200 38.800 429.000 ;
        RECT 39.600 428.800 40.400 430.400 ;
        RECT 41.200 428.800 42.000 430.400 ;
        RECT 42.800 430.300 43.600 430.400 ;
        RECT 44.800 430.300 45.400 431.800 ;
        RECT 42.800 429.700 45.400 430.300 ;
        RECT 42.800 429.600 43.600 429.700 ;
        RECT 44.800 428.400 45.400 429.700 ;
        RECT 46.000 428.800 46.800 430.400 ;
        RECT 50.600 428.400 51.200 431.800 ;
        RECT 52.200 429.800 52.800 431.800 ;
        RECT 55.600 431.600 56.200 435.000 ;
        RECT 59.800 432.800 60.600 439.800 ;
        RECT 69.000 438.400 69.800 439.800 ;
        RECT 68.400 437.600 69.800 438.400 ;
        RECT 69.000 432.800 69.800 437.600 ;
        RECT 73.200 435.000 74.000 439.000 ;
        RECT 59.800 432.200 61.400 432.800 ;
        RECT 55.600 431.000 59.400 431.600 ;
        RECT 51.800 429.000 52.800 429.800 ;
        RECT 21.200 427.200 22.000 427.600 ;
        RECT 12.200 425.400 13.000 425.600 ;
        RECT 6.000 424.200 6.800 425.000 ;
        RECT 10.200 424.800 13.000 425.400 ;
        RECT 14.000 424.800 14.800 425.600 ;
        RECT 10.200 424.200 10.800 424.800 ;
        RECT 15.600 424.200 16.400 425.000 ;
        RECT 5.400 423.600 6.800 424.200 ;
        RECT 5.400 422.200 6.600 423.600 ;
        RECT 10.000 422.200 10.800 424.200 ;
        RECT 14.400 423.600 16.400 424.200 ;
        RECT 14.400 422.200 15.200 423.600 ;
        RECT 18.800 422.200 19.600 427.000 ;
        RECT 20.600 426.200 24.200 426.600 ;
        RECT 25.200 426.200 25.800 427.600 ;
        RECT 27.000 426.200 27.600 427.600 ;
        RECT 30.800 427.200 31.600 427.600 ;
        RECT 36.200 427.000 36.800 427.600 ;
        RECT 37.800 427.800 38.800 428.200 ;
        RECT 37.800 427.200 42.000 427.800 ;
        RECT 42.800 427.600 45.400 428.400 ;
        RECT 47.600 428.200 48.400 428.400 ;
        RECT 46.800 427.600 48.400 428.200 ;
        RECT 50.600 427.600 51.600 428.400 ;
        RECT 36.200 426.600 37.000 427.000 ;
        RECT 28.600 426.200 32.200 426.600 ;
        RECT 20.400 426.000 24.400 426.200 ;
        RECT 20.400 422.200 21.200 426.000 ;
        RECT 23.600 422.200 24.400 426.000 ;
        RECT 25.200 422.200 26.000 426.200 ;
        RECT 26.800 422.200 27.600 426.200 ;
        RECT 28.400 426.000 32.400 426.200 ;
        RECT 36.200 426.000 37.800 426.600 ;
        RECT 28.400 422.200 29.200 426.000 ;
        RECT 31.600 422.200 32.400 426.000 ;
        RECT 37.000 423.000 37.800 426.000 ;
        RECT 41.400 425.000 42.000 427.200 ;
        RECT 43.000 426.200 43.600 427.600 ;
        RECT 46.800 427.200 47.600 427.600 ;
        RECT 44.600 426.200 48.200 426.600 ;
        RECT 50.600 426.200 51.200 427.600 ;
        RECT 52.200 427.400 52.800 429.000 ;
        RECT 53.800 429.600 54.800 430.400 ;
        RECT 53.800 428.800 54.600 429.600 ;
        RECT 55.600 428.800 56.400 430.400 ;
        RECT 57.200 428.800 58.000 430.400 ;
        RECT 58.800 429.000 59.400 431.000 ;
        RECT 58.800 428.200 60.200 429.000 ;
        RECT 60.800 428.400 61.400 432.200 ;
        RECT 68.200 432.200 69.800 432.800 ;
        RECT 62.000 430.300 62.800 431.200 ;
        RECT 63.600 430.300 64.400 430.400 ;
        RECT 62.000 429.700 64.400 430.300 ;
        RECT 62.000 429.600 62.800 429.700 ;
        RECT 63.600 429.600 64.400 429.700 ;
        RECT 66.800 429.600 67.600 431.200 ;
        RECT 68.200 428.400 68.800 432.200 ;
        RECT 73.400 431.600 74.000 435.000 ;
        RECT 77.400 432.400 78.200 439.800 ;
        RECT 78.800 433.600 79.600 434.400 ;
        RECT 79.000 432.400 79.600 433.600 ;
        RECT 82.000 433.600 82.800 434.400 ;
        RECT 82.000 432.400 82.600 433.600 ;
        RECT 83.400 432.400 84.200 439.800 ;
        RECT 77.400 431.800 78.400 432.400 ;
        RECT 79.000 431.800 80.400 432.400 ;
        RECT 70.200 431.000 74.000 431.600 ;
        RECT 70.200 429.000 70.800 431.000 ;
        RECT 60.800 428.300 62.800 428.400 ;
        RECT 65.200 428.300 66.000 428.400 ;
        RECT 58.800 427.800 59.800 428.200 ;
        RECT 52.200 426.800 54.800 427.400 ;
        RECT 41.200 423.000 42.000 425.000 ;
        RECT 42.800 422.200 43.600 426.200 ;
        RECT 44.400 426.000 48.400 426.200 ;
        RECT 44.400 422.200 45.200 426.000 ;
        RECT 47.600 422.200 48.400 426.000 ;
        RECT 50.600 425.600 51.600 426.200 ;
        RECT 50.800 422.200 51.600 425.600 ;
        RECT 54.000 422.200 54.800 426.800 ;
        RECT 55.600 427.200 59.800 427.800 ;
        RECT 60.800 427.700 66.000 428.300 ;
        RECT 60.800 427.600 62.800 427.700 ;
        RECT 65.200 427.600 66.000 427.700 ;
        RECT 66.800 427.600 68.800 428.400 ;
        RECT 69.400 428.200 70.800 429.000 ;
        RECT 71.600 428.800 72.400 430.400 ;
        RECT 73.200 428.800 74.000 430.400 ;
        RECT 76.400 428.800 77.200 430.400 ;
        RECT 77.800 430.300 78.400 431.800 ;
        RECT 79.600 431.600 80.400 431.800 ;
        RECT 81.200 431.800 82.600 432.400 ;
        RECT 81.200 431.600 82.000 431.800 ;
        RECT 83.200 431.600 85.200 432.400 ;
        RECT 81.300 430.300 81.900 431.600 ;
        RECT 77.800 429.700 81.900 430.300 ;
        RECT 77.800 428.400 78.400 429.700 ;
        RECT 83.200 428.400 83.800 431.600 ;
        RECT 87.600 431.200 88.400 439.800 ;
        RECT 91.800 435.800 93.000 439.800 ;
        RECT 96.400 435.800 97.200 439.800 ;
        RECT 100.800 436.400 101.600 439.800 ;
        RECT 100.800 435.800 102.800 436.400 ;
        RECT 92.400 435.000 93.200 435.800 ;
        RECT 96.600 435.200 97.200 435.800 ;
        RECT 95.800 434.600 99.400 435.200 ;
        RECT 102.000 435.000 102.800 435.800 ;
        RECT 95.800 434.400 96.600 434.600 ;
        RECT 98.600 434.400 99.400 434.600 ;
        RECT 91.600 433.200 93.000 434.000 ;
        RECT 92.400 432.200 93.000 433.200 ;
        RECT 94.600 433.000 96.800 433.600 ;
        RECT 94.600 432.800 95.400 433.000 ;
        RECT 92.400 431.600 94.800 432.200 ;
        RECT 87.600 430.600 91.800 431.200 ;
        RECT 84.400 428.800 85.200 430.400 ;
        RECT 55.600 425.000 56.200 427.200 ;
        RECT 60.800 427.000 61.400 427.600 ;
        RECT 60.600 426.600 61.400 427.000 ;
        RECT 59.800 426.000 61.400 426.600 ;
        RECT 68.200 427.000 68.800 427.600 ;
        RECT 69.800 427.800 70.800 428.200 ;
        RECT 74.800 428.200 75.600 428.400 ;
        RECT 69.800 427.200 74.000 427.800 ;
        RECT 74.800 427.600 76.400 428.200 ;
        RECT 77.800 427.600 80.400 428.400 ;
        RECT 81.200 427.600 83.800 428.400 ;
        RECT 86.000 428.200 86.800 428.400 ;
        RECT 85.200 427.600 86.800 428.200 ;
        RECT 75.600 427.200 76.400 427.600 ;
        RECT 68.200 426.600 69.000 427.000 ;
        RECT 68.200 426.000 69.800 426.600 ;
        RECT 55.600 423.000 56.400 425.000 ;
        RECT 59.800 423.000 60.600 426.000 ;
        RECT 69.000 423.000 69.800 426.000 ;
        RECT 73.400 425.000 74.000 427.200 ;
        RECT 75.000 426.200 78.600 426.600 ;
        RECT 79.600 426.200 80.200 427.600 ;
        RECT 81.400 426.200 82.000 427.600 ;
        RECT 85.200 427.200 86.000 427.600 ;
        RECT 87.600 427.200 88.400 430.600 ;
        RECT 91.000 430.400 91.800 430.600 ;
        RECT 94.200 430.300 94.800 431.600 ;
        RECT 96.200 431.800 96.800 433.000 ;
        RECT 97.400 433.000 98.200 433.200 ;
        RECT 102.000 433.000 102.800 433.200 ;
        RECT 97.400 432.400 102.800 433.000 ;
        RECT 96.200 431.400 101.000 431.800 ;
        RECT 105.200 431.400 106.000 439.800 ;
        RECT 115.400 432.800 116.200 439.800 ;
        RECT 119.600 435.000 120.400 439.000 ;
        RECT 96.200 431.200 106.000 431.400 ;
        RECT 114.600 432.200 116.200 432.800 ;
        RECT 100.200 431.000 106.000 431.200 ;
        RECT 100.400 430.800 106.000 431.000 ;
        RECT 95.600 430.300 96.400 430.400 ;
        RECT 89.400 429.800 90.200 430.000 ;
        RECT 89.400 429.200 93.200 429.800 ;
        RECT 94.100 429.700 96.400 430.300 ;
        RECT 92.400 429.000 93.200 429.200 ;
        RECT 94.200 428.400 94.800 429.700 ;
        RECT 95.600 429.600 96.400 429.700 ;
        RECT 98.800 430.200 99.600 430.400 ;
        RECT 106.800 430.300 107.600 430.400 ;
        RECT 113.200 430.300 114.000 431.200 ;
        RECT 98.800 429.600 103.800 430.200 ;
        RECT 106.800 429.700 114.000 430.300 ;
        RECT 106.800 429.600 107.600 429.700 ;
        RECT 113.200 429.600 114.000 429.700 ;
        RECT 103.000 429.400 103.800 429.600 ;
        RECT 101.400 428.400 102.200 428.600 ;
        RECT 114.600 428.400 115.200 432.200 ;
        RECT 119.800 431.600 120.400 435.000 ;
        RECT 121.200 432.400 122.000 439.800 ;
        RECT 124.400 432.800 125.200 439.800 ;
        RECT 129.200 432.800 130.000 439.800 ;
        RECT 121.200 431.800 123.800 432.400 ;
        RECT 124.400 431.800 125.400 432.800 ;
        RECT 116.600 431.000 120.400 431.600 ;
        RECT 116.600 429.000 117.200 431.000 ;
        RECT 94.200 427.800 105.200 428.400 ;
        RECT 94.600 427.600 95.400 427.800 ;
        RECT 98.800 427.600 99.600 427.800 ;
        RECT 87.600 426.600 91.400 427.200 ;
        RECT 83.000 426.200 86.600 426.600 ;
        RECT 73.200 423.000 74.000 425.000 ;
        RECT 74.800 426.000 78.800 426.200 ;
        RECT 74.800 422.200 75.600 426.000 ;
        RECT 78.000 422.200 78.800 426.000 ;
        RECT 79.600 422.200 80.400 426.200 ;
        RECT 81.200 422.200 82.000 426.200 ;
        RECT 82.800 426.000 86.800 426.200 ;
        RECT 82.800 422.200 83.600 426.000 ;
        RECT 86.000 422.200 86.800 426.000 ;
        RECT 87.600 422.200 88.400 426.600 ;
        RECT 90.600 426.400 91.400 426.600 ;
        RECT 100.400 425.600 101.000 427.800 ;
        RECT 103.600 427.600 105.200 427.800 ;
        RECT 108.400 428.300 109.200 428.400 ;
        RECT 113.200 428.300 115.200 428.400 ;
        RECT 108.400 427.700 115.200 428.300 ;
        RECT 115.800 428.200 117.200 429.000 ;
        RECT 118.000 428.800 118.800 430.400 ;
        RECT 119.600 428.800 120.400 430.400 ;
        RECT 121.200 429.600 122.200 430.400 ;
        RECT 121.400 428.800 122.200 429.600 ;
        RECT 123.200 429.800 123.800 431.800 ;
        RECT 123.200 429.000 124.200 429.800 ;
        RECT 108.400 427.600 109.200 427.700 ;
        RECT 113.200 427.600 115.200 427.700 ;
        RECT 114.600 427.000 115.200 427.600 ;
        RECT 116.200 427.800 117.200 428.200 ;
        RECT 116.200 427.200 120.400 427.800 ;
        RECT 123.200 427.400 123.800 429.000 ;
        RECT 124.800 428.400 125.400 431.800 ;
        RECT 129.000 431.800 130.000 432.800 ;
        RECT 132.400 432.400 133.200 439.800 ;
        RECT 130.600 431.800 133.200 432.400 ;
        RECT 134.000 432.400 134.800 439.800 ;
        RECT 137.200 432.800 138.000 439.800 ;
        RECT 134.000 431.800 136.600 432.400 ;
        RECT 137.200 431.800 138.200 432.800 ;
        RECT 129.000 428.400 129.600 431.800 ;
        RECT 130.600 429.800 131.200 431.800 ;
        RECT 130.200 429.000 131.200 429.800 ;
        RECT 124.400 428.300 125.400 428.400 ;
        RECT 126.000 428.300 126.800 428.400 ;
        RECT 124.400 427.700 126.800 428.300 ;
        RECT 124.400 427.600 125.400 427.700 ;
        RECT 126.000 427.600 126.800 427.700 ;
        RECT 129.000 427.600 130.000 428.400 ;
        RECT 98.600 425.400 99.400 425.600 ;
        RECT 92.400 424.200 93.200 425.000 ;
        RECT 96.600 424.800 99.400 425.400 ;
        RECT 100.400 424.800 101.200 425.600 ;
        RECT 96.600 424.200 97.200 424.800 ;
        RECT 102.000 424.200 102.800 425.000 ;
        RECT 91.800 423.600 93.200 424.200 ;
        RECT 91.800 422.200 93.000 423.600 ;
        RECT 96.400 422.200 97.200 424.200 ;
        RECT 100.800 423.600 102.800 424.200 ;
        RECT 100.800 422.200 101.600 423.600 ;
        RECT 105.200 422.200 106.000 427.000 ;
        RECT 114.600 426.600 115.400 427.000 ;
        RECT 114.600 426.000 116.200 426.600 ;
        RECT 115.400 423.000 116.200 426.000 ;
        RECT 119.800 425.000 120.400 427.200 ;
        RECT 119.600 423.000 120.400 425.000 ;
        RECT 121.200 426.800 123.800 427.400 ;
        RECT 121.200 422.200 122.000 426.800 ;
        RECT 124.800 426.200 125.400 427.600 ;
        RECT 124.400 425.600 125.400 426.200 ;
        RECT 129.000 426.200 129.600 427.600 ;
        RECT 130.600 427.400 131.200 429.000 ;
        RECT 132.200 429.600 133.200 430.400 ;
        RECT 134.000 429.600 135.000 430.400 ;
        RECT 132.200 428.800 133.000 429.600 ;
        RECT 134.200 428.800 135.000 429.600 ;
        RECT 136.000 429.800 136.600 431.800 ;
        RECT 136.000 429.000 137.000 429.800 ;
        RECT 136.000 427.400 136.600 429.000 ;
        RECT 137.600 428.400 138.200 431.800 ;
        RECT 137.200 427.600 138.200 428.400 ;
        RECT 130.600 426.800 133.200 427.400 ;
        RECT 129.000 425.600 130.000 426.200 ;
        RECT 124.400 422.200 125.200 425.600 ;
        RECT 129.200 422.200 130.000 425.600 ;
        RECT 132.400 422.200 133.200 426.800 ;
        RECT 134.000 426.800 136.600 427.400 ;
        RECT 134.000 422.200 134.800 426.800 ;
        RECT 137.600 426.200 138.200 427.600 ;
        RECT 137.200 425.600 138.200 426.200 ;
        RECT 140.400 431.200 141.200 439.800 ;
        RECT 144.600 435.800 145.800 439.800 ;
        RECT 149.200 435.800 150.000 439.800 ;
        RECT 153.600 436.400 154.400 439.800 ;
        RECT 153.600 435.800 155.600 436.400 ;
        RECT 145.200 435.000 146.000 435.800 ;
        RECT 149.400 435.200 150.000 435.800 ;
        RECT 148.600 434.600 152.200 435.200 ;
        RECT 154.800 435.000 155.600 435.800 ;
        RECT 148.600 434.400 149.400 434.600 ;
        RECT 151.400 434.400 152.200 434.600 ;
        RECT 144.400 433.200 145.800 434.000 ;
        RECT 145.200 432.200 145.800 433.200 ;
        RECT 147.400 433.000 149.600 433.600 ;
        RECT 147.400 432.800 148.200 433.000 ;
        RECT 145.200 431.600 147.600 432.200 ;
        RECT 140.400 430.600 144.600 431.200 ;
        RECT 140.400 427.200 141.200 430.600 ;
        RECT 143.800 430.400 144.600 430.600 ;
        RECT 142.200 429.800 143.000 430.000 ;
        RECT 142.200 429.200 146.000 429.800 ;
        RECT 145.200 429.000 146.000 429.200 ;
        RECT 147.000 428.400 147.600 431.600 ;
        RECT 149.000 431.800 149.600 433.000 ;
        RECT 150.200 433.000 151.000 433.200 ;
        RECT 154.800 433.000 155.600 433.200 ;
        RECT 150.200 432.400 155.600 433.000 ;
        RECT 149.000 431.400 153.800 431.800 ;
        RECT 158.000 431.400 158.800 439.800 ;
        RECT 160.400 433.600 161.200 434.400 ;
        RECT 160.400 432.400 161.000 433.600 ;
        RECT 161.800 432.400 162.600 439.800 ;
        RECT 168.200 434.400 169.000 439.800 ;
        RECT 172.400 435.000 173.200 439.000 ;
        RECT 166.800 433.600 167.600 434.400 ;
        RECT 168.200 433.600 170.000 434.400 ;
        RECT 166.800 432.400 167.400 433.600 ;
        RECT 168.200 432.400 169.000 433.600 ;
        RECT 159.600 431.800 161.000 432.400 ;
        RECT 161.600 431.800 162.600 432.400 ;
        RECT 166.000 431.800 167.400 432.400 ;
        RECT 168.000 431.800 169.000 432.400 ;
        RECT 159.600 431.600 160.400 431.800 ;
        RECT 149.000 431.200 158.800 431.400 ;
        RECT 153.000 431.000 158.800 431.200 ;
        RECT 153.200 430.800 158.800 431.000 ;
        RECT 151.600 430.200 152.400 430.400 ;
        RECT 159.600 430.300 160.400 430.400 ;
        RECT 161.600 430.300 162.200 431.800 ;
        RECT 166.000 431.600 166.800 431.800 ;
        RECT 151.600 429.600 156.600 430.200 ;
        RECT 159.600 429.700 162.200 430.300 ;
        RECT 159.600 429.600 160.400 429.700 ;
        RECT 155.800 429.400 156.600 429.600 ;
        RECT 154.200 428.400 155.000 428.600 ;
        RECT 161.600 428.400 162.200 429.700 ;
        RECT 162.800 428.800 163.600 430.400 ;
        RECT 168.000 428.400 168.600 431.800 ;
        RECT 172.400 431.600 173.000 435.000 ;
        RECT 176.600 432.800 177.400 439.800 ;
        RECT 184.200 438.400 185.000 439.800 ;
        RECT 184.200 437.600 186.000 438.400 ;
        RECT 182.800 433.600 183.600 434.400 ;
        RECT 176.600 432.200 178.200 432.800 ;
        RECT 182.800 432.400 183.400 433.600 ;
        RECT 184.200 432.400 185.000 437.600 ;
        RECT 177.200 431.600 178.200 432.200 ;
        RECT 182.000 431.800 183.400 432.400 ;
        RECT 184.000 431.800 185.000 432.400 ;
        RECT 188.400 432.400 189.200 439.800 ;
        RECT 191.600 432.800 192.400 439.800 ;
        RECT 188.400 431.800 191.000 432.400 ;
        RECT 191.600 431.800 192.600 432.800 ;
        RECT 182.000 431.600 182.800 431.800 ;
        RECT 172.400 431.000 176.200 431.600 ;
        RECT 169.200 428.800 170.000 430.400 ;
        RECT 172.400 428.800 173.200 430.400 ;
        RECT 174.000 428.800 174.800 430.400 ;
        RECT 175.600 429.000 176.200 431.000 ;
        RECT 147.000 427.800 158.000 428.400 ;
        RECT 147.400 427.600 148.200 427.800 ;
        RECT 153.200 427.600 154.000 427.800 ;
        RECT 156.400 427.600 158.000 427.800 ;
        RECT 159.600 427.600 162.200 428.400 ;
        RECT 164.400 428.200 165.200 428.400 ;
        RECT 163.600 427.600 165.200 428.200 ;
        RECT 166.000 427.600 168.600 428.400 ;
        RECT 170.800 428.200 171.600 428.400 ;
        RECT 170.000 427.600 171.600 428.200 ;
        RECT 175.600 428.200 177.000 429.000 ;
        RECT 177.600 428.400 178.200 431.600 ;
        RECT 178.800 429.600 179.600 431.200 ;
        RECT 184.000 428.400 184.600 431.800 ;
        RECT 185.200 428.800 186.000 430.400 ;
        RECT 188.400 429.600 189.400 430.400 ;
        RECT 188.600 428.800 189.400 429.600 ;
        RECT 190.400 429.800 191.000 431.800 ;
        RECT 190.400 429.000 191.400 429.800 ;
        RECT 175.600 427.800 176.600 428.200 ;
        RECT 140.400 426.600 144.200 427.200 ;
        RECT 137.200 422.200 138.000 425.600 ;
        RECT 140.400 422.200 141.200 426.600 ;
        RECT 143.400 426.400 144.200 426.600 ;
        RECT 153.200 425.600 153.800 427.600 ;
        RECT 151.400 425.400 152.200 425.600 ;
        RECT 145.200 424.200 146.000 425.000 ;
        RECT 149.400 424.800 152.200 425.400 ;
        RECT 153.200 424.800 154.000 425.600 ;
        RECT 149.400 424.200 150.000 424.800 ;
        RECT 154.800 424.200 155.600 425.000 ;
        RECT 144.600 423.600 146.000 424.200 ;
        RECT 144.600 422.200 145.800 423.600 ;
        RECT 149.200 422.200 150.000 424.200 ;
        RECT 153.600 423.600 155.600 424.200 ;
        RECT 153.600 422.200 154.400 423.600 ;
        RECT 158.000 422.200 158.800 427.000 ;
        RECT 159.800 426.200 160.400 427.600 ;
        RECT 163.600 427.200 164.400 427.600 ;
        RECT 161.400 426.200 165.000 426.600 ;
        RECT 166.200 426.200 166.800 427.600 ;
        RECT 170.000 427.200 170.800 427.600 ;
        RECT 172.400 427.200 176.600 427.800 ;
        RECT 177.600 427.600 179.600 428.400 ;
        RECT 182.000 427.600 184.600 428.400 ;
        RECT 186.800 428.200 187.600 428.400 ;
        RECT 186.000 427.600 187.600 428.200 ;
        RECT 167.800 426.200 171.400 426.600 ;
        RECT 159.600 422.200 160.400 426.200 ;
        RECT 161.200 426.000 165.200 426.200 ;
        RECT 161.200 422.200 162.000 426.000 ;
        RECT 164.400 422.200 165.200 426.000 ;
        RECT 166.000 422.200 166.800 426.200 ;
        RECT 167.600 426.000 171.600 426.200 ;
        RECT 167.600 422.200 168.400 426.000 ;
        RECT 170.800 422.200 171.600 426.000 ;
        RECT 172.400 425.000 173.000 427.200 ;
        RECT 177.600 427.000 178.200 427.600 ;
        RECT 177.400 426.600 178.200 427.000 ;
        RECT 176.600 426.000 178.200 426.600 ;
        RECT 182.200 426.200 182.800 427.600 ;
        RECT 186.000 427.200 186.800 427.600 ;
        RECT 190.400 427.400 191.000 429.000 ;
        RECT 192.000 428.400 192.600 431.800 ;
        RECT 191.600 427.600 192.600 428.400 ;
        RECT 188.400 426.800 191.000 427.400 ;
        RECT 183.800 426.200 187.400 426.600 ;
        RECT 172.400 423.000 173.200 425.000 ;
        RECT 176.600 423.000 177.400 426.000 ;
        RECT 182.000 422.200 182.800 426.200 ;
        RECT 183.600 426.000 187.600 426.200 ;
        RECT 183.600 422.200 184.400 426.000 ;
        RECT 186.800 422.200 187.600 426.000 ;
        RECT 188.400 422.200 189.200 426.800 ;
        RECT 192.000 426.200 192.600 427.600 ;
        RECT 191.600 425.600 192.600 426.200 ;
        RECT 194.800 431.200 195.600 439.800 ;
        RECT 199.000 435.800 200.200 439.800 ;
        RECT 203.600 435.800 204.400 439.800 ;
        RECT 208.000 436.400 208.800 439.800 ;
        RECT 208.000 435.800 210.000 436.400 ;
        RECT 199.600 435.000 200.400 435.800 ;
        RECT 203.800 435.200 204.400 435.800 ;
        RECT 203.000 434.600 206.600 435.200 ;
        RECT 209.200 435.000 210.000 435.800 ;
        RECT 203.000 434.400 203.800 434.600 ;
        RECT 205.800 434.400 206.600 434.600 ;
        RECT 198.800 433.200 200.200 434.000 ;
        RECT 199.600 432.200 200.200 433.200 ;
        RECT 201.800 433.000 204.000 433.600 ;
        RECT 201.800 432.800 202.600 433.000 ;
        RECT 199.600 431.600 202.000 432.200 ;
        RECT 194.800 430.600 199.000 431.200 ;
        RECT 194.800 427.200 195.600 430.600 ;
        RECT 198.200 430.400 199.000 430.600 ;
        RECT 201.400 430.400 202.000 431.600 ;
        RECT 203.400 431.800 204.000 433.000 ;
        RECT 204.600 433.000 205.400 433.200 ;
        RECT 209.200 433.000 210.000 433.200 ;
        RECT 204.600 432.400 210.000 433.000 ;
        RECT 203.400 431.400 208.200 431.800 ;
        RECT 212.400 431.400 213.200 439.800 ;
        RECT 216.600 432.600 217.400 439.800 ;
        RECT 215.600 431.800 217.400 432.600 ;
        RECT 203.400 431.200 213.200 431.400 ;
        RECT 207.400 431.000 213.200 431.200 ;
        RECT 207.600 430.800 213.200 431.000 ;
        RECT 196.600 429.800 197.400 430.000 ;
        RECT 196.600 429.200 200.400 429.800 ;
        RECT 201.200 429.600 202.000 430.400 ;
        RECT 206.000 430.200 206.800 430.400 ;
        RECT 206.000 429.600 211.000 430.200 ;
        RECT 199.600 429.000 200.400 429.200 ;
        RECT 201.400 428.400 202.000 429.600 ;
        RECT 210.200 429.400 211.000 429.600 ;
        RECT 208.600 428.400 209.400 428.600 ;
        RECT 215.800 428.400 216.400 431.800 ;
        RECT 217.200 429.600 218.000 431.200 ;
        RECT 201.400 427.800 212.400 428.400 ;
        RECT 201.800 427.600 202.600 427.800 ;
        RECT 194.800 426.600 198.600 427.200 ;
        RECT 191.600 422.200 192.400 425.600 ;
        RECT 194.800 422.200 195.600 426.600 ;
        RECT 197.800 426.400 198.600 426.600 ;
        RECT 207.600 425.600 208.200 427.800 ;
        RECT 210.800 427.600 212.400 427.800 ;
        RECT 215.600 427.600 216.400 428.400 ;
        RECT 205.800 425.400 206.600 425.600 ;
        RECT 199.600 424.200 200.400 425.000 ;
        RECT 203.800 424.800 206.600 425.400 ;
        RECT 207.600 424.800 208.400 425.600 ;
        RECT 203.800 424.200 204.400 424.800 ;
        RECT 209.200 424.200 210.000 425.000 ;
        RECT 199.000 423.600 200.400 424.200 ;
        RECT 199.000 422.200 200.200 423.600 ;
        RECT 203.600 422.200 204.400 424.200 ;
        RECT 208.000 423.600 210.000 424.200 ;
        RECT 208.000 422.200 208.800 423.600 ;
        RECT 212.400 422.200 213.200 427.000 ;
        RECT 214.000 424.800 214.800 426.400 ;
        RECT 215.800 424.400 216.400 427.600 ;
        RECT 217.200 426.300 218.000 426.400 ;
        RECT 218.800 426.300 219.600 439.800 ;
        RECT 222.000 431.800 222.800 439.800 ;
        RECT 223.600 432.400 224.400 439.800 ;
        RECT 226.800 432.400 227.600 439.800 ;
        RECT 229.000 432.400 229.800 439.800 ;
        RECT 223.600 431.800 227.600 432.400 ;
        RECT 228.400 431.800 229.800 432.400 ;
        RECT 222.200 430.400 222.800 431.800 ;
        RECT 228.400 431.600 229.200 431.800 ;
        RECT 226.000 430.400 226.800 430.800 ;
        RECT 228.400 430.400 229.000 431.600 ;
        RECT 233.200 431.200 234.000 439.800 ;
        RECT 235.400 432.600 236.200 439.800 ;
        RECT 235.400 431.800 237.200 432.600 ;
        RECT 241.200 432.000 242.000 439.800 ;
        RECT 244.400 435.200 245.200 439.800 ;
        RECT 230.000 430.800 234.000 431.200 ;
        RECT 229.800 430.600 234.000 430.800 ;
        RECT 222.000 429.800 224.400 430.400 ;
        RECT 226.000 429.800 227.600 430.400 ;
        RECT 222.000 429.600 222.800 429.800 ;
        RECT 220.400 428.300 221.200 428.400 ;
        RECT 220.400 427.700 222.700 428.300 ;
        RECT 220.400 427.600 221.200 427.700 ;
        RECT 222.100 426.400 222.700 427.700 ;
        RECT 217.200 425.700 219.600 426.300 ;
        RECT 217.200 425.600 218.000 425.700 ;
        RECT 215.600 422.200 216.400 424.400 ;
        RECT 218.800 422.200 219.600 425.700 ;
        RECT 220.400 424.800 221.200 426.400 ;
        RECT 222.000 425.600 222.800 426.400 ;
        RECT 223.800 426.200 224.400 429.800 ;
        RECT 226.800 429.600 227.600 429.800 ;
        RECT 228.400 429.600 229.200 430.400 ;
        RECT 229.800 430.000 230.600 430.600 ;
        RECT 225.200 427.600 226.000 429.200 ;
        RECT 222.200 424.800 223.000 425.600 ;
        RECT 223.600 422.200 224.400 426.200 ;
        RECT 228.400 426.200 229.000 429.600 ;
        RECT 229.800 427.000 230.400 430.000 ;
        RECT 234.800 429.600 235.600 431.200 ;
        RECT 231.200 428.400 232.000 429.200 ;
        RECT 236.400 428.400 237.000 431.800 ;
        RECT 241.000 431.200 242.000 432.000 ;
        RECT 242.600 434.600 245.200 435.200 ;
        RECT 242.600 433.000 243.200 434.600 ;
        RECT 247.600 434.400 248.400 439.800 ;
        RECT 250.800 437.000 251.600 439.800 ;
        RECT 252.400 437.000 253.200 439.800 ;
        RECT 254.000 437.000 254.800 439.800 ;
        RECT 249.000 434.400 253.200 435.200 ;
        RECT 245.800 433.600 248.400 434.400 ;
        RECT 255.600 433.600 256.400 439.800 ;
        RECT 258.800 435.000 259.600 439.800 ;
        RECT 262.000 435.000 262.800 439.800 ;
        RECT 263.600 437.000 264.400 439.800 ;
        RECT 265.200 437.000 266.000 439.800 ;
        RECT 268.400 435.200 269.200 439.800 ;
        RECT 271.600 436.400 272.400 439.800 ;
        RECT 271.600 435.800 272.600 436.400 ;
        RECT 272.000 435.200 272.600 435.800 ;
        RECT 267.200 434.400 271.400 435.200 ;
        RECT 272.000 434.600 274.000 435.200 ;
        RECT 258.800 433.600 261.400 434.400 ;
        RECT 262.000 433.800 267.800 434.400 ;
        RECT 270.800 434.000 271.400 434.400 ;
        RECT 250.800 433.000 251.600 433.200 ;
        RECT 242.600 432.400 251.600 433.000 ;
        RECT 254.000 433.000 254.800 433.200 ;
        RECT 262.000 433.000 262.600 433.800 ;
        RECT 268.400 433.200 269.800 433.800 ;
        RECT 270.800 433.200 272.400 434.000 ;
        RECT 254.000 432.400 262.600 433.000 ;
        RECT 263.600 433.000 269.800 433.200 ;
        RECT 263.600 432.600 269.000 433.000 ;
        RECT 263.600 432.400 264.400 432.600 ;
        RECT 231.400 427.600 232.400 428.400 ;
        RECT 236.400 427.600 237.200 428.400 ;
        RECT 229.800 426.400 232.200 427.000 ;
        RECT 228.400 422.200 229.200 426.200 ;
        RECT 231.600 424.200 232.200 426.400 ;
        RECT 233.200 426.300 234.000 426.400 ;
        RECT 234.800 426.300 235.600 426.400 ;
        RECT 233.200 425.700 235.600 426.300 ;
        RECT 233.200 424.800 234.000 425.700 ;
        RECT 234.800 425.600 235.600 425.700 ;
        RECT 236.400 424.400 237.000 427.600 ;
        RECT 241.000 426.800 241.800 431.200 ;
        RECT 242.600 430.600 243.200 432.400 ;
        RECT 242.400 430.000 243.200 430.600 ;
        RECT 249.200 430.000 272.600 430.600 ;
        RECT 242.400 428.000 243.000 430.000 ;
        RECT 249.200 429.400 250.000 430.000 ;
        RECT 260.400 429.600 261.200 430.000 ;
        RECT 266.800 429.600 267.600 430.000 ;
        RECT 270.000 429.600 270.800 430.000 ;
        RECT 271.800 429.800 272.600 430.000 ;
        RECT 243.600 428.600 247.400 429.400 ;
        RECT 242.400 427.400 243.600 428.000 ;
        RECT 238.000 424.800 238.800 426.400 ;
        RECT 241.000 426.000 242.000 426.800 ;
        RECT 231.600 422.200 232.400 424.200 ;
        RECT 236.400 422.200 237.200 424.400 ;
        RECT 241.200 422.200 242.000 426.000 ;
        RECT 242.800 422.200 243.600 427.400 ;
        RECT 246.600 427.400 247.400 428.600 ;
        RECT 246.600 426.800 248.400 427.400 ;
        RECT 247.600 426.200 248.400 426.800 ;
        RECT 252.400 426.400 253.200 429.200 ;
        RECT 255.600 428.600 258.800 429.400 ;
        RECT 262.600 428.600 264.600 429.400 ;
        RECT 273.200 429.000 274.000 434.600 ;
        RECT 279.600 431.600 280.400 434.400 ;
        RECT 255.200 427.800 256.000 428.000 ;
        RECT 255.200 427.200 259.600 427.800 ;
        RECT 258.800 427.000 259.600 427.200 ;
        RECT 260.400 426.800 261.200 428.400 ;
        RECT 247.600 425.400 250.000 426.200 ;
        RECT 252.400 425.600 253.400 426.400 ;
        RECT 256.400 425.600 258.000 426.400 ;
        RECT 258.800 426.200 259.600 426.400 ;
        RECT 262.600 426.200 263.400 428.600 ;
        RECT 265.200 428.200 274.000 429.000 ;
        RECT 268.600 426.800 271.600 427.600 ;
        RECT 268.600 426.200 269.400 426.800 ;
        RECT 258.800 425.600 263.400 426.200 ;
        RECT 249.200 422.200 250.000 425.400 ;
        RECT 266.800 425.400 269.400 426.200 ;
        RECT 250.800 422.200 251.600 425.000 ;
        RECT 252.400 422.200 253.200 425.000 ;
        RECT 254.000 422.200 254.800 425.000 ;
        RECT 255.600 422.200 256.400 425.000 ;
        RECT 258.800 422.200 259.600 425.000 ;
        RECT 262.000 422.200 262.800 425.000 ;
        RECT 263.600 422.200 264.400 425.000 ;
        RECT 265.200 422.200 266.000 425.000 ;
        RECT 266.800 422.200 267.600 425.400 ;
        RECT 273.200 422.200 274.000 428.200 ;
        RECT 281.200 426.200 282.000 439.800 ;
        RECT 286.000 431.200 286.800 439.800 ;
        RECT 289.200 431.200 290.000 439.800 ;
        RECT 292.400 431.200 293.200 439.800 ;
        RECT 295.600 431.200 296.400 439.800 ;
        RECT 301.400 438.400 302.200 439.800 ;
        RECT 300.400 437.600 302.200 438.400 ;
        RECT 301.400 432.400 302.200 437.600 ;
        RECT 307.400 438.400 308.200 439.800 ;
        RECT 307.400 437.600 309.200 438.400 ;
        RECT 302.800 433.600 303.600 434.400 ;
        RECT 303.000 432.400 303.600 433.600 ;
        RECT 306.000 433.600 306.800 434.400 ;
        RECT 306.000 432.400 306.600 433.600 ;
        RECT 307.400 432.400 308.200 437.600 ;
        RECT 301.400 431.800 302.400 432.400 ;
        RECT 303.000 431.800 304.400 432.400 ;
        RECT 284.400 430.400 286.800 431.200 ;
        RECT 287.800 430.400 290.000 431.200 ;
        RECT 291.000 430.400 293.200 431.200 ;
        RECT 294.600 430.400 296.400 431.200 ;
        RECT 282.800 426.800 283.600 428.400 ;
        RECT 284.400 427.600 285.200 430.400 ;
        RECT 287.800 429.000 288.600 430.400 ;
        RECT 291.000 429.000 291.800 430.400 ;
        RECT 294.600 429.000 295.400 430.400 ;
        RECT 286.000 428.200 288.600 429.000 ;
        RECT 289.400 428.200 291.800 429.000 ;
        RECT 292.800 428.200 295.400 429.000 ;
        RECT 296.200 428.200 298.000 429.000 ;
        RECT 300.400 428.800 301.200 430.400 ;
        RECT 301.800 428.400 302.400 431.800 ;
        RECT 303.600 431.600 304.400 431.800 ;
        RECT 305.200 431.800 306.600 432.400 ;
        RECT 307.200 431.800 308.200 432.400 ;
        RECT 305.200 431.600 306.000 431.800 ;
        RECT 307.200 428.400 307.800 431.800 ;
        RECT 308.400 428.800 309.200 430.400 ;
        RECT 287.800 427.600 288.600 428.200 ;
        RECT 291.000 427.600 291.800 428.200 ;
        RECT 294.600 427.600 295.400 428.200 ;
        RECT 297.200 427.600 298.000 428.200 ;
        RECT 298.800 428.200 299.600 428.400 ;
        RECT 298.800 427.600 300.400 428.200 ;
        RECT 301.800 427.600 304.400 428.400 ;
        RECT 305.200 427.600 307.800 428.400 ;
        RECT 310.000 428.300 310.800 428.400 ;
        RECT 311.600 428.300 312.400 439.800 ;
        RECT 317.400 432.600 318.200 439.800 ;
        RECT 316.400 431.800 318.200 432.600 ;
        RECT 320.200 432.600 321.000 439.800 ;
        RECT 320.200 431.800 322.000 432.600 ;
        RECT 313.200 430.300 314.000 430.400 ;
        RECT 316.600 430.300 317.200 431.800 ;
        RECT 313.200 429.700 317.200 430.300 ;
        RECT 313.200 429.600 314.000 429.700 ;
        RECT 316.600 428.400 317.200 429.700 ;
        RECT 318.000 429.600 318.800 431.200 ;
        RECT 319.600 429.600 320.400 431.200 ;
        RECT 310.000 428.200 312.400 428.300 ;
        RECT 309.200 427.700 312.400 428.200 ;
        RECT 309.200 427.600 310.800 427.700 ;
        RECT 284.400 426.800 286.800 427.600 ;
        RECT 287.800 426.800 290.000 427.600 ;
        RECT 291.000 426.800 293.200 427.600 ;
        RECT 294.600 426.800 296.400 427.600 ;
        RECT 299.600 427.200 300.400 427.600 ;
        RECT 280.200 425.600 282.000 426.200 ;
        RECT 280.200 422.200 281.000 425.600 ;
        RECT 286.000 422.200 286.800 426.800 ;
        RECT 289.200 422.200 290.000 426.800 ;
        RECT 292.400 422.200 293.200 426.800 ;
        RECT 295.600 422.200 296.400 426.800 ;
        RECT 299.000 426.200 302.600 426.600 ;
        RECT 303.600 426.200 304.200 427.600 ;
        RECT 305.400 426.200 306.000 427.600 ;
        RECT 309.200 427.200 310.000 427.600 ;
        RECT 307.000 426.200 310.600 426.600 ;
        RECT 298.800 426.000 302.800 426.200 ;
        RECT 298.800 422.200 299.600 426.000 ;
        RECT 302.000 422.200 302.800 426.000 ;
        RECT 303.600 422.200 304.400 426.200 ;
        RECT 305.200 422.200 306.000 426.200 ;
        RECT 306.800 426.000 310.800 426.200 ;
        RECT 306.800 422.200 307.600 426.000 ;
        RECT 310.000 422.200 310.800 426.000 ;
        RECT 311.600 422.200 312.400 427.700 ;
        RECT 316.400 427.600 317.200 428.400 ;
        RECT 313.200 424.800 314.000 426.400 ;
        RECT 314.800 424.800 315.600 426.400 ;
        RECT 316.600 424.200 317.200 427.600 ;
        RECT 316.400 422.200 317.200 424.200 ;
        RECT 321.200 428.400 321.800 431.800 ;
        RECT 321.200 427.600 322.000 428.400 ;
        RECT 324.400 428.300 325.200 428.400 ;
        RECT 322.900 427.700 325.200 428.300 ;
        RECT 321.200 426.400 321.800 427.600 ;
        RECT 322.900 426.400 323.500 427.700 ;
        RECT 324.400 426.800 325.200 427.700 ;
        RECT 326.000 428.300 326.800 439.800 ;
        RECT 327.600 431.600 328.400 433.200 ;
        RECT 329.200 428.300 330.000 428.400 ;
        RECT 326.000 427.700 330.000 428.300 ;
        RECT 321.200 425.600 322.000 426.400 ;
        RECT 321.200 424.200 321.800 425.600 ;
        RECT 322.800 424.800 323.600 426.400 ;
        RECT 326.000 426.200 326.800 427.700 ;
        RECT 329.200 426.800 330.000 427.700 ;
        RECT 330.800 426.200 331.600 439.800 ;
        RECT 332.400 431.600 333.200 433.200 ;
        RECT 332.400 428.300 333.200 428.400 ;
        RECT 334.000 428.300 334.800 428.400 ;
        RECT 332.400 427.700 334.800 428.300 ;
        RECT 332.400 427.600 333.200 427.700 ;
        RECT 334.000 426.800 334.800 427.700 ;
        RECT 335.600 428.300 336.400 439.800 ;
        RECT 339.800 432.400 340.600 439.800 ;
        RECT 341.200 433.600 342.800 434.400 ;
        RECT 341.400 432.400 342.000 433.600 ;
        RECT 339.800 431.800 340.800 432.400 ;
        RECT 341.400 431.800 342.800 432.400 ;
        RECT 346.200 431.800 348.200 439.800 ;
        RECT 340.200 430.400 340.800 431.800 ;
        RECT 342.000 431.600 342.800 431.800 ;
        RECT 337.200 430.300 338.000 430.400 ;
        RECT 338.800 430.300 339.600 430.400 ;
        RECT 337.200 429.700 339.600 430.300 ;
        RECT 337.200 429.600 338.000 429.700 ;
        RECT 338.800 428.800 339.600 429.700 ;
        RECT 340.200 429.600 341.200 430.400 ;
        RECT 340.200 428.400 340.800 429.600 ;
        RECT 337.200 428.300 338.000 428.400 ;
        RECT 335.600 428.200 338.000 428.300 ;
        RECT 335.600 427.700 338.800 428.200 ;
        RECT 326.000 425.600 327.800 426.200 ;
        RECT 330.800 425.600 332.600 426.200 ;
        RECT 321.200 422.200 322.000 424.200 ;
        RECT 327.000 422.200 327.800 425.600 ;
        RECT 331.800 422.200 332.600 425.600 ;
        RECT 335.600 422.200 336.400 427.700 ;
        RECT 337.200 427.600 338.800 427.700 ;
        RECT 340.200 427.600 342.800 428.400 ;
        RECT 343.600 427.600 344.400 429.200 ;
        RECT 345.200 428.800 346.000 430.400 ;
        RECT 347.000 428.400 347.600 431.800 ;
        RECT 348.400 428.800 349.200 430.400 ;
        RECT 346.800 428.200 347.600 428.400 ;
        RECT 350.000 428.200 350.800 428.400 ;
        RECT 345.200 427.600 347.600 428.200 ;
        RECT 349.200 427.600 350.800 428.200 ;
        RECT 338.000 427.200 338.800 427.600 ;
        RECT 337.400 426.200 341.000 426.600 ;
        RECT 342.000 426.200 342.600 427.600 ;
        RECT 345.200 426.200 345.800 427.600 ;
        RECT 349.200 427.200 350.000 427.600 ;
        RECT 347.000 426.200 350.600 426.600 ;
        RECT 337.200 426.000 341.200 426.200 ;
        RECT 337.200 422.200 338.000 426.000 ;
        RECT 340.400 422.200 341.200 426.000 ;
        RECT 342.000 422.200 342.800 426.200 ;
        RECT 343.600 422.800 344.400 426.200 ;
        RECT 345.200 423.400 346.000 426.200 ;
        RECT 346.800 426.000 350.800 426.200 ;
        RECT 346.800 422.800 347.600 426.000 ;
        RECT 343.600 422.200 347.600 422.800 ;
        RECT 350.000 422.200 350.800 426.000 ;
        RECT 351.600 422.200 352.400 439.800 ;
        RECT 357.400 431.800 359.400 439.800 ;
        RECT 362.800 435.800 363.600 439.800 ;
        RECT 363.000 435.600 363.600 435.800 ;
        RECT 366.000 435.800 366.800 439.800 ;
        RECT 366.000 435.600 366.600 435.800 ;
        RECT 363.000 435.000 366.600 435.600 ;
        RECT 363.000 432.400 363.600 435.000 ;
        RECT 364.400 432.800 365.200 434.400 ;
        RECT 354.800 427.600 355.600 429.200 ;
        RECT 356.400 428.800 357.200 430.400 ;
        RECT 358.200 428.400 358.800 431.800 ;
        RECT 362.800 431.600 363.600 432.400 ;
        RECT 359.600 428.800 360.400 430.400 ;
        RECT 363.000 428.400 363.600 431.600 ;
        RECT 367.600 430.800 368.400 432.400 ;
        RECT 365.200 429.600 366.800 430.400 ;
        RECT 358.000 428.200 358.800 428.400 ;
        RECT 361.200 428.200 362.000 428.400 ;
        RECT 356.400 427.600 358.800 428.200 ;
        RECT 360.400 427.600 362.000 428.200 ;
        RECT 363.000 428.200 364.600 428.400 ;
        RECT 363.000 427.800 364.800 428.200 ;
        RECT 353.200 424.800 354.000 426.400 ;
        RECT 356.400 426.200 357.000 427.600 ;
        RECT 360.400 427.200 361.200 427.600 ;
        RECT 358.200 426.200 361.800 426.600 ;
        RECT 354.800 422.800 355.600 426.200 ;
        RECT 356.400 423.400 357.200 426.200 ;
        RECT 358.000 426.000 362.000 426.200 ;
        RECT 358.000 422.800 358.800 426.000 ;
        RECT 354.800 422.200 358.800 422.800 ;
        RECT 361.200 422.200 362.000 426.000 ;
        RECT 364.000 422.200 364.800 427.800 ;
        RECT 369.200 422.200 370.000 439.800 ;
        RECT 372.400 435.800 373.200 439.800 ;
        RECT 372.600 435.600 373.200 435.800 ;
        RECT 375.600 435.800 376.400 439.800 ;
        RECT 375.600 435.600 376.200 435.800 ;
        RECT 372.600 435.000 376.200 435.600 ;
        RECT 372.600 432.400 373.200 435.000 ;
        RECT 374.000 432.800 374.800 434.400 ;
        RECT 372.400 431.600 373.200 432.400 ;
        RECT 372.600 428.400 373.200 431.600 ;
        RECT 377.200 430.800 378.000 432.400 ;
        RECT 378.800 431.800 379.600 439.800 ;
        RECT 382.000 435.800 382.800 439.800 ;
        RECT 378.800 430.400 379.400 431.800 ;
        RECT 382.000 431.600 382.600 435.800 ;
        RECT 380.200 431.000 382.600 431.600 ;
        RECT 385.200 431.800 386.000 439.800 ;
        RECT 388.400 432.400 389.200 439.800 ;
        RECT 390.000 433.600 391.600 434.400 ;
        RECT 390.800 432.400 391.400 433.600 ;
        RECT 392.200 432.400 393.000 439.800 ;
        RECT 387.000 431.800 389.200 432.400 ;
        RECT 390.000 431.800 391.400 432.400 ;
        RECT 392.000 431.800 393.000 432.400 ;
        RECT 374.800 429.600 376.400 430.400 ;
        RECT 378.800 429.600 379.600 430.400 ;
        RECT 372.600 428.200 374.200 428.400 ;
        RECT 372.600 427.800 374.400 428.200 ;
        RECT 370.800 424.800 371.600 426.400 ;
        RECT 373.600 422.200 374.400 427.800 ;
        RECT 378.800 426.200 379.400 429.600 ;
        RECT 380.200 427.600 380.800 431.000 ;
        RECT 382.000 429.600 382.800 430.400 ;
        RECT 385.200 429.600 385.800 431.800 ;
        RECT 387.000 431.200 387.600 431.800 ;
        RECT 390.000 431.600 390.800 431.800 ;
        RECT 386.400 430.400 387.600 431.200 ;
        RECT 382.000 428.800 382.600 429.600 ;
        RECT 381.600 428.200 382.600 428.800 ;
        RECT 381.600 428.000 382.400 428.200 ;
        RECT 383.600 427.600 384.400 429.200 ;
        RECT 380.000 427.400 380.800 427.600 ;
        RECT 380.000 427.000 383.000 427.400 ;
        RECT 380.000 426.800 384.200 427.000 ;
        RECT 382.400 426.400 384.200 426.800 ;
        RECT 383.600 426.200 384.200 426.400 ;
        RECT 378.800 425.200 380.200 426.200 ;
        RECT 379.400 424.400 380.200 425.200 ;
        RECT 378.800 423.600 380.200 424.400 ;
        RECT 379.400 422.200 380.200 423.600 ;
        RECT 383.600 422.200 384.400 426.200 ;
        RECT 385.200 422.200 386.000 429.600 ;
        RECT 387.000 427.400 387.600 430.400 ;
        RECT 388.400 428.800 389.200 430.400 ;
        RECT 392.000 428.400 392.600 431.800 ;
        RECT 393.200 428.800 394.000 430.400 ;
        RECT 390.000 427.600 392.600 428.400 ;
        RECT 394.800 428.200 395.600 428.400 ;
        RECT 394.000 427.600 395.600 428.200 ;
        RECT 387.000 426.800 389.200 427.400 ;
        RECT 388.400 422.200 389.200 426.800 ;
        RECT 390.200 426.200 390.800 427.600 ;
        RECT 394.000 427.200 394.800 427.600 ;
        RECT 396.400 426.800 397.200 428.400 ;
        RECT 391.800 426.200 395.400 426.600 ;
        RECT 398.000 426.200 398.800 439.800 ;
        RECT 407.600 436.400 408.400 439.800 ;
        RECT 407.400 435.800 408.400 436.400 ;
        RECT 407.400 435.200 408.000 435.800 ;
        RECT 410.800 435.200 411.600 439.800 ;
        RECT 414.000 437.000 414.800 439.800 ;
        RECT 415.600 437.000 416.400 439.800 ;
        RECT 406.000 434.600 408.000 435.200 ;
        RECT 399.600 431.600 400.400 433.200 ;
        RECT 406.000 429.000 406.800 434.600 ;
        RECT 408.600 434.400 412.800 435.200 ;
        RECT 417.200 435.000 418.000 439.800 ;
        RECT 420.400 435.000 421.200 439.800 ;
        RECT 408.600 434.000 409.200 434.400 ;
        RECT 407.600 433.200 409.200 434.000 ;
        RECT 412.200 433.800 418.000 434.400 ;
        RECT 410.200 433.200 411.600 433.800 ;
        RECT 410.200 433.000 416.400 433.200 ;
        RECT 411.000 432.600 416.400 433.000 ;
        RECT 415.600 432.400 416.400 432.600 ;
        RECT 417.400 433.000 418.000 433.800 ;
        RECT 418.600 433.600 421.200 434.400 ;
        RECT 423.600 433.600 424.400 439.800 ;
        RECT 425.200 437.000 426.000 439.800 ;
        RECT 426.800 437.000 427.600 439.800 ;
        RECT 428.400 437.000 429.200 439.800 ;
        RECT 426.800 434.400 431.000 435.200 ;
        RECT 431.600 434.400 432.400 439.800 ;
        RECT 434.800 435.200 435.600 439.800 ;
        RECT 434.800 434.600 437.400 435.200 ;
        RECT 431.600 433.600 434.200 434.400 ;
        RECT 425.200 433.000 426.000 433.200 ;
        RECT 417.400 432.400 426.000 433.000 ;
        RECT 428.400 433.000 429.200 433.200 ;
        RECT 436.800 433.000 437.400 434.600 ;
        RECT 428.400 432.400 437.400 433.000 ;
        RECT 436.800 430.600 437.400 432.400 ;
        RECT 438.000 432.000 438.800 439.800 ;
        RECT 438.000 431.200 439.000 432.000 ;
        RECT 407.400 430.000 430.800 430.600 ;
        RECT 436.800 430.000 437.600 430.600 ;
        RECT 407.400 429.800 408.400 430.000 ;
        RECT 407.600 429.600 408.400 429.800 ;
        RECT 412.400 429.600 413.200 430.000 ;
        RECT 430.000 429.400 430.800 430.000 ;
        RECT 406.000 428.200 414.800 429.000 ;
        RECT 415.400 428.600 417.400 429.400 ;
        RECT 421.200 428.600 424.400 429.400 ;
        RECT 390.000 422.200 390.800 426.200 ;
        RECT 391.600 426.000 395.600 426.200 ;
        RECT 391.600 422.200 392.400 426.000 ;
        RECT 394.800 422.200 395.600 426.000 ;
        RECT 398.000 425.600 399.800 426.200 ;
        RECT 399.000 422.200 399.800 425.600 ;
        RECT 406.000 422.200 406.800 428.200 ;
        RECT 408.400 426.800 411.400 427.600 ;
        RECT 410.600 426.200 411.400 426.800 ;
        RECT 416.600 426.200 417.400 428.600 ;
        RECT 418.800 426.800 419.600 428.400 ;
        RECT 424.000 427.800 424.800 428.000 ;
        RECT 420.400 427.200 424.800 427.800 ;
        RECT 420.400 427.000 421.200 427.200 ;
        RECT 426.800 426.400 427.600 429.200 ;
        RECT 432.600 428.600 436.400 429.400 ;
        RECT 432.600 427.400 433.400 428.600 ;
        RECT 437.000 428.000 437.600 430.000 ;
        RECT 420.400 426.200 421.200 426.400 ;
        RECT 410.600 425.400 413.200 426.200 ;
        RECT 416.600 425.600 421.200 426.200 ;
        RECT 422.000 425.600 423.600 426.400 ;
        RECT 426.600 425.600 427.600 426.400 ;
        RECT 431.600 426.800 433.400 427.400 ;
        RECT 436.400 427.400 437.600 428.000 ;
        RECT 431.600 426.200 432.400 426.800 ;
        RECT 412.400 422.200 413.200 425.400 ;
        RECT 430.000 425.400 432.400 426.200 ;
        RECT 414.000 422.200 414.800 425.000 ;
        RECT 415.600 422.200 416.400 425.000 ;
        RECT 417.200 422.200 418.000 425.000 ;
        RECT 420.400 422.200 421.200 425.000 ;
        RECT 423.600 422.200 424.400 425.000 ;
        RECT 425.200 422.200 426.000 425.000 ;
        RECT 426.800 422.200 427.600 425.000 ;
        RECT 428.400 422.200 429.200 425.000 ;
        RECT 430.000 422.200 430.800 425.400 ;
        RECT 436.400 422.200 437.200 427.400 ;
        RECT 438.200 426.800 439.000 431.200 ;
        RECT 438.000 426.000 439.000 426.800 ;
        RECT 438.000 422.200 438.800 426.000 ;
        RECT 441.200 422.200 442.000 439.800 ;
        RECT 446.000 432.800 446.800 439.800 ;
        RECT 445.800 431.800 446.800 432.800 ;
        RECT 449.200 432.400 450.000 439.800 ;
        RECT 447.400 431.800 450.000 432.400 ;
        RECT 445.800 428.400 446.400 431.800 ;
        RECT 447.400 429.800 448.000 431.800 ;
        RECT 452.400 431.200 453.200 439.800 ;
        RECT 455.600 431.200 456.400 439.800 ;
        RECT 458.800 431.200 459.600 439.800 ;
        RECT 462.000 431.200 462.800 439.800 ;
        RECT 466.800 436.400 467.600 439.800 ;
        RECT 466.600 435.800 467.600 436.400 ;
        RECT 466.600 435.200 467.200 435.800 ;
        RECT 470.000 435.200 470.800 439.800 ;
        RECT 473.200 437.000 474.000 439.800 ;
        RECT 474.800 437.000 475.600 439.800 ;
        RECT 450.800 430.400 453.200 431.200 ;
        RECT 454.200 430.400 456.400 431.200 ;
        RECT 457.400 430.400 459.600 431.200 ;
        RECT 461.000 430.400 462.800 431.200 ;
        RECT 465.200 434.600 467.200 435.200 ;
        RECT 447.000 429.000 448.000 429.800 ;
        RECT 445.800 428.300 446.800 428.400 ;
        RECT 442.900 427.700 446.800 428.300 ;
        RECT 442.900 426.400 443.500 427.700 ;
        RECT 445.800 427.600 446.800 427.700 ;
        RECT 442.800 424.800 443.600 426.400 ;
        RECT 445.800 426.200 446.400 427.600 ;
        RECT 447.400 427.400 448.000 429.000 ;
        RECT 449.000 429.600 450.000 430.400 ;
        RECT 449.000 428.800 449.800 429.600 ;
        RECT 450.800 427.600 451.600 430.400 ;
        RECT 454.200 429.000 455.000 430.400 ;
        RECT 457.400 429.000 458.200 430.400 ;
        RECT 461.000 429.000 461.800 430.400 ;
        RECT 465.200 429.000 466.000 434.600 ;
        RECT 467.800 434.400 472.000 435.200 ;
        RECT 476.400 435.000 477.200 439.800 ;
        RECT 479.600 435.000 480.400 439.800 ;
        RECT 467.800 434.000 468.400 434.400 ;
        RECT 466.800 433.200 468.400 434.000 ;
        RECT 471.400 433.800 477.200 434.400 ;
        RECT 469.400 433.200 470.800 433.800 ;
        RECT 469.400 433.000 475.600 433.200 ;
        RECT 470.200 432.600 475.600 433.000 ;
        RECT 474.800 432.400 475.600 432.600 ;
        RECT 476.600 433.000 477.200 433.800 ;
        RECT 477.800 433.600 480.400 434.400 ;
        RECT 482.800 433.600 483.600 439.800 ;
        RECT 484.400 437.000 485.200 439.800 ;
        RECT 486.000 437.000 486.800 439.800 ;
        RECT 487.600 437.000 488.400 439.800 ;
        RECT 486.000 434.400 490.200 435.200 ;
        RECT 490.800 434.400 491.600 439.800 ;
        RECT 494.000 435.200 494.800 439.800 ;
        RECT 494.000 434.600 496.600 435.200 ;
        RECT 490.800 433.600 493.400 434.400 ;
        RECT 484.400 433.000 485.200 433.200 ;
        RECT 476.600 432.400 485.200 433.000 ;
        RECT 487.600 433.000 488.400 433.200 ;
        RECT 496.000 433.000 496.600 434.600 ;
        RECT 487.600 432.400 496.600 433.000 ;
        RECT 496.000 430.600 496.600 432.400 ;
        RECT 497.200 432.300 498.000 439.800 ;
        RECT 501.200 433.600 502.000 434.400 ;
        RECT 501.200 432.400 501.800 433.600 ;
        RECT 502.600 432.400 503.400 439.800 ;
        RECT 500.400 432.300 501.800 432.400 ;
        RECT 497.200 431.800 501.800 432.300 ;
        RECT 502.400 431.800 503.400 432.400 ;
        RECT 497.200 431.700 501.200 431.800 ;
        RECT 497.200 431.200 498.200 431.700 ;
        RECT 500.400 431.600 501.200 431.700 ;
        RECT 466.600 430.000 490.000 430.600 ;
        RECT 496.000 430.000 496.800 430.600 ;
        RECT 466.600 429.800 467.400 430.000 ;
        RECT 468.400 429.600 469.200 430.000 ;
        RECT 471.600 429.600 472.400 430.000 ;
        RECT 489.200 429.400 490.000 430.000 ;
        RECT 452.400 428.200 455.000 429.000 ;
        RECT 455.800 428.200 458.200 429.000 ;
        RECT 459.200 428.200 461.800 429.000 ;
        RECT 462.600 428.200 464.400 429.000 ;
        RECT 454.200 427.600 455.000 428.200 ;
        RECT 457.400 427.600 458.200 428.200 ;
        RECT 461.000 427.600 461.800 428.200 ;
        RECT 463.600 427.600 464.400 428.200 ;
        RECT 465.200 428.200 474.000 429.000 ;
        RECT 474.600 428.600 476.600 429.400 ;
        RECT 480.400 428.600 483.600 429.400 ;
        RECT 447.400 426.800 450.000 427.400 ;
        RECT 450.800 426.800 453.200 427.600 ;
        RECT 454.200 426.800 456.400 427.600 ;
        RECT 457.400 426.800 459.600 427.600 ;
        RECT 461.000 426.800 462.800 427.600 ;
        RECT 445.800 425.600 446.800 426.200 ;
        RECT 446.000 422.200 446.800 425.600 ;
        RECT 449.200 422.200 450.000 426.800 ;
        RECT 452.400 422.200 453.200 426.800 ;
        RECT 455.600 422.200 456.400 426.800 ;
        RECT 458.800 422.200 459.600 426.800 ;
        RECT 462.000 422.200 462.800 426.800 ;
        RECT 465.200 422.200 466.000 428.200 ;
        RECT 467.600 426.800 470.600 427.600 ;
        RECT 469.800 426.200 470.600 426.800 ;
        RECT 475.800 426.200 476.600 428.600 ;
        RECT 478.000 426.800 478.800 428.400 ;
        RECT 483.200 427.800 484.000 428.000 ;
        RECT 479.600 427.200 484.000 427.800 ;
        RECT 479.600 427.000 480.400 427.200 ;
        RECT 486.000 426.400 486.800 429.200 ;
        RECT 491.800 428.600 495.600 429.400 ;
        RECT 491.800 427.400 492.600 428.600 ;
        RECT 496.200 428.000 496.800 430.000 ;
        RECT 479.600 426.200 480.400 426.400 ;
        RECT 469.800 425.400 472.400 426.200 ;
        RECT 475.800 425.600 480.400 426.200 ;
        RECT 481.200 425.600 482.800 426.400 ;
        RECT 485.800 425.600 486.800 426.400 ;
        RECT 490.800 426.800 492.600 427.400 ;
        RECT 495.600 427.400 496.800 428.000 ;
        RECT 490.800 426.200 491.600 426.800 ;
        RECT 471.600 422.200 472.400 425.400 ;
        RECT 489.200 425.400 491.600 426.200 ;
        RECT 473.200 422.200 474.000 425.000 ;
        RECT 474.800 422.200 475.600 425.000 ;
        RECT 476.400 422.200 477.200 425.000 ;
        RECT 479.600 422.200 480.400 425.000 ;
        RECT 482.800 422.200 483.600 425.000 ;
        RECT 484.400 422.200 485.200 425.000 ;
        RECT 486.000 422.200 486.800 425.000 ;
        RECT 487.600 422.200 488.400 425.000 ;
        RECT 489.200 422.200 490.000 425.400 ;
        RECT 495.600 422.200 496.400 427.400 ;
        RECT 497.400 426.800 498.200 431.200 ;
        RECT 498.800 430.300 499.600 430.400 ;
        RECT 502.400 430.300 503.000 431.800 ;
        RECT 508.400 431.200 509.200 439.800 ;
        RECT 511.600 431.200 512.400 439.800 ;
        RECT 514.800 431.200 515.600 439.800 ;
        RECT 518.000 431.200 518.800 439.800 ;
        RECT 522.800 432.800 523.600 439.800 ;
        RECT 522.600 431.800 523.600 432.800 ;
        RECT 526.000 432.400 526.800 439.800 ;
        RECT 530.200 438.400 531.000 439.800 ;
        RECT 529.200 437.600 531.000 438.400 ;
        RECT 524.200 431.800 526.800 432.400 ;
        RECT 530.200 432.400 531.000 437.600 ;
        RECT 531.600 433.600 532.400 434.400 ;
        RECT 531.800 432.400 532.400 433.600 ;
        RECT 530.200 431.800 531.200 432.400 ;
        RECT 531.800 431.800 533.200 432.400 ;
        RECT 508.400 430.400 510.200 431.200 ;
        RECT 511.600 430.400 513.800 431.200 ;
        RECT 514.800 430.400 517.000 431.200 ;
        RECT 518.000 430.400 520.400 431.200 ;
        RECT 498.800 429.700 503.000 430.300 ;
        RECT 498.800 429.600 499.600 429.700 ;
        RECT 502.400 428.400 503.000 429.700 ;
        RECT 503.600 428.800 504.400 430.400 ;
        RECT 509.400 429.000 510.200 430.400 ;
        RECT 513.000 429.000 513.800 430.400 ;
        RECT 516.200 429.000 517.000 430.400 ;
        RECT 500.400 427.600 503.000 428.400 ;
        RECT 505.200 428.200 506.000 428.400 ;
        RECT 504.400 427.600 506.000 428.200 ;
        RECT 506.800 428.200 508.600 429.000 ;
        RECT 509.400 428.200 512.000 429.000 ;
        RECT 513.000 428.200 515.400 429.000 ;
        RECT 516.200 428.200 518.800 429.000 ;
        RECT 506.800 427.600 507.600 428.200 ;
        RECT 509.400 427.600 510.200 428.200 ;
        RECT 513.000 427.600 513.800 428.200 ;
        RECT 516.200 427.600 517.000 428.200 ;
        RECT 519.600 427.600 520.400 430.400 ;
        RECT 497.200 426.300 498.200 426.800 ;
        RECT 498.800 426.300 499.600 426.400 ;
        RECT 497.200 425.700 499.600 426.300 ;
        RECT 500.600 426.200 501.200 427.600 ;
        RECT 504.400 427.200 505.200 427.600 ;
        RECT 508.400 426.800 510.200 427.600 ;
        RECT 511.600 426.800 513.800 427.600 ;
        RECT 514.800 426.800 517.000 427.600 ;
        RECT 518.000 426.800 520.400 427.600 ;
        RECT 522.600 428.400 523.200 431.800 ;
        RECT 524.200 429.800 524.800 431.800 ;
        RECT 523.800 429.000 524.800 429.800 ;
        RECT 522.600 427.600 523.600 428.400 ;
        RECT 502.200 426.200 505.800 426.600 ;
        RECT 497.200 422.200 498.000 425.700 ;
        RECT 498.800 425.600 499.600 425.700 ;
        RECT 500.400 422.200 501.200 426.200 ;
        RECT 502.000 426.000 506.000 426.200 ;
        RECT 502.000 422.200 502.800 426.000 ;
        RECT 505.200 422.200 506.000 426.000 ;
        RECT 508.400 422.200 509.200 426.800 ;
        RECT 511.600 422.200 512.400 426.800 ;
        RECT 514.800 422.200 515.600 426.800 ;
        RECT 518.000 422.200 518.800 426.800 ;
        RECT 522.600 426.200 523.200 427.600 ;
        RECT 524.200 427.400 524.800 429.000 ;
        RECT 525.800 429.600 526.800 430.400 ;
        RECT 525.800 428.800 526.600 429.600 ;
        RECT 529.200 428.800 530.000 430.400 ;
        RECT 530.600 428.400 531.200 431.800 ;
        RECT 532.400 431.600 533.200 431.800 ;
        RECT 534.000 431.200 534.800 439.800 ;
        RECT 538.200 438.400 539.000 439.800 ;
        RECT 538.200 437.600 539.600 438.400 ;
        RECT 538.200 432.400 539.000 437.600 ;
        RECT 540.400 432.400 541.200 439.800 ;
        RECT 543.600 432.800 544.400 439.800 ;
        RECT 549.000 438.400 549.800 439.800 ;
        RECT 549.000 437.600 550.800 438.400 ;
        RECT 547.600 433.600 548.400 434.400 ;
        RECT 538.200 431.800 539.600 432.400 ;
        RECT 540.400 431.800 543.000 432.400 ;
        RECT 543.600 431.800 544.600 432.800 ;
        RECT 547.600 432.400 548.200 433.600 ;
        RECT 549.000 432.400 549.800 437.600 ;
        RECT 534.000 430.800 538.000 431.200 ;
        RECT 534.000 430.600 538.200 430.800 ;
        RECT 537.400 430.000 538.200 430.600 ;
        RECT 539.000 430.400 539.600 431.800 ;
        RECT 536.000 428.400 536.800 429.200 ;
        RECT 527.600 428.200 528.400 428.400 ;
        RECT 527.600 427.600 529.200 428.200 ;
        RECT 530.600 427.600 533.200 428.400 ;
        RECT 535.600 427.600 536.600 428.400 ;
        RECT 524.200 426.800 526.800 427.400 ;
        RECT 528.400 427.200 529.200 427.600 ;
        RECT 522.600 425.600 523.600 426.200 ;
        RECT 522.800 422.200 523.600 425.600 ;
        RECT 526.000 422.200 526.800 426.800 ;
        RECT 527.800 426.200 531.400 426.600 ;
        RECT 532.400 426.200 533.000 427.600 ;
        RECT 537.600 427.000 538.200 430.000 ;
        RECT 538.800 429.600 539.600 430.400 ;
        RECT 540.400 429.600 541.400 430.400 ;
        RECT 535.800 426.400 538.200 427.000 ;
        RECT 527.600 426.000 531.600 426.200 ;
        RECT 527.600 422.200 528.400 426.000 ;
        RECT 530.800 422.200 531.600 426.000 ;
        RECT 532.400 422.200 533.200 426.200 ;
        RECT 534.000 424.800 534.800 426.400 ;
        RECT 535.800 424.200 536.400 426.400 ;
        RECT 539.000 426.200 539.600 429.600 ;
        RECT 540.600 428.800 541.400 429.600 ;
        RECT 542.400 429.800 543.000 431.800 ;
        RECT 542.400 429.000 543.400 429.800 ;
        RECT 542.400 427.400 543.000 429.000 ;
        RECT 544.000 428.400 544.600 431.800 ;
        RECT 546.800 431.800 548.200 432.400 ;
        RECT 548.800 431.800 549.800 432.400 ;
        RECT 554.800 432.000 555.600 439.800 ;
        RECT 558.000 435.200 558.800 439.800 ;
        RECT 546.800 431.600 547.600 431.800 ;
        RECT 548.800 428.400 549.400 431.800 ;
        RECT 554.600 431.200 555.600 432.000 ;
        RECT 556.200 434.600 558.800 435.200 ;
        RECT 556.200 433.000 556.800 434.600 ;
        RECT 561.200 434.400 562.000 439.800 ;
        RECT 564.400 437.000 565.200 439.800 ;
        RECT 566.000 437.000 566.800 439.800 ;
        RECT 567.600 437.000 568.400 439.800 ;
        RECT 562.600 434.400 566.800 435.200 ;
        RECT 559.400 433.600 562.000 434.400 ;
        RECT 569.200 433.600 570.000 439.800 ;
        RECT 572.400 435.000 573.200 439.800 ;
        RECT 575.600 435.000 576.400 439.800 ;
        RECT 577.200 437.000 578.000 439.800 ;
        RECT 578.800 437.000 579.600 439.800 ;
        RECT 582.000 435.200 582.800 439.800 ;
        RECT 585.200 436.400 586.000 439.800 ;
        RECT 585.200 435.800 586.200 436.400 ;
        RECT 585.600 435.200 586.200 435.800 ;
        RECT 580.800 434.400 585.000 435.200 ;
        RECT 585.600 434.600 587.600 435.200 ;
        RECT 572.400 433.600 575.000 434.400 ;
        RECT 575.600 433.800 581.400 434.400 ;
        RECT 584.400 434.000 585.000 434.400 ;
        RECT 564.400 433.000 565.200 433.200 ;
        RECT 556.200 432.400 565.200 433.000 ;
        RECT 567.600 433.000 568.400 433.200 ;
        RECT 575.600 433.000 576.200 433.800 ;
        RECT 582.000 433.200 583.400 433.800 ;
        RECT 584.400 433.200 586.000 434.000 ;
        RECT 567.600 432.400 576.200 433.000 ;
        RECT 577.200 433.000 583.400 433.200 ;
        RECT 577.200 432.600 582.600 433.000 ;
        RECT 577.200 432.400 578.000 432.600 ;
        RECT 550.000 428.800 550.800 430.400 ;
        RECT 543.600 427.600 544.600 428.400 ;
        RECT 546.800 427.600 549.400 428.400 ;
        RECT 551.600 428.200 552.400 428.400 ;
        RECT 550.800 427.600 552.400 428.200 ;
        RECT 535.600 422.200 536.400 424.200 ;
        RECT 538.800 422.200 539.600 426.200 ;
        RECT 540.400 426.800 543.000 427.400 ;
        RECT 540.400 422.200 541.200 426.800 ;
        RECT 544.000 426.200 544.600 427.600 ;
        RECT 547.000 426.200 547.600 427.600 ;
        RECT 550.800 427.200 551.600 427.600 ;
        RECT 554.600 426.800 555.400 431.200 ;
        RECT 556.200 430.600 556.800 432.400 ;
        RECT 580.200 431.800 581.000 432.000 ;
        RECT 583.600 431.800 584.400 432.400 ;
        RECT 557.400 431.200 584.400 431.800 ;
        RECT 557.400 431.000 558.200 431.200 ;
        RECT 556.000 430.000 556.800 430.600 ;
        RECT 556.000 428.000 556.600 430.000 ;
        RECT 557.200 428.600 561.000 429.400 ;
        RECT 556.000 427.400 557.200 428.000 ;
        RECT 548.600 426.200 552.200 426.600 ;
        RECT 543.600 425.600 544.600 426.200 ;
        RECT 543.600 422.200 544.400 425.600 ;
        RECT 546.800 422.200 547.600 426.200 ;
        RECT 548.400 426.000 552.400 426.200 ;
        RECT 554.600 426.000 555.600 426.800 ;
        RECT 548.400 422.200 549.200 426.000 ;
        RECT 551.600 422.200 552.400 426.000 ;
        RECT 554.800 422.200 555.600 426.000 ;
        RECT 556.400 422.200 557.200 427.400 ;
        RECT 560.200 427.400 561.000 428.600 ;
        RECT 560.200 426.800 562.000 427.400 ;
        RECT 561.200 426.200 562.000 426.800 ;
        RECT 566.000 426.400 566.800 429.200 ;
        RECT 569.200 428.600 572.400 429.400 ;
        RECT 576.200 428.600 578.200 429.400 ;
        RECT 586.800 429.000 587.600 434.600 ;
        RECT 593.200 432.400 594.000 439.800 ;
        RECT 596.400 432.800 597.200 439.800 ;
        RECT 593.200 431.800 595.800 432.400 ;
        RECT 593.200 429.600 594.200 430.400 ;
        RECT 568.800 427.800 569.600 428.000 ;
        RECT 568.800 427.200 573.200 427.800 ;
        RECT 572.400 427.000 573.200 427.200 ;
        RECT 574.000 426.800 574.800 428.400 ;
        RECT 561.200 425.400 563.600 426.200 ;
        RECT 566.000 425.600 567.000 426.400 ;
        RECT 570.000 425.600 571.600 426.400 ;
        RECT 572.400 426.200 573.200 426.400 ;
        RECT 576.200 426.200 577.000 428.600 ;
        RECT 578.800 428.200 587.600 429.000 ;
        RECT 593.400 428.800 594.200 429.600 ;
        RECT 595.200 429.800 595.800 431.800 ;
        RECT 596.400 431.600 597.400 432.800 ;
        RECT 601.200 432.000 602.000 439.800 ;
        RECT 604.400 435.200 605.200 439.800 ;
        RECT 595.200 429.000 596.200 429.800 ;
        RECT 582.200 426.800 585.200 427.600 ;
        RECT 582.200 426.200 583.000 426.800 ;
        RECT 572.400 425.600 577.000 426.200 ;
        RECT 562.800 422.200 563.600 425.400 ;
        RECT 580.400 425.400 583.000 426.200 ;
        RECT 564.400 422.200 565.200 425.000 ;
        RECT 566.000 422.200 566.800 425.000 ;
        RECT 567.600 422.200 568.400 425.000 ;
        RECT 569.200 422.200 570.000 425.000 ;
        RECT 572.400 422.200 573.200 425.000 ;
        RECT 575.600 422.200 576.400 425.000 ;
        RECT 577.200 422.200 578.000 425.000 ;
        RECT 578.800 422.200 579.600 425.000 ;
        RECT 580.400 422.200 581.200 425.400 ;
        RECT 586.800 422.200 587.600 428.200 ;
        RECT 595.200 427.400 595.800 429.000 ;
        RECT 596.800 428.400 597.400 431.600 ;
        RECT 596.400 427.600 597.400 428.400 ;
        RECT 593.200 426.800 595.800 427.400 ;
        RECT 593.200 422.200 594.000 426.800 ;
        RECT 596.800 426.200 597.400 427.600 ;
        RECT 596.400 425.600 597.400 426.200 ;
        RECT 601.000 431.200 602.000 432.000 ;
        RECT 602.600 434.600 605.200 435.200 ;
        RECT 602.600 433.000 603.200 434.600 ;
        RECT 607.600 434.400 608.400 439.800 ;
        RECT 610.800 437.000 611.600 439.800 ;
        RECT 612.400 437.000 613.200 439.800 ;
        RECT 614.000 437.000 614.800 439.800 ;
        RECT 609.000 434.400 613.200 435.200 ;
        RECT 605.800 433.600 608.400 434.400 ;
        RECT 615.600 433.600 616.400 439.800 ;
        RECT 618.800 435.000 619.600 439.800 ;
        RECT 622.000 435.000 622.800 439.800 ;
        RECT 623.600 437.000 624.400 439.800 ;
        RECT 625.200 437.000 626.000 439.800 ;
        RECT 628.400 435.200 629.200 439.800 ;
        RECT 631.600 436.400 632.400 439.800 ;
        RECT 631.600 435.800 632.600 436.400 ;
        RECT 632.000 435.200 632.600 435.800 ;
        RECT 627.200 434.400 631.400 435.200 ;
        RECT 632.000 434.600 634.000 435.200 ;
        RECT 618.800 433.600 621.400 434.400 ;
        RECT 622.000 433.800 627.800 434.400 ;
        RECT 630.800 434.000 631.400 434.400 ;
        RECT 610.800 433.000 611.600 433.200 ;
        RECT 602.600 432.400 611.600 433.000 ;
        RECT 614.000 433.000 614.800 433.200 ;
        RECT 622.000 433.000 622.600 433.800 ;
        RECT 628.400 433.200 629.800 433.800 ;
        RECT 630.800 433.200 632.400 434.000 ;
        RECT 614.000 432.400 622.600 433.000 ;
        RECT 623.600 433.000 629.800 433.200 ;
        RECT 623.600 432.600 629.000 433.000 ;
        RECT 623.600 432.400 624.400 432.600 ;
        RECT 601.000 426.800 601.800 431.200 ;
        RECT 602.600 430.600 603.200 432.400 ;
        RECT 602.400 430.000 603.200 430.600 ;
        RECT 609.200 430.000 632.600 430.600 ;
        RECT 602.400 428.000 603.000 430.000 ;
        RECT 609.200 429.400 610.000 430.000 ;
        RECT 626.800 429.600 627.600 430.000 ;
        RECT 631.600 429.800 632.600 430.000 ;
        RECT 631.600 429.600 632.400 429.800 ;
        RECT 603.600 428.600 607.400 429.400 ;
        RECT 602.400 427.400 603.600 428.000 ;
        RECT 601.000 426.000 602.000 426.800 ;
        RECT 596.400 422.200 597.200 425.600 ;
        RECT 601.200 422.200 602.000 426.000 ;
        RECT 602.800 422.200 603.600 427.400 ;
        RECT 606.600 427.400 607.400 428.600 ;
        RECT 606.600 426.800 608.400 427.400 ;
        RECT 607.600 426.200 608.400 426.800 ;
        RECT 612.400 426.400 613.200 429.200 ;
        RECT 615.600 428.600 618.800 429.400 ;
        RECT 622.600 428.600 624.600 429.400 ;
        RECT 633.200 429.000 634.000 434.600 ;
        RECT 636.400 431.200 637.200 439.800 ;
        RECT 639.600 431.200 640.400 439.800 ;
        RECT 642.800 431.200 643.600 439.800 ;
        RECT 646.000 431.200 646.800 439.800 ;
        RECT 650.800 432.000 651.600 439.800 ;
        RECT 654.000 435.200 654.800 439.800 ;
        RECT 615.200 427.800 616.000 428.000 ;
        RECT 615.200 427.200 619.600 427.800 ;
        RECT 618.800 427.000 619.600 427.200 ;
        RECT 620.400 426.800 621.200 428.400 ;
        RECT 607.600 425.400 610.000 426.200 ;
        RECT 612.400 425.600 613.400 426.400 ;
        RECT 616.400 425.600 618.000 426.400 ;
        RECT 618.800 426.200 619.600 426.400 ;
        RECT 622.600 426.200 623.400 428.600 ;
        RECT 625.200 428.200 634.000 429.000 ;
        RECT 628.600 426.800 631.600 427.600 ;
        RECT 628.600 426.200 629.400 426.800 ;
        RECT 618.800 425.600 623.400 426.200 ;
        RECT 609.200 422.200 610.000 425.400 ;
        RECT 626.800 425.400 629.400 426.200 ;
        RECT 610.800 422.200 611.600 425.000 ;
        RECT 612.400 422.200 613.200 425.000 ;
        RECT 614.000 422.200 614.800 425.000 ;
        RECT 615.600 422.200 616.400 425.000 ;
        RECT 618.800 422.200 619.600 425.000 ;
        RECT 622.000 422.200 622.800 425.000 ;
        RECT 623.600 422.200 624.400 425.000 ;
        RECT 625.200 422.200 626.000 425.000 ;
        RECT 626.800 422.200 627.600 425.400 ;
        RECT 633.200 422.200 634.000 428.200 ;
        RECT 634.800 430.400 637.200 431.200 ;
        RECT 638.200 430.400 640.400 431.200 ;
        RECT 641.400 430.400 643.600 431.200 ;
        RECT 645.000 430.400 646.800 431.200 ;
        RECT 650.600 431.200 651.600 432.000 ;
        RECT 652.200 434.600 654.800 435.200 ;
        RECT 652.200 433.000 652.800 434.600 ;
        RECT 657.200 434.400 658.000 439.800 ;
        RECT 660.400 437.000 661.200 439.800 ;
        RECT 662.000 437.000 662.800 439.800 ;
        RECT 663.600 437.000 664.400 439.800 ;
        RECT 658.600 434.400 662.800 435.200 ;
        RECT 655.400 433.600 658.000 434.400 ;
        RECT 665.200 433.600 666.000 439.800 ;
        RECT 668.400 435.000 669.200 439.800 ;
        RECT 671.600 435.000 672.400 439.800 ;
        RECT 673.200 437.000 674.000 439.800 ;
        RECT 674.800 437.000 675.600 439.800 ;
        RECT 678.000 435.200 678.800 439.800 ;
        RECT 681.200 436.400 682.000 439.800 ;
        RECT 681.200 435.800 682.200 436.400 ;
        RECT 681.600 435.200 682.200 435.800 ;
        RECT 676.800 434.400 681.000 435.200 ;
        RECT 681.600 434.600 683.600 435.200 ;
        RECT 668.400 433.600 671.000 434.400 ;
        RECT 671.600 433.800 677.400 434.400 ;
        RECT 680.400 434.000 681.000 434.400 ;
        RECT 660.400 433.000 661.200 433.200 ;
        RECT 652.200 432.400 661.200 433.000 ;
        RECT 663.600 433.000 664.400 433.200 ;
        RECT 671.600 433.000 672.200 433.800 ;
        RECT 678.000 433.200 679.400 433.800 ;
        RECT 680.400 433.200 682.000 434.000 ;
        RECT 663.600 432.400 672.200 433.000 ;
        RECT 673.200 433.000 679.400 433.200 ;
        RECT 673.200 432.600 678.600 433.000 ;
        RECT 673.200 432.400 674.000 432.600 ;
        RECT 634.800 427.600 635.600 430.400 ;
        RECT 638.200 429.000 639.000 430.400 ;
        RECT 641.400 429.000 642.200 430.400 ;
        RECT 645.000 429.000 645.800 430.400 ;
        RECT 636.400 428.200 639.000 429.000 ;
        RECT 639.800 428.200 642.200 429.000 ;
        RECT 643.200 428.200 645.800 429.000 ;
        RECT 646.600 428.200 648.400 429.000 ;
        RECT 638.200 427.600 639.000 428.200 ;
        RECT 641.400 427.600 642.200 428.200 ;
        RECT 645.000 427.600 645.800 428.200 ;
        RECT 647.600 427.600 648.400 428.200 ;
        RECT 634.800 426.800 637.200 427.600 ;
        RECT 638.200 426.800 640.400 427.600 ;
        RECT 641.400 426.800 643.600 427.600 ;
        RECT 645.000 426.800 646.800 427.600 ;
        RECT 636.400 422.200 637.200 426.800 ;
        RECT 639.600 422.200 640.400 426.800 ;
        RECT 642.800 422.200 643.600 426.800 ;
        RECT 646.000 422.200 646.800 426.800 ;
        RECT 650.600 426.800 651.400 431.200 ;
        RECT 652.200 430.600 652.800 432.400 ;
        RECT 652.000 430.000 652.800 430.600 ;
        RECT 658.800 430.000 682.200 430.600 ;
        RECT 652.000 428.000 652.600 430.000 ;
        RECT 658.800 429.400 659.600 430.000 ;
        RECT 676.400 429.600 677.200 430.000 ;
        RECT 681.400 429.800 682.200 430.000 ;
        RECT 653.200 428.600 657.000 429.400 ;
        RECT 652.000 427.400 653.200 428.000 ;
        RECT 650.600 426.000 651.600 426.800 ;
        RECT 650.800 422.200 651.600 426.000 ;
        RECT 652.400 422.200 653.200 427.400 ;
        RECT 656.200 427.400 657.000 428.600 ;
        RECT 656.200 426.800 658.000 427.400 ;
        RECT 657.200 426.200 658.000 426.800 ;
        RECT 662.000 426.400 662.800 429.200 ;
        RECT 665.200 428.600 668.400 429.400 ;
        RECT 672.200 428.600 674.200 429.400 ;
        RECT 682.800 429.000 683.600 434.600 ;
        RECT 664.800 427.800 665.600 428.000 ;
        RECT 664.800 427.200 669.200 427.800 ;
        RECT 668.400 427.000 669.200 427.200 ;
        RECT 670.000 426.800 670.800 428.400 ;
        RECT 657.200 425.400 659.600 426.200 ;
        RECT 662.000 425.600 663.000 426.400 ;
        RECT 666.000 425.600 667.600 426.400 ;
        RECT 668.400 426.200 669.200 426.400 ;
        RECT 672.200 426.200 673.000 428.600 ;
        RECT 674.800 428.200 683.600 429.000 ;
        RECT 678.200 426.800 681.200 427.600 ;
        RECT 678.200 426.200 679.000 426.800 ;
        RECT 668.400 425.600 673.000 426.200 ;
        RECT 658.800 422.200 659.600 425.400 ;
        RECT 676.400 425.400 679.000 426.200 ;
        RECT 660.400 422.200 661.200 425.000 ;
        RECT 662.000 422.200 662.800 425.000 ;
        RECT 663.600 422.200 664.400 425.000 ;
        RECT 665.200 422.200 666.000 425.000 ;
        RECT 668.400 422.200 669.200 425.000 ;
        RECT 671.600 422.200 672.400 425.000 ;
        RECT 673.200 422.200 674.000 425.000 ;
        RECT 674.800 422.200 675.600 425.000 ;
        RECT 676.400 422.200 677.200 425.400 ;
        RECT 682.800 422.200 683.600 428.200 ;
        RECT 1.200 415.000 2.000 419.800 ;
        RECT 5.600 418.400 6.400 419.800 ;
        RECT 4.400 417.800 6.400 418.400 ;
        RECT 10.000 417.800 10.800 419.800 ;
        RECT 14.200 418.400 15.400 419.800 ;
        RECT 14.000 417.800 15.400 418.400 ;
        RECT 4.400 417.000 5.200 417.800 ;
        RECT 10.000 417.200 10.600 417.800 ;
        RECT 6.000 416.400 6.800 417.200 ;
        RECT 7.800 416.600 10.600 417.200 ;
        RECT 14.000 417.000 14.800 417.800 ;
        RECT 7.800 416.400 8.600 416.600 ;
        RECT 2.000 414.200 3.600 414.400 ;
        RECT 6.200 414.200 6.800 416.400 ;
        RECT 15.800 415.400 16.600 415.600 ;
        RECT 18.800 415.400 19.600 419.800 ;
        RECT 20.400 416.000 21.200 419.800 ;
        RECT 23.600 416.000 24.400 419.800 ;
        RECT 20.400 415.800 24.400 416.000 ;
        RECT 25.200 415.800 26.000 419.800 ;
        RECT 30.600 416.000 31.400 419.000 ;
        RECT 34.800 417.000 35.600 419.000 ;
        RECT 20.600 415.400 24.200 415.800 ;
        RECT 15.800 414.800 19.600 415.400 ;
        RECT 11.800 414.200 12.600 414.400 ;
        RECT 2.000 413.600 13.000 414.200 ;
        RECT 5.000 413.400 5.800 413.600 ;
        RECT 3.400 412.400 4.200 412.600 ;
        RECT 12.400 412.400 13.000 413.600 ;
        RECT 14.000 412.800 14.800 413.000 ;
        RECT 3.400 411.800 8.400 412.400 ;
        RECT 7.600 411.600 8.400 411.800 ;
        RECT 12.400 411.600 13.200 412.400 ;
        RECT 14.000 412.200 17.800 412.800 ;
        RECT 17.000 412.000 17.800 412.200 ;
        RECT 1.200 411.000 6.800 411.200 ;
        RECT 1.200 410.800 7.000 411.000 ;
        RECT 1.200 410.600 11.000 410.800 ;
        RECT 1.200 402.200 2.000 410.600 ;
        RECT 6.200 410.200 11.000 410.600 ;
        RECT 4.400 409.000 9.800 409.600 ;
        RECT 4.400 408.800 5.200 409.000 ;
        RECT 9.000 408.800 9.800 409.000 ;
        RECT 10.400 409.000 11.000 410.200 ;
        RECT 12.400 410.400 13.000 411.600 ;
        RECT 15.400 411.400 16.200 411.600 ;
        RECT 18.800 411.400 19.600 414.800 ;
        RECT 21.200 414.400 22.000 414.800 ;
        RECT 25.200 414.400 25.800 415.800 ;
        RECT 29.800 415.400 31.400 416.000 ;
        RECT 29.800 415.000 30.600 415.400 ;
        RECT 29.800 414.400 30.400 415.000 ;
        RECT 35.000 414.800 35.600 417.000 ;
        RECT 20.400 413.800 22.000 414.400 ;
        RECT 20.400 413.600 21.200 413.800 ;
        RECT 23.400 413.600 26.000 414.400 ;
        RECT 26.800 414.300 27.600 414.400 ;
        RECT 28.400 414.300 30.400 414.400 ;
        RECT 26.800 413.700 30.400 414.300 ;
        RECT 31.400 414.200 35.600 414.800 ;
        RECT 36.400 415.200 37.200 419.800 ;
        RECT 39.600 416.400 40.400 419.800 ;
        RECT 39.600 415.800 40.600 416.400 ;
        RECT 42.800 416.000 43.600 419.800 ;
        RECT 46.000 416.000 46.800 419.800 ;
        RECT 42.800 415.800 46.800 416.000 ;
        RECT 47.600 415.800 48.400 419.800 ;
        RECT 49.200 415.800 50.000 419.800 ;
        RECT 50.800 416.000 51.600 419.800 ;
        RECT 54.000 416.000 54.800 419.800 ;
        RECT 59.400 416.000 60.200 419.000 ;
        RECT 63.600 417.000 64.400 419.000 ;
        RECT 50.800 415.800 54.800 416.000 ;
        RECT 36.400 414.600 39.000 415.200 ;
        RECT 31.400 413.800 32.400 414.200 ;
        RECT 26.800 413.600 27.600 413.700 ;
        RECT 28.400 413.600 30.400 413.700 ;
        RECT 22.000 411.600 22.800 413.200 ;
        RECT 23.400 412.400 24.000 413.600 ;
        RECT 23.400 411.600 24.400 412.400 ;
        RECT 26.800 412.300 27.600 412.400 ;
        RECT 28.400 412.300 29.200 412.400 ;
        RECT 26.800 411.700 29.200 412.300 ;
        RECT 26.800 411.600 27.600 411.700 ;
        RECT 15.400 410.800 19.600 411.400 ;
        RECT 12.400 409.800 14.800 410.400 ;
        RECT 11.800 409.000 12.600 409.200 ;
        RECT 10.400 408.400 12.600 409.000 ;
        RECT 14.200 408.800 14.800 409.800 ;
        RECT 14.200 408.000 15.600 408.800 ;
        RECT 7.800 407.400 8.600 407.600 ;
        RECT 10.600 407.400 11.400 407.600 ;
        RECT 4.400 406.200 5.200 407.000 ;
        RECT 7.800 406.800 11.400 407.400 ;
        RECT 10.000 406.200 10.600 406.800 ;
        RECT 14.000 406.200 14.800 407.000 ;
        RECT 4.400 405.600 6.400 406.200 ;
        RECT 5.600 402.200 6.400 405.600 ;
        RECT 10.000 402.200 10.800 406.200 ;
        RECT 14.200 402.200 15.400 406.200 ;
        RECT 18.800 402.200 19.600 410.800 ;
        RECT 23.400 410.200 24.000 411.600 ;
        RECT 28.400 410.800 29.200 411.700 ;
        RECT 25.200 410.200 26.000 410.400 ;
        RECT 23.000 409.600 24.000 410.200 ;
        RECT 24.600 409.600 26.000 410.200 ;
        RECT 29.800 409.800 30.400 413.600 ;
        RECT 31.000 413.000 32.400 413.800 ;
        RECT 31.800 411.000 32.400 413.000 ;
        RECT 33.200 411.600 34.000 413.200 ;
        RECT 34.800 411.600 35.600 413.200 ;
        RECT 36.600 412.400 37.400 413.200 ;
        RECT 36.400 411.600 37.400 412.400 ;
        RECT 38.400 413.000 39.000 414.600 ;
        RECT 40.000 414.400 40.600 415.800 ;
        RECT 43.000 415.400 46.600 415.800 ;
        RECT 43.600 414.400 44.400 414.800 ;
        RECT 47.600 414.400 48.200 415.800 ;
        RECT 49.400 414.400 50.000 415.800 ;
        RECT 51.000 415.400 54.600 415.800 ;
        RECT 58.600 415.400 60.200 416.000 ;
        RECT 58.600 415.000 59.400 415.400 ;
        RECT 53.200 414.400 54.000 414.800 ;
        RECT 58.600 414.400 59.200 415.000 ;
        RECT 63.800 414.800 64.400 417.000 ;
        RECT 65.200 415.600 66.000 417.200 ;
        RECT 39.600 414.300 40.600 414.400 ;
        RECT 39.600 413.700 41.900 414.300 ;
        RECT 39.600 413.600 40.600 413.700 ;
        RECT 38.400 412.200 39.400 413.000 ;
        RECT 31.800 410.400 35.600 411.000 ;
        RECT 23.000 402.200 23.800 409.600 ;
        RECT 24.600 408.400 25.200 409.600 ;
        RECT 29.800 409.200 31.400 409.800 ;
        RECT 24.400 407.600 25.200 408.400 ;
        RECT 30.600 402.200 31.400 409.200 ;
        RECT 35.000 407.000 35.600 410.400 ;
        RECT 38.400 410.200 39.000 412.200 ;
        RECT 40.000 410.200 40.600 413.600 ;
        RECT 41.300 412.300 41.900 413.700 ;
        RECT 42.800 413.800 44.400 414.400 ;
        RECT 42.800 413.600 43.600 413.800 ;
        RECT 45.800 413.600 48.400 414.400 ;
        RECT 49.200 413.600 51.800 414.400 ;
        RECT 53.200 414.300 54.800 414.400 ;
        RECT 55.600 414.300 56.400 414.400 ;
        RECT 53.200 413.800 56.400 414.300 ;
        RECT 54.000 413.700 56.400 413.800 ;
        RECT 54.000 413.600 54.800 413.700 ;
        RECT 55.600 413.600 56.400 413.700 ;
        RECT 57.200 413.600 59.200 414.400 ;
        RECT 60.200 414.200 64.400 414.800 ;
        RECT 60.200 413.800 61.200 414.200 ;
        RECT 44.400 412.300 45.200 413.200 ;
        RECT 41.300 411.700 45.200 412.300 ;
        RECT 44.400 411.600 45.200 411.700 ;
        RECT 45.800 412.300 46.400 413.600 ;
        RECT 45.800 411.700 49.900 412.300 ;
        RECT 45.800 410.200 46.400 411.700 ;
        RECT 49.300 410.400 49.900 411.700 ;
        RECT 47.600 410.200 48.400 410.400 ;
        RECT 34.800 403.000 35.600 407.000 ;
        RECT 36.400 409.600 39.000 410.200 ;
        RECT 36.400 402.200 37.200 409.600 ;
        RECT 39.600 409.200 40.600 410.200 ;
        RECT 45.400 409.600 46.400 410.200 ;
        RECT 47.000 409.600 48.400 410.200 ;
        RECT 49.200 410.200 50.000 410.400 ;
        RECT 51.200 410.200 51.800 413.600 ;
        RECT 52.400 411.600 53.200 413.200 ;
        RECT 58.600 412.400 59.200 413.600 ;
        RECT 59.800 413.000 61.200 413.800 ;
        RECT 57.200 410.800 58.000 412.400 ;
        RECT 58.600 411.600 59.600 412.400 ;
        RECT 49.200 409.600 50.600 410.200 ;
        RECT 51.200 409.600 52.200 410.200 ;
        RECT 39.600 402.200 40.400 409.200 ;
        RECT 45.400 402.200 46.200 409.600 ;
        RECT 47.000 408.400 47.600 409.600 ;
        RECT 46.800 407.600 47.600 408.400 ;
        RECT 50.000 408.400 50.600 409.600 ;
        RECT 50.000 407.600 50.800 408.400 ;
        RECT 51.400 402.200 52.200 409.600 ;
        RECT 58.600 409.800 59.200 411.600 ;
        RECT 60.600 411.000 61.200 413.000 ;
        RECT 62.000 411.600 62.800 413.200 ;
        RECT 63.600 411.600 64.400 413.200 ;
        RECT 60.600 410.400 64.400 411.000 ;
        RECT 58.600 409.200 60.200 409.800 ;
        RECT 59.400 402.200 60.200 409.200 ;
        RECT 63.800 407.000 64.400 410.400 ;
        RECT 63.600 403.000 64.400 407.000 ;
        RECT 66.800 402.200 67.600 419.800 ;
        RECT 68.400 415.400 69.200 419.800 ;
        RECT 72.600 418.400 73.800 419.800 ;
        RECT 72.600 417.800 74.000 418.400 ;
        RECT 77.200 417.800 78.000 419.800 ;
        RECT 81.600 418.400 82.400 419.800 ;
        RECT 81.600 417.800 83.600 418.400 ;
        RECT 73.200 417.000 74.000 417.800 ;
        RECT 77.400 417.200 78.000 417.800 ;
        RECT 77.400 416.600 80.200 417.200 ;
        RECT 79.400 416.400 80.200 416.600 ;
        RECT 81.200 416.400 82.000 417.200 ;
        RECT 82.800 417.000 83.600 417.800 ;
        RECT 71.400 415.400 72.200 415.600 ;
        RECT 68.400 414.800 72.200 415.400 ;
        RECT 68.400 411.400 69.200 414.800 ;
        RECT 75.400 414.200 76.200 414.400 ;
        RECT 81.200 414.200 81.800 416.400 ;
        RECT 86.000 415.000 86.800 419.800 ;
        RECT 87.600 415.600 88.400 417.200 ;
        RECT 84.400 414.200 86.000 414.400 ;
        RECT 75.000 413.600 86.000 414.200 ;
        RECT 73.200 412.800 74.000 413.000 ;
        RECT 70.200 412.200 74.000 412.800 ;
        RECT 70.200 412.000 71.000 412.200 ;
        RECT 71.800 411.400 72.600 411.600 ;
        RECT 68.400 410.800 72.600 411.400 ;
        RECT 68.400 402.200 69.200 410.800 ;
        RECT 75.000 410.400 75.600 413.600 ;
        RECT 82.200 413.400 83.000 413.600 ;
        RECT 83.800 412.400 84.600 412.600 ;
        RECT 79.600 411.800 84.600 412.400 ;
        RECT 79.600 411.600 80.400 411.800 ;
        RECT 81.200 411.000 86.800 411.200 ;
        RECT 81.000 410.800 86.800 411.000 ;
        RECT 73.200 409.800 75.600 410.400 ;
        RECT 77.000 410.600 86.800 410.800 ;
        RECT 77.000 410.200 81.800 410.600 ;
        RECT 73.200 408.800 73.800 409.800 ;
        RECT 72.400 408.000 73.800 408.800 ;
        RECT 75.400 409.000 76.200 409.200 ;
        RECT 77.000 409.000 77.600 410.200 ;
        RECT 75.400 408.400 77.600 409.000 ;
        RECT 78.200 409.000 83.600 409.600 ;
        RECT 78.200 408.800 79.000 409.000 ;
        RECT 82.800 408.800 83.600 409.000 ;
        RECT 76.600 407.400 77.400 407.600 ;
        RECT 79.400 407.400 80.200 407.600 ;
        RECT 73.200 406.200 74.000 407.000 ;
        RECT 76.600 406.800 80.200 407.400 ;
        RECT 77.400 406.200 78.000 406.800 ;
        RECT 82.800 406.200 83.600 407.000 ;
        RECT 72.600 402.200 73.800 406.200 ;
        RECT 77.200 402.200 78.000 406.200 ;
        RECT 81.600 405.600 83.600 406.200 ;
        RECT 81.600 402.200 82.400 405.600 ;
        RECT 86.000 402.200 86.800 410.600 ;
        RECT 89.200 402.200 90.000 419.800 ;
        RECT 94.400 414.200 95.200 419.800 ;
        RECT 97.200 415.000 98.000 419.800 ;
        RECT 101.600 418.400 102.400 419.800 ;
        RECT 100.400 417.800 102.400 418.400 ;
        RECT 106.000 417.800 106.800 419.800 ;
        RECT 110.200 418.400 111.400 419.800 ;
        RECT 110.000 417.800 111.400 418.400 ;
        RECT 100.400 417.000 101.200 417.800 ;
        RECT 106.000 417.200 106.600 417.800 ;
        RECT 102.000 416.400 102.800 417.200 ;
        RECT 103.800 416.600 106.600 417.200 ;
        RECT 110.000 417.000 110.800 417.800 ;
        RECT 103.800 416.400 104.600 416.600 ;
        RECT 98.000 414.200 99.600 414.400 ;
        RECT 102.200 414.200 102.800 416.400 ;
        RECT 111.800 415.400 112.600 415.600 ;
        RECT 114.800 415.400 115.600 419.800 ;
        RECT 121.200 415.800 122.000 419.800 ;
        RECT 122.800 416.000 123.600 419.800 ;
        RECT 126.000 416.000 126.800 419.800 ;
        RECT 122.800 415.800 126.800 416.000 ;
        RECT 111.800 414.800 115.600 415.400 ;
        RECT 107.800 414.200 108.600 414.400 ;
        RECT 94.400 413.800 96.200 414.200 ;
        RECT 94.600 413.600 96.200 413.800 ;
        RECT 98.000 413.600 109.000 414.200 ;
        RECT 92.400 411.600 94.000 412.400 ;
        RECT 90.800 409.600 91.600 411.200 ;
        RECT 95.600 410.400 96.200 413.600 ;
        RECT 101.000 413.400 101.800 413.600 ;
        RECT 99.400 412.400 100.200 412.600 ;
        RECT 99.400 411.800 104.400 412.400 ;
        RECT 103.600 411.600 104.400 411.800 ;
        RECT 97.200 411.000 102.800 411.200 ;
        RECT 97.200 410.800 103.000 411.000 ;
        RECT 97.200 410.600 107.000 410.800 ;
        RECT 95.600 409.600 96.400 410.400 ;
        RECT 94.000 407.600 94.800 409.200 ;
        RECT 95.600 407.000 96.200 409.600 ;
        RECT 92.600 406.400 96.200 407.000 ;
        RECT 92.600 406.200 93.200 406.400 ;
        RECT 92.400 402.200 93.200 406.200 ;
        RECT 95.600 406.200 96.200 406.400 ;
        RECT 95.600 402.200 96.400 406.200 ;
        RECT 97.200 402.200 98.000 410.600 ;
        RECT 102.200 410.200 107.000 410.600 ;
        RECT 100.400 409.000 105.800 409.600 ;
        RECT 100.400 408.800 101.200 409.000 ;
        RECT 105.000 408.800 105.800 409.000 ;
        RECT 106.400 409.000 107.000 410.200 ;
        RECT 108.400 410.400 109.000 413.600 ;
        RECT 110.000 412.800 110.800 413.000 ;
        RECT 110.000 412.200 113.800 412.800 ;
        RECT 113.000 412.000 113.800 412.200 ;
        RECT 111.400 411.400 112.200 411.600 ;
        RECT 114.800 411.400 115.600 414.800 ;
        RECT 121.400 414.400 122.000 415.800 ;
        RECT 123.000 415.400 126.600 415.800 ;
        RECT 125.200 414.400 126.000 414.800 ;
        RECT 116.400 414.300 117.200 414.400 ;
        RECT 121.200 414.300 123.800 414.400 ;
        RECT 116.400 413.700 123.800 414.300 ;
        RECT 125.200 413.800 126.800 414.400 ;
        RECT 131.200 414.200 132.000 419.800 ;
        RECT 134.000 417.000 134.800 419.000 ;
        RECT 134.000 414.800 134.600 417.000 ;
        RECT 138.200 416.400 139.000 419.000 ;
        RECT 137.200 416.000 139.000 416.400 ;
        RECT 137.200 415.600 139.800 416.000 ;
        RECT 138.200 415.400 139.800 415.600 ;
        RECT 139.000 415.000 139.800 415.400 ;
        RECT 134.000 414.200 138.200 414.800 ;
        RECT 131.200 413.800 133.000 414.200 ;
        RECT 116.400 413.600 117.200 413.700 ;
        RECT 121.200 413.600 123.800 413.700 ;
        RECT 126.000 413.600 126.800 413.800 ;
        RECT 131.400 413.600 133.000 413.800 ;
        RECT 111.400 410.800 115.600 411.400 ;
        RECT 108.400 409.800 110.800 410.400 ;
        RECT 107.800 409.000 108.600 409.200 ;
        RECT 106.400 408.400 108.600 409.000 ;
        RECT 110.200 408.800 110.800 409.800 ;
        RECT 110.200 408.000 111.600 408.800 ;
        RECT 103.800 407.400 104.600 407.600 ;
        RECT 106.600 407.400 107.400 407.600 ;
        RECT 100.400 406.200 101.200 407.000 ;
        RECT 103.800 406.800 107.400 407.400 ;
        RECT 106.000 406.200 106.600 406.800 ;
        RECT 110.000 406.200 110.800 407.000 ;
        RECT 100.400 405.600 102.400 406.200 ;
        RECT 101.600 402.200 102.400 405.600 ;
        RECT 106.000 402.200 106.800 406.200 ;
        RECT 110.200 402.200 111.400 406.200 ;
        RECT 114.800 404.300 115.600 410.800 ;
        RECT 121.200 410.200 122.000 410.400 ;
        RECT 123.200 410.200 123.800 413.600 ;
        RECT 124.400 411.600 125.200 413.200 ;
        RECT 129.200 411.600 130.800 412.400 ;
        RECT 121.200 409.600 122.600 410.200 ;
        RECT 123.200 409.600 124.200 410.200 ;
        RECT 127.600 409.600 128.400 411.200 ;
        RECT 132.400 410.400 133.000 413.600 ;
        RECT 137.200 413.800 138.200 414.200 ;
        RECT 139.200 414.400 139.800 415.000 ;
        RECT 134.000 411.600 134.800 413.200 ;
        RECT 135.600 411.600 136.400 413.200 ;
        RECT 137.200 413.000 138.600 413.800 ;
        RECT 139.200 413.600 141.200 414.400 ;
        RECT 137.200 411.000 137.800 413.000 ;
        RECT 134.000 410.400 137.800 411.000 ;
        RECT 132.400 409.600 133.200 410.400 ;
        RECT 122.000 408.400 122.600 409.600 ;
        RECT 122.000 407.600 122.800 408.400 ;
        RECT 119.600 404.300 120.400 404.400 ;
        RECT 114.800 403.700 120.400 404.300 ;
        RECT 114.800 402.200 115.600 403.700 ;
        RECT 119.600 403.600 120.400 403.700 ;
        RECT 123.400 402.200 124.200 409.600 ;
        RECT 127.600 408.300 128.400 408.400 ;
        RECT 130.800 408.300 131.600 409.200 ;
        RECT 127.600 407.700 131.600 408.300 ;
        RECT 127.600 407.600 128.400 407.700 ;
        RECT 130.800 407.600 131.600 407.700 ;
        RECT 132.400 407.000 133.000 409.600 ;
        RECT 129.400 406.400 133.000 407.000 ;
        RECT 129.400 406.200 130.000 406.400 ;
        RECT 129.200 402.200 130.000 406.200 ;
        RECT 132.400 406.200 133.000 406.400 ;
        RECT 134.000 407.000 134.600 410.400 ;
        RECT 139.200 409.800 139.800 413.600 ;
        RECT 140.400 410.800 141.200 412.400 ;
        RECT 138.200 409.200 139.800 409.800 ;
        RECT 132.400 402.200 133.200 406.200 ;
        RECT 134.000 403.000 134.800 407.000 ;
        RECT 138.200 402.200 139.000 409.200 ;
        RECT 143.600 402.200 144.400 419.800 ;
        RECT 145.200 415.600 146.000 417.200 ;
        RECT 148.000 414.200 148.800 419.800 ;
        RECT 147.000 413.800 148.800 414.200 ;
        RECT 147.000 413.600 148.600 413.800 ;
        RECT 147.000 410.400 147.600 413.600 ;
        RECT 149.200 411.600 150.800 412.400 ;
        RECT 146.800 409.600 147.600 410.400 ;
        RECT 151.600 409.600 152.400 411.200 ;
        RECT 147.000 407.000 147.600 409.600 ;
        RECT 148.400 407.600 149.200 409.200 ;
        RECT 153.200 408.300 154.000 419.800 ;
        RECT 154.800 415.600 155.600 417.200 ;
        RECT 156.400 415.200 157.200 419.800 ;
        RECT 159.600 416.400 160.400 419.800 ;
        RECT 159.600 415.800 160.600 416.400 ;
        RECT 162.800 416.000 163.600 419.800 ;
        RECT 166.000 416.000 166.800 419.800 ;
        RECT 162.800 415.800 166.800 416.000 ;
        RECT 167.600 415.800 168.400 419.800 ;
        RECT 169.200 417.000 170.000 419.000 ;
        RECT 156.400 414.600 159.000 415.200 ;
        RECT 156.600 412.400 157.400 413.200 ;
        RECT 154.800 412.300 155.600 412.400 ;
        RECT 156.400 412.300 157.400 412.400 ;
        RECT 154.800 411.700 157.400 412.300 ;
        RECT 154.800 411.600 155.600 411.700 ;
        RECT 156.400 411.600 157.400 411.700 ;
        RECT 158.400 413.000 159.000 414.600 ;
        RECT 160.000 414.400 160.600 415.800 ;
        RECT 163.000 415.400 166.600 415.800 ;
        RECT 163.600 414.400 164.400 414.800 ;
        RECT 167.600 414.400 168.200 415.800 ;
        RECT 169.200 414.800 169.800 417.000 ;
        RECT 173.400 416.000 174.200 419.000 ;
        RECT 178.800 416.000 179.600 419.800 ;
        RECT 182.000 416.000 182.800 419.800 ;
        RECT 173.400 415.400 175.000 416.000 ;
        RECT 178.800 415.800 182.800 416.000 ;
        RECT 183.600 415.800 184.400 419.800 ;
        RECT 185.200 415.800 186.000 419.800 ;
        RECT 186.800 416.000 187.600 419.800 ;
        RECT 190.000 416.000 190.800 419.800 ;
        RECT 193.200 416.000 194.000 419.800 ;
        RECT 186.800 415.800 190.800 416.000 ;
        RECT 179.000 415.400 182.600 415.800 ;
        RECT 174.200 415.000 175.000 415.400 ;
        RECT 159.600 414.300 160.600 414.400 ;
        RECT 159.600 413.700 161.900 414.300 ;
        RECT 159.600 413.600 160.600 413.700 ;
        RECT 158.400 412.200 159.400 413.000 ;
        RECT 158.400 410.200 159.000 412.200 ;
        RECT 160.000 410.200 160.600 413.600 ;
        RECT 161.300 412.300 161.900 413.700 ;
        RECT 162.800 413.800 164.400 414.400 ;
        RECT 162.800 413.600 163.600 413.800 ;
        RECT 165.800 413.600 168.400 414.400 ;
        RECT 169.200 414.200 173.400 414.800 ;
        RECT 172.400 413.800 173.400 414.200 ;
        RECT 174.400 414.400 175.000 415.000 ;
        RECT 179.600 414.400 180.400 414.800 ;
        RECT 183.600 414.400 184.200 415.800 ;
        RECT 185.400 414.400 186.000 415.800 ;
        RECT 187.000 415.400 190.600 415.800 ;
        RECT 193.000 415.200 194.000 416.000 ;
        RECT 189.200 414.400 190.000 414.800 ;
        RECT 164.400 412.300 165.200 413.200 ;
        RECT 161.300 411.700 165.200 412.300 ;
        RECT 164.400 411.600 165.200 411.700 ;
        RECT 165.800 410.200 166.400 413.600 ;
        RECT 169.200 411.600 170.000 413.200 ;
        RECT 170.800 411.600 171.600 413.200 ;
        RECT 172.400 413.000 173.800 413.800 ;
        RECT 174.400 413.600 176.400 414.400 ;
        RECT 178.800 413.800 180.400 414.400 ;
        RECT 178.800 413.600 179.600 413.800 ;
        RECT 181.800 413.600 184.400 414.400 ;
        RECT 185.200 413.600 187.800 414.400 ;
        RECT 189.200 413.800 190.800 414.400 ;
        RECT 190.000 413.600 190.800 413.800 ;
        RECT 172.400 411.000 173.000 413.000 ;
        RECT 169.200 410.400 173.000 411.000 ;
        RECT 174.400 410.400 175.000 413.600 ;
        RECT 175.600 412.300 176.400 412.400 ;
        RECT 178.800 412.300 179.600 412.400 ;
        RECT 175.600 411.700 179.600 412.300 ;
        RECT 175.600 410.800 176.400 411.700 ;
        RECT 178.800 411.600 179.600 411.700 ;
        RECT 180.400 411.600 181.200 413.200 ;
        RECT 181.800 412.300 182.400 413.600 ;
        RECT 181.800 411.700 185.900 412.300 ;
        RECT 167.600 410.200 168.400 410.400 ;
        RECT 156.400 409.600 159.000 410.200 ;
        RECT 154.800 408.300 155.600 408.400 ;
        RECT 153.200 407.700 155.600 408.300 ;
        RECT 147.000 406.400 150.600 407.000 ;
        RECT 147.000 406.200 147.600 406.400 ;
        RECT 146.800 402.200 147.600 406.200 ;
        RECT 150.000 406.200 150.600 406.400 ;
        RECT 150.000 402.200 150.800 406.200 ;
        RECT 153.200 402.200 154.000 407.700 ;
        RECT 154.800 407.600 155.600 407.700 ;
        RECT 156.400 402.200 157.200 409.600 ;
        RECT 159.600 409.200 160.600 410.200 ;
        RECT 165.400 409.600 166.400 410.200 ;
        RECT 167.000 409.600 168.400 410.200 ;
        RECT 159.600 402.200 160.400 409.200 ;
        RECT 165.400 402.200 166.200 409.600 ;
        RECT 167.000 408.400 167.600 409.600 ;
        RECT 166.800 407.600 167.600 408.400 ;
        RECT 169.200 407.000 169.800 410.400 ;
        RECT 174.000 409.800 175.000 410.400 ;
        RECT 181.800 410.200 182.400 411.700 ;
        RECT 185.300 410.400 185.900 411.700 ;
        RECT 183.600 410.200 184.400 410.400 ;
        RECT 173.400 409.200 175.000 409.800 ;
        RECT 181.400 409.600 182.400 410.200 ;
        RECT 183.000 409.600 184.400 410.200 ;
        RECT 185.200 410.200 186.000 410.400 ;
        RECT 187.200 410.200 187.800 413.600 ;
        RECT 188.400 411.600 189.200 413.200 ;
        RECT 193.000 410.800 193.800 415.200 ;
        RECT 194.800 414.600 195.600 419.800 ;
        RECT 201.200 416.600 202.000 419.800 ;
        RECT 202.800 417.000 203.600 419.800 ;
        RECT 204.400 417.000 205.200 419.800 ;
        RECT 206.000 417.000 206.800 419.800 ;
        RECT 207.600 417.000 208.400 419.800 ;
        RECT 210.800 417.000 211.600 419.800 ;
        RECT 214.000 417.000 214.800 419.800 ;
        RECT 215.600 417.000 216.400 419.800 ;
        RECT 217.200 417.000 218.000 419.800 ;
        RECT 199.600 415.800 202.000 416.600 ;
        RECT 218.800 416.600 219.600 419.800 ;
        RECT 199.600 415.200 200.400 415.800 ;
        RECT 194.400 414.000 195.600 414.600 ;
        RECT 198.600 414.600 200.400 415.200 ;
        RECT 204.400 415.600 205.400 416.400 ;
        RECT 208.400 415.600 210.000 416.400 ;
        RECT 210.800 415.800 215.400 416.400 ;
        RECT 218.800 415.800 221.400 416.600 ;
        RECT 210.800 415.600 211.600 415.800 ;
        RECT 194.400 412.000 195.000 414.000 ;
        RECT 198.600 413.400 199.400 414.600 ;
        RECT 195.600 412.600 199.400 413.400 ;
        RECT 204.400 412.800 205.200 415.600 ;
        RECT 210.800 414.800 211.600 415.000 ;
        RECT 207.200 414.200 211.600 414.800 ;
        RECT 207.200 414.000 208.000 414.200 ;
        RECT 212.400 413.600 213.200 415.200 ;
        RECT 214.600 413.400 215.400 415.800 ;
        RECT 220.600 415.200 221.400 415.800 ;
        RECT 220.600 414.400 223.600 415.200 ;
        RECT 225.200 413.800 226.000 419.800 ;
        RECT 229.400 418.400 230.200 419.800 ;
        RECT 228.400 417.600 230.200 418.400 ;
        RECT 229.400 416.400 230.200 417.600 ;
        RECT 228.400 415.800 230.200 416.400 ;
        RECT 232.200 416.400 233.000 419.800 ;
        RECT 232.200 415.800 234.000 416.400 ;
        RECT 236.400 415.800 237.200 419.800 ;
        RECT 240.600 416.800 241.400 419.800 ;
        RECT 240.600 415.800 242.000 416.800 ;
        RECT 242.800 416.000 243.600 419.800 ;
        RECT 246.000 416.000 246.800 419.800 ;
        RECT 242.800 415.800 246.800 416.000 ;
        RECT 247.600 415.800 248.400 419.800 ;
        RECT 249.800 418.400 250.600 419.800 ;
        RECT 249.200 417.600 250.600 418.400 ;
        RECT 249.800 416.400 250.600 417.600 ;
        RECT 249.800 415.800 251.600 416.400 ;
        RECT 254.000 415.800 254.800 419.800 ;
        RECT 255.600 416.000 256.400 419.800 ;
        RECT 258.800 416.000 259.600 419.800 ;
        RECT 255.600 415.800 259.600 416.000 ;
        RECT 207.600 412.600 210.800 413.400 ;
        RECT 214.600 412.600 216.600 413.400 ;
        RECT 217.200 413.000 226.000 413.800 ;
        RECT 226.800 413.600 227.600 415.200 ;
        RECT 201.200 412.000 202.000 412.600 ;
        RECT 218.800 412.000 219.600 412.400 ;
        RECT 223.800 412.000 224.600 412.200 ;
        RECT 194.400 411.400 195.200 412.000 ;
        RECT 201.200 411.400 224.600 412.000 ;
        RECT 185.200 409.600 186.600 410.200 ;
        RECT 187.200 409.600 188.200 410.200 ;
        RECT 193.000 410.000 194.000 410.800 ;
        RECT 169.200 403.000 170.000 407.000 ;
        RECT 173.400 402.200 174.200 409.200 ;
        RECT 181.400 402.200 182.200 409.600 ;
        RECT 183.000 408.400 183.600 409.600 ;
        RECT 182.800 407.600 183.600 408.400 ;
        RECT 186.000 408.400 186.600 409.600 ;
        RECT 186.000 407.600 186.800 408.400 ;
        RECT 187.400 402.200 188.200 409.600 ;
        RECT 193.200 402.200 194.000 410.000 ;
        RECT 194.600 409.600 195.200 411.400 ;
        RECT 194.600 409.000 203.600 409.600 ;
        RECT 194.600 407.400 195.200 409.000 ;
        RECT 202.800 408.800 203.600 409.000 ;
        RECT 206.000 409.000 214.600 409.600 ;
        RECT 206.000 408.800 206.800 409.000 ;
        RECT 197.800 407.600 200.400 408.400 ;
        RECT 194.600 406.800 197.200 407.400 ;
        RECT 196.400 402.200 197.200 406.800 ;
        RECT 199.600 402.200 200.400 407.600 ;
        RECT 201.000 406.800 205.200 407.600 ;
        RECT 202.800 402.200 203.600 405.000 ;
        RECT 204.400 402.200 205.200 405.000 ;
        RECT 206.000 402.200 206.800 405.000 ;
        RECT 207.600 402.200 208.400 408.400 ;
        RECT 210.800 407.600 213.400 408.400 ;
        RECT 214.000 408.200 214.600 409.000 ;
        RECT 215.600 409.400 216.400 409.600 ;
        RECT 215.600 409.000 221.000 409.400 ;
        RECT 215.600 408.800 221.800 409.000 ;
        RECT 220.400 408.200 221.800 408.800 ;
        RECT 214.000 407.600 219.800 408.200 ;
        RECT 222.800 408.000 224.400 408.800 ;
        RECT 222.800 407.600 223.400 408.000 ;
        RECT 210.800 402.200 211.600 407.000 ;
        RECT 214.000 402.200 214.800 407.000 ;
        RECT 219.200 406.800 223.400 407.600 ;
        RECT 225.200 407.400 226.000 413.000 ;
        RECT 224.000 406.800 226.000 407.400 ;
        RECT 215.600 402.200 216.400 405.000 ;
        RECT 217.200 402.200 218.000 405.000 ;
        RECT 220.400 402.200 221.200 406.800 ;
        RECT 224.000 406.200 224.600 406.800 ;
        RECT 223.600 405.600 224.600 406.200 ;
        RECT 223.600 402.200 224.400 405.600 ;
        RECT 228.400 402.200 229.200 415.800 ;
        RECT 233.200 412.300 234.000 415.800 ;
        RECT 236.600 415.600 237.200 415.800 ;
        RECT 236.600 415.200 238.400 415.600 ;
        RECT 234.800 413.600 235.600 415.200 ;
        RECT 236.600 415.000 240.800 415.200 ;
        RECT 237.800 414.600 240.800 415.000 ;
        RECT 240.000 414.400 240.800 414.600 ;
        RECT 236.400 412.800 237.200 414.400 ;
        RECT 238.400 413.800 239.200 414.000 ;
        RECT 238.200 413.200 239.200 413.800 ;
        RECT 238.200 412.400 238.800 413.200 ;
        RECT 230.100 411.700 234.000 412.300 ;
        RECT 230.100 410.400 230.700 411.700 ;
        RECT 230.000 408.800 230.800 410.400 ;
        RECT 231.600 408.800 232.400 410.400 ;
        RECT 233.200 402.200 234.000 411.700 ;
        RECT 238.000 411.600 238.800 412.400 ;
        RECT 240.000 411.000 240.600 414.400 ;
        RECT 241.400 412.400 242.000 415.800 ;
        RECT 243.000 415.400 246.600 415.800 ;
        RECT 243.600 414.400 244.400 414.800 ;
        RECT 247.600 414.400 248.200 415.800 ;
        RECT 242.800 413.800 244.400 414.400 ;
        RECT 242.800 413.600 243.600 413.800 ;
        RECT 245.800 413.600 248.400 414.400 ;
        RECT 241.200 412.300 242.000 412.400 ;
        RECT 242.900 412.300 243.500 413.600 ;
        RECT 241.200 411.700 243.500 412.300 ;
        RECT 241.200 411.600 242.000 411.700 ;
        RECT 244.400 411.600 245.200 413.200 ;
        RECT 245.800 412.300 246.400 413.600 ;
        RECT 245.800 411.700 249.900 412.300 ;
        RECT 238.200 410.400 240.600 411.000 ;
        RECT 238.200 406.200 238.800 410.400 ;
        RECT 241.400 410.200 242.000 411.600 ;
        RECT 245.800 410.200 246.400 411.700 ;
        RECT 249.300 410.400 249.900 411.700 ;
        RECT 247.600 410.200 248.400 410.400 ;
        RECT 238.000 402.200 238.800 406.200 ;
        RECT 241.200 402.200 242.000 410.200 ;
        RECT 245.400 409.600 246.400 410.200 ;
        RECT 247.000 409.600 248.400 410.200 ;
        RECT 245.400 402.200 246.200 409.600 ;
        RECT 247.000 408.400 247.600 409.600 ;
        RECT 249.200 408.800 250.000 410.400 ;
        RECT 246.800 407.600 247.600 408.400 ;
        RECT 250.800 402.200 251.600 415.800 ;
        RECT 252.400 414.300 253.200 415.200 ;
        RECT 254.200 414.400 254.800 415.800 ;
        RECT 255.800 415.400 259.400 415.800 ;
        RECT 258.000 414.400 258.800 414.800 ;
        RECT 254.000 414.300 256.600 414.400 ;
        RECT 252.400 413.700 256.600 414.300 ;
        RECT 258.000 413.800 259.600 414.400 ;
        RECT 252.400 413.600 253.200 413.700 ;
        RECT 254.000 413.600 256.600 413.700 ;
        RECT 258.800 413.600 259.600 413.800 ;
        RECT 265.200 413.800 266.000 419.800 ;
        RECT 271.600 416.600 272.400 419.800 ;
        RECT 273.200 417.000 274.000 419.800 ;
        RECT 274.800 417.000 275.600 419.800 ;
        RECT 276.400 417.000 277.200 419.800 ;
        RECT 279.600 417.000 280.400 419.800 ;
        RECT 282.800 417.000 283.600 419.800 ;
        RECT 284.400 417.000 285.200 419.800 ;
        RECT 286.000 417.000 286.800 419.800 ;
        RECT 287.600 417.000 288.400 419.800 ;
        RECT 269.800 415.800 272.400 416.600 ;
        RECT 289.200 416.600 290.000 419.800 ;
        RECT 275.800 415.800 280.400 416.400 ;
        RECT 269.800 415.200 270.600 415.800 ;
        RECT 267.600 414.400 270.600 415.200 ;
        RECT 252.400 410.300 253.200 410.400 ;
        RECT 254.000 410.300 254.800 410.400 ;
        RECT 252.400 410.200 254.800 410.300 ;
        RECT 256.000 410.200 256.600 413.600 ;
        RECT 257.200 411.600 258.000 413.200 ;
        RECT 265.200 413.000 274.000 413.800 ;
        RECT 275.800 413.400 276.600 415.800 ;
        RECT 279.600 415.600 280.400 415.800 ;
        RECT 281.200 415.600 282.800 416.400 ;
        RECT 285.800 415.600 286.800 416.400 ;
        RECT 289.200 415.800 291.600 416.600 ;
        RECT 278.000 413.600 278.800 415.200 ;
        RECT 279.600 414.800 280.400 415.000 ;
        RECT 279.600 414.200 284.000 414.800 ;
        RECT 283.200 414.000 284.000 414.200 ;
        RECT 252.400 409.700 255.400 410.200 ;
        RECT 252.400 409.600 253.200 409.700 ;
        RECT 254.000 409.600 255.400 409.700 ;
        RECT 256.000 409.600 257.000 410.200 ;
        RECT 254.800 408.400 255.400 409.600 ;
        RECT 254.800 407.600 255.600 408.400 ;
        RECT 256.200 402.200 257.000 409.600 ;
        RECT 265.200 407.400 266.000 413.000 ;
        RECT 274.600 412.600 276.600 413.400 ;
        RECT 280.400 412.600 283.600 413.400 ;
        RECT 286.000 412.800 286.800 415.600 ;
        RECT 290.800 415.200 291.600 415.800 ;
        RECT 290.800 414.600 292.600 415.200 ;
        RECT 291.800 413.400 292.600 414.600 ;
        RECT 295.600 414.600 296.400 419.800 ;
        RECT 297.200 416.000 298.000 419.800 ;
        RECT 301.000 416.400 301.800 419.800 ;
        RECT 297.200 415.200 298.200 416.000 ;
        RECT 301.000 415.800 302.800 416.400 ;
        RECT 295.600 414.000 296.800 414.600 ;
        RECT 291.800 412.600 295.600 413.400 ;
        RECT 296.200 412.000 296.800 414.000 ;
        RECT 296.000 411.400 296.800 412.000 ;
        RECT 294.600 410.800 295.400 411.000 ;
        RECT 268.400 410.200 295.400 410.800 ;
        RECT 268.400 409.600 269.200 410.200 ;
        RECT 271.800 410.000 272.600 410.200 ;
        RECT 296.000 409.600 296.600 411.400 ;
        RECT 297.400 410.800 298.200 415.200 ;
        RECT 274.800 409.400 275.600 409.600 ;
        RECT 270.200 409.000 275.600 409.400 ;
        RECT 269.400 408.800 275.600 409.000 ;
        RECT 276.600 409.000 285.200 409.600 ;
        RECT 266.800 408.000 268.400 408.800 ;
        RECT 269.400 408.200 270.800 408.800 ;
        RECT 276.600 408.200 277.200 409.000 ;
        RECT 284.400 408.800 285.200 409.000 ;
        RECT 287.600 409.000 296.600 409.600 ;
        RECT 287.600 408.800 288.400 409.000 ;
        RECT 267.800 407.600 268.400 408.000 ;
        RECT 271.400 407.600 277.200 408.200 ;
        RECT 277.800 407.600 280.400 408.400 ;
        RECT 265.200 406.800 267.200 407.400 ;
        RECT 267.800 406.800 272.000 407.600 ;
        RECT 266.600 406.200 267.200 406.800 ;
        RECT 266.600 405.600 267.600 406.200 ;
        RECT 266.800 402.200 267.600 405.600 ;
        RECT 270.000 402.200 270.800 406.800 ;
        RECT 273.200 402.200 274.000 405.000 ;
        RECT 274.800 402.200 275.600 405.000 ;
        RECT 276.400 402.200 277.200 407.000 ;
        RECT 279.600 402.200 280.400 407.000 ;
        RECT 282.800 402.200 283.600 408.400 ;
        RECT 290.800 407.600 293.400 408.400 ;
        RECT 286.000 406.800 290.200 407.600 ;
        RECT 284.400 402.200 285.200 405.000 ;
        RECT 286.000 402.200 286.800 405.000 ;
        RECT 287.600 402.200 288.400 405.000 ;
        RECT 290.800 402.200 291.600 407.600 ;
        RECT 296.000 407.400 296.600 409.000 ;
        RECT 294.000 406.800 296.600 407.400 ;
        RECT 297.200 410.000 298.200 410.800 ;
        RECT 294.000 402.200 294.800 406.800 ;
        RECT 297.200 402.200 298.000 410.000 ;
        RECT 300.400 408.800 301.200 410.400 ;
        RECT 302.000 410.300 302.800 415.800 ;
        RECT 303.600 414.300 304.400 415.200 ;
        RECT 305.200 414.300 306.000 419.800 ;
        RECT 311.000 418.400 311.800 419.800 ;
        RECT 310.000 417.600 311.800 418.400 ;
        RECT 306.800 415.600 307.600 417.200 ;
        RECT 311.000 416.400 311.800 417.600 ;
        RECT 310.000 415.800 311.800 416.400 ;
        RECT 314.800 417.800 315.600 419.800 ;
        RECT 303.600 413.700 306.000 414.300 ;
        RECT 303.600 413.600 304.400 413.700 ;
        RECT 303.600 410.300 304.400 410.400 ;
        RECT 302.000 409.700 304.400 410.300 ;
        RECT 302.000 402.200 302.800 409.700 ;
        RECT 303.600 409.600 304.400 409.700 ;
        RECT 305.200 402.200 306.000 413.700 ;
        RECT 308.400 413.600 309.200 415.200 ;
        RECT 310.000 402.200 310.800 415.800 ;
        RECT 314.800 414.400 315.400 417.800 ;
        RECT 319.600 417.600 320.400 419.800 ;
        RECT 316.400 415.600 317.200 417.200 ;
        RECT 319.600 414.400 320.200 417.600 ;
        RECT 321.200 415.600 322.000 417.200 ;
        RECT 322.800 415.800 323.600 419.800 ;
        RECT 324.400 416.000 325.200 419.800 ;
        RECT 327.600 416.000 328.400 419.800 ;
        RECT 329.400 416.400 330.200 417.200 ;
        RECT 324.400 415.800 328.400 416.000 ;
        RECT 323.000 414.400 323.600 415.800 ;
        RECT 324.600 415.400 328.200 415.800 ;
        RECT 329.200 415.600 330.000 416.400 ;
        RECT 330.800 415.800 331.600 419.800 ;
        RECT 336.200 416.400 337.000 419.800 ;
        RECT 336.200 415.800 338.000 416.400 ;
        RECT 340.400 415.800 341.200 419.800 ;
        RECT 342.000 416.000 342.800 419.800 ;
        RECT 345.200 416.000 346.000 419.800 ;
        RECT 347.000 416.400 347.800 417.200 ;
        RECT 342.000 415.800 346.000 416.000 ;
        RECT 326.800 414.400 327.600 414.800 ;
        RECT 314.800 413.600 315.600 414.400 ;
        RECT 319.600 413.600 320.400 414.400 ;
        RECT 322.800 413.600 325.400 414.400 ;
        RECT 326.800 413.800 328.400 414.400 ;
        RECT 327.600 413.600 328.400 413.800 ;
        RECT 313.200 412.300 314.000 412.400 ;
        RECT 311.700 411.700 314.000 412.300 ;
        RECT 311.700 410.400 312.300 411.700 ;
        RECT 313.200 410.800 314.000 411.700 ;
        RECT 314.800 412.300 315.400 413.600 ;
        RECT 318.000 412.300 318.800 412.400 ;
        RECT 314.800 411.700 318.800 412.300 ;
        RECT 311.600 408.800 312.400 410.400 ;
        RECT 314.800 410.200 315.400 411.700 ;
        RECT 318.000 410.800 318.800 411.700 ;
        RECT 319.600 410.200 320.200 413.600 ;
        RECT 322.800 410.200 323.600 410.400 ;
        RECT 324.800 410.200 325.400 413.600 ;
        RECT 326.000 411.600 326.800 413.200 ;
        RECT 329.200 412.200 330.000 412.400 ;
        RECT 331.000 412.200 331.600 415.800 ;
        RECT 332.400 412.800 333.200 414.400 ;
        RECT 334.000 412.200 334.800 412.400 ;
        RECT 329.200 411.600 331.600 412.200 ;
        RECT 333.200 411.600 334.800 412.200 ;
        RECT 329.400 410.200 330.000 411.600 ;
        RECT 333.200 411.200 334.000 411.600 ;
        RECT 313.800 409.400 315.600 410.200 ;
        RECT 318.600 409.400 320.400 410.200 ;
        RECT 322.800 409.600 324.200 410.200 ;
        RECT 324.800 409.600 325.800 410.200 ;
        RECT 313.800 402.200 314.600 409.400 ;
        RECT 318.600 402.200 319.400 409.400 ;
        RECT 323.600 408.400 324.200 409.600 ;
        RECT 323.600 407.600 324.400 408.400 ;
        RECT 325.000 402.200 325.800 409.600 ;
        RECT 329.200 402.200 330.000 410.200 ;
        RECT 330.800 409.600 334.800 410.200 ;
        RECT 330.800 402.200 331.600 409.600 ;
        RECT 334.000 402.200 334.800 409.600 ;
        RECT 335.600 408.800 336.400 410.400 ;
        RECT 337.200 402.200 338.000 415.800 ;
        RECT 338.800 413.600 339.600 415.200 ;
        RECT 340.600 414.400 341.200 415.800 ;
        RECT 342.200 415.400 345.800 415.800 ;
        RECT 346.800 415.600 347.600 416.400 ;
        RECT 348.400 415.800 349.200 419.800 ;
        RECT 354.800 417.800 355.600 419.800 ;
        RECT 344.400 414.400 345.200 414.800 ;
        RECT 340.400 413.600 343.000 414.400 ;
        RECT 344.400 414.300 346.000 414.400 ;
        RECT 346.800 414.300 347.600 414.400 ;
        RECT 344.400 413.800 347.600 414.300 ;
        RECT 345.200 413.700 347.600 413.800 ;
        RECT 345.200 413.600 346.000 413.700 ;
        RECT 346.800 413.600 347.600 413.700 ;
        RECT 338.900 412.300 339.500 413.600 ;
        RECT 340.400 412.300 341.200 412.400 ;
        RECT 338.900 411.700 341.200 412.300 ;
        RECT 340.400 411.600 341.200 411.700 ;
        RECT 338.800 410.300 339.600 410.400 ;
        RECT 340.400 410.300 341.200 410.400 ;
        RECT 338.800 410.200 341.200 410.300 ;
        RECT 342.400 410.200 343.000 413.600 ;
        RECT 343.600 411.600 344.400 413.200 ;
        RECT 346.800 412.200 347.600 412.400 ;
        RECT 348.600 412.200 349.200 415.800 ;
        RECT 353.200 415.600 354.000 417.200 ;
        RECT 355.000 414.400 355.600 417.800 ;
        RECT 360.600 416.400 361.400 419.800 ;
        RECT 359.600 415.800 361.400 416.400 ;
        RECT 350.000 412.800 350.800 414.400 ;
        RECT 354.800 413.600 355.600 414.400 ;
        RECT 358.000 413.600 358.800 415.200 ;
        RECT 351.600 412.200 352.400 412.400 ;
        RECT 346.800 411.600 349.200 412.200 ;
        RECT 350.800 411.600 352.400 412.200 ;
        RECT 353.200 412.300 354.000 412.400 ;
        RECT 355.000 412.300 355.600 413.600 ;
        RECT 353.200 411.700 355.600 412.300 ;
        RECT 353.200 411.600 354.000 411.700 ;
        RECT 347.000 410.200 347.600 411.600 ;
        RECT 350.800 411.200 351.600 411.600 ;
        RECT 355.000 410.200 355.600 411.700 ;
        RECT 356.400 410.800 357.200 412.400 ;
        RECT 338.800 409.700 341.800 410.200 ;
        RECT 338.800 409.600 339.600 409.700 ;
        RECT 340.400 409.600 341.800 409.700 ;
        RECT 342.400 409.600 343.400 410.200 ;
        RECT 341.200 408.400 341.800 409.600 ;
        RECT 341.200 407.600 342.000 408.400 ;
        RECT 342.600 402.200 343.400 409.600 ;
        RECT 346.800 402.200 347.600 410.200 ;
        RECT 348.400 409.600 352.400 410.200 ;
        RECT 348.400 402.200 349.200 409.600 ;
        RECT 351.600 402.200 352.400 409.600 ;
        RECT 354.800 409.400 356.600 410.200 ;
        RECT 355.800 402.200 356.600 409.400 ;
        RECT 359.600 402.200 360.400 415.800 ;
        RECT 364.000 414.200 364.800 419.800 ;
        RECT 363.000 413.800 364.800 414.200 ;
        RECT 372.800 414.200 373.600 419.800 ;
        RECT 376.800 414.200 377.600 419.800 ;
        RECT 372.800 413.800 374.600 414.200 ;
        RECT 363.000 413.600 364.600 413.800 ;
        RECT 373.000 413.600 374.600 413.800 ;
        RECT 363.000 410.400 363.600 413.600 ;
        RECT 365.200 411.600 366.800 412.400 ;
        RECT 370.800 411.600 372.400 412.400 ;
        RECT 361.200 408.800 362.000 410.400 ;
        RECT 362.800 409.600 363.600 410.400 ;
        RECT 367.600 409.600 368.400 411.200 ;
        RECT 369.200 409.600 370.000 411.200 ;
        RECT 374.000 410.400 374.600 413.600 ;
        RECT 375.800 413.800 377.600 414.200 ;
        RECT 375.800 413.600 377.400 413.800 ;
        RECT 375.800 410.400 376.400 413.600 ;
        RECT 378.000 411.600 379.600 412.400 ;
        RECT 374.000 409.600 374.800 410.400 ;
        RECT 375.600 409.600 376.400 410.400 ;
        RECT 380.400 409.600 381.200 411.200 ;
        RECT 363.000 407.000 363.600 409.600 ;
        RECT 364.400 407.600 365.200 409.200 ;
        RECT 367.700 408.300 368.300 409.600 ;
        RECT 370.800 408.300 371.600 408.400 ;
        RECT 367.700 407.700 371.600 408.300 ;
        RECT 370.800 407.600 371.600 407.700 ;
        RECT 372.400 407.600 373.200 409.200 ;
        RECT 374.000 407.000 374.600 409.600 ;
        RECT 363.000 406.400 366.600 407.000 ;
        RECT 371.000 406.400 374.600 407.000 ;
        RECT 363.000 406.200 363.600 406.400 ;
        RECT 362.800 402.200 363.600 406.200 ;
        RECT 366.000 406.200 366.600 406.400 ;
        RECT 366.000 402.200 366.800 406.200 ;
        RECT 370.800 402.200 371.600 406.400 ;
        RECT 374.000 406.200 374.600 406.400 ;
        RECT 375.800 407.000 376.400 409.600 ;
        RECT 377.200 407.600 378.000 409.200 ;
        RECT 375.800 406.400 379.400 407.000 ;
        RECT 375.800 406.200 376.400 406.400 ;
        RECT 374.000 402.200 374.800 406.200 ;
        RECT 375.600 402.200 376.400 406.200 ;
        RECT 378.800 402.200 379.600 406.400 ;
        RECT 382.000 402.200 382.800 419.800 ;
        RECT 387.800 415.800 389.400 419.800 ;
        RECT 383.600 413.600 384.400 415.200 ;
        RECT 386.800 413.600 387.600 414.400 ;
        RECT 387.000 413.200 387.600 413.600 ;
        RECT 387.000 412.400 387.800 413.200 ;
        RECT 388.400 412.400 389.000 415.800 ;
        RECT 390.000 412.800 390.800 414.400 ;
        RECT 396.800 414.200 397.600 419.800 ;
        RECT 399.800 416.400 400.600 417.200 ;
        RECT 399.600 415.600 400.400 416.400 ;
        RECT 401.200 415.600 402.000 419.800 ;
        RECT 396.800 413.800 398.600 414.200 ;
        RECT 397.000 413.600 398.600 413.800 ;
        RECT 385.200 410.800 386.000 412.400 ;
        RECT 388.400 411.600 389.200 412.400 ;
        RECT 391.600 412.200 392.400 412.400 ;
        RECT 390.800 411.600 392.400 412.200 ;
        RECT 394.800 411.600 396.400 412.400 ;
        RECT 388.400 411.400 389.000 411.600 ;
        RECT 387.000 410.800 389.000 411.400 ;
        RECT 390.800 411.200 391.600 411.600 ;
        RECT 387.000 410.200 387.600 410.800 ;
        RECT 385.200 402.800 386.000 410.200 ;
        RECT 386.800 403.400 387.600 410.200 ;
        RECT 388.400 409.600 392.400 410.200 ;
        RECT 393.200 409.600 394.000 411.200 ;
        RECT 398.000 410.400 398.600 413.600 ;
        RECT 399.600 412.200 400.400 412.400 ;
        RECT 401.400 412.200 402.000 415.600 ;
        RECT 407.600 417.800 408.400 419.800 ;
        RECT 407.600 414.400 408.200 417.800 ;
        RECT 409.200 415.600 410.000 417.200 ;
        RECT 417.200 416.000 418.000 419.800 ;
        RECT 417.000 415.200 418.000 416.000 ;
        RECT 402.800 412.800 403.600 414.400 ;
        RECT 407.600 414.300 408.400 414.400 ;
        RECT 404.500 413.700 408.400 414.300 ;
        RECT 404.500 412.400 405.100 413.700 ;
        RECT 407.600 413.600 408.400 413.700 ;
        RECT 404.400 412.200 405.200 412.400 ;
        RECT 399.600 411.600 402.000 412.200 ;
        RECT 403.600 411.600 405.200 412.200 ;
        RECT 398.000 409.600 398.800 410.400 ;
        RECT 399.800 410.200 400.400 411.600 ;
        RECT 403.600 411.200 404.400 411.600 ;
        RECT 406.000 410.800 406.800 412.400 ;
        RECT 407.600 410.200 408.200 413.600 ;
        RECT 417.000 410.800 417.800 415.200 ;
        RECT 418.800 414.600 419.600 419.800 ;
        RECT 425.200 416.600 426.000 419.800 ;
        RECT 426.800 417.000 427.600 419.800 ;
        RECT 428.400 417.000 429.200 419.800 ;
        RECT 430.000 417.000 430.800 419.800 ;
        RECT 431.600 417.000 432.400 419.800 ;
        RECT 434.800 417.000 435.600 419.800 ;
        RECT 438.000 417.000 438.800 419.800 ;
        RECT 439.600 417.000 440.400 419.800 ;
        RECT 441.200 417.000 442.000 419.800 ;
        RECT 423.600 415.800 426.000 416.600 ;
        RECT 442.800 416.600 443.600 419.800 ;
        RECT 423.600 415.200 424.400 415.800 ;
        RECT 418.400 414.000 419.600 414.600 ;
        RECT 422.600 414.600 424.400 415.200 ;
        RECT 428.400 415.600 429.400 416.400 ;
        RECT 432.400 415.600 434.000 416.400 ;
        RECT 434.800 415.800 439.400 416.400 ;
        RECT 442.800 415.800 445.400 416.600 ;
        RECT 434.800 415.600 435.600 415.800 ;
        RECT 418.400 412.000 419.000 414.000 ;
        RECT 422.600 413.400 423.400 414.600 ;
        RECT 419.600 412.600 423.400 413.400 ;
        RECT 428.400 412.800 429.200 415.600 ;
        RECT 434.800 414.800 435.600 415.000 ;
        RECT 431.200 414.200 435.600 414.800 ;
        RECT 431.200 414.000 432.000 414.200 ;
        RECT 436.400 413.600 437.200 415.200 ;
        RECT 438.600 413.400 439.400 415.800 ;
        RECT 444.600 415.200 445.400 415.800 ;
        RECT 444.600 414.400 447.600 415.200 ;
        RECT 449.200 413.800 450.000 419.800 ;
        RECT 431.600 412.600 434.800 413.400 ;
        RECT 438.600 412.600 440.600 413.400 ;
        RECT 441.200 413.000 450.000 413.800 ;
        RECT 425.200 412.000 426.000 412.600 ;
        RECT 442.800 412.000 443.600 412.400 ;
        RECT 447.600 412.200 448.400 412.400 ;
        RECT 447.600 412.000 448.600 412.200 ;
        RECT 418.400 411.400 419.200 412.000 ;
        RECT 425.200 411.400 448.600 412.000 ;
        RECT 388.400 402.800 389.200 409.600 ;
        RECT 385.200 402.200 389.200 402.800 ;
        RECT 391.600 402.200 392.400 409.600 ;
        RECT 396.400 407.600 397.200 409.200 ;
        RECT 398.000 407.000 398.600 409.600 ;
        RECT 395.000 406.400 398.600 407.000 ;
        RECT 395.000 406.200 395.600 406.400 ;
        RECT 394.800 402.200 395.600 406.200 ;
        RECT 398.000 406.200 398.600 406.400 ;
        RECT 398.000 402.200 398.800 406.200 ;
        RECT 399.600 402.200 400.400 410.200 ;
        RECT 401.200 409.600 405.200 410.200 ;
        RECT 401.200 402.200 402.000 409.600 ;
        RECT 404.400 402.200 405.200 409.600 ;
        RECT 406.600 409.400 408.400 410.200 ;
        RECT 417.000 410.000 418.000 410.800 ;
        RECT 406.600 404.400 407.400 409.400 ;
        RECT 412.400 408.300 413.200 408.400 ;
        RECT 417.200 408.300 418.000 410.000 ;
        RECT 412.400 407.700 418.000 408.300 ;
        RECT 412.400 407.600 413.200 407.700 ;
        RECT 406.000 403.600 407.400 404.400 ;
        RECT 406.600 402.200 407.400 403.600 ;
        RECT 417.200 402.200 418.000 407.700 ;
        RECT 418.600 409.600 419.200 411.400 ;
        RECT 418.600 409.000 427.600 409.600 ;
        RECT 418.600 407.400 419.200 409.000 ;
        RECT 426.800 408.800 427.600 409.000 ;
        RECT 430.000 409.000 438.600 409.600 ;
        RECT 430.000 408.800 430.800 409.000 ;
        RECT 421.800 407.600 424.400 408.400 ;
        RECT 418.600 406.800 421.200 407.400 ;
        RECT 420.400 402.200 421.200 406.800 ;
        RECT 423.600 402.200 424.400 407.600 ;
        RECT 425.000 406.800 429.200 407.600 ;
        RECT 426.800 402.200 427.600 405.000 ;
        RECT 428.400 402.200 429.200 405.000 ;
        RECT 430.000 402.200 430.800 405.000 ;
        RECT 431.600 402.200 432.400 408.400 ;
        RECT 434.800 407.600 437.400 408.400 ;
        RECT 438.000 408.200 438.600 409.000 ;
        RECT 439.600 409.400 440.400 409.600 ;
        RECT 439.600 409.000 445.000 409.400 ;
        RECT 439.600 408.800 445.800 409.000 ;
        RECT 444.400 408.200 445.800 408.800 ;
        RECT 438.000 407.600 443.800 408.200 ;
        RECT 446.800 408.000 448.400 408.800 ;
        RECT 446.800 407.600 447.400 408.000 ;
        RECT 434.800 402.200 435.600 407.000 ;
        RECT 438.000 402.200 438.800 407.000 ;
        RECT 443.200 406.800 447.400 407.600 ;
        RECT 449.200 407.400 450.000 413.000 ;
        RECT 448.000 406.800 450.000 407.400 ;
        RECT 450.800 413.800 451.600 419.800 ;
        RECT 457.200 416.600 458.000 419.800 ;
        RECT 458.800 417.000 459.600 419.800 ;
        RECT 460.400 417.000 461.200 419.800 ;
        RECT 462.000 417.000 462.800 419.800 ;
        RECT 465.200 417.000 466.000 419.800 ;
        RECT 468.400 417.000 469.200 419.800 ;
        RECT 470.000 417.000 470.800 419.800 ;
        RECT 471.600 417.000 472.400 419.800 ;
        RECT 473.200 417.000 474.000 419.800 ;
        RECT 455.400 415.800 458.000 416.600 ;
        RECT 474.800 416.600 475.600 419.800 ;
        RECT 461.400 415.800 466.000 416.400 ;
        RECT 455.400 415.200 456.200 415.800 ;
        RECT 453.200 414.400 456.200 415.200 ;
        RECT 450.800 413.000 459.600 413.800 ;
        RECT 461.400 413.400 462.200 415.800 ;
        RECT 465.200 415.600 466.000 415.800 ;
        RECT 466.800 415.600 468.400 416.400 ;
        RECT 471.400 415.600 472.400 416.400 ;
        RECT 474.800 415.800 477.200 416.600 ;
        RECT 463.600 413.600 464.400 415.200 ;
        RECT 465.200 414.800 466.000 415.000 ;
        RECT 465.200 414.200 469.600 414.800 ;
        RECT 468.800 414.000 469.600 414.200 ;
        RECT 450.800 407.400 451.600 413.000 ;
        RECT 460.200 412.600 462.200 413.400 ;
        RECT 466.000 412.600 469.200 413.400 ;
        RECT 471.600 412.800 472.400 415.600 ;
        RECT 476.400 415.200 477.200 415.800 ;
        RECT 476.400 414.600 478.200 415.200 ;
        RECT 477.400 413.400 478.200 414.600 ;
        RECT 481.200 414.600 482.000 419.800 ;
        RECT 482.800 416.000 483.600 419.800 ;
        RECT 486.000 416.000 486.800 419.800 ;
        RECT 489.200 416.000 490.000 419.800 ;
        RECT 482.800 415.200 483.800 416.000 ;
        RECT 486.000 415.800 490.000 416.000 ;
        RECT 490.800 415.800 491.600 419.800 ;
        RECT 492.400 415.800 493.200 419.800 ;
        RECT 494.000 416.000 494.800 419.800 ;
        RECT 497.200 416.000 498.000 419.800 ;
        RECT 494.000 415.800 498.000 416.000 ;
        RECT 486.200 415.400 489.800 415.800 ;
        RECT 481.200 414.000 482.400 414.600 ;
        RECT 477.400 412.600 481.200 413.400 ;
        RECT 452.200 412.000 453.000 412.200 ;
        RECT 454.000 412.000 454.800 412.400 ;
        RECT 455.600 412.000 456.400 412.400 ;
        RECT 457.200 412.000 458.000 412.400 ;
        RECT 474.800 412.000 475.600 412.600 ;
        RECT 481.800 412.000 482.400 414.000 ;
        RECT 452.200 411.400 475.600 412.000 ;
        RECT 481.600 411.400 482.400 412.000 ;
        RECT 481.600 409.600 482.200 411.400 ;
        RECT 483.000 410.800 483.800 415.200 ;
        RECT 486.800 414.400 487.600 414.800 ;
        RECT 490.800 414.400 491.400 415.800 ;
        RECT 492.600 414.400 493.200 415.800 ;
        RECT 494.200 415.400 497.800 415.800 ;
        RECT 496.400 414.400 497.200 414.800 ;
        RECT 486.000 413.800 487.600 414.400 ;
        RECT 486.000 413.600 486.800 413.800 ;
        RECT 489.000 413.600 491.600 414.400 ;
        RECT 492.400 413.600 495.000 414.400 ;
        RECT 496.400 414.300 498.000 414.400 ;
        RECT 498.800 414.300 499.600 419.800 ;
        RECT 500.400 415.600 501.200 417.200 ;
        RECT 502.000 416.000 502.800 419.800 ;
        RECT 505.200 416.000 506.000 419.800 ;
        RECT 502.000 415.800 506.000 416.000 ;
        RECT 506.800 415.800 507.600 419.800 ;
        RECT 510.000 416.000 510.800 419.800 ;
        RECT 502.200 415.400 505.800 415.800 ;
        RECT 502.800 414.400 503.600 414.800 ;
        RECT 506.800 414.400 507.400 415.800 ;
        RECT 509.800 415.200 510.800 416.000 ;
        RECT 496.400 413.800 499.600 414.300 ;
        RECT 497.200 413.700 499.600 413.800 ;
        RECT 497.200 413.600 498.000 413.700 ;
        RECT 487.600 411.600 488.400 413.200 ;
        RECT 489.000 412.400 489.600 413.600 ;
        RECT 489.000 411.600 490.000 412.400 ;
        RECT 460.400 409.400 461.200 409.600 ;
        RECT 455.800 409.000 461.200 409.400 ;
        RECT 455.000 408.800 461.200 409.000 ;
        RECT 462.200 409.000 470.800 409.600 ;
        RECT 452.400 408.000 454.000 408.800 ;
        RECT 455.000 408.200 456.400 408.800 ;
        RECT 462.200 408.200 462.800 409.000 ;
        RECT 470.000 408.800 470.800 409.000 ;
        RECT 473.200 409.000 482.200 409.600 ;
        RECT 473.200 408.800 474.000 409.000 ;
        RECT 453.400 407.600 454.000 408.000 ;
        RECT 457.000 407.600 462.800 408.200 ;
        RECT 463.400 407.600 466.000 408.400 ;
        RECT 450.800 406.800 452.800 407.400 ;
        RECT 453.400 406.800 457.600 407.600 ;
        RECT 439.600 402.200 440.400 405.000 ;
        RECT 441.200 402.200 442.000 405.000 ;
        RECT 444.400 402.200 445.200 406.800 ;
        RECT 448.000 406.200 448.600 406.800 ;
        RECT 447.600 405.600 448.600 406.200 ;
        RECT 452.200 406.200 452.800 406.800 ;
        RECT 452.200 405.600 453.200 406.200 ;
        RECT 447.600 402.200 448.400 405.600 ;
        RECT 452.400 402.200 453.200 405.600 ;
        RECT 455.600 402.200 456.400 406.800 ;
        RECT 458.800 402.200 459.600 405.000 ;
        RECT 460.400 402.200 461.200 405.000 ;
        RECT 462.000 402.200 462.800 407.000 ;
        RECT 465.200 402.200 466.000 407.000 ;
        RECT 468.400 402.200 469.200 408.400 ;
        RECT 476.400 407.600 479.000 408.400 ;
        RECT 471.600 406.800 475.800 407.600 ;
        RECT 470.000 402.200 470.800 405.000 ;
        RECT 471.600 402.200 472.400 405.000 ;
        RECT 473.200 402.200 474.000 405.000 ;
        RECT 476.400 402.200 477.200 407.600 ;
        RECT 481.600 407.400 482.200 409.000 ;
        RECT 479.600 406.800 482.200 407.400 ;
        RECT 482.800 410.000 483.800 410.800 ;
        RECT 489.000 410.200 489.600 411.600 ;
        RECT 490.800 410.200 491.600 410.400 ;
        RECT 479.600 402.200 480.400 406.800 ;
        RECT 482.800 402.200 483.600 410.000 ;
        RECT 488.600 409.600 489.600 410.200 ;
        RECT 490.200 409.600 491.600 410.200 ;
        RECT 492.400 410.200 493.200 410.400 ;
        RECT 494.400 410.200 495.000 413.600 ;
        RECT 495.600 411.600 496.400 413.200 ;
        RECT 492.400 409.600 493.800 410.200 ;
        RECT 494.400 409.600 495.400 410.200 ;
        RECT 488.600 402.200 489.400 409.600 ;
        RECT 490.200 408.400 490.800 409.600 ;
        RECT 490.000 407.600 490.800 408.400 ;
        RECT 493.200 408.400 493.800 409.600 ;
        RECT 493.200 407.600 494.000 408.400 ;
        RECT 494.600 402.200 495.400 409.600 ;
        RECT 498.800 402.200 499.600 413.700 ;
        RECT 502.000 413.800 503.600 414.400 ;
        RECT 502.000 413.600 502.800 413.800 ;
        RECT 505.000 413.600 507.600 414.400 ;
        RECT 503.600 411.600 504.400 413.200 ;
        RECT 505.000 410.200 505.600 413.600 ;
        RECT 509.800 410.800 510.600 415.200 ;
        RECT 511.600 414.600 512.400 419.800 ;
        RECT 518.000 416.600 518.800 419.800 ;
        RECT 519.600 417.000 520.400 419.800 ;
        RECT 521.200 417.000 522.000 419.800 ;
        RECT 522.800 417.000 523.600 419.800 ;
        RECT 524.400 417.000 525.200 419.800 ;
        RECT 527.600 417.000 528.400 419.800 ;
        RECT 530.800 417.000 531.600 419.800 ;
        RECT 532.400 417.000 533.200 419.800 ;
        RECT 534.000 417.000 534.800 419.800 ;
        RECT 516.400 415.800 518.800 416.600 ;
        RECT 535.600 416.600 536.400 419.800 ;
        RECT 516.400 415.200 517.200 415.800 ;
        RECT 511.200 414.000 512.400 414.600 ;
        RECT 515.400 414.600 517.200 415.200 ;
        RECT 521.200 415.600 522.200 416.400 ;
        RECT 525.200 415.600 526.800 416.400 ;
        RECT 527.600 415.800 532.200 416.400 ;
        RECT 535.600 415.800 538.200 416.600 ;
        RECT 527.600 415.600 528.400 415.800 ;
        RECT 511.200 412.000 511.800 414.000 ;
        RECT 515.400 413.400 516.200 414.600 ;
        RECT 512.400 412.600 516.200 413.400 ;
        RECT 521.200 412.800 522.000 415.600 ;
        RECT 527.600 414.800 528.400 415.000 ;
        RECT 524.000 414.200 528.400 414.800 ;
        RECT 524.000 414.000 524.800 414.200 ;
        RECT 529.200 413.600 530.000 415.200 ;
        RECT 531.400 413.400 532.200 415.800 ;
        RECT 537.400 415.200 538.200 415.800 ;
        RECT 537.400 414.400 540.400 415.200 ;
        RECT 542.000 413.800 542.800 419.800 ;
        RECT 545.200 416.400 546.000 419.800 ;
        RECT 524.400 412.600 527.600 413.400 ;
        RECT 531.400 412.600 533.400 413.400 ;
        RECT 534.000 413.000 542.800 413.800 ;
        RECT 518.000 412.000 518.800 412.600 ;
        RECT 535.600 412.000 536.400 412.400 ;
        RECT 540.400 412.200 541.200 412.400 ;
        RECT 540.400 412.000 541.400 412.200 ;
        RECT 511.200 411.400 512.000 412.000 ;
        RECT 518.000 411.400 541.400 412.000 ;
        RECT 506.800 410.200 507.600 410.400 ;
        RECT 504.600 409.600 505.600 410.200 ;
        RECT 506.200 409.600 507.600 410.200 ;
        RECT 509.800 410.000 510.800 410.800 ;
        RECT 504.600 402.200 505.400 409.600 ;
        RECT 506.200 408.400 506.800 409.600 ;
        RECT 506.000 407.600 506.800 408.400 ;
        RECT 510.000 402.200 510.800 410.000 ;
        RECT 511.400 409.600 512.000 411.400 ;
        RECT 511.400 409.000 520.400 409.600 ;
        RECT 511.400 407.400 512.000 409.000 ;
        RECT 519.600 408.800 520.400 409.000 ;
        RECT 522.800 409.000 531.400 409.600 ;
        RECT 522.800 408.800 523.600 409.000 ;
        RECT 514.600 407.600 517.200 408.400 ;
        RECT 511.400 406.800 514.000 407.400 ;
        RECT 513.200 402.200 514.000 406.800 ;
        RECT 516.400 402.200 517.200 407.600 ;
        RECT 517.800 406.800 522.000 407.600 ;
        RECT 519.600 402.200 520.400 405.000 ;
        RECT 521.200 402.200 522.000 405.000 ;
        RECT 522.800 402.200 523.600 405.000 ;
        RECT 524.400 402.200 525.200 408.400 ;
        RECT 527.600 407.600 530.200 408.400 ;
        RECT 530.800 408.200 531.400 409.000 ;
        RECT 532.400 409.400 533.200 409.600 ;
        RECT 532.400 409.000 537.800 409.400 ;
        RECT 532.400 408.800 538.600 409.000 ;
        RECT 537.200 408.200 538.600 408.800 ;
        RECT 530.800 407.600 536.600 408.200 ;
        RECT 539.600 408.000 541.200 408.800 ;
        RECT 539.600 407.600 540.200 408.000 ;
        RECT 527.600 402.200 528.400 407.000 ;
        RECT 530.800 402.200 531.600 407.000 ;
        RECT 536.000 406.800 540.200 407.600 ;
        RECT 542.000 407.400 542.800 413.000 ;
        RECT 545.000 415.800 546.000 416.400 ;
        RECT 545.000 414.400 545.600 415.800 ;
        RECT 548.400 415.200 549.200 419.800 ;
        RECT 550.000 416.000 550.800 419.800 ;
        RECT 553.200 416.000 554.000 419.800 ;
        RECT 550.000 415.800 554.000 416.000 ;
        RECT 554.800 415.800 555.600 419.800 ;
        RECT 550.200 415.400 553.800 415.800 ;
        RECT 546.600 414.600 549.200 415.200 ;
        RECT 545.000 413.600 546.000 414.400 ;
        RECT 545.000 410.200 545.600 413.600 ;
        RECT 546.600 413.000 547.200 414.600 ;
        RECT 550.800 414.400 551.600 414.800 ;
        RECT 554.800 414.400 555.400 415.800 ;
        RECT 550.000 413.800 551.600 414.400 ;
        RECT 550.000 413.600 550.800 413.800 ;
        RECT 553.000 413.600 555.600 414.400 ;
        RECT 546.200 412.200 547.200 413.000 ;
        RECT 546.600 410.200 547.200 412.200 ;
        RECT 548.200 412.400 549.000 413.200 ;
        RECT 548.200 411.600 549.200 412.400 ;
        RECT 551.600 411.600 552.400 413.200 ;
        RECT 553.000 410.200 553.600 413.600 ;
        RECT 554.800 410.200 555.600 410.400 ;
        RECT 545.000 409.200 546.000 410.200 ;
        RECT 546.600 409.600 549.200 410.200 ;
        RECT 540.800 406.800 542.800 407.400 ;
        RECT 532.400 402.200 533.200 405.000 ;
        RECT 534.000 402.200 534.800 405.000 ;
        RECT 537.200 402.200 538.000 406.800 ;
        RECT 540.800 406.200 541.400 406.800 ;
        RECT 540.400 405.600 541.400 406.200 ;
        RECT 540.400 402.200 541.200 405.600 ;
        RECT 545.200 402.200 546.000 409.200 ;
        RECT 548.400 402.200 549.200 409.600 ;
        RECT 552.600 409.600 553.600 410.200 ;
        RECT 554.200 409.600 555.600 410.200 ;
        RECT 552.600 402.200 553.400 409.600 ;
        RECT 554.200 408.400 554.800 409.600 ;
        RECT 554.000 407.600 554.800 408.400 ;
        RECT 556.400 402.200 557.200 419.800 ;
        RECT 558.000 415.600 558.800 417.200 ;
        RECT 559.600 415.800 560.400 419.800 ;
        RECT 561.200 416.000 562.000 419.800 ;
        RECT 564.400 416.000 565.200 419.800 ;
        RECT 561.200 415.800 565.200 416.000 ;
        RECT 566.000 416.000 566.800 419.800 ;
        RECT 569.200 416.000 570.000 419.800 ;
        RECT 566.000 415.800 570.000 416.000 ;
        RECT 570.800 415.800 571.600 419.800 ;
        RECT 578.800 416.000 579.600 419.800 ;
        RECT 559.800 414.400 560.400 415.800 ;
        RECT 561.400 415.400 565.000 415.800 ;
        RECT 566.200 415.400 569.800 415.800 ;
        RECT 563.600 414.400 564.400 414.800 ;
        RECT 566.800 414.400 567.600 414.800 ;
        RECT 570.800 414.400 571.400 415.800 ;
        RECT 578.600 415.200 579.600 416.000 ;
        RECT 559.600 413.600 562.200 414.400 ;
        RECT 563.600 413.800 565.200 414.400 ;
        RECT 564.400 413.600 565.200 413.800 ;
        RECT 566.000 413.800 567.600 414.400 ;
        RECT 566.000 413.600 566.800 413.800 ;
        RECT 569.000 413.600 571.600 414.400 ;
        RECT 559.600 410.200 560.400 410.400 ;
        RECT 561.600 410.200 562.200 413.600 ;
        RECT 562.800 411.600 563.600 413.200 ;
        RECT 567.600 411.600 568.400 413.200 ;
        RECT 569.000 410.200 569.600 413.600 ;
        RECT 578.600 410.800 579.400 415.200 ;
        RECT 580.400 414.600 581.200 419.800 ;
        RECT 586.800 416.600 587.600 419.800 ;
        RECT 588.400 417.000 589.200 419.800 ;
        RECT 590.000 417.000 590.800 419.800 ;
        RECT 591.600 417.000 592.400 419.800 ;
        RECT 593.200 417.000 594.000 419.800 ;
        RECT 596.400 417.000 597.200 419.800 ;
        RECT 599.600 417.000 600.400 419.800 ;
        RECT 601.200 417.000 602.000 419.800 ;
        RECT 602.800 417.000 603.600 419.800 ;
        RECT 585.200 415.800 587.600 416.600 ;
        RECT 604.400 416.600 605.200 419.800 ;
        RECT 585.200 415.200 586.000 415.800 ;
        RECT 580.000 414.000 581.200 414.600 ;
        RECT 584.200 414.600 586.000 415.200 ;
        RECT 590.000 415.600 591.000 416.400 ;
        RECT 594.000 415.600 595.600 416.400 ;
        RECT 596.400 415.800 601.000 416.400 ;
        RECT 604.400 415.800 607.000 416.600 ;
        RECT 596.400 415.600 597.200 415.800 ;
        RECT 580.000 412.000 580.600 414.000 ;
        RECT 584.200 413.400 585.000 414.600 ;
        RECT 581.200 412.600 585.000 413.400 ;
        RECT 590.000 412.800 590.800 415.600 ;
        RECT 596.400 414.800 597.200 415.000 ;
        RECT 592.800 414.200 597.200 414.800 ;
        RECT 592.800 414.000 593.600 414.200 ;
        RECT 598.000 413.600 598.800 415.200 ;
        RECT 600.200 413.400 601.000 415.800 ;
        RECT 606.200 415.200 607.000 415.800 ;
        RECT 606.200 414.400 609.200 415.200 ;
        RECT 610.800 413.800 611.600 419.800 ;
        RECT 612.400 415.800 613.200 419.800 ;
        RECT 616.800 418.400 618.400 419.800 ;
        RECT 616.800 417.600 619.600 418.400 ;
        RECT 616.800 416.200 618.400 417.600 ;
        RECT 612.400 415.200 614.600 415.800 ;
        RECT 615.600 415.400 617.200 415.600 ;
        RECT 613.800 415.000 614.600 415.200 ;
        RECT 615.200 414.800 617.200 415.400 ;
        RECT 615.200 414.400 615.800 414.800 ;
        RECT 593.200 412.600 596.400 413.400 ;
        RECT 600.200 412.600 602.200 413.400 ;
        RECT 602.800 413.000 611.600 413.800 ;
        RECT 612.400 413.800 615.800 414.400 ;
        RECT 612.400 413.600 614.000 413.800 ;
        RECT 586.800 412.000 587.600 412.600 ;
        RECT 604.400 412.000 605.200 412.400 ;
        RECT 609.200 412.200 610.000 412.400 ;
        RECT 609.200 412.000 610.200 412.200 ;
        RECT 580.000 411.400 580.800 412.000 ;
        RECT 586.800 411.400 610.200 412.000 ;
        RECT 570.800 410.200 571.600 410.400 ;
        RECT 559.600 409.600 561.000 410.200 ;
        RECT 561.600 409.600 562.600 410.200 ;
        RECT 560.400 408.400 561.000 409.600 ;
        RECT 560.400 407.600 561.200 408.400 ;
        RECT 561.800 402.200 562.600 409.600 ;
        RECT 568.600 409.600 569.600 410.200 ;
        RECT 570.200 409.600 571.600 410.200 ;
        RECT 578.600 410.000 579.600 410.800 ;
        RECT 568.600 402.200 569.400 409.600 ;
        RECT 570.200 408.400 570.800 409.600 ;
        RECT 570.000 407.600 570.800 408.400 ;
        RECT 575.600 408.300 576.400 408.400 ;
        RECT 578.800 408.300 579.600 410.000 ;
        RECT 575.600 407.700 579.600 408.300 ;
        RECT 575.600 407.600 576.400 407.700 ;
        RECT 578.800 402.200 579.600 407.700 ;
        RECT 580.200 409.600 580.800 411.400 ;
        RECT 580.200 409.000 589.200 409.600 ;
        RECT 580.200 407.400 580.800 409.000 ;
        RECT 588.400 408.800 589.200 409.000 ;
        RECT 591.600 409.000 600.200 409.600 ;
        RECT 591.600 408.800 592.400 409.000 ;
        RECT 583.400 407.600 586.000 408.400 ;
        RECT 580.200 406.800 582.800 407.400 ;
        RECT 582.000 402.200 582.800 406.800 ;
        RECT 585.200 402.200 586.000 407.600 ;
        RECT 586.600 406.800 590.800 407.600 ;
        RECT 588.400 402.200 589.200 405.000 ;
        RECT 590.000 402.200 590.800 405.000 ;
        RECT 591.600 402.200 592.400 405.000 ;
        RECT 593.200 402.200 594.000 408.400 ;
        RECT 596.400 407.600 599.000 408.400 ;
        RECT 599.600 408.200 600.200 409.000 ;
        RECT 601.200 409.400 602.000 409.600 ;
        RECT 601.200 409.000 606.600 409.400 ;
        RECT 601.200 408.800 607.400 409.000 ;
        RECT 606.000 408.200 607.400 408.800 ;
        RECT 599.600 407.600 605.400 408.200 ;
        RECT 608.400 408.000 610.000 408.800 ;
        RECT 608.400 407.600 609.000 408.000 ;
        RECT 596.400 402.200 597.200 407.000 ;
        RECT 599.600 402.200 600.400 407.000 ;
        RECT 604.800 406.800 609.000 407.600 ;
        RECT 610.800 407.400 611.600 413.000 ;
        RECT 616.400 413.400 617.200 414.200 ;
        RECT 616.400 412.800 617.000 413.400 ;
        RECT 614.400 412.200 617.000 412.800 ;
        RECT 617.800 412.800 618.400 416.200 ;
        RECT 622.000 415.800 622.800 419.800 ;
        RECT 624.200 416.400 625.000 419.800 ;
        RECT 624.200 415.800 626.000 416.400 ;
        RECT 619.000 414.800 619.800 415.600 ;
        RECT 620.400 415.200 622.800 415.800 ;
        RECT 620.400 415.000 621.200 415.200 ;
        RECT 619.200 414.400 619.800 414.800 ;
        RECT 619.200 413.600 620.000 414.400 ;
        RECT 621.200 413.600 622.800 414.400 ;
        RECT 617.800 412.400 618.800 412.800 ;
        RECT 617.800 412.200 619.600 412.400 ;
        RECT 614.400 412.000 615.200 412.200 ;
        RECT 618.200 411.600 619.600 412.200 ;
        RECT 622.000 412.300 622.800 412.400 ;
        RECT 625.200 412.300 626.000 415.800 ;
        RECT 626.800 413.600 627.600 415.200 ;
        RECT 628.400 413.600 629.200 415.200 ;
        RECT 630.000 414.300 630.800 419.800 ;
        RECT 631.600 416.000 632.400 419.800 ;
        RECT 634.800 416.000 635.600 419.800 ;
        RECT 631.600 415.800 635.600 416.000 ;
        RECT 636.400 415.800 637.200 419.800 ;
        RECT 638.000 415.800 638.800 419.800 ;
        RECT 642.400 418.400 644.000 419.800 ;
        RECT 642.400 417.600 645.200 418.400 ;
        RECT 642.400 416.200 644.000 417.600 ;
        RECT 631.800 415.400 635.400 415.800 ;
        RECT 632.400 414.400 633.200 414.800 ;
        RECT 636.400 414.400 637.000 415.800 ;
        RECT 638.000 415.200 640.200 415.800 ;
        RECT 641.200 415.400 642.800 415.600 ;
        RECT 639.400 415.000 640.200 415.200 ;
        RECT 640.800 414.800 642.800 415.400 ;
        RECT 640.800 414.400 641.400 414.800 ;
        RECT 631.600 414.300 633.200 414.400 ;
        RECT 630.000 413.800 633.200 414.300 ;
        RECT 630.000 413.700 632.400 413.800 ;
        RECT 622.000 411.700 626.000 412.300 ;
        RECT 622.000 411.600 622.800 411.700 ;
        RECT 616.600 411.400 617.400 411.600 ;
        RECT 614.000 410.800 617.400 411.400 ;
        RECT 614.000 410.200 614.600 410.800 ;
        RECT 618.200 410.200 618.800 411.600 ;
        RECT 609.600 406.800 611.600 407.400 ;
        RECT 612.400 409.600 614.600 410.200 ;
        RECT 601.200 402.200 602.000 405.000 ;
        RECT 602.800 402.200 603.600 405.000 ;
        RECT 606.000 402.200 606.800 406.800 ;
        RECT 609.600 406.200 610.200 406.800 ;
        RECT 609.200 405.600 610.200 406.200 ;
        RECT 609.200 402.200 610.000 405.600 ;
        RECT 612.400 402.200 613.200 409.600 ;
        RECT 613.800 409.400 614.600 409.600 ;
        RECT 616.800 409.600 618.800 410.200 ;
        RECT 620.400 409.600 622.800 410.200 ;
        RECT 616.800 402.200 618.400 409.600 ;
        RECT 620.400 409.400 621.200 409.600 ;
        RECT 622.000 402.200 622.800 409.600 ;
        RECT 623.600 408.800 624.400 410.400 ;
        RECT 625.200 402.200 626.000 411.700 ;
        RECT 630.000 402.200 630.800 413.700 ;
        RECT 631.600 413.600 632.400 413.700 ;
        RECT 634.600 413.600 637.200 414.400 ;
        RECT 638.000 413.800 641.400 414.400 ;
        RECT 638.000 413.600 639.600 413.800 ;
        RECT 633.200 411.600 634.000 413.200 ;
        RECT 634.600 410.200 635.200 413.600 ;
        RECT 642.000 413.400 642.800 414.200 ;
        RECT 642.000 412.800 642.600 413.400 ;
        RECT 640.000 412.200 642.600 412.800 ;
        RECT 643.400 412.800 644.000 416.200 ;
        RECT 647.600 415.800 648.400 419.800 ;
        RECT 650.800 416.000 651.600 419.800 ;
        RECT 644.600 414.800 645.400 415.600 ;
        RECT 646.000 415.200 648.400 415.800 ;
        RECT 650.600 415.200 651.600 416.000 ;
        RECT 646.000 415.000 646.800 415.200 ;
        RECT 644.800 414.400 645.400 414.800 ;
        RECT 644.800 413.600 645.600 414.400 ;
        RECT 646.800 413.600 648.400 414.400 ;
        RECT 643.400 412.400 644.400 412.800 ;
        RECT 643.400 412.200 645.200 412.400 ;
        RECT 640.000 412.000 640.800 412.200 ;
        RECT 643.800 411.600 645.200 412.200 ;
        RECT 642.200 411.400 643.000 411.600 ;
        RECT 639.600 410.800 643.000 411.400 ;
        RECT 636.400 410.200 637.200 410.400 ;
        RECT 639.600 410.200 640.200 410.800 ;
        RECT 643.800 410.200 644.400 411.600 ;
        RECT 650.600 410.800 651.400 415.200 ;
        RECT 652.400 414.600 653.200 419.800 ;
        RECT 658.800 416.600 659.600 419.800 ;
        RECT 660.400 417.000 661.200 419.800 ;
        RECT 662.000 417.000 662.800 419.800 ;
        RECT 663.600 417.000 664.400 419.800 ;
        RECT 665.200 417.000 666.000 419.800 ;
        RECT 668.400 417.000 669.200 419.800 ;
        RECT 671.600 417.000 672.400 419.800 ;
        RECT 673.200 417.000 674.000 419.800 ;
        RECT 674.800 417.000 675.600 419.800 ;
        RECT 657.200 415.800 659.600 416.600 ;
        RECT 676.400 416.600 677.200 419.800 ;
        RECT 657.200 415.200 658.000 415.800 ;
        RECT 652.000 414.000 653.200 414.600 ;
        RECT 656.200 414.600 658.000 415.200 ;
        RECT 662.000 415.600 663.000 416.400 ;
        RECT 666.000 415.600 667.600 416.400 ;
        RECT 668.400 415.800 673.000 416.400 ;
        RECT 676.400 415.800 679.000 416.600 ;
        RECT 668.400 415.600 669.200 415.800 ;
        RECT 652.000 412.000 652.600 414.000 ;
        RECT 656.200 413.400 657.000 414.600 ;
        RECT 653.200 412.600 657.000 413.400 ;
        RECT 662.000 412.800 662.800 415.600 ;
        RECT 668.400 414.800 669.200 415.000 ;
        RECT 664.800 414.200 669.200 414.800 ;
        RECT 664.800 414.000 665.600 414.200 ;
        RECT 670.000 413.600 670.800 415.200 ;
        RECT 672.200 413.400 673.000 415.800 ;
        RECT 678.200 415.200 679.000 415.800 ;
        RECT 678.200 414.400 681.200 415.200 ;
        RECT 682.800 413.800 683.600 419.800 ;
        RECT 665.200 412.600 668.400 413.400 ;
        RECT 672.200 412.600 674.200 413.400 ;
        RECT 674.800 413.000 683.600 413.800 ;
        RECT 658.800 412.000 659.600 412.600 ;
        RECT 676.400 412.000 677.200 412.400 ;
        RECT 679.600 412.000 680.400 412.400 ;
        RECT 681.400 412.000 682.200 412.200 ;
        RECT 652.000 411.400 652.800 412.000 ;
        RECT 658.800 411.400 682.200 412.000 ;
        RECT 634.200 409.600 635.200 410.200 ;
        RECT 635.800 409.600 637.200 410.200 ;
        RECT 638.000 409.600 640.200 410.200 ;
        RECT 634.200 404.400 635.000 409.600 ;
        RECT 635.800 408.400 636.400 409.600 ;
        RECT 635.600 407.600 636.400 408.400 ;
        RECT 633.200 403.600 635.000 404.400 ;
        RECT 634.200 402.200 635.000 403.600 ;
        RECT 638.000 402.200 638.800 409.600 ;
        RECT 639.400 409.400 640.200 409.600 ;
        RECT 642.400 409.600 644.400 410.200 ;
        RECT 646.000 409.600 648.400 410.200 ;
        RECT 650.600 410.000 651.600 410.800 ;
        RECT 642.400 402.200 644.000 409.600 ;
        RECT 646.000 409.400 646.800 409.600 ;
        RECT 647.600 402.200 648.400 409.600 ;
        RECT 650.800 402.200 651.600 410.000 ;
        RECT 652.200 409.600 652.800 411.400 ;
        RECT 652.200 409.000 661.200 409.600 ;
        RECT 652.200 407.400 652.800 409.000 ;
        RECT 660.400 408.800 661.200 409.000 ;
        RECT 663.600 409.000 672.200 409.600 ;
        RECT 663.600 408.800 664.400 409.000 ;
        RECT 655.400 407.600 658.000 408.400 ;
        RECT 652.200 406.800 654.800 407.400 ;
        RECT 654.000 402.200 654.800 406.800 ;
        RECT 657.200 402.200 658.000 407.600 ;
        RECT 658.600 406.800 662.800 407.600 ;
        RECT 660.400 402.200 661.200 405.000 ;
        RECT 662.000 402.200 662.800 405.000 ;
        RECT 663.600 402.200 664.400 405.000 ;
        RECT 665.200 402.200 666.000 408.400 ;
        RECT 668.400 407.600 671.000 408.400 ;
        RECT 671.600 408.200 672.200 409.000 ;
        RECT 673.200 409.400 674.000 409.600 ;
        RECT 673.200 409.000 678.600 409.400 ;
        RECT 673.200 408.800 679.400 409.000 ;
        RECT 678.000 408.200 679.400 408.800 ;
        RECT 671.600 407.600 677.400 408.200 ;
        RECT 680.400 408.000 682.000 408.800 ;
        RECT 680.400 407.600 681.000 408.000 ;
        RECT 668.400 402.200 669.200 407.000 ;
        RECT 671.600 402.200 672.400 407.000 ;
        RECT 676.800 406.800 681.000 407.600 ;
        RECT 682.800 407.400 683.600 413.000 ;
        RECT 681.600 406.800 683.600 407.400 ;
        RECT 673.200 402.200 674.000 405.000 ;
        RECT 674.800 402.200 675.600 405.000 ;
        RECT 678.000 402.200 678.800 406.800 ;
        RECT 681.600 406.200 682.200 406.800 ;
        RECT 681.200 405.600 682.200 406.200 ;
        RECT 681.200 402.200 682.000 405.600 ;
        RECT 4.400 392.400 5.200 399.800 ;
        RECT 3.000 391.800 5.200 392.400 ;
        RECT 3.000 391.200 3.600 391.800 ;
        RECT 2.400 390.400 3.600 391.200 ;
        RECT 6.000 391.400 6.800 399.800 ;
        RECT 10.400 396.400 11.200 399.800 ;
        RECT 9.200 395.800 11.200 396.400 ;
        RECT 14.800 395.800 15.600 399.800 ;
        RECT 19.000 395.800 20.200 399.800 ;
        RECT 9.200 395.000 10.000 395.800 ;
        RECT 14.800 395.200 15.400 395.800 ;
        RECT 12.600 394.600 16.200 395.200 ;
        RECT 18.800 395.000 19.600 395.800 ;
        RECT 12.600 394.400 13.400 394.600 ;
        RECT 15.400 394.400 16.200 394.600 ;
        RECT 9.200 393.000 10.000 393.200 ;
        RECT 13.800 393.000 14.600 393.200 ;
        RECT 9.200 392.400 14.600 393.000 ;
        RECT 15.200 393.000 17.400 393.600 ;
        RECT 15.200 391.800 15.800 393.000 ;
        RECT 16.600 392.800 17.400 393.000 ;
        RECT 19.000 393.200 20.400 394.000 ;
        RECT 19.000 392.200 19.600 393.200 ;
        RECT 11.000 391.400 15.800 391.800 ;
        RECT 6.000 391.200 15.800 391.400 ;
        RECT 17.200 391.600 19.600 392.200 ;
        RECT 6.000 391.000 11.800 391.200 ;
        RECT 6.000 390.800 11.600 391.000 ;
        RECT 3.000 387.400 3.600 390.400 ;
        RECT 4.400 388.800 5.200 390.400 ;
        RECT 12.400 390.300 13.200 390.400 ;
        RECT 14.000 390.300 14.800 390.400 ;
        RECT 12.400 390.200 14.800 390.300 ;
        RECT 8.200 389.700 14.800 390.200 ;
        RECT 8.200 389.600 13.200 389.700 ;
        RECT 14.000 389.600 14.800 389.700 ;
        RECT 8.200 389.400 9.000 389.600 ;
        RECT 9.800 388.400 10.600 388.600 ;
        RECT 17.200 388.400 17.800 391.600 ;
        RECT 23.600 391.200 24.400 399.800 ;
        RECT 27.400 398.400 28.200 399.800 ;
        RECT 27.400 397.600 29.200 398.400 ;
        RECT 26.000 393.600 26.800 394.400 ;
        RECT 26.000 392.400 26.600 393.600 ;
        RECT 27.400 392.400 28.200 397.600 ;
        RECT 33.200 392.800 34.000 399.800 ;
        RECT 25.200 391.800 26.600 392.400 ;
        RECT 27.200 391.800 28.200 392.400 ;
        RECT 33.000 391.800 34.000 392.800 ;
        RECT 36.400 392.400 37.200 399.800 ;
        RECT 34.600 391.800 37.200 392.400 ;
        RECT 40.600 392.400 41.400 399.800 ;
        RECT 46.600 394.400 47.400 399.800 ;
        RECT 42.000 393.600 42.800 394.400 ;
        RECT 42.200 392.400 42.800 393.600 ;
        RECT 45.200 393.600 46.000 394.400 ;
        RECT 46.600 393.600 48.400 394.400 ;
        RECT 45.200 392.400 45.800 393.600 ;
        RECT 46.600 392.400 47.400 393.600 ;
        RECT 54.600 392.800 55.400 399.800 ;
        RECT 58.800 395.000 59.600 399.000 ;
        RECT 64.200 398.400 65.000 399.800 ;
        RECT 63.600 397.600 65.000 398.400 ;
        RECT 40.600 391.800 41.600 392.400 ;
        RECT 42.200 391.800 43.600 392.400 ;
        RECT 25.200 391.600 26.000 391.800 ;
        RECT 20.200 390.600 24.400 391.200 ;
        RECT 20.200 390.400 21.000 390.600 ;
        RECT 21.800 389.800 22.600 390.000 ;
        RECT 18.800 389.200 22.600 389.800 ;
        RECT 18.800 389.000 19.600 389.200 ;
        RECT 6.800 387.800 17.800 388.400 ;
        RECT 6.800 387.600 8.400 387.800 ;
        RECT 3.000 386.800 5.200 387.400 ;
        RECT 4.400 382.200 5.200 386.800 ;
        RECT 6.000 382.200 6.800 387.000 ;
        RECT 11.000 385.600 11.600 387.800 ;
        RECT 12.400 387.600 13.200 387.800 ;
        RECT 16.600 387.600 17.400 387.800 ;
        RECT 23.600 387.200 24.400 390.600 ;
        RECT 27.200 388.400 27.800 391.800 ;
        RECT 28.400 390.300 29.200 390.400 ;
        RECT 28.400 389.700 32.300 390.300 ;
        RECT 28.400 388.800 29.200 389.700 ;
        RECT 25.200 387.600 27.800 388.400 ;
        RECT 30.000 388.200 30.800 388.400 ;
        RECT 29.200 387.600 30.800 388.200 ;
        RECT 31.700 388.300 32.300 389.700 ;
        RECT 33.000 388.400 33.600 391.800 ;
        RECT 34.600 389.800 35.200 391.800 ;
        RECT 34.200 389.000 35.200 389.800 ;
        RECT 33.000 388.300 34.000 388.400 ;
        RECT 31.700 387.700 34.000 388.300 ;
        RECT 33.000 387.600 34.000 387.700 ;
        RECT 20.600 386.600 24.400 387.200 ;
        RECT 20.600 386.400 21.400 386.600 ;
        RECT 9.200 384.200 10.000 385.000 ;
        RECT 10.800 384.800 11.600 385.600 ;
        RECT 12.600 385.400 13.400 385.600 ;
        RECT 12.600 384.800 15.400 385.400 ;
        RECT 14.800 384.200 15.400 384.800 ;
        RECT 18.800 384.200 19.600 385.000 ;
        RECT 9.200 383.600 11.200 384.200 ;
        RECT 10.400 382.200 11.200 383.600 ;
        RECT 14.800 382.200 15.600 384.200 ;
        RECT 18.800 383.600 20.200 384.200 ;
        RECT 19.000 382.200 20.200 383.600 ;
        RECT 23.600 382.200 24.400 386.600 ;
        RECT 25.400 386.200 26.000 387.600 ;
        RECT 29.200 387.200 30.000 387.600 ;
        RECT 27.000 386.200 30.600 386.600 ;
        RECT 33.000 386.200 33.600 387.600 ;
        RECT 34.600 387.400 35.200 389.000 ;
        RECT 36.200 389.600 37.200 390.400 ;
        RECT 36.200 388.800 37.000 389.600 ;
        RECT 39.600 388.800 40.400 390.400 ;
        RECT 41.000 390.300 41.600 391.800 ;
        RECT 42.800 391.600 43.600 391.800 ;
        RECT 44.400 391.800 45.800 392.400 ;
        RECT 46.400 391.800 47.400 392.400 ;
        RECT 53.800 392.200 55.400 392.800 ;
        RECT 44.400 391.600 45.200 391.800 ;
        RECT 44.500 390.300 45.100 391.600 ;
        RECT 41.000 389.700 45.100 390.300 ;
        RECT 41.000 388.400 41.600 389.700 ;
        RECT 46.400 388.400 47.000 391.800 ;
        RECT 47.600 388.800 48.400 390.400 ;
        RECT 49.200 390.300 50.000 390.400 ;
        RECT 52.400 390.300 53.200 391.200 ;
        RECT 49.200 389.700 53.200 390.300 ;
        RECT 49.200 389.600 50.000 389.700 ;
        RECT 52.400 389.600 53.200 389.700 ;
        RECT 53.800 388.400 54.400 392.200 ;
        RECT 59.000 391.600 59.600 395.000 ;
        RECT 64.200 392.800 65.000 397.600 ;
        RECT 68.400 395.000 69.200 399.000 ;
        RECT 55.800 391.000 59.600 391.600 ;
        RECT 63.400 392.200 65.000 392.800 ;
        RECT 55.800 389.000 56.400 391.000 ;
        RECT 38.000 388.200 38.800 388.400 ;
        RECT 38.000 387.600 39.600 388.200 ;
        RECT 41.000 387.600 43.600 388.400 ;
        RECT 44.400 387.600 47.000 388.400 ;
        RECT 49.200 388.300 50.000 388.400 ;
        RECT 50.800 388.300 51.600 388.400 ;
        RECT 49.200 388.200 51.600 388.300 ;
        RECT 48.400 387.700 51.600 388.200 ;
        RECT 48.400 387.600 50.000 387.700 ;
        RECT 50.800 387.600 51.600 387.700 ;
        RECT 52.400 387.600 54.400 388.400 ;
        RECT 55.000 388.200 56.400 389.000 ;
        RECT 57.200 388.800 58.000 390.400 ;
        RECT 58.800 388.800 59.600 390.400 ;
        RECT 60.400 390.300 61.200 390.400 ;
        RECT 62.000 390.300 62.800 391.200 ;
        RECT 60.400 389.700 62.800 390.300 ;
        RECT 60.400 389.600 61.200 389.700 ;
        RECT 62.000 389.600 62.800 389.700 ;
        RECT 63.400 388.400 64.000 392.200 ;
        RECT 68.600 391.600 69.200 395.000 ;
        RECT 65.400 391.000 69.200 391.600 ;
        RECT 65.400 389.000 66.000 391.000 ;
        RECT 34.600 386.800 37.200 387.400 ;
        RECT 38.800 387.200 39.600 387.600 ;
        RECT 25.200 382.200 26.000 386.200 ;
        RECT 26.800 386.000 30.800 386.200 ;
        RECT 26.800 382.200 27.600 386.000 ;
        RECT 30.000 382.200 30.800 386.000 ;
        RECT 33.000 385.600 34.000 386.200 ;
        RECT 33.200 382.200 34.000 385.600 ;
        RECT 36.400 382.200 37.200 386.800 ;
        RECT 38.200 386.200 41.800 386.600 ;
        RECT 42.800 386.200 43.400 387.600 ;
        RECT 44.600 386.200 45.200 387.600 ;
        RECT 48.400 387.200 49.200 387.600 ;
        RECT 53.800 387.000 54.400 387.600 ;
        RECT 55.400 387.800 56.400 388.200 ;
        RECT 55.400 387.200 59.600 387.800 ;
        RECT 62.000 387.600 64.000 388.400 ;
        RECT 64.600 388.200 66.000 389.000 ;
        RECT 66.800 388.800 67.600 390.400 ;
        RECT 68.400 388.800 69.200 390.400 ;
        RECT 53.800 386.600 54.600 387.000 ;
        RECT 46.200 386.200 49.800 386.600 ;
        RECT 38.000 386.000 42.000 386.200 ;
        RECT 38.000 382.200 38.800 386.000 ;
        RECT 41.200 382.200 42.000 386.000 ;
        RECT 42.800 382.200 43.600 386.200 ;
        RECT 44.400 382.200 45.200 386.200 ;
        RECT 46.000 386.000 50.000 386.200 ;
        RECT 53.800 386.000 55.400 386.600 ;
        RECT 46.000 382.200 46.800 386.000 ;
        RECT 49.200 382.200 50.000 386.000 ;
        RECT 54.600 383.000 55.400 386.000 ;
        RECT 59.000 385.000 59.600 387.200 ;
        RECT 63.400 387.000 64.000 387.600 ;
        RECT 65.000 387.800 66.000 388.200 ;
        RECT 65.000 387.200 69.200 387.800 ;
        RECT 63.400 386.600 64.200 387.000 ;
        RECT 63.400 386.000 65.000 386.600 ;
        RECT 58.800 383.000 59.600 385.000 ;
        RECT 64.200 383.000 65.000 386.000 ;
        RECT 68.600 385.000 69.200 387.200 ;
        RECT 68.400 383.000 69.200 385.000 ;
        RECT 70.000 384.800 70.800 386.400 ;
        RECT 71.600 382.200 72.400 399.800 ;
        RECT 74.800 392.800 75.600 399.800 ;
        RECT 74.600 391.800 75.600 392.800 ;
        RECT 78.000 392.400 78.800 399.800 ;
        RECT 76.200 391.800 78.800 392.400 ;
        RECT 74.600 388.400 75.200 391.800 ;
        RECT 76.200 389.800 76.800 391.800 ;
        RECT 75.800 389.000 76.800 389.800 ;
        RECT 74.600 387.600 75.600 388.400 ;
        RECT 74.600 386.200 75.200 387.600 ;
        RECT 76.200 387.400 76.800 389.000 ;
        RECT 77.800 389.600 78.800 390.400 ;
        RECT 77.800 388.800 78.600 389.600 ;
        RECT 76.200 386.800 78.800 387.400 ;
        RECT 79.600 386.800 80.400 388.400 ;
        RECT 74.600 385.600 75.600 386.200 ;
        RECT 74.800 382.200 75.600 385.600 ;
        RECT 78.000 382.200 78.800 386.800 ;
        RECT 81.200 386.200 82.000 399.800 ;
        RECT 82.800 391.600 83.600 393.200 ;
        RECT 84.400 392.400 85.200 399.800 ;
        RECT 87.600 392.800 88.400 399.800 ;
        RECT 91.600 393.600 92.400 394.400 ;
        RECT 84.400 391.800 87.000 392.400 ;
        RECT 87.600 391.800 88.600 392.800 ;
        RECT 91.600 392.400 92.200 393.600 ;
        RECT 93.000 392.400 93.800 399.800 ;
        RECT 98.800 392.800 99.600 399.800 ;
        RECT 84.400 389.600 85.400 390.400 ;
        RECT 84.600 388.800 85.400 389.600 ;
        RECT 86.400 389.800 87.000 391.800 ;
        RECT 86.400 389.000 87.400 389.800 ;
        RECT 86.400 387.400 87.000 389.000 ;
        RECT 88.000 388.400 88.600 391.800 ;
        RECT 90.800 391.800 92.200 392.400 ;
        RECT 92.800 391.800 93.800 392.400 ;
        RECT 98.600 391.800 99.600 392.800 ;
        RECT 102.000 392.400 102.800 399.800 ;
        RECT 100.200 391.800 102.800 392.400 ;
        RECT 106.200 392.400 107.000 399.800 ;
        RECT 107.600 393.600 108.400 394.400 ;
        RECT 107.800 392.400 108.400 393.600 ;
        RECT 117.400 392.600 118.200 399.800 ;
        RECT 122.200 398.400 123.000 399.800 ;
        RECT 121.200 397.600 123.000 398.400 ;
        RECT 106.200 391.800 107.200 392.400 ;
        RECT 107.800 391.800 109.200 392.400 ;
        RECT 116.400 391.800 118.200 392.600 ;
        RECT 122.200 392.400 123.000 397.600 ;
        RECT 123.600 393.600 124.400 394.400 ;
        RECT 123.800 392.400 124.400 393.600 ;
        RECT 126.800 393.600 127.600 394.400 ;
        RECT 126.800 392.400 127.400 393.600 ;
        RECT 128.200 392.400 129.000 399.800 ;
        RECT 132.400 395.600 133.200 399.800 ;
        RECT 135.600 395.800 136.400 399.800 ;
        RECT 135.600 395.600 136.200 395.800 ;
        RECT 132.600 395.000 136.200 395.600 ;
        RECT 132.600 392.400 133.200 395.000 ;
        RECT 134.000 392.800 134.800 394.400 ;
        RECT 139.600 393.600 140.400 394.400 ;
        RECT 139.600 392.400 140.200 393.600 ;
        RECT 141.000 392.400 141.800 399.800 ;
        RECT 122.200 391.800 123.200 392.400 ;
        RECT 123.800 391.800 125.200 392.400 ;
        RECT 90.800 391.600 91.600 391.800 ;
        RECT 92.800 388.400 93.400 391.800 ;
        RECT 94.000 390.300 94.800 390.400 ;
        RECT 97.200 390.300 98.000 390.400 ;
        RECT 94.000 389.700 98.000 390.300 ;
        RECT 94.000 388.800 94.800 389.700 ;
        RECT 97.200 389.600 98.000 389.700 ;
        RECT 98.600 388.400 99.200 391.800 ;
        RECT 100.200 389.800 100.800 391.800 ;
        RECT 99.800 389.000 100.800 389.800 ;
        RECT 87.600 387.600 88.600 388.400 ;
        RECT 90.800 387.600 93.400 388.400 ;
        RECT 95.600 388.200 96.400 388.400 ;
        RECT 94.800 387.600 96.400 388.200 ;
        RECT 98.600 387.600 99.600 388.400 ;
        RECT 84.400 386.800 87.000 387.400 ;
        RECT 81.200 385.600 83.000 386.200 ;
        RECT 82.200 382.200 83.000 385.600 ;
        RECT 84.400 382.200 85.200 386.800 ;
        RECT 88.000 386.200 88.600 387.600 ;
        RECT 91.000 386.200 91.600 387.600 ;
        RECT 94.800 387.200 95.600 387.600 ;
        RECT 92.600 386.200 96.200 386.600 ;
        RECT 98.600 386.200 99.200 387.600 ;
        RECT 100.200 387.400 100.800 389.000 ;
        RECT 101.800 390.300 102.800 390.400 ;
        RECT 103.600 390.300 104.400 390.400 ;
        RECT 101.800 389.700 104.400 390.300 ;
        RECT 101.800 389.600 102.800 389.700 ;
        RECT 103.600 389.600 104.400 389.700 ;
        RECT 101.800 388.800 102.600 389.600 ;
        RECT 105.200 388.800 106.000 390.400 ;
        RECT 106.600 388.400 107.200 391.800 ;
        RECT 108.400 391.600 109.200 391.800 ;
        RECT 108.400 390.300 109.200 390.400 ;
        RECT 116.600 390.300 117.200 391.800 ;
        RECT 108.400 389.700 117.200 390.300 ;
        RECT 108.400 389.600 109.200 389.700 ;
        RECT 116.600 388.400 117.200 389.700 ;
        RECT 118.000 389.600 118.800 391.200 ;
        RECT 121.200 388.800 122.000 390.400 ;
        RECT 122.600 388.400 123.200 391.800 ;
        RECT 124.400 391.600 125.200 391.800 ;
        RECT 126.000 391.800 127.400 392.400 ;
        RECT 128.000 391.800 129.000 392.400 ;
        RECT 126.000 391.600 126.800 391.800 ;
        RECT 128.000 388.400 128.600 391.800 ;
        RECT 132.400 391.600 133.200 392.400 ;
        RECT 135.600 392.300 136.400 392.400 ;
        RECT 137.200 392.300 138.000 392.400 ;
        RECT 135.600 391.700 138.000 392.300 ;
        RECT 135.600 391.600 136.400 391.700 ;
        RECT 129.200 388.800 130.000 390.400 ;
        RECT 132.600 388.400 133.200 391.600 ;
        RECT 137.200 390.800 138.000 391.700 ;
        RECT 138.800 391.800 140.200 392.400 ;
        RECT 138.800 391.600 139.600 391.800 ;
        RECT 140.800 391.600 142.800 392.400 ;
        RECT 145.200 391.600 146.000 393.200 ;
        RECT 146.800 392.300 147.600 399.800 ;
        RECT 150.800 393.600 151.600 394.400 ;
        RECT 150.800 392.400 151.400 393.600 ;
        RECT 152.200 392.400 153.000 399.800 ;
        RECT 150.000 392.300 151.400 392.400 ;
        RECT 146.800 391.800 151.400 392.300 ;
        RECT 152.000 391.800 153.000 392.400 ;
        RECT 156.400 395.000 157.200 399.000 ;
        RECT 146.800 391.700 150.800 391.800 ;
        RECT 134.800 389.600 136.400 390.400 ;
        RECT 140.800 388.400 141.400 391.600 ;
        RECT 142.000 390.300 142.800 390.400 ;
        RECT 143.600 390.300 144.400 390.400 ;
        RECT 142.000 389.700 144.400 390.300 ;
        RECT 142.000 388.800 142.800 389.700 ;
        RECT 143.600 389.600 144.400 389.700 ;
        RECT 103.600 388.200 104.400 388.400 ;
        RECT 103.600 387.600 105.200 388.200 ;
        RECT 106.600 387.600 109.200 388.400 ;
        RECT 116.400 387.600 117.200 388.400 ;
        RECT 119.600 388.200 120.400 388.400 ;
        RECT 119.600 387.600 121.200 388.200 ;
        RECT 122.600 387.600 125.200 388.400 ;
        RECT 126.000 387.600 128.600 388.400 ;
        RECT 130.800 388.200 131.600 388.400 ;
        RECT 130.000 387.600 131.600 388.200 ;
        RECT 132.600 388.200 134.200 388.400 ;
        RECT 132.600 387.800 134.400 388.200 ;
        RECT 100.200 386.800 102.800 387.400 ;
        RECT 104.400 387.200 105.200 387.600 ;
        RECT 87.600 385.600 88.600 386.200 ;
        RECT 87.600 382.200 88.400 385.600 ;
        RECT 90.800 382.200 91.600 386.200 ;
        RECT 92.400 386.000 96.400 386.200 ;
        RECT 92.400 382.200 93.200 386.000 ;
        RECT 95.600 382.200 96.400 386.000 ;
        RECT 98.600 385.600 99.600 386.200 ;
        RECT 98.800 382.200 99.600 385.600 ;
        RECT 102.000 382.200 102.800 386.800 ;
        RECT 103.800 386.200 107.400 386.600 ;
        RECT 108.400 386.200 109.000 387.600 ;
        RECT 103.600 386.000 107.600 386.200 ;
        RECT 103.600 382.200 104.400 386.000 ;
        RECT 106.800 382.200 107.600 386.000 ;
        RECT 108.400 384.300 109.200 386.200 ;
        RECT 114.800 384.800 115.600 386.400 ;
        RECT 116.600 384.400 117.200 387.600 ;
        RECT 120.400 387.200 121.200 387.600 ;
        RECT 119.800 386.200 123.400 386.600 ;
        RECT 124.400 386.200 125.000 387.600 ;
        RECT 126.200 386.200 126.800 387.600 ;
        RECT 130.000 387.200 130.800 387.600 ;
        RECT 127.800 386.200 131.400 386.600 ;
        RECT 111.600 384.300 112.400 384.400 ;
        RECT 108.400 383.700 112.400 384.300 ;
        RECT 108.400 382.200 109.200 383.700 ;
        RECT 111.600 383.600 112.400 383.700 ;
        RECT 116.400 382.200 117.200 384.400 ;
        RECT 119.600 386.000 123.600 386.200 ;
        RECT 119.600 382.200 120.400 386.000 ;
        RECT 122.800 382.200 123.600 386.000 ;
        RECT 124.400 382.200 125.200 386.200 ;
        RECT 126.000 382.200 126.800 386.200 ;
        RECT 127.600 386.000 131.600 386.200 ;
        RECT 127.600 382.200 128.400 386.000 ;
        RECT 130.800 382.200 131.600 386.000 ;
        RECT 133.600 382.200 134.400 387.800 ;
        RECT 138.800 387.600 141.400 388.400 ;
        RECT 143.600 388.200 144.400 388.400 ;
        RECT 142.800 387.600 144.400 388.200 ;
        RECT 139.000 386.200 139.600 387.600 ;
        RECT 142.800 387.200 143.600 387.600 ;
        RECT 140.600 386.200 144.200 386.600 ;
        RECT 146.800 386.200 147.600 391.700 ;
        RECT 150.000 391.600 150.800 391.700 ;
        RECT 148.400 390.300 149.200 390.400 ;
        RECT 152.000 390.300 152.600 391.800 ;
        RECT 156.400 391.600 157.000 395.000 ;
        RECT 160.600 392.800 161.400 399.800 ;
        RECT 160.600 392.200 162.200 392.800 ;
        RECT 156.400 391.000 160.200 391.600 ;
        RECT 148.400 389.700 152.600 390.300 ;
        RECT 148.400 389.600 149.200 389.700 ;
        RECT 152.000 388.400 152.600 389.700 ;
        RECT 153.200 388.800 154.000 390.400 ;
        RECT 156.400 388.800 157.200 390.400 ;
        RECT 158.000 388.800 158.800 390.400 ;
        RECT 159.600 389.000 160.200 391.000 ;
        RECT 148.400 386.800 149.200 388.400 ;
        RECT 150.000 387.600 152.600 388.400 ;
        RECT 154.800 388.200 155.600 388.400 ;
        RECT 154.000 387.600 155.600 388.200 ;
        RECT 159.600 388.200 161.000 389.000 ;
        RECT 161.600 388.400 162.200 392.200 ;
        RECT 168.600 392.400 169.400 399.800 ;
        RECT 170.000 393.600 170.800 394.400 ;
        RECT 170.200 392.400 170.800 393.600 ;
        RECT 173.200 393.600 174.000 394.400 ;
        RECT 173.200 392.400 173.800 393.600 ;
        RECT 174.600 392.400 175.400 399.800 ;
        RECT 168.600 391.800 169.600 392.400 ;
        RECT 170.200 391.800 171.600 392.400 ;
        RECT 162.800 389.600 163.600 391.200 ;
        RECT 167.600 390.300 168.400 390.400 ;
        RECT 164.500 389.700 168.400 390.300 ;
        RECT 161.600 388.300 163.600 388.400 ;
        RECT 164.500 388.300 165.100 389.700 ;
        RECT 167.600 388.800 168.400 389.700 ;
        RECT 169.000 388.400 169.600 391.800 ;
        RECT 170.800 391.600 171.600 391.800 ;
        RECT 172.400 391.800 173.800 392.400 ;
        RECT 174.400 391.800 175.400 392.400 ;
        RECT 178.800 395.000 179.600 399.000 ;
        RECT 172.400 391.600 173.200 391.800 ;
        RECT 170.900 390.300 171.500 391.600 ;
        RECT 174.400 390.300 175.000 391.800 ;
        RECT 178.800 391.600 179.400 395.000 ;
        RECT 183.000 392.800 183.800 399.800 ;
        RECT 183.000 392.200 184.600 392.800 ;
        RECT 178.800 391.000 182.600 391.600 ;
        RECT 170.900 389.700 175.000 390.300 ;
        RECT 174.400 388.400 175.000 389.700 ;
        RECT 175.600 388.800 176.400 390.400 ;
        RECT 178.800 388.800 179.600 390.400 ;
        RECT 180.400 388.800 181.200 390.400 ;
        RECT 182.000 389.000 182.600 391.000 ;
        RECT 159.600 387.800 160.600 388.200 ;
        RECT 150.200 386.200 150.800 387.600 ;
        RECT 154.000 387.200 154.800 387.600 ;
        RECT 156.400 387.200 160.600 387.800 ;
        RECT 161.600 387.700 165.100 388.300 ;
        RECT 166.000 388.200 166.800 388.400 ;
        RECT 161.600 387.600 163.600 387.700 ;
        RECT 166.000 387.600 167.600 388.200 ;
        RECT 169.000 387.600 171.600 388.400 ;
        RECT 172.400 387.600 175.000 388.400 ;
        RECT 177.200 388.200 178.000 388.400 ;
        RECT 176.400 387.600 178.000 388.200 ;
        RECT 182.000 388.200 183.400 389.000 ;
        RECT 184.000 388.400 184.600 392.200 ;
        RECT 191.000 392.400 191.800 399.800 ;
        RECT 192.400 393.600 193.200 394.400 ;
        RECT 192.600 392.400 193.200 393.600 ;
        RECT 197.400 392.400 198.200 399.800 ;
        RECT 198.800 393.600 199.600 394.400 ;
        RECT 199.000 392.400 199.600 393.600 ;
        RECT 191.000 391.800 192.000 392.400 ;
        RECT 192.600 391.800 194.000 392.400 ;
        RECT 197.400 391.800 198.400 392.400 ;
        RECT 199.000 391.800 200.400 392.400 ;
        RECT 185.200 389.600 186.000 391.200 ;
        RECT 188.400 390.300 189.200 390.400 ;
        RECT 190.000 390.300 190.800 390.400 ;
        RECT 188.400 389.700 190.800 390.300 ;
        RECT 188.400 389.600 189.200 389.700 ;
        RECT 190.000 388.800 190.800 389.700 ;
        RECT 191.400 390.300 192.000 391.800 ;
        RECT 193.200 391.600 194.000 391.800 ;
        RECT 194.800 390.300 195.600 390.400 ;
        RECT 191.400 389.700 195.600 390.300 ;
        RECT 191.400 388.400 192.000 389.700 ;
        RECT 194.800 389.600 195.600 389.700 ;
        RECT 196.400 388.800 197.200 390.400 ;
        RECT 197.800 388.400 198.400 391.800 ;
        RECT 199.600 391.600 200.400 391.800 ;
        RECT 201.200 391.200 202.000 399.800 ;
        RECT 205.400 395.800 206.600 399.800 ;
        RECT 210.000 395.800 210.800 399.800 ;
        RECT 214.400 396.400 215.200 399.800 ;
        RECT 214.400 395.800 216.400 396.400 ;
        RECT 206.000 395.000 206.800 395.800 ;
        RECT 210.200 395.200 210.800 395.800 ;
        RECT 209.400 394.600 213.000 395.200 ;
        RECT 215.600 395.000 216.400 395.800 ;
        RECT 209.400 394.400 210.200 394.600 ;
        RECT 212.200 394.400 213.000 394.600 ;
        RECT 205.200 393.200 206.600 394.000 ;
        RECT 206.000 392.200 206.600 393.200 ;
        RECT 208.200 393.000 210.400 393.600 ;
        RECT 208.200 392.800 209.000 393.000 ;
        RECT 206.000 391.600 208.400 392.200 ;
        RECT 201.200 390.600 205.400 391.200 ;
        RECT 184.000 388.300 186.000 388.400 ;
        RECT 186.800 388.300 187.600 388.400 ;
        RECT 182.000 387.800 183.000 388.200 ;
        RECT 151.800 386.200 155.400 386.600 ;
        RECT 138.800 382.200 139.600 386.200 ;
        RECT 140.400 386.000 144.400 386.200 ;
        RECT 140.400 382.200 141.200 386.000 ;
        RECT 143.600 382.200 144.400 386.000 ;
        RECT 145.800 385.600 147.600 386.200 ;
        RECT 145.800 382.200 146.600 385.600 ;
        RECT 150.000 382.200 150.800 386.200 ;
        RECT 151.600 386.000 155.600 386.200 ;
        RECT 151.600 382.200 152.400 386.000 ;
        RECT 154.800 382.200 155.600 386.000 ;
        RECT 156.400 385.000 157.000 387.200 ;
        RECT 161.600 387.000 162.200 387.600 ;
        RECT 166.800 387.200 167.600 387.600 ;
        RECT 161.400 386.600 162.200 387.000 ;
        RECT 160.600 386.000 162.200 386.600 ;
        RECT 166.200 386.200 169.800 386.600 ;
        RECT 170.800 386.200 171.400 387.600 ;
        RECT 172.600 386.200 173.200 387.600 ;
        RECT 176.400 387.200 177.200 387.600 ;
        RECT 178.800 387.200 183.000 387.800 ;
        RECT 184.000 387.700 187.600 388.300 ;
        RECT 184.000 387.600 186.000 387.700 ;
        RECT 186.800 387.600 187.600 387.700 ;
        RECT 188.400 388.200 189.200 388.400 ;
        RECT 188.400 387.600 190.000 388.200 ;
        RECT 191.400 387.600 194.000 388.400 ;
        RECT 194.800 388.200 195.600 388.400 ;
        RECT 194.800 387.600 196.400 388.200 ;
        RECT 197.800 387.600 200.400 388.400 ;
        RECT 174.200 386.200 177.800 386.600 ;
        RECT 166.000 386.000 170.000 386.200 ;
        RECT 156.400 383.000 157.200 385.000 ;
        RECT 160.600 383.000 161.400 386.000 ;
        RECT 166.000 382.200 166.800 386.000 ;
        RECT 169.200 382.200 170.000 386.000 ;
        RECT 170.800 382.200 171.600 386.200 ;
        RECT 172.400 382.200 173.200 386.200 ;
        RECT 174.000 386.000 178.000 386.200 ;
        RECT 174.000 382.200 174.800 386.000 ;
        RECT 177.200 382.200 178.000 386.000 ;
        RECT 178.800 385.000 179.400 387.200 ;
        RECT 184.000 387.000 184.600 387.600 ;
        RECT 189.200 387.200 190.000 387.600 ;
        RECT 183.800 386.600 184.600 387.000 ;
        RECT 183.000 386.000 184.600 386.600 ;
        RECT 188.600 386.200 192.200 386.600 ;
        RECT 193.200 386.200 193.800 387.600 ;
        RECT 195.600 387.200 196.400 387.600 ;
        RECT 195.000 386.200 198.600 386.600 ;
        RECT 199.600 386.200 200.200 387.600 ;
        RECT 201.200 387.200 202.000 390.600 ;
        RECT 204.600 390.400 205.400 390.600 ;
        RECT 207.800 390.300 208.400 391.600 ;
        RECT 209.800 391.800 210.400 393.000 ;
        RECT 211.000 393.000 211.800 393.200 ;
        RECT 215.600 393.000 216.400 393.200 ;
        RECT 211.000 392.400 216.400 393.000 ;
        RECT 209.800 391.400 214.600 391.800 ;
        RECT 218.800 391.400 219.600 399.800 ;
        RECT 220.400 392.400 221.200 399.800 ;
        RECT 224.800 394.400 226.400 399.800 ;
        RECT 224.800 393.600 227.600 394.400 ;
        RECT 222.200 392.400 223.000 392.600 ;
        RECT 220.400 391.800 223.000 392.400 ;
        RECT 224.800 391.800 226.400 393.600 ;
        RECT 228.400 392.400 229.200 392.600 ;
        RECT 230.000 392.400 230.800 399.800 ;
        RECT 228.400 391.800 230.800 392.400 ;
        RECT 231.600 395.000 232.400 399.000 ;
        RECT 209.800 391.200 219.600 391.400 ;
        RECT 213.800 391.000 219.600 391.200 ;
        RECT 214.000 390.800 219.600 391.000 ;
        RECT 223.400 390.400 224.200 390.600 ;
        RECT 225.400 390.400 226.000 391.800 ;
        RECT 231.600 391.600 232.200 395.000 ;
        RECT 235.800 392.800 236.600 399.800 ;
        RECT 241.200 395.000 242.000 399.000 ;
        RECT 245.400 398.400 246.200 399.800 ;
        RECT 245.400 397.600 246.800 398.400 ;
        RECT 235.800 392.200 237.400 392.800 ;
        RECT 231.600 391.000 235.400 391.600 ;
        RECT 209.200 390.300 210.000 390.400 ;
        RECT 203.000 389.800 203.800 390.000 ;
        RECT 203.000 389.200 206.800 389.800 ;
        RECT 207.700 389.700 210.000 390.300 ;
        RECT 206.000 389.000 206.800 389.200 ;
        RECT 207.800 388.400 208.400 389.700 ;
        RECT 209.200 389.600 210.000 389.700 ;
        RECT 210.800 390.300 211.600 390.400 ;
        RECT 212.400 390.300 213.200 390.400 ;
        RECT 210.800 390.200 213.200 390.300 ;
        RECT 210.800 389.700 217.400 390.200 ;
        RECT 210.800 389.600 211.600 389.700 ;
        RECT 212.400 389.600 217.400 389.700 ;
        RECT 222.600 389.800 224.200 390.400 ;
        RECT 222.600 389.600 223.400 389.800 ;
        RECT 225.200 389.600 226.000 390.400 ;
        RECT 216.600 389.400 217.400 389.600 ;
        RECT 224.000 388.600 224.800 388.800 ;
        RECT 215.000 388.400 215.800 388.600 ;
        RECT 222.000 388.400 224.800 388.600 ;
        RECT 207.800 387.800 218.800 388.400 ;
        RECT 208.200 387.600 209.000 387.800 ;
        RECT 201.200 386.600 205.000 387.200 ;
        RECT 188.400 386.000 192.400 386.200 ;
        RECT 178.800 383.000 179.600 385.000 ;
        RECT 183.000 383.000 183.800 386.000 ;
        RECT 188.400 382.200 189.200 386.000 ;
        RECT 191.600 382.200 192.400 386.000 ;
        RECT 193.200 382.200 194.000 386.200 ;
        RECT 194.800 386.000 198.800 386.200 ;
        RECT 194.800 382.200 195.600 386.000 ;
        RECT 198.000 382.200 198.800 386.000 ;
        RECT 199.600 382.200 200.400 386.200 ;
        RECT 201.200 382.200 202.000 386.600 ;
        RECT 204.200 386.400 205.000 386.600 ;
        RECT 214.000 385.600 214.600 387.800 ;
        RECT 217.200 387.600 218.800 387.800 ;
        RECT 220.400 388.000 224.800 388.400 ;
        RECT 225.400 388.400 226.000 389.600 ;
        RECT 231.600 388.800 232.400 390.400 ;
        RECT 233.200 388.800 234.000 390.400 ;
        RECT 234.800 389.000 235.400 391.000 ;
        RECT 220.400 387.800 222.600 388.000 ;
        RECT 225.400 387.800 226.400 388.400 ;
        RECT 220.400 387.600 222.000 387.800 ;
        RECT 212.200 385.400 213.000 385.600 ;
        RECT 206.000 384.200 206.800 385.000 ;
        RECT 210.200 384.800 213.000 385.400 ;
        RECT 214.000 384.800 214.800 385.600 ;
        RECT 210.200 384.200 210.800 384.800 ;
        RECT 215.600 384.200 216.400 385.000 ;
        RECT 205.400 383.600 206.800 384.200 ;
        RECT 205.400 382.200 206.600 383.600 ;
        RECT 210.000 382.200 210.800 384.200 ;
        RECT 214.400 383.600 216.400 384.200 ;
        RECT 214.400 382.200 215.200 383.600 ;
        RECT 218.800 382.200 219.600 387.000 ;
        RECT 222.200 386.800 223.000 387.000 ;
        RECT 220.400 386.200 223.000 386.800 ;
        RECT 223.600 386.400 225.200 387.200 ;
        RECT 220.400 382.200 221.200 386.200 ;
        RECT 225.800 385.800 226.400 387.800 ;
        RECT 227.200 387.600 228.000 388.400 ;
        RECT 229.200 387.600 230.800 388.400 ;
        RECT 234.800 388.200 236.200 389.000 ;
        RECT 236.800 388.400 237.400 392.200 ;
        RECT 241.200 391.600 241.800 395.000 ;
        RECT 245.400 392.800 246.200 397.600 ;
        RECT 245.400 392.200 247.000 392.800 ;
        RECT 238.000 389.600 238.800 391.200 ;
        RECT 241.200 391.000 245.000 391.600 ;
        RECT 241.200 388.800 242.000 390.400 ;
        RECT 242.800 388.800 243.600 390.400 ;
        RECT 244.400 389.000 245.000 391.000 ;
        RECT 236.800 388.300 238.800 388.400 ;
        RECT 239.600 388.300 240.400 388.400 ;
        RECT 234.800 387.800 235.800 388.200 ;
        RECT 227.200 387.200 227.800 387.600 ;
        RECT 227.000 386.400 227.800 387.200 ;
        RECT 231.600 387.200 235.800 387.800 ;
        RECT 236.800 387.700 240.400 388.300 ;
        RECT 244.400 388.200 245.800 389.000 ;
        RECT 246.400 388.400 247.000 392.200 ;
        RECT 250.800 392.400 251.600 399.800 ;
        RECT 254.000 392.800 254.800 399.800 ;
        RECT 250.800 391.800 253.400 392.400 ;
        RECT 254.000 391.800 255.000 392.800 ;
        RECT 247.600 389.600 248.400 391.200 ;
        RECT 250.800 389.600 251.800 390.400 ;
        RECT 251.000 388.800 251.800 389.600 ;
        RECT 252.800 389.800 253.400 391.800 ;
        RECT 252.800 389.000 253.800 389.800 ;
        RECT 244.400 387.800 245.400 388.200 ;
        RECT 236.800 387.600 238.800 387.700 ;
        RECT 239.600 387.600 240.400 387.700 ;
        RECT 228.400 386.800 229.200 387.000 ;
        RECT 228.400 386.200 230.800 386.800 ;
        RECT 224.800 382.200 226.400 385.800 ;
        RECT 230.000 382.200 230.800 386.200 ;
        RECT 231.600 385.000 232.200 387.200 ;
        RECT 236.800 387.000 237.400 387.600 ;
        RECT 236.600 386.600 237.400 387.000 ;
        RECT 235.800 386.000 237.400 386.600 ;
        RECT 241.200 387.200 245.400 387.800 ;
        RECT 246.400 387.600 248.400 388.400 ;
        RECT 231.600 383.000 232.400 385.000 ;
        RECT 235.800 383.000 236.600 386.000 ;
        RECT 241.200 385.000 241.800 387.200 ;
        RECT 246.400 387.000 247.000 387.600 ;
        RECT 252.800 387.400 253.400 389.000 ;
        RECT 254.400 388.400 255.000 391.800 ;
        RECT 258.800 391.200 259.600 399.800 ;
        RECT 262.000 391.200 262.800 399.800 ;
        RECT 273.800 398.400 274.600 399.800 ;
        RECT 273.800 397.600 275.600 398.400 ;
        RECT 273.800 392.800 274.600 397.600 ;
        RECT 278.000 395.000 278.800 399.000 ;
        RECT 281.200 396.400 282.000 399.800 ;
        RECT 281.000 395.800 282.000 396.400 ;
        RECT 281.000 395.200 281.600 395.800 ;
        RECT 284.400 395.200 285.200 399.800 ;
        RECT 287.600 397.000 288.400 399.800 ;
        RECT 289.200 397.000 290.000 399.800 ;
        RECT 273.000 392.200 274.600 392.800 ;
        RECT 258.800 390.400 262.800 391.200 ;
        RECT 254.000 387.600 255.000 388.400 ;
        RECT 262.000 387.600 262.800 390.400 ;
        RECT 271.600 389.600 272.400 391.200 ;
        RECT 273.000 388.400 273.600 392.200 ;
        RECT 278.200 391.600 278.800 395.000 ;
        RECT 275.000 391.000 278.800 391.600 ;
        RECT 279.600 394.600 281.600 395.200 ;
        RECT 275.000 389.000 275.600 391.000 ;
        RECT 271.600 387.600 273.600 388.400 ;
        RECT 274.200 388.200 275.600 389.000 ;
        RECT 276.400 388.800 277.200 390.400 ;
        RECT 278.000 388.800 278.800 390.400 ;
        RECT 279.600 389.000 280.400 394.600 ;
        RECT 282.200 394.400 286.400 395.200 ;
        RECT 290.800 395.000 291.600 399.800 ;
        RECT 294.000 395.000 294.800 399.800 ;
        RECT 282.200 394.000 282.800 394.400 ;
        RECT 281.200 393.200 282.800 394.000 ;
        RECT 285.800 393.800 291.600 394.400 ;
        RECT 283.800 393.200 285.200 393.800 ;
        RECT 283.800 393.000 290.000 393.200 ;
        RECT 284.600 392.600 290.000 393.000 ;
        RECT 289.200 392.400 290.000 392.600 ;
        RECT 291.000 393.000 291.600 393.800 ;
        RECT 292.200 393.600 294.800 394.400 ;
        RECT 297.200 393.600 298.000 399.800 ;
        RECT 298.800 397.000 299.600 399.800 ;
        RECT 300.400 397.000 301.200 399.800 ;
        RECT 302.000 397.000 302.800 399.800 ;
        RECT 300.400 394.400 304.600 395.200 ;
        RECT 305.200 394.400 306.000 399.800 ;
        RECT 308.400 395.200 309.200 399.800 ;
        RECT 308.400 394.600 311.000 395.200 ;
        RECT 305.200 393.600 307.800 394.400 ;
        RECT 298.800 393.000 299.600 393.200 ;
        RECT 291.000 392.400 299.600 393.000 ;
        RECT 302.000 393.000 302.800 393.200 ;
        RECT 310.400 393.000 311.000 394.600 ;
        RECT 302.000 392.400 311.000 393.000 ;
        RECT 310.400 390.600 311.000 392.400 ;
        RECT 311.600 392.000 312.400 399.800 ;
        RECT 313.200 392.300 314.000 392.400 ;
        RECT 314.800 392.300 315.600 393.200 ;
        RECT 311.600 391.200 312.600 392.000 ;
        RECT 313.200 391.700 315.600 392.300 ;
        RECT 313.200 391.600 314.000 391.700 ;
        RECT 314.800 391.600 315.600 391.700 ;
        RECT 281.000 390.000 304.400 390.600 ;
        RECT 310.400 390.000 311.200 390.600 ;
        RECT 281.000 389.800 281.800 390.000 ;
        RECT 284.400 389.600 285.200 390.000 ;
        RECT 286.000 389.600 286.800 390.000 ;
        RECT 303.600 389.400 304.400 390.000 ;
        RECT 246.200 386.600 247.000 387.000 ;
        RECT 245.400 386.000 247.000 386.600 ;
        RECT 250.800 386.800 253.400 387.400 ;
        RECT 241.200 383.000 242.000 385.000 ;
        RECT 245.400 383.000 246.200 386.000 ;
        RECT 250.800 382.200 251.600 386.800 ;
        RECT 254.400 386.200 255.000 387.600 ;
        RECT 254.000 385.600 255.000 386.200 ;
        RECT 258.800 386.800 262.800 387.600 ;
        RECT 254.000 382.200 254.800 385.600 ;
        RECT 258.800 382.200 259.600 386.800 ;
        RECT 262.000 382.200 262.800 386.800 ;
        RECT 273.000 387.000 273.600 387.600 ;
        RECT 274.600 387.800 275.600 388.200 ;
        RECT 279.600 388.200 288.400 389.000 ;
        RECT 289.000 388.600 291.000 389.400 ;
        RECT 294.800 388.600 298.000 389.400 ;
        RECT 274.600 387.200 278.800 387.800 ;
        RECT 273.000 386.600 273.800 387.000 ;
        RECT 273.000 386.000 274.600 386.600 ;
        RECT 273.800 383.000 274.600 386.000 ;
        RECT 278.200 385.000 278.800 387.200 ;
        RECT 278.000 383.000 278.800 385.000 ;
        RECT 279.600 382.200 280.400 388.200 ;
        RECT 282.000 386.800 285.000 387.600 ;
        RECT 284.200 386.200 285.000 386.800 ;
        RECT 290.200 386.200 291.000 388.600 ;
        RECT 292.400 386.800 293.200 388.400 ;
        RECT 297.600 387.800 298.400 388.000 ;
        RECT 294.000 387.200 298.400 387.800 ;
        RECT 294.000 387.000 294.800 387.200 ;
        RECT 300.400 386.400 301.200 389.200 ;
        RECT 306.200 388.600 310.000 389.400 ;
        RECT 306.200 387.400 307.000 388.600 ;
        RECT 310.600 388.000 311.200 390.000 ;
        RECT 294.000 386.200 294.800 386.400 ;
        RECT 284.200 385.400 286.800 386.200 ;
        RECT 290.200 385.600 294.800 386.200 ;
        RECT 295.600 385.600 297.200 386.400 ;
        RECT 300.200 385.600 301.200 386.400 ;
        RECT 305.200 386.800 307.000 387.400 ;
        RECT 310.000 387.400 311.200 388.000 ;
        RECT 311.800 390.300 312.600 391.200 ;
        RECT 314.800 390.300 315.600 390.400 ;
        RECT 311.800 389.700 315.600 390.300 ;
        RECT 305.200 386.200 306.000 386.800 ;
        RECT 286.000 382.200 286.800 385.400 ;
        RECT 303.600 385.400 306.000 386.200 ;
        RECT 287.600 382.200 288.400 385.000 ;
        RECT 289.200 382.200 290.000 385.000 ;
        RECT 290.800 382.200 291.600 385.000 ;
        RECT 294.000 382.200 294.800 385.000 ;
        RECT 297.200 382.200 298.000 385.000 ;
        RECT 298.800 382.200 299.600 385.000 ;
        RECT 300.400 382.200 301.200 385.000 ;
        RECT 302.000 382.200 302.800 385.000 ;
        RECT 303.600 382.200 304.400 385.400 ;
        RECT 310.000 382.200 310.800 387.400 ;
        RECT 311.800 386.800 312.600 389.700 ;
        RECT 314.800 389.600 315.600 389.700 ;
        RECT 311.600 386.000 312.600 386.800 ;
        RECT 316.400 386.200 317.200 399.800 ;
        RECT 322.200 392.400 323.000 399.800 ;
        RECT 323.600 393.600 324.400 394.400 ;
        RECT 323.800 392.400 324.400 393.600 ;
        RECT 322.200 391.800 323.200 392.400 ;
        RECT 323.800 391.800 325.200 392.400 ;
        RECT 321.200 388.800 322.000 390.400 ;
        RECT 322.600 388.400 323.200 391.800 ;
        RECT 324.400 391.600 325.200 391.800 ;
        RECT 326.000 391.600 326.800 393.200 ;
        RECT 327.600 392.300 328.400 399.800 ;
        RECT 333.000 398.400 333.800 399.800 ;
        RECT 333.000 397.600 334.800 398.400 ;
        RECT 331.600 393.600 332.400 394.400 ;
        RECT 331.600 392.400 332.200 393.600 ;
        RECT 333.000 392.400 333.800 397.600 ;
        RECT 338.000 393.600 338.800 394.400 ;
        RECT 338.000 392.400 338.600 393.600 ;
        RECT 339.400 392.400 340.200 399.800 ;
        RECT 330.800 392.300 332.200 392.400 ;
        RECT 327.600 391.800 332.200 392.300 ;
        RECT 332.800 391.800 333.800 392.400 ;
        RECT 337.200 391.800 338.600 392.400 ;
        RECT 339.200 391.800 340.200 392.400 ;
        RECT 343.600 391.800 344.400 399.800 ;
        RECT 345.200 392.400 346.000 399.800 ;
        RECT 348.400 392.400 349.200 399.800 ;
        RECT 345.200 391.800 349.200 392.400 ;
        RECT 352.600 391.800 354.600 399.800 ;
        RECT 360.600 392.600 361.400 399.800 ;
        RECT 359.600 391.800 361.400 392.600 ;
        RECT 327.600 391.700 331.600 391.800 ;
        RECT 318.000 386.800 318.800 388.400 ;
        RECT 319.600 388.200 320.400 388.400 ;
        RECT 319.600 387.600 321.200 388.200 ;
        RECT 322.600 387.600 325.200 388.400 ;
        RECT 320.400 387.200 321.200 387.600 ;
        RECT 319.800 386.200 323.400 386.600 ;
        RECT 324.400 386.400 325.000 387.600 ;
        RECT 311.600 382.200 312.400 386.000 ;
        RECT 315.400 385.600 317.200 386.200 ;
        RECT 319.600 386.000 323.600 386.200 ;
        RECT 315.400 384.400 316.200 385.600 ;
        RECT 314.800 383.600 316.200 384.400 ;
        RECT 315.400 382.200 316.200 383.600 ;
        RECT 319.600 382.200 320.400 386.000 ;
        RECT 322.800 382.200 323.600 386.000 ;
        RECT 324.400 382.200 325.200 386.400 ;
        RECT 327.600 386.200 328.400 391.700 ;
        RECT 330.800 391.600 331.600 391.700 ;
        RECT 332.800 388.400 333.400 391.800 ;
        RECT 337.200 391.600 338.000 391.800 ;
        RECT 334.000 388.800 334.800 390.400 ;
        RECT 339.200 388.400 339.800 391.800 ;
        RECT 343.800 390.400 344.400 391.800 ;
        RECT 347.600 390.400 348.400 390.800 ;
        RECT 340.400 388.800 341.200 390.400 ;
        RECT 343.600 389.800 346.000 390.400 ;
        RECT 347.600 389.800 349.200 390.400 ;
        RECT 343.600 389.600 344.400 389.800 ;
        RECT 329.200 386.800 330.000 388.400 ;
        RECT 330.800 387.600 333.400 388.400 ;
        RECT 335.600 388.200 336.400 388.400 ;
        RECT 334.800 387.600 336.400 388.200 ;
        RECT 337.200 387.600 339.800 388.400 ;
        RECT 342.000 388.300 342.800 388.400 ;
        RECT 343.600 388.300 344.400 388.400 ;
        RECT 342.000 388.200 344.400 388.300 ;
        RECT 341.200 387.700 344.400 388.200 ;
        RECT 341.200 387.600 342.800 387.700 ;
        RECT 343.600 387.600 344.400 387.700 ;
        RECT 331.000 386.200 331.600 387.600 ;
        RECT 334.800 387.200 335.600 387.600 ;
        RECT 332.600 386.200 336.200 386.600 ;
        RECT 337.400 386.200 338.000 387.600 ;
        RECT 341.200 387.200 342.000 387.600 ;
        RECT 339.000 386.200 342.600 386.600 ;
        RECT 326.600 385.600 328.400 386.200 ;
        RECT 326.600 382.200 327.400 385.600 ;
        RECT 330.800 382.200 331.600 386.200 ;
        RECT 332.400 386.000 336.400 386.200 ;
        RECT 332.400 382.200 333.200 386.000 ;
        RECT 335.600 382.200 336.400 386.000 ;
        RECT 337.200 382.200 338.000 386.200 ;
        RECT 338.800 386.000 342.800 386.200 ;
        RECT 338.800 382.200 339.600 386.000 ;
        RECT 342.000 382.200 342.800 386.000 ;
        RECT 343.600 385.600 344.400 386.400 ;
        RECT 345.400 386.200 346.000 389.800 ;
        RECT 348.400 389.600 349.200 389.800 ;
        RECT 346.800 387.600 347.600 389.200 ;
        RECT 350.000 387.600 350.800 389.200 ;
        RECT 351.600 388.800 352.400 390.400 ;
        RECT 353.400 388.400 354.000 391.800 ;
        RECT 354.800 390.300 355.600 390.400 ;
        RECT 358.000 390.300 358.800 390.400 ;
        RECT 354.800 389.700 358.800 390.300 ;
        RECT 354.800 388.800 355.600 389.700 ;
        RECT 358.000 389.600 358.800 389.700 ;
        RECT 359.800 388.400 360.400 391.800 ;
        RECT 362.800 391.600 363.600 399.800 ;
        RECT 364.400 392.400 365.200 399.800 ;
        RECT 367.600 392.400 368.400 399.800 ;
        RECT 364.400 391.800 368.400 392.400 ;
        RECT 369.200 391.600 370.000 393.200 ;
        RECT 361.200 389.600 362.000 391.200 ;
        RECT 363.000 390.400 363.600 391.600 ;
        RECT 366.800 390.400 367.600 390.800 ;
        RECT 362.800 389.800 365.200 390.400 ;
        RECT 366.800 390.300 368.400 390.400 ;
        RECT 369.200 390.300 370.000 390.400 ;
        RECT 366.800 389.800 370.000 390.300 ;
        RECT 362.800 389.600 363.600 389.800 ;
        RECT 353.200 388.200 354.000 388.400 ;
        RECT 356.400 388.300 357.200 388.400 ;
        RECT 356.400 388.200 358.700 388.300 ;
        RECT 351.600 387.600 354.000 388.200 ;
        RECT 355.600 387.700 358.700 388.200 ;
        RECT 355.600 387.600 357.200 387.700 ;
        RECT 351.600 386.200 352.200 387.600 ;
        RECT 355.600 387.200 356.400 387.600 ;
        RECT 353.400 386.200 357.000 386.600 ;
        RECT 358.100 386.400 358.700 387.700 ;
        RECT 359.600 387.600 360.400 388.400 ;
        RECT 359.800 386.400 360.400 387.600 ;
        RECT 343.800 384.800 344.600 385.600 ;
        RECT 345.200 382.200 346.000 386.200 ;
        RECT 350.000 382.800 350.800 386.200 ;
        RECT 351.600 383.400 352.400 386.200 ;
        RECT 353.200 386.000 357.200 386.200 ;
        RECT 353.200 382.800 354.000 386.000 ;
        RECT 350.000 382.200 354.000 382.800 ;
        RECT 356.400 382.200 357.200 386.000 ;
        RECT 358.000 384.800 358.800 386.400 ;
        RECT 359.600 385.600 360.400 386.400 ;
        RECT 362.800 385.600 363.600 386.400 ;
        RECT 364.600 386.200 365.200 389.800 ;
        RECT 367.600 389.700 370.000 389.800 ;
        RECT 367.600 389.600 368.400 389.700 ;
        RECT 369.200 389.600 370.000 389.700 ;
        RECT 366.000 388.300 366.800 389.200 ;
        RECT 370.800 388.300 371.600 399.800 ;
        RECT 375.600 395.800 376.400 399.800 ;
        RECT 375.800 395.600 376.400 395.800 ;
        RECT 378.800 395.800 379.600 399.800 ;
        RECT 378.800 395.600 379.400 395.800 ;
        RECT 375.800 395.000 379.400 395.600 ;
        RECT 377.200 392.800 378.000 394.400 ;
        RECT 378.800 392.400 379.400 395.000 ;
        RECT 374.000 390.800 374.800 392.400 ;
        RECT 378.800 391.600 379.600 392.400 ;
        RECT 375.600 389.600 377.200 390.400 ;
        RECT 378.800 388.400 379.400 391.600 ;
        RECT 366.000 387.700 371.600 388.300 ;
        RECT 366.000 387.600 366.800 387.700 ;
        RECT 370.800 386.200 371.600 387.700 ;
        RECT 372.400 386.800 373.200 388.400 ;
        RECT 377.800 388.200 379.400 388.400 ;
        RECT 377.600 387.800 379.400 388.200 ;
        RECT 359.800 384.200 360.400 385.600 ;
        RECT 363.000 384.800 363.800 385.600 ;
        RECT 359.600 382.200 360.400 384.200 ;
        RECT 364.400 382.200 365.200 386.200 ;
        RECT 369.800 385.600 371.600 386.200 ;
        RECT 369.800 382.200 370.600 385.600 ;
        RECT 377.600 382.200 378.400 387.800 ;
        RECT 380.400 386.800 381.200 388.400 ;
        RECT 382.000 386.200 382.800 399.800 ;
        RECT 386.800 396.400 387.600 399.800 ;
        RECT 386.600 395.800 387.600 396.400 ;
        RECT 386.600 395.200 387.200 395.800 ;
        RECT 390.000 395.200 390.800 399.800 ;
        RECT 393.200 397.000 394.000 399.800 ;
        RECT 394.800 397.000 395.600 399.800 ;
        RECT 385.200 394.600 387.200 395.200 ;
        RECT 383.600 391.600 384.400 393.200 ;
        RECT 385.200 389.000 386.000 394.600 ;
        RECT 387.800 394.400 392.000 395.200 ;
        RECT 396.400 395.000 397.200 399.800 ;
        RECT 399.600 395.000 400.400 399.800 ;
        RECT 387.800 394.000 388.400 394.400 ;
        RECT 386.800 393.200 388.400 394.000 ;
        RECT 391.400 393.800 397.200 394.400 ;
        RECT 389.400 393.200 390.800 393.800 ;
        RECT 389.400 393.000 395.600 393.200 ;
        RECT 390.200 392.600 395.600 393.000 ;
        RECT 394.800 392.400 395.600 392.600 ;
        RECT 396.600 393.000 397.200 393.800 ;
        RECT 397.800 393.600 400.400 394.400 ;
        RECT 402.800 393.600 403.600 399.800 ;
        RECT 404.400 397.000 405.200 399.800 ;
        RECT 406.000 397.000 406.800 399.800 ;
        RECT 407.600 397.000 408.400 399.800 ;
        RECT 406.000 394.400 410.200 395.200 ;
        RECT 410.800 394.400 411.600 399.800 ;
        RECT 414.000 395.200 414.800 399.800 ;
        RECT 414.000 394.600 416.600 395.200 ;
        RECT 410.800 393.600 413.400 394.400 ;
        RECT 404.400 393.000 405.200 393.200 ;
        RECT 396.600 392.400 405.200 393.000 ;
        RECT 407.600 393.000 408.400 393.200 ;
        RECT 416.000 393.000 416.600 394.600 ;
        RECT 407.600 392.400 416.600 393.000 ;
        RECT 416.000 390.600 416.600 392.400 ;
        RECT 417.200 392.000 418.000 399.800 ;
        RECT 425.200 395.000 426.000 399.000 ;
        RECT 417.200 391.200 418.200 392.000 ;
        RECT 386.600 390.000 410.000 390.600 ;
        RECT 416.000 390.000 416.800 390.600 ;
        RECT 386.600 389.800 387.400 390.000 ;
        RECT 388.400 389.600 389.200 390.000 ;
        RECT 391.600 389.600 392.400 390.000 ;
        RECT 409.200 389.400 410.000 390.000 ;
        RECT 385.200 388.200 394.000 389.000 ;
        RECT 394.600 388.600 396.600 389.400 ;
        RECT 400.400 388.600 403.600 389.400 ;
        RECT 382.000 385.600 383.800 386.200 ;
        RECT 383.000 382.200 383.800 385.600 ;
        RECT 385.200 382.200 386.000 388.200 ;
        RECT 387.600 386.800 390.600 387.600 ;
        RECT 389.800 386.200 390.600 386.800 ;
        RECT 395.800 386.200 396.600 388.600 ;
        RECT 398.000 386.800 398.800 388.400 ;
        RECT 403.200 387.800 404.000 388.000 ;
        RECT 399.600 387.200 404.000 387.800 ;
        RECT 399.600 387.000 400.400 387.200 ;
        RECT 406.000 386.400 406.800 389.200 ;
        RECT 411.800 388.600 415.600 389.400 ;
        RECT 411.800 387.400 412.600 388.600 ;
        RECT 416.200 388.000 416.800 390.000 ;
        RECT 399.600 386.200 400.400 386.400 ;
        RECT 389.800 385.400 392.400 386.200 ;
        RECT 395.800 385.600 400.400 386.200 ;
        RECT 401.200 385.600 402.800 386.400 ;
        RECT 405.800 385.600 406.800 386.400 ;
        RECT 410.800 386.800 412.600 387.400 ;
        RECT 415.600 387.400 416.800 388.000 ;
        RECT 417.400 390.300 418.200 391.200 ;
        RECT 425.200 391.600 425.800 395.000 ;
        RECT 429.400 392.800 430.200 399.800 ;
        RECT 436.400 392.800 437.200 399.800 ;
        RECT 429.400 392.200 431.000 392.800 ;
        RECT 425.200 391.000 429.000 391.600 ;
        RECT 425.200 390.300 426.000 390.400 ;
        RECT 417.400 389.700 426.000 390.300 ;
        RECT 410.800 386.200 411.600 386.800 ;
        RECT 391.600 382.200 392.400 385.400 ;
        RECT 409.200 385.400 411.600 386.200 ;
        RECT 393.200 382.200 394.000 385.000 ;
        RECT 394.800 382.200 395.600 385.000 ;
        RECT 396.400 382.200 397.200 385.000 ;
        RECT 399.600 382.200 400.400 385.000 ;
        RECT 402.800 382.200 403.600 385.000 ;
        RECT 404.400 382.200 405.200 385.000 ;
        RECT 406.000 382.200 406.800 385.000 ;
        RECT 407.600 382.200 408.400 385.000 ;
        RECT 409.200 382.200 410.000 385.400 ;
        RECT 415.600 382.200 416.400 387.400 ;
        RECT 417.400 386.800 418.200 389.700 ;
        RECT 425.200 388.800 426.000 389.700 ;
        RECT 426.800 388.800 427.600 390.400 ;
        RECT 428.400 389.000 429.000 391.000 ;
        RECT 428.400 388.200 429.800 389.000 ;
        RECT 430.400 388.400 431.000 392.200 ;
        RECT 436.200 391.800 437.200 392.800 ;
        RECT 439.600 392.400 440.400 399.800 ;
        RECT 437.800 391.800 440.400 392.400 ;
        RECT 443.800 392.400 444.600 399.800 ;
        RECT 445.200 394.300 446.000 394.400 ;
        RECT 449.200 394.300 450.000 399.800 ;
        RECT 452.400 395.200 453.200 399.800 ;
        RECT 445.200 393.700 450.000 394.300 ;
        RECT 445.200 393.600 446.000 393.700 ;
        RECT 445.400 392.400 446.000 393.600 ;
        RECT 443.800 391.800 444.800 392.400 ;
        RECT 445.400 391.800 446.800 392.400 ;
        RECT 449.200 392.000 450.000 393.700 ;
        RECT 431.600 389.600 432.400 391.200 ;
        RECT 436.200 388.400 436.800 391.800 ;
        RECT 437.800 389.800 438.400 391.800 ;
        RECT 437.400 389.000 438.400 389.800 ;
        RECT 428.400 387.800 429.400 388.200 ;
        RECT 417.200 386.000 418.200 386.800 ;
        RECT 425.200 387.200 429.400 387.800 ;
        RECT 430.400 387.600 432.400 388.400 ;
        RECT 436.200 387.600 437.200 388.400 ;
        RECT 417.200 382.200 418.000 386.000 ;
        RECT 425.200 385.000 425.800 387.200 ;
        RECT 430.400 387.000 431.000 387.600 ;
        RECT 430.200 386.600 431.000 387.000 ;
        RECT 429.400 386.400 431.000 386.600 ;
        RECT 428.400 386.000 431.000 386.400 ;
        RECT 436.200 386.200 436.800 387.600 ;
        RECT 437.800 387.400 438.400 389.000 ;
        RECT 439.400 389.600 440.400 390.400 ;
        RECT 439.400 388.800 440.200 389.600 ;
        RECT 442.800 388.800 443.600 390.400 ;
        RECT 444.200 388.400 444.800 391.800 ;
        RECT 446.000 391.600 446.800 391.800 ;
        RECT 449.000 391.200 450.000 392.000 ;
        RECT 450.600 394.600 453.200 395.200 ;
        RECT 450.600 393.000 451.200 394.600 ;
        RECT 455.600 394.400 456.400 399.800 ;
        RECT 458.800 397.000 459.600 399.800 ;
        RECT 460.400 397.000 461.200 399.800 ;
        RECT 462.000 397.000 462.800 399.800 ;
        RECT 457.000 394.400 461.200 395.200 ;
        RECT 453.800 393.600 456.400 394.400 ;
        RECT 463.600 393.600 464.400 399.800 ;
        RECT 466.800 395.000 467.600 399.800 ;
        RECT 470.000 395.000 470.800 399.800 ;
        RECT 471.600 397.000 472.400 399.800 ;
        RECT 473.200 397.000 474.000 399.800 ;
        RECT 476.400 395.200 477.200 399.800 ;
        RECT 479.600 396.400 480.400 399.800 ;
        RECT 479.600 395.800 480.600 396.400 ;
        RECT 480.000 395.200 480.600 395.800 ;
        RECT 475.200 394.400 479.400 395.200 ;
        RECT 480.000 394.600 482.000 395.200 ;
        RECT 466.800 393.600 469.400 394.400 ;
        RECT 470.000 393.800 475.800 394.400 ;
        RECT 478.800 394.000 479.400 394.400 ;
        RECT 458.800 393.000 459.600 393.200 ;
        RECT 450.600 392.400 459.600 393.000 ;
        RECT 462.000 393.000 462.800 393.200 ;
        RECT 470.000 393.000 470.600 393.800 ;
        RECT 476.400 393.200 477.800 393.800 ;
        RECT 478.800 393.200 480.400 394.000 ;
        RECT 462.000 392.400 470.600 393.000 ;
        RECT 471.600 393.000 477.800 393.200 ;
        RECT 471.600 392.600 477.000 393.000 ;
        RECT 471.600 392.400 472.400 392.600 ;
        RECT 441.200 388.200 442.000 388.400 ;
        RECT 444.200 388.300 446.800 388.400 ;
        RECT 447.600 388.300 448.400 388.400 ;
        RECT 441.200 387.600 442.800 388.200 ;
        RECT 444.200 387.700 448.400 388.300 ;
        RECT 444.200 387.600 446.800 387.700 ;
        RECT 447.600 387.600 448.400 387.700 ;
        RECT 437.800 386.800 440.400 387.400 ;
        RECT 442.000 387.200 442.800 387.600 ;
        RECT 428.400 385.600 430.200 386.000 ;
        RECT 436.200 385.600 437.200 386.200 ;
        RECT 425.200 383.000 426.000 385.000 ;
        RECT 429.400 383.000 430.200 385.600 ;
        RECT 436.400 382.200 437.200 385.600 ;
        RECT 439.600 382.200 440.400 386.800 ;
        RECT 441.400 386.200 445.000 386.600 ;
        RECT 446.000 386.200 446.600 387.600 ;
        RECT 449.000 386.800 449.800 391.200 ;
        RECT 450.600 390.600 451.200 392.400 ;
        RECT 450.400 390.000 451.200 390.600 ;
        RECT 457.200 390.000 480.600 390.600 ;
        RECT 450.400 388.000 451.000 390.000 ;
        RECT 457.200 389.400 458.000 390.000 ;
        RECT 474.800 389.600 475.600 390.000 ;
        RECT 478.000 389.600 478.800 390.000 ;
        RECT 479.800 389.800 480.600 390.000 ;
        RECT 451.600 388.600 455.400 389.400 ;
        RECT 450.400 387.400 451.600 388.000 ;
        RECT 441.200 386.000 445.200 386.200 ;
        RECT 441.200 382.200 442.000 386.000 ;
        RECT 444.400 382.200 445.200 386.000 ;
        RECT 446.000 382.200 446.800 386.200 ;
        RECT 449.000 386.000 450.000 386.800 ;
        RECT 449.200 382.200 450.000 386.000 ;
        RECT 450.800 382.200 451.600 387.400 ;
        RECT 454.600 387.400 455.400 388.600 ;
        RECT 454.600 386.800 456.400 387.400 ;
        RECT 455.600 386.200 456.400 386.800 ;
        RECT 460.400 386.400 461.200 389.200 ;
        RECT 463.600 388.600 466.800 389.400 ;
        RECT 470.600 388.600 472.600 389.400 ;
        RECT 481.200 389.000 482.000 394.600 ;
        RECT 463.200 387.800 464.000 388.000 ;
        RECT 463.200 387.200 467.600 387.800 ;
        RECT 466.800 387.000 467.600 387.200 ;
        RECT 468.400 386.800 469.200 388.400 ;
        RECT 455.600 385.400 458.000 386.200 ;
        RECT 460.400 385.600 461.400 386.400 ;
        RECT 464.400 385.600 466.000 386.400 ;
        RECT 466.800 386.200 467.600 386.400 ;
        RECT 470.600 386.200 471.400 388.600 ;
        RECT 473.200 388.200 482.000 389.000 ;
        RECT 476.600 386.800 479.600 387.600 ;
        RECT 476.600 386.200 477.400 386.800 ;
        RECT 466.800 385.600 471.400 386.200 ;
        RECT 457.200 382.200 458.000 385.400 ;
        RECT 474.800 385.400 477.400 386.200 ;
        RECT 458.800 382.200 459.600 385.000 ;
        RECT 460.400 382.200 461.200 385.000 ;
        RECT 462.000 382.200 462.800 385.000 ;
        RECT 463.600 382.200 464.400 385.000 ;
        RECT 466.800 382.200 467.600 385.000 ;
        RECT 470.000 382.200 470.800 385.000 ;
        RECT 471.600 382.200 472.400 385.000 ;
        RECT 473.200 382.200 474.000 385.000 ;
        RECT 474.800 382.200 475.600 385.400 ;
        RECT 481.200 382.200 482.000 388.200 ;
        RECT 482.800 386.800 483.600 388.400 ;
        RECT 484.400 386.200 485.200 399.800 ;
        RECT 486.000 391.600 486.800 393.200 ;
        RECT 487.600 391.600 488.400 394.400 ;
        RECT 489.200 386.200 490.000 399.800 ;
        RECT 494.000 391.200 494.800 399.800 ;
        RECT 497.200 391.200 498.000 399.800 ;
        RECT 500.400 391.600 501.200 394.400 ;
        RECT 494.000 390.400 498.000 391.200 ;
        RECT 490.800 386.800 491.600 388.400 ;
        RECT 497.200 387.600 498.000 390.400 ;
        RECT 494.000 386.800 498.000 387.600 ;
        RECT 484.400 385.600 486.200 386.200 ;
        RECT 485.400 384.400 486.200 385.600 ;
        RECT 488.200 385.600 490.000 386.200 ;
        RECT 488.200 384.400 489.000 385.600 ;
        RECT 484.400 383.600 486.200 384.400 ;
        RECT 487.600 383.600 489.000 384.400 ;
        RECT 485.400 382.200 486.200 383.600 ;
        RECT 488.200 382.200 489.000 383.600 ;
        RECT 494.000 382.200 494.800 386.800 ;
        RECT 497.200 382.200 498.000 386.800 ;
        RECT 502.000 386.200 502.800 399.800 ;
        RECT 506.000 393.600 506.800 394.400 ;
        RECT 506.000 392.400 506.600 393.600 ;
        RECT 507.400 392.400 508.200 399.800 ;
        RECT 512.400 393.600 513.200 394.400 ;
        RECT 512.400 392.400 513.000 393.600 ;
        RECT 513.800 392.400 514.600 399.800 ;
        RECT 520.200 398.400 521.000 399.800 ;
        RECT 520.200 397.600 522.000 398.400 ;
        RECT 518.800 393.600 519.600 394.400 ;
        RECT 518.800 392.400 519.400 393.600 ;
        RECT 520.200 392.400 521.000 397.600 ;
        RECT 526.000 392.800 526.800 399.800 ;
        RECT 503.600 392.300 504.400 392.400 ;
        RECT 505.200 392.300 506.600 392.400 ;
        RECT 503.600 391.800 506.600 392.300 ;
        RECT 507.200 391.800 508.200 392.400 ;
        RECT 511.600 391.800 513.000 392.400 ;
        RECT 513.600 391.800 514.600 392.400 ;
        RECT 518.000 391.800 519.400 392.400 ;
        RECT 520.000 391.800 521.000 392.400 ;
        RECT 525.800 391.800 526.800 392.800 ;
        RECT 529.200 392.400 530.000 399.800 ;
        RECT 527.400 391.800 530.000 392.400 ;
        RECT 503.600 391.700 506.000 391.800 ;
        RECT 503.600 391.600 504.400 391.700 ;
        RECT 505.200 391.600 506.000 391.700 ;
        RECT 507.200 390.400 507.800 391.800 ;
        RECT 511.600 391.600 512.400 391.800 ;
        RECT 506.800 389.600 507.800 390.400 ;
        RECT 507.200 388.400 507.800 389.600 ;
        RECT 508.400 388.800 509.200 390.400 ;
        RECT 510.000 390.300 510.800 390.400 ;
        RECT 513.600 390.300 514.200 391.800 ;
        RECT 518.000 391.600 518.800 391.800 ;
        RECT 510.000 389.700 514.200 390.300 ;
        RECT 510.000 389.600 510.800 389.700 ;
        RECT 513.600 388.400 514.200 389.700 ;
        RECT 514.800 388.800 515.600 390.400 ;
        RECT 520.000 388.400 520.600 391.800 ;
        RECT 521.200 388.800 522.000 390.400 ;
        RECT 525.800 388.400 526.400 391.800 ;
        RECT 527.400 389.800 528.000 391.800 ;
        RECT 530.800 391.600 531.600 394.400 ;
        RECT 527.000 389.000 528.000 389.800 ;
        RECT 503.600 386.800 504.400 388.400 ;
        RECT 505.200 387.600 507.800 388.400 ;
        RECT 510.000 388.200 510.800 388.400 ;
        RECT 509.200 387.600 510.800 388.200 ;
        RECT 511.600 387.600 514.200 388.400 ;
        RECT 516.400 388.200 517.200 388.400 ;
        RECT 515.600 387.600 517.200 388.200 ;
        RECT 518.000 387.600 520.600 388.400 ;
        RECT 522.800 388.200 523.600 388.400 ;
        RECT 522.000 387.600 523.600 388.200 ;
        RECT 525.800 387.600 526.800 388.400 ;
        RECT 505.400 386.200 506.000 387.600 ;
        RECT 509.200 387.200 510.000 387.600 ;
        RECT 507.000 386.200 510.600 386.600 ;
        RECT 511.800 386.200 512.400 387.600 ;
        RECT 515.600 387.200 516.400 387.600 ;
        RECT 513.400 386.200 517.000 386.600 ;
        RECT 518.200 386.200 518.800 387.600 ;
        RECT 522.000 387.200 522.800 387.600 ;
        RECT 519.800 386.200 523.400 386.600 ;
        RECT 525.800 386.200 526.400 387.600 ;
        RECT 527.400 387.400 528.000 389.000 ;
        RECT 529.000 389.600 530.000 390.400 ;
        RECT 529.000 388.800 529.800 389.600 ;
        RECT 527.400 386.800 530.000 387.400 ;
        RECT 501.000 385.600 502.800 386.200 ;
        RECT 501.000 384.400 501.800 385.600 ;
        RECT 500.400 383.600 501.800 384.400 ;
        RECT 501.000 382.200 501.800 383.600 ;
        RECT 505.200 382.200 506.000 386.200 ;
        RECT 506.800 386.000 510.800 386.200 ;
        RECT 506.800 382.200 507.600 386.000 ;
        RECT 510.000 382.200 510.800 386.000 ;
        RECT 511.600 382.200 512.400 386.200 ;
        RECT 513.200 386.000 517.200 386.200 ;
        RECT 513.200 382.200 514.000 386.000 ;
        RECT 516.400 382.200 517.200 386.000 ;
        RECT 518.000 382.200 518.800 386.200 ;
        RECT 519.600 386.000 523.600 386.200 ;
        RECT 519.600 382.200 520.400 386.000 ;
        RECT 522.800 382.200 523.600 386.000 ;
        RECT 525.800 385.600 526.800 386.200 ;
        RECT 526.000 382.200 526.800 385.600 ;
        RECT 529.200 382.200 530.000 386.800 ;
        RECT 532.400 386.200 533.200 399.800 ;
        RECT 538.200 392.400 539.000 399.800 ;
        RECT 539.600 393.600 540.400 394.400 ;
        RECT 539.800 392.400 540.400 393.600 ;
        RECT 542.800 393.600 543.600 394.400 ;
        RECT 542.800 392.400 543.400 393.600 ;
        RECT 544.200 392.400 545.000 399.800 ;
        RECT 538.200 391.800 539.200 392.400 ;
        RECT 539.800 391.800 541.200 392.400 ;
        RECT 537.200 388.800 538.000 390.400 ;
        RECT 538.600 390.300 539.200 391.800 ;
        RECT 540.400 391.600 541.200 391.800 ;
        RECT 542.000 391.800 543.400 392.400 ;
        RECT 542.000 391.600 542.800 391.800 ;
        RECT 544.000 391.600 546.000 392.400 ;
        RECT 542.100 390.300 542.700 391.600 ;
        RECT 538.600 389.700 542.700 390.300 ;
        RECT 538.600 388.400 539.200 389.700 ;
        RECT 544.000 388.400 544.600 391.600 ;
        RECT 548.400 391.400 549.200 399.800 ;
        RECT 552.800 396.400 553.600 399.800 ;
        RECT 551.600 395.800 553.600 396.400 ;
        RECT 557.200 395.800 558.000 399.800 ;
        RECT 561.400 395.800 562.600 399.800 ;
        RECT 551.600 395.000 552.400 395.800 ;
        RECT 557.200 395.200 557.800 395.800 ;
        RECT 555.000 394.600 558.600 395.200 ;
        RECT 561.200 395.000 562.000 395.800 ;
        RECT 555.000 394.400 555.800 394.600 ;
        RECT 557.800 394.400 558.600 394.600 ;
        RECT 551.600 393.000 552.400 393.200 ;
        RECT 556.200 393.000 557.000 393.200 ;
        RECT 551.600 392.400 557.000 393.000 ;
        RECT 557.600 393.000 559.800 393.600 ;
        RECT 557.600 391.800 558.200 393.000 ;
        RECT 559.000 392.800 559.800 393.000 ;
        RECT 561.400 393.200 562.800 394.000 ;
        RECT 561.400 392.200 562.000 393.200 ;
        RECT 553.400 391.400 558.200 391.800 ;
        RECT 548.400 391.200 558.200 391.400 ;
        RECT 559.600 391.600 562.000 392.200 ;
        RECT 548.400 391.000 554.200 391.200 ;
        RECT 548.400 390.800 554.000 391.000 ;
        RECT 545.200 390.300 546.000 390.400 ;
        RECT 546.800 390.300 547.600 390.400 ;
        RECT 545.200 389.700 547.600 390.300 ;
        RECT 554.800 390.200 555.600 390.400 ;
        RECT 545.200 388.800 546.000 389.700 ;
        RECT 546.800 389.600 547.600 389.700 ;
        RECT 550.600 389.600 555.600 390.200 ;
        RECT 550.600 389.400 551.400 389.600 ;
        RECT 552.200 388.400 553.000 388.600 ;
        RECT 559.600 388.400 560.200 391.600 ;
        RECT 566.000 391.200 566.800 399.800 ;
        RECT 562.600 390.600 566.800 391.200 ;
        RECT 562.600 390.400 563.400 390.600 ;
        RECT 564.200 389.800 565.000 390.000 ;
        RECT 561.200 389.200 565.000 389.800 ;
        RECT 561.200 389.000 562.000 389.200 ;
        RECT 534.000 386.800 534.800 388.400 ;
        RECT 535.600 388.200 536.400 388.400 ;
        RECT 535.600 387.600 537.200 388.200 ;
        RECT 538.600 387.600 541.200 388.400 ;
        RECT 542.000 387.600 544.600 388.400 ;
        RECT 546.800 388.200 547.600 388.400 ;
        RECT 546.000 387.600 547.600 388.200 ;
        RECT 549.200 387.800 560.200 388.400 ;
        RECT 549.200 387.600 550.800 387.800 ;
        RECT 536.400 387.200 537.200 387.600 ;
        RECT 535.800 386.200 539.400 386.600 ;
        RECT 540.400 386.200 541.000 387.600 ;
        RECT 542.200 386.200 542.800 387.600 ;
        RECT 546.000 387.200 546.800 387.600 ;
        RECT 543.800 386.200 547.400 386.600 ;
        RECT 531.400 385.600 533.200 386.200 ;
        RECT 535.600 386.000 539.600 386.200 ;
        RECT 531.400 384.400 532.200 385.600 ;
        RECT 530.800 383.600 532.200 384.400 ;
        RECT 531.400 382.200 532.200 383.600 ;
        RECT 535.600 382.200 536.400 386.000 ;
        RECT 538.800 382.200 539.600 386.000 ;
        RECT 540.400 382.200 541.200 386.200 ;
        RECT 542.000 382.200 542.800 386.200 ;
        RECT 543.600 386.000 547.600 386.200 ;
        RECT 543.600 382.200 544.400 386.000 ;
        RECT 546.800 382.200 547.600 386.000 ;
        RECT 548.400 382.200 549.200 387.000 ;
        RECT 553.400 385.600 554.000 387.800 ;
        RECT 556.400 387.600 557.200 387.800 ;
        RECT 559.000 387.600 559.800 387.800 ;
        RECT 564.400 387.200 565.200 388.400 ;
        RECT 566.000 387.200 566.800 390.600 ;
        RECT 563.000 386.600 566.800 387.200 ;
        RECT 563.000 386.400 563.800 386.600 ;
        RECT 551.600 384.200 552.400 385.000 ;
        RECT 553.200 384.800 554.000 385.600 ;
        RECT 555.000 385.400 555.800 385.600 ;
        RECT 555.000 384.800 557.800 385.400 ;
        RECT 557.200 384.200 557.800 384.800 ;
        RECT 561.200 384.200 562.000 385.000 ;
        RECT 551.600 383.600 553.600 384.200 ;
        RECT 552.800 382.200 553.600 383.600 ;
        RECT 557.200 382.200 558.000 384.200 ;
        RECT 561.200 383.600 562.600 384.200 ;
        RECT 561.400 382.200 562.600 383.600 ;
        RECT 566.000 382.200 566.800 386.600 ;
        RECT 567.600 382.200 568.400 399.800 ;
        RECT 575.600 391.600 576.400 394.400 ;
        RECT 569.200 384.800 570.000 386.400 ;
        RECT 577.200 386.200 578.000 399.800 ;
        RECT 582.600 398.400 583.400 399.800 ;
        RECT 582.600 397.600 584.400 398.400 ;
        RECT 581.200 393.600 582.000 394.400 ;
        RECT 581.200 392.400 581.800 393.600 ;
        RECT 582.600 392.400 583.400 397.600 ;
        RECT 580.400 391.800 581.800 392.400 ;
        RECT 582.400 391.800 583.400 392.400 ;
        RECT 580.400 391.600 581.200 391.800 ;
        RECT 582.400 388.400 583.000 391.800 ;
        RECT 586.800 391.400 587.600 399.800 ;
        RECT 591.200 396.400 592.000 399.800 ;
        RECT 590.000 395.800 592.000 396.400 ;
        RECT 595.600 395.800 596.400 399.800 ;
        RECT 599.800 395.800 601.000 399.800 ;
        RECT 590.000 395.000 590.800 395.800 ;
        RECT 595.600 395.200 596.200 395.800 ;
        RECT 593.400 394.600 597.000 395.200 ;
        RECT 599.600 395.000 600.400 395.800 ;
        RECT 593.400 394.400 594.200 394.600 ;
        RECT 596.200 394.400 597.000 394.600 ;
        RECT 590.000 393.000 590.800 393.200 ;
        RECT 594.600 393.000 595.400 393.200 ;
        RECT 590.000 392.400 595.400 393.000 ;
        RECT 596.000 393.000 598.200 393.600 ;
        RECT 596.000 391.800 596.600 393.000 ;
        RECT 597.400 392.800 598.200 393.000 ;
        RECT 599.800 393.200 601.200 394.000 ;
        RECT 599.800 392.200 600.400 393.200 ;
        RECT 591.800 391.400 596.600 391.800 ;
        RECT 586.800 391.200 596.600 391.400 ;
        RECT 598.000 391.600 600.400 392.200 ;
        RECT 586.800 391.000 592.600 391.200 ;
        RECT 586.800 390.800 592.400 391.000 ;
        RECT 583.600 388.800 584.400 390.400 ;
        RECT 593.200 390.200 594.000 390.400 ;
        RECT 589.000 389.600 594.000 390.200 ;
        RECT 589.000 389.400 589.800 389.600 ;
        RECT 591.600 389.400 592.400 389.600 ;
        RECT 590.600 388.400 591.400 388.600 ;
        RECT 598.000 388.400 598.600 391.600 ;
        RECT 604.400 391.200 605.200 399.800 ;
        RECT 606.000 395.800 606.800 399.800 ;
        RECT 606.200 395.600 606.800 395.800 ;
        RECT 609.200 395.800 610.000 399.800 ;
        RECT 609.200 395.600 609.800 395.800 ;
        RECT 606.200 395.000 609.800 395.600 ;
        RECT 606.200 392.400 606.800 395.000 ;
        RECT 607.600 392.800 608.400 394.400 ;
        RECT 615.000 392.400 615.800 399.800 ;
        RECT 616.400 393.600 617.200 394.400 ;
        RECT 616.600 392.400 617.200 393.600 ;
        RECT 606.000 391.600 606.800 392.400 ;
        RECT 601.000 390.600 605.200 391.200 ;
        RECT 601.000 390.400 601.800 390.600 ;
        RECT 602.600 389.800 603.400 390.000 ;
        RECT 599.600 389.200 603.400 389.800 ;
        RECT 599.600 389.000 600.400 389.200 ;
        RECT 578.800 386.800 579.600 388.400 ;
        RECT 580.400 387.600 583.000 388.400 ;
        RECT 585.200 388.200 586.000 388.400 ;
        RECT 584.400 387.600 586.000 388.200 ;
        RECT 587.600 387.800 598.600 388.400 ;
        RECT 587.600 387.600 589.200 387.800 ;
        RECT 580.600 386.200 581.200 387.600 ;
        RECT 584.400 387.200 585.200 387.600 ;
        RECT 582.200 386.200 585.800 386.600 ;
        RECT 576.200 385.600 578.000 386.200 ;
        RECT 570.800 384.300 571.600 384.400 ;
        RECT 576.200 384.300 577.000 385.600 ;
        RECT 570.800 383.700 577.000 384.300 ;
        RECT 570.800 383.600 571.600 383.700 ;
        RECT 576.200 382.200 577.000 383.700 ;
        RECT 580.400 382.200 581.200 386.200 ;
        RECT 582.000 386.000 586.000 386.200 ;
        RECT 582.000 382.200 582.800 386.000 ;
        RECT 585.200 382.200 586.000 386.000 ;
        RECT 586.800 382.200 587.600 387.000 ;
        RECT 591.800 385.600 592.400 387.800 ;
        RECT 596.400 387.600 598.200 387.800 ;
        RECT 604.400 387.200 605.200 390.600 ;
        RECT 606.200 388.400 606.800 391.600 ;
        RECT 610.800 390.800 611.600 392.400 ;
        RECT 615.000 391.800 616.000 392.400 ;
        RECT 616.600 391.800 618.000 392.400 ;
        RECT 608.400 389.600 610.000 390.400 ;
        RECT 614.000 388.800 614.800 390.400 ;
        RECT 615.400 388.400 616.000 391.800 ;
        RECT 617.200 391.600 618.000 391.800 ;
        RECT 618.800 391.600 619.600 393.200 ;
        RECT 617.300 390.300 617.900 391.600 ;
        RECT 620.400 390.300 621.200 399.800 ;
        RECT 617.300 389.700 621.200 390.300 ;
        RECT 606.200 388.200 607.800 388.400 ;
        RECT 612.400 388.200 613.200 388.400 ;
        RECT 615.400 388.300 618.000 388.400 ;
        RECT 618.800 388.300 619.600 388.400 ;
        RECT 606.200 387.800 608.000 388.200 ;
        RECT 601.400 386.600 605.200 387.200 ;
        RECT 601.400 386.400 602.200 386.600 ;
        RECT 590.000 384.200 590.800 385.000 ;
        RECT 591.600 384.800 592.400 385.600 ;
        RECT 593.400 385.400 594.200 385.600 ;
        RECT 593.400 384.800 596.200 385.400 ;
        RECT 595.600 384.200 596.200 384.800 ;
        RECT 599.600 384.200 600.400 385.000 ;
        RECT 590.000 383.600 592.000 384.200 ;
        RECT 591.200 382.200 592.000 383.600 ;
        RECT 595.600 382.200 596.400 384.200 ;
        RECT 599.600 383.600 601.000 384.200 ;
        RECT 599.800 382.200 601.000 383.600 ;
        RECT 604.400 382.200 605.200 386.600 ;
        RECT 607.200 382.200 608.000 387.800 ;
        RECT 612.400 387.600 614.000 388.200 ;
        RECT 615.400 387.700 619.600 388.300 ;
        RECT 615.400 387.600 618.000 387.700 ;
        RECT 618.800 387.600 619.600 387.700 ;
        RECT 613.200 387.200 614.000 387.600 ;
        RECT 612.600 386.200 616.200 386.600 ;
        RECT 617.200 386.200 617.800 387.600 ;
        RECT 620.400 386.200 621.200 389.700 ;
        RECT 623.600 391.200 624.400 399.800 ;
        RECT 627.800 395.800 629.000 399.800 ;
        RECT 632.400 395.800 633.200 399.800 ;
        RECT 636.800 396.400 637.600 399.800 ;
        RECT 636.800 395.800 638.800 396.400 ;
        RECT 628.400 395.000 629.200 395.800 ;
        RECT 632.600 395.200 633.200 395.800 ;
        RECT 631.800 394.600 635.400 395.200 ;
        RECT 638.000 395.000 638.800 395.800 ;
        RECT 631.800 394.400 632.600 394.600 ;
        RECT 634.600 394.400 635.400 394.600 ;
        RECT 627.600 393.200 629.000 394.000 ;
        RECT 628.400 392.200 629.000 393.200 ;
        RECT 630.600 393.000 632.800 393.600 ;
        RECT 630.600 392.800 631.400 393.000 ;
        RECT 628.400 391.600 630.800 392.200 ;
        RECT 623.600 390.600 627.800 391.200 ;
        RECT 622.000 386.800 622.800 388.400 ;
        RECT 623.600 387.200 624.400 390.600 ;
        RECT 627.000 390.400 627.800 390.600 ;
        RECT 625.400 389.800 626.200 390.000 ;
        RECT 625.400 389.200 629.200 389.800 ;
        RECT 628.400 389.000 629.200 389.200 ;
        RECT 630.200 388.400 630.800 391.600 ;
        RECT 632.200 391.800 632.800 393.000 ;
        RECT 633.400 393.000 634.200 393.200 ;
        RECT 638.000 393.000 638.800 393.200 ;
        RECT 633.400 392.400 638.800 393.000 ;
        RECT 632.200 391.400 637.000 391.800 ;
        RECT 641.200 391.400 642.000 399.800 ;
        RECT 643.600 393.600 644.400 394.400 ;
        RECT 643.600 392.400 644.200 393.600 ;
        RECT 645.000 392.400 645.800 399.800 ;
        RECT 650.800 396.400 651.600 399.800 ;
        RECT 650.600 395.800 651.600 396.400 ;
        RECT 650.600 395.200 651.200 395.800 ;
        RECT 654.000 395.200 654.800 399.800 ;
        RECT 657.200 397.000 658.000 399.800 ;
        RECT 658.800 397.000 659.600 399.800 ;
        RECT 642.800 391.800 644.200 392.400 ;
        RECT 644.800 391.800 645.800 392.400 ;
        RECT 649.200 394.600 651.200 395.200 ;
        RECT 642.800 391.600 643.600 391.800 ;
        RECT 632.200 391.200 642.000 391.400 ;
        RECT 636.200 391.000 642.000 391.200 ;
        RECT 636.400 390.800 642.000 391.000 ;
        RECT 634.800 390.200 635.600 390.400 ;
        RECT 634.800 389.600 639.800 390.200 ;
        RECT 636.400 389.400 637.200 389.600 ;
        RECT 639.000 389.400 639.800 389.600 ;
        RECT 637.400 388.400 638.200 388.600 ;
        RECT 644.800 388.400 645.400 391.800 ;
        RECT 646.000 388.800 646.800 390.400 ;
        RECT 649.200 389.000 650.000 394.600 ;
        RECT 651.800 394.400 656.000 395.200 ;
        RECT 660.400 395.000 661.200 399.800 ;
        RECT 663.600 395.000 664.400 399.800 ;
        RECT 651.800 394.000 652.400 394.400 ;
        RECT 650.800 393.200 652.400 394.000 ;
        RECT 655.400 393.800 661.200 394.400 ;
        RECT 653.400 393.200 654.800 393.800 ;
        RECT 653.400 393.000 659.600 393.200 ;
        RECT 654.200 392.600 659.600 393.000 ;
        RECT 658.800 392.400 659.600 392.600 ;
        RECT 660.600 393.000 661.200 393.800 ;
        RECT 661.800 393.600 664.400 394.400 ;
        RECT 666.800 393.600 667.600 399.800 ;
        RECT 668.400 397.000 669.200 399.800 ;
        RECT 670.000 397.000 670.800 399.800 ;
        RECT 671.600 397.000 672.400 399.800 ;
        RECT 670.000 394.400 674.200 395.200 ;
        RECT 674.800 394.400 675.600 399.800 ;
        RECT 678.000 395.200 678.800 399.800 ;
        RECT 678.000 394.600 680.600 395.200 ;
        RECT 674.800 393.600 677.400 394.400 ;
        RECT 668.400 393.000 669.200 393.200 ;
        RECT 660.600 392.400 669.200 393.000 ;
        RECT 671.600 393.000 672.400 393.200 ;
        RECT 680.000 393.000 680.600 394.600 ;
        RECT 671.600 392.400 680.600 393.000 ;
        RECT 680.000 390.600 680.600 392.400 ;
        RECT 681.200 392.000 682.000 399.800 ;
        RECT 681.200 391.200 682.200 392.000 ;
        RECT 650.600 390.000 674.000 390.600 ;
        RECT 680.000 390.000 680.800 390.600 ;
        RECT 650.600 389.800 651.400 390.000 ;
        RECT 654.000 389.600 654.800 390.000 ;
        RECT 655.600 389.600 656.400 390.000 ;
        RECT 673.200 389.400 674.000 390.000 ;
        RECT 630.200 387.800 641.200 388.400 ;
        RECT 630.600 387.600 631.400 387.800 ;
        RECT 612.400 386.000 616.400 386.200 ;
        RECT 612.400 382.200 613.200 386.000 ;
        RECT 615.600 382.200 616.400 386.000 ;
        RECT 617.200 382.200 618.000 386.200 ;
        RECT 619.400 385.600 621.200 386.200 ;
        RECT 623.600 386.600 627.400 387.200 ;
        RECT 619.400 382.200 620.200 385.600 ;
        RECT 623.600 382.200 624.400 386.600 ;
        RECT 626.600 386.400 627.400 386.600 ;
        RECT 636.400 385.600 637.000 387.800 ;
        RECT 639.600 387.600 641.200 387.800 ;
        RECT 642.800 387.600 645.400 388.400 ;
        RECT 647.600 388.200 648.400 388.400 ;
        RECT 646.800 387.600 648.400 388.200 ;
        RECT 649.200 388.200 658.000 389.000 ;
        RECT 658.600 388.600 660.600 389.400 ;
        RECT 664.400 388.600 667.600 389.400 ;
        RECT 634.600 385.400 635.400 385.600 ;
        RECT 628.400 384.200 629.200 385.000 ;
        RECT 632.600 384.800 635.400 385.400 ;
        RECT 636.400 384.800 637.200 385.600 ;
        RECT 632.600 384.200 633.200 384.800 ;
        RECT 638.000 384.200 638.800 385.000 ;
        RECT 627.800 383.600 629.200 384.200 ;
        RECT 627.800 382.200 629.000 383.600 ;
        RECT 632.400 382.200 633.200 384.200 ;
        RECT 636.800 383.600 638.800 384.200 ;
        RECT 636.800 382.200 637.600 383.600 ;
        RECT 641.200 382.200 642.000 387.000 ;
        RECT 643.000 386.200 643.600 387.600 ;
        RECT 646.800 387.200 647.600 387.600 ;
        RECT 644.600 386.200 648.200 386.600 ;
        RECT 642.800 382.200 643.600 386.200 ;
        RECT 644.400 386.000 648.400 386.200 ;
        RECT 644.400 382.200 645.200 386.000 ;
        RECT 647.600 382.200 648.400 386.000 ;
        RECT 649.200 382.200 650.000 388.200 ;
        RECT 651.600 386.800 654.600 387.600 ;
        RECT 653.800 386.200 654.600 386.800 ;
        RECT 659.800 386.200 660.600 388.600 ;
        RECT 662.000 386.800 662.800 388.400 ;
        RECT 667.200 387.800 668.000 388.000 ;
        RECT 663.600 387.200 668.000 387.800 ;
        RECT 663.600 387.000 664.400 387.200 ;
        RECT 670.000 386.400 670.800 389.200 ;
        RECT 675.800 388.600 679.600 389.400 ;
        RECT 675.800 387.400 676.600 388.600 ;
        RECT 680.200 388.000 680.800 390.000 ;
        RECT 663.600 386.200 664.400 386.400 ;
        RECT 653.800 385.400 656.400 386.200 ;
        RECT 659.800 385.600 664.400 386.200 ;
        RECT 665.200 385.600 666.800 386.400 ;
        RECT 669.800 385.600 670.800 386.400 ;
        RECT 674.800 386.800 676.600 387.400 ;
        RECT 679.600 387.400 680.800 388.000 ;
        RECT 674.800 386.200 675.600 386.800 ;
        RECT 655.600 382.200 656.400 385.400 ;
        RECT 673.200 385.400 675.600 386.200 ;
        RECT 657.200 382.200 658.000 385.000 ;
        RECT 658.800 382.200 659.600 385.000 ;
        RECT 660.400 382.200 661.200 385.000 ;
        RECT 663.600 382.200 664.400 385.000 ;
        RECT 666.800 382.200 667.600 385.000 ;
        RECT 668.400 382.200 669.200 385.000 ;
        RECT 670.000 382.200 670.800 385.000 ;
        RECT 671.600 382.200 672.400 385.000 ;
        RECT 673.200 382.200 674.000 385.400 ;
        RECT 679.600 382.200 680.400 387.400 ;
        RECT 681.400 386.800 682.200 391.200 ;
        RECT 681.200 386.000 682.200 386.800 ;
        RECT 681.200 382.200 682.000 386.000 ;
        RECT 1.200 375.000 2.000 379.800 ;
        RECT 5.600 378.400 6.400 379.800 ;
        RECT 4.400 377.800 6.400 378.400 ;
        RECT 10.000 377.800 10.800 379.800 ;
        RECT 14.200 378.400 15.400 379.800 ;
        RECT 14.000 377.800 15.400 378.400 ;
        RECT 4.400 377.000 5.200 377.800 ;
        RECT 10.000 377.200 10.600 377.800 ;
        RECT 6.000 376.400 6.800 377.200 ;
        RECT 7.800 376.600 10.600 377.200 ;
        RECT 14.000 377.000 14.800 377.800 ;
        RECT 7.800 376.400 8.600 376.600 ;
        RECT 2.000 374.200 3.600 374.400 ;
        RECT 6.200 374.200 6.800 376.400 ;
        RECT 15.800 375.400 16.600 375.600 ;
        RECT 18.800 375.400 19.600 379.800 ;
        RECT 20.400 375.600 21.200 377.200 ;
        RECT 15.800 374.800 19.600 375.400 ;
        RECT 11.800 374.200 12.600 374.400 ;
        RECT 2.000 373.600 13.000 374.200 ;
        RECT 5.000 373.400 5.800 373.600 ;
        RECT 3.400 372.400 4.200 372.600 ;
        RECT 12.400 372.400 13.000 373.600 ;
        RECT 14.000 372.800 14.800 373.000 ;
        RECT 3.400 371.800 8.400 372.400 ;
        RECT 7.600 371.600 8.400 371.800 ;
        RECT 12.400 371.600 13.200 372.400 ;
        RECT 14.000 372.200 17.800 372.800 ;
        RECT 17.000 372.000 17.800 372.200 ;
        RECT 1.200 371.000 6.800 371.200 ;
        RECT 1.200 370.800 7.000 371.000 ;
        RECT 1.200 370.600 11.000 370.800 ;
        RECT 1.200 362.200 2.000 370.600 ;
        RECT 6.200 370.200 11.000 370.600 ;
        RECT 4.400 369.000 9.800 369.600 ;
        RECT 4.400 368.800 5.200 369.000 ;
        RECT 9.000 368.800 9.800 369.000 ;
        RECT 10.400 369.000 11.000 370.200 ;
        RECT 12.400 370.400 13.000 371.600 ;
        RECT 15.400 371.400 16.200 371.600 ;
        RECT 18.800 371.400 19.600 374.800 ;
        RECT 15.400 370.800 19.600 371.400 ;
        RECT 12.400 369.800 14.800 370.400 ;
        RECT 11.800 369.000 12.600 369.200 ;
        RECT 10.400 368.400 12.600 369.000 ;
        RECT 14.200 368.800 14.800 369.800 ;
        RECT 14.200 368.000 15.600 368.800 ;
        RECT 7.800 367.400 8.600 367.600 ;
        RECT 10.600 367.400 11.400 367.600 ;
        RECT 4.400 366.200 5.200 367.000 ;
        RECT 7.800 366.800 11.400 367.400 ;
        RECT 10.000 366.200 10.600 366.800 ;
        RECT 14.000 366.200 14.800 367.000 ;
        RECT 4.400 365.600 6.400 366.200 ;
        RECT 5.600 362.200 6.400 365.600 ;
        RECT 10.000 362.200 10.800 366.200 ;
        RECT 14.200 362.200 15.400 366.200 ;
        RECT 18.800 362.200 19.600 370.800 ;
        RECT 22.000 362.200 22.800 379.800 ;
        RECT 23.600 376.000 24.400 379.800 ;
        RECT 26.800 376.000 27.600 379.800 ;
        RECT 23.600 375.800 27.600 376.000 ;
        RECT 28.400 375.800 29.200 379.800 ;
        RECT 30.000 375.800 30.800 379.800 ;
        RECT 31.600 376.000 32.400 379.800 ;
        RECT 34.800 376.000 35.600 379.800 ;
        RECT 40.200 376.000 41.000 379.000 ;
        RECT 44.400 377.000 45.200 379.000 ;
        RECT 31.600 375.800 35.600 376.000 ;
        RECT 23.800 375.400 27.400 375.800 ;
        RECT 24.400 374.400 25.200 374.800 ;
        RECT 28.400 374.400 29.000 375.800 ;
        RECT 30.200 374.400 30.800 375.800 ;
        RECT 31.800 375.400 35.400 375.800 ;
        RECT 39.400 375.400 41.000 376.000 ;
        RECT 39.400 375.000 40.200 375.400 ;
        RECT 34.000 374.400 34.800 374.800 ;
        RECT 39.400 374.400 40.000 375.000 ;
        RECT 44.600 374.800 45.200 377.000 ;
        RECT 49.800 376.000 50.600 379.000 ;
        RECT 54.000 377.000 54.800 379.000 ;
        RECT 23.600 373.800 25.200 374.400 ;
        RECT 23.600 373.600 24.400 373.800 ;
        RECT 26.600 373.600 29.200 374.400 ;
        RECT 30.000 373.600 32.600 374.400 ;
        RECT 34.000 374.300 35.600 374.400 ;
        RECT 36.400 374.300 37.200 374.400 ;
        RECT 34.000 373.800 37.200 374.300 ;
        RECT 34.800 373.700 37.200 373.800 ;
        RECT 34.800 373.600 35.600 373.700 ;
        RECT 36.400 373.600 37.200 373.700 ;
        RECT 38.000 373.600 40.000 374.400 ;
        RECT 41.000 374.200 45.200 374.800 ;
        RECT 49.000 375.400 50.600 376.000 ;
        RECT 49.000 375.000 49.800 375.400 ;
        RECT 49.000 374.400 49.600 375.000 ;
        RECT 54.200 374.800 54.800 377.000 ;
        RECT 55.600 375.600 56.400 377.200 ;
        RECT 46.000 374.300 46.800 374.400 ;
        RECT 47.600 374.300 49.600 374.400 ;
        RECT 41.000 373.800 42.000 374.200 ;
        RECT 25.200 371.600 26.000 373.200 ;
        RECT 26.600 372.300 27.200 373.600 ;
        RECT 26.600 371.700 30.700 372.300 ;
        RECT 26.600 370.200 27.200 371.700 ;
        RECT 30.100 370.400 30.700 371.700 ;
        RECT 28.400 370.200 29.200 370.400 ;
        RECT 26.200 369.600 27.200 370.200 ;
        RECT 27.800 369.600 29.200 370.200 ;
        RECT 30.000 370.200 30.800 370.400 ;
        RECT 32.000 370.200 32.600 373.600 ;
        RECT 33.200 371.600 34.000 373.200 ;
        RECT 34.800 372.300 35.600 372.400 ;
        RECT 38.000 372.300 38.800 372.400 ;
        RECT 34.800 371.700 38.800 372.300 ;
        RECT 34.800 371.600 35.600 371.700 ;
        RECT 38.000 370.800 38.800 371.700 ;
        RECT 30.000 369.600 31.400 370.200 ;
        RECT 32.000 369.600 33.000 370.200 ;
        RECT 26.200 362.200 27.000 369.600 ;
        RECT 27.800 368.400 28.400 369.600 ;
        RECT 27.600 367.600 28.400 368.400 ;
        RECT 30.800 368.400 31.400 369.600 ;
        RECT 30.800 367.600 31.600 368.400 ;
        RECT 32.200 362.200 33.000 369.600 ;
        RECT 39.400 369.800 40.000 373.600 ;
        RECT 40.600 373.000 42.000 373.800 ;
        RECT 46.000 373.700 49.600 374.300 ;
        RECT 50.600 374.200 54.800 374.800 ;
        RECT 50.600 373.800 51.600 374.200 ;
        RECT 46.000 373.600 46.800 373.700 ;
        RECT 47.600 373.600 49.600 373.700 ;
        RECT 41.400 371.000 42.000 373.000 ;
        RECT 42.800 371.600 43.600 373.200 ;
        RECT 44.400 371.600 45.200 373.200 ;
        RECT 41.400 370.400 45.200 371.000 ;
        RECT 47.600 370.800 48.400 372.400 ;
        RECT 39.400 369.200 41.000 369.800 ;
        RECT 40.200 364.400 41.000 369.200 ;
        RECT 44.600 367.000 45.200 370.400 ;
        RECT 49.000 369.800 49.600 373.600 ;
        RECT 50.200 373.000 51.600 373.800 ;
        RECT 51.000 371.000 51.600 373.000 ;
        RECT 52.400 371.600 53.200 373.200 ;
        RECT 54.000 371.600 54.800 373.200 ;
        RECT 51.000 370.400 54.800 371.000 ;
        RECT 49.000 369.200 50.600 369.800 ;
        RECT 39.600 363.600 41.000 364.400 ;
        RECT 40.200 362.200 41.000 363.600 ;
        RECT 44.400 363.000 45.200 367.000 ;
        RECT 49.800 362.200 50.600 369.200 ;
        RECT 54.200 367.000 54.800 370.400 ;
        RECT 54.000 363.000 54.800 367.000 ;
        RECT 57.200 362.200 58.000 379.800 ;
        RECT 58.800 375.800 59.600 379.800 ;
        RECT 60.400 376.000 61.200 379.800 ;
        RECT 63.600 376.000 64.400 379.800 ;
        RECT 67.800 376.400 68.600 379.800 ;
        RECT 60.400 375.800 64.400 376.000 ;
        RECT 66.800 375.800 68.600 376.400 ;
        RECT 59.000 374.400 59.600 375.800 ;
        RECT 60.600 375.400 64.200 375.800 ;
        RECT 62.800 374.400 63.600 374.800 ;
        RECT 58.800 373.600 61.400 374.400 ;
        RECT 62.800 373.800 64.400 374.400 ;
        RECT 63.600 373.600 64.400 373.800 ;
        RECT 65.200 373.600 66.000 375.200 ;
        RECT 58.800 370.200 59.600 370.400 ;
        RECT 60.800 370.200 61.400 373.600 ;
        RECT 62.000 371.600 62.800 373.200 ;
        RECT 58.800 369.600 60.200 370.200 ;
        RECT 60.800 369.600 61.800 370.200 ;
        RECT 59.600 368.400 60.200 369.600 ;
        RECT 61.000 368.400 61.800 369.600 ;
        RECT 59.600 367.600 60.400 368.400 ;
        RECT 61.000 367.600 62.800 368.400 ;
        RECT 61.000 362.200 61.800 367.600 ;
        RECT 66.800 362.200 67.600 375.800 ;
        RECT 70.000 375.600 70.800 377.200 ;
        RECT 68.400 370.300 69.200 370.400 ;
        RECT 70.000 370.300 70.800 370.400 ;
        RECT 68.400 369.700 70.800 370.300 ;
        RECT 68.400 368.800 69.200 369.700 ;
        RECT 70.000 369.600 70.800 369.700 ;
        RECT 71.600 362.200 72.400 379.800 ;
        RECT 73.200 376.000 74.000 379.800 ;
        RECT 76.400 376.000 77.200 379.800 ;
        RECT 73.200 375.800 77.200 376.000 ;
        RECT 78.000 375.800 78.800 379.800 ;
        RECT 73.400 375.400 77.000 375.800 ;
        RECT 74.000 374.400 74.800 374.800 ;
        RECT 78.000 374.400 78.600 375.800 ;
        RECT 79.600 375.600 80.400 377.200 ;
        RECT 73.200 373.800 74.800 374.400 ;
        RECT 73.200 373.600 74.000 373.800 ;
        RECT 76.200 373.600 78.800 374.400 ;
        RECT 73.200 372.300 74.000 372.400 ;
        RECT 74.800 372.300 75.600 373.200 ;
        RECT 73.200 371.700 75.600 372.300 ;
        RECT 73.200 371.600 74.000 371.700 ;
        RECT 74.800 371.600 75.600 371.700 ;
        RECT 76.200 372.300 76.800 373.600 ;
        RECT 79.600 372.300 80.400 372.400 ;
        RECT 76.200 371.700 80.400 372.300 ;
        RECT 76.200 370.200 76.800 371.700 ;
        RECT 79.600 371.600 80.400 371.700 ;
        RECT 78.000 370.200 78.800 370.400 ;
        RECT 75.800 369.600 76.800 370.200 ;
        RECT 77.400 369.600 78.800 370.200 ;
        RECT 75.800 362.200 76.600 369.600 ;
        RECT 77.400 368.400 78.000 369.600 ;
        RECT 77.200 367.600 78.000 368.400 ;
        RECT 79.600 368.300 80.400 368.400 ;
        RECT 81.200 368.300 82.000 379.800 ;
        RECT 82.800 375.200 83.600 379.800 ;
        RECT 86.000 376.400 86.800 379.800 ;
        RECT 86.000 375.800 87.000 376.400 ;
        RECT 89.200 376.000 90.000 379.800 ;
        RECT 92.400 376.000 93.200 379.800 ;
        RECT 89.200 375.800 93.200 376.000 ;
        RECT 94.000 375.800 94.800 379.800 ;
        RECT 95.600 376.000 96.400 379.800 ;
        RECT 98.800 376.000 99.600 379.800 ;
        RECT 95.600 375.800 99.600 376.000 ;
        RECT 100.400 375.800 101.200 379.800 ;
        RECT 102.000 376.000 102.800 379.800 ;
        RECT 105.200 376.000 106.000 379.800 ;
        RECT 102.000 375.800 106.000 376.000 ;
        RECT 106.800 375.800 107.600 379.800 ;
        RECT 82.800 374.600 85.400 375.200 ;
        RECT 83.000 372.400 83.800 373.200 ;
        RECT 82.800 371.600 83.800 372.400 ;
        RECT 84.800 373.000 85.400 374.600 ;
        RECT 86.400 374.400 87.000 375.800 ;
        RECT 89.400 375.400 93.000 375.800 ;
        RECT 90.000 374.400 90.800 374.800 ;
        RECT 94.000 374.400 94.600 375.800 ;
        RECT 95.800 375.400 99.400 375.800 ;
        RECT 96.400 374.400 97.200 374.800 ;
        RECT 100.400 374.400 101.000 375.800 ;
        RECT 102.200 375.400 105.800 375.800 ;
        RECT 102.800 374.400 103.600 374.800 ;
        RECT 106.800 374.400 107.400 375.800 ;
        RECT 86.000 373.600 87.000 374.400 ;
        RECT 89.200 373.800 90.800 374.400 ;
        RECT 89.200 373.600 90.000 373.800 ;
        RECT 92.200 373.600 94.800 374.400 ;
        RECT 95.600 373.800 97.200 374.400 ;
        RECT 98.600 374.300 101.200 374.400 ;
        RECT 102.000 374.300 103.600 374.400 ;
        RECT 98.600 373.800 103.600 374.300 ;
        RECT 95.600 373.600 96.400 373.800 ;
        RECT 98.600 373.700 102.800 373.800 ;
        RECT 98.600 373.600 101.200 373.700 ;
        RECT 102.000 373.600 102.800 373.700 ;
        RECT 105.000 373.600 107.600 374.400 ;
        RECT 116.800 374.200 117.600 379.800 ;
        RECT 119.600 375.800 120.400 379.800 ;
        RECT 121.200 376.000 122.000 379.800 ;
        RECT 124.400 376.000 125.200 379.800 ;
        RECT 121.200 375.800 125.200 376.000 ;
        RECT 119.800 374.400 120.400 375.800 ;
        RECT 121.400 375.400 125.000 375.800 ;
        RECT 126.000 375.200 126.800 379.800 ;
        RECT 129.200 376.400 130.000 379.800 ;
        RECT 134.000 377.800 134.800 379.800 ;
        RECT 134.000 376.400 134.600 377.800 ;
        RECT 129.200 375.800 130.200 376.400 ;
        RECT 123.600 374.400 124.400 374.800 ;
        RECT 126.000 374.600 128.600 375.200 ;
        RECT 116.800 373.800 118.600 374.200 ;
        RECT 117.000 373.600 118.600 373.800 ;
        RECT 119.600 373.600 122.200 374.400 ;
        RECT 123.600 373.800 125.200 374.400 ;
        RECT 124.400 373.600 125.200 373.800 ;
        RECT 84.800 372.200 85.800 373.000 ;
        RECT 84.800 370.200 85.400 372.200 ;
        RECT 86.400 370.200 87.000 373.600 ;
        RECT 90.800 371.600 91.600 373.200 ;
        RECT 92.200 370.200 92.800 373.600 ;
        RECT 97.200 371.600 98.000 373.200 ;
        RECT 94.000 370.200 94.800 370.400 ;
        RECT 98.600 370.200 99.200 373.600 ;
        RECT 103.600 371.600 104.400 373.200 ;
        RECT 100.400 370.200 101.200 370.400 ;
        RECT 105.000 370.200 105.600 373.600 ;
        RECT 114.800 371.600 116.400 372.400 ;
        RECT 106.800 370.300 107.600 370.400 ;
        RECT 108.400 370.300 109.200 370.400 ;
        RECT 106.800 370.200 109.200 370.300 ;
        RECT 79.600 367.700 82.000 368.300 ;
        RECT 79.600 367.600 80.400 367.700 ;
        RECT 81.200 362.200 82.000 367.700 ;
        RECT 82.800 369.600 85.400 370.200 ;
        RECT 82.800 362.200 83.600 369.600 ;
        RECT 86.000 369.200 87.000 370.200 ;
        RECT 91.800 369.600 92.800 370.200 ;
        RECT 93.400 369.600 94.800 370.200 ;
        RECT 98.200 369.600 99.200 370.200 ;
        RECT 99.800 369.600 101.200 370.200 ;
        RECT 104.600 369.600 105.600 370.200 ;
        RECT 106.200 369.700 109.200 370.200 ;
        RECT 106.200 369.600 107.600 369.700 ;
        RECT 108.400 369.600 109.200 369.700 ;
        RECT 113.200 369.600 114.000 371.200 ;
        RECT 118.000 370.400 118.600 373.600 ;
        RECT 118.000 369.600 118.800 370.400 ;
        RECT 119.600 370.200 120.400 370.400 ;
        RECT 121.600 370.200 122.200 373.600 ;
        RECT 122.800 371.600 123.600 373.200 ;
        RECT 126.200 372.400 127.000 373.200 ;
        RECT 126.000 371.600 127.000 372.400 ;
        RECT 128.000 373.000 128.600 374.600 ;
        RECT 129.600 374.400 130.200 375.800 ;
        RECT 129.200 373.600 130.200 374.400 ;
        RECT 128.000 372.200 129.000 373.000 ;
        RECT 128.000 370.200 128.600 372.200 ;
        RECT 129.600 370.200 130.200 373.600 ;
        RECT 134.000 375.600 134.800 376.400 ;
        RECT 135.600 375.600 136.400 377.200 ;
        RECT 137.200 375.800 138.000 379.800 ;
        RECT 138.800 376.000 139.600 379.800 ;
        RECT 142.000 376.000 142.800 379.800 ;
        RECT 138.800 375.800 142.800 376.000 ;
        RECT 134.000 374.400 134.600 375.600 ;
        RECT 137.400 374.400 138.000 375.800 ;
        RECT 139.000 375.400 142.600 375.800 ;
        RECT 141.200 374.400 142.000 374.800 ;
        RECT 134.000 373.600 134.800 374.400 ;
        RECT 137.200 373.600 139.800 374.400 ;
        RECT 141.200 373.800 142.800 374.400 ;
        RECT 142.000 373.600 142.800 373.800 ;
        RECT 132.400 370.800 133.200 372.400 ;
        RECT 134.000 370.200 134.600 373.600 ;
        RECT 137.200 370.200 138.000 370.400 ;
        RECT 139.200 370.200 139.800 373.600 ;
        RECT 140.400 371.600 141.200 373.200 ;
        RECT 119.600 369.600 121.000 370.200 ;
        RECT 121.600 369.600 122.600 370.200 ;
        RECT 86.000 362.200 86.800 369.200 ;
        RECT 91.800 364.400 92.600 369.600 ;
        RECT 93.400 368.400 94.000 369.600 ;
        RECT 93.200 367.600 94.000 368.400 ;
        RECT 90.800 363.600 92.600 364.400 ;
        RECT 91.800 362.200 92.600 363.600 ;
        RECT 98.200 362.200 99.000 369.600 ;
        RECT 99.800 368.400 100.400 369.600 ;
        RECT 99.600 367.600 100.400 368.400 ;
        RECT 104.600 364.400 105.400 369.600 ;
        RECT 106.200 368.400 106.800 369.600 ;
        RECT 106.000 367.600 106.800 368.400 ;
        RECT 116.400 367.600 117.200 369.200 ;
        RECT 118.000 367.000 118.600 369.600 ;
        RECT 120.400 368.400 121.000 369.600 ;
        RECT 120.400 367.600 121.200 368.400 ;
        RECT 115.000 366.400 118.600 367.000 ;
        RECT 103.600 363.600 105.400 364.400 ;
        RECT 104.600 362.200 105.400 363.600 ;
        RECT 114.800 362.200 115.600 366.400 ;
        RECT 118.000 366.200 118.600 366.400 ;
        RECT 121.800 366.400 122.600 369.600 ;
        RECT 126.000 369.600 128.600 370.200 ;
        RECT 118.000 362.200 118.800 366.200 ;
        RECT 121.800 365.600 123.600 366.400 ;
        RECT 121.800 362.200 122.600 365.600 ;
        RECT 126.000 362.200 126.800 369.600 ;
        RECT 129.200 369.200 130.200 370.200 ;
        RECT 133.000 369.400 134.800 370.200 ;
        RECT 137.200 369.600 138.600 370.200 ;
        RECT 139.200 369.600 140.200 370.200 ;
        RECT 129.200 362.200 130.000 369.200 ;
        RECT 133.000 362.200 133.800 369.400 ;
        RECT 138.000 368.400 138.600 369.600 ;
        RECT 138.000 367.600 138.800 368.400 ;
        RECT 139.400 362.200 140.200 369.600 ;
        RECT 143.600 362.200 144.400 379.800 ;
        RECT 145.200 375.600 146.000 377.200 ;
        RECT 145.200 368.300 146.000 368.400 ;
        RECT 146.800 368.300 147.600 379.800 ;
        RECT 148.400 375.600 149.200 377.200 ;
        RECT 145.200 367.700 147.600 368.300 ;
        RECT 145.200 367.600 146.000 367.700 ;
        RECT 146.800 362.200 147.600 367.700 ;
        RECT 150.000 375.400 150.800 379.800 ;
        RECT 154.200 378.400 155.400 379.800 ;
        RECT 154.200 377.800 155.600 378.400 ;
        RECT 158.800 377.800 159.600 379.800 ;
        RECT 163.200 378.400 164.000 379.800 ;
        RECT 163.200 377.800 165.200 378.400 ;
        RECT 154.800 377.000 155.600 377.800 ;
        RECT 159.000 377.200 159.600 377.800 ;
        RECT 159.000 376.600 161.800 377.200 ;
        RECT 161.000 376.400 161.800 376.600 ;
        RECT 162.800 376.400 163.600 377.200 ;
        RECT 164.400 377.000 165.200 377.800 ;
        RECT 153.000 375.400 153.800 375.600 ;
        RECT 150.000 374.800 153.800 375.400 ;
        RECT 150.000 371.400 150.800 374.800 ;
        RECT 162.800 374.400 163.400 376.400 ;
        RECT 167.600 375.000 168.400 379.800 ;
        RECT 169.200 375.200 170.000 379.800 ;
        RECT 172.400 376.400 173.200 379.800 ;
        RECT 176.200 376.400 177.000 379.800 ;
        RECT 172.400 375.800 173.400 376.400 ;
        RECT 176.200 375.800 178.000 376.400 ;
        RECT 169.200 374.600 171.800 375.200 ;
        RECT 157.000 374.200 157.800 374.400 ;
        RECT 162.800 374.200 163.600 374.400 ;
        RECT 166.000 374.200 167.600 374.400 ;
        RECT 156.600 373.600 167.600 374.200 ;
        RECT 154.800 372.800 155.600 373.000 ;
        RECT 151.800 372.200 155.600 372.800 ;
        RECT 151.800 372.000 152.600 372.200 ;
        RECT 153.400 371.400 154.200 371.600 ;
        RECT 150.000 370.800 154.200 371.400 ;
        RECT 150.000 362.200 150.800 370.800 ;
        RECT 156.600 370.400 157.200 373.600 ;
        RECT 163.800 373.400 164.600 373.600 ;
        RECT 165.400 372.400 166.200 372.600 ;
        RECT 169.400 372.400 170.200 373.200 ;
        RECT 161.200 371.800 166.200 372.400 ;
        RECT 161.200 371.600 162.000 371.800 ;
        RECT 169.200 371.600 170.200 372.400 ;
        RECT 171.200 373.000 171.800 374.600 ;
        RECT 172.800 374.400 173.400 375.800 ;
        RECT 172.400 374.300 173.400 374.400 ;
        RECT 175.600 374.300 176.400 374.400 ;
        RECT 172.400 373.700 176.400 374.300 ;
        RECT 172.400 373.600 173.400 373.700 ;
        RECT 175.600 373.600 176.400 373.700 ;
        RECT 171.200 372.200 172.200 373.000 ;
        RECT 162.800 371.000 168.400 371.200 ;
        RECT 162.600 370.800 168.400 371.000 ;
        RECT 154.800 369.800 157.200 370.400 ;
        RECT 158.600 370.600 168.400 370.800 ;
        RECT 158.600 370.200 163.400 370.600 ;
        RECT 154.800 368.800 155.400 369.800 ;
        RECT 154.000 368.000 155.400 368.800 ;
        RECT 157.000 369.000 157.800 369.200 ;
        RECT 158.600 369.000 159.200 370.200 ;
        RECT 157.000 368.400 159.200 369.000 ;
        RECT 159.800 369.000 165.200 369.600 ;
        RECT 159.800 368.800 160.600 369.000 ;
        RECT 164.400 368.800 165.200 369.000 ;
        RECT 158.200 367.400 159.000 367.600 ;
        RECT 161.000 367.400 161.800 367.600 ;
        RECT 154.800 366.200 155.600 367.000 ;
        RECT 158.200 366.800 161.800 367.400 ;
        RECT 159.000 366.200 159.600 366.800 ;
        RECT 164.400 366.200 165.200 367.000 ;
        RECT 154.200 362.200 155.400 366.200 ;
        RECT 158.800 362.200 159.600 366.200 ;
        RECT 163.200 365.600 165.200 366.200 ;
        RECT 163.200 362.200 164.000 365.600 ;
        RECT 167.600 362.200 168.400 370.600 ;
        RECT 171.200 370.200 171.800 372.200 ;
        RECT 172.800 370.200 173.400 373.600 ;
        RECT 174.000 372.300 174.800 372.400 ;
        RECT 174.000 371.700 176.300 372.300 ;
        RECT 174.000 371.600 174.800 371.700 ;
        RECT 175.700 370.400 176.300 371.700 ;
        RECT 169.200 369.600 171.800 370.200 ;
        RECT 169.200 362.200 170.000 369.600 ;
        RECT 172.400 369.200 173.400 370.200 ;
        RECT 172.400 362.200 173.200 369.200 ;
        RECT 175.600 368.800 176.400 370.400 ;
        RECT 177.200 362.200 178.000 375.800 ;
        RECT 178.800 373.600 179.600 375.200 ;
        RECT 180.400 373.800 181.200 379.800 ;
        RECT 186.800 376.600 187.600 379.800 ;
        RECT 188.400 377.000 189.200 379.800 ;
        RECT 190.000 377.000 190.800 379.800 ;
        RECT 191.600 377.000 192.400 379.800 ;
        RECT 194.800 377.000 195.600 379.800 ;
        RECT 198.000 377.000 198.800 379.800 ;
        RECT 199.600 377.000 200.400 379.800 ;
        RECT 201.200 377.000 202.000 379.800 ;
        RECT 202.800 377.000 203.600 379.800 ;
        RECT 185.000 375.800 187.600 376.600 ;
        RECT 204.400 376.600 205.200 379.800 ;
        RECT 191.000 375.800 195.600 376.400 ;
        RECT 185.000 375.200 185.800 375.800 ;
        RECT 182.800 374.400 185.800 375.200 ;
        RECT 180.400 373.000 189.200 373.800 ;
        RECT 191.000 373.400 191.800 375.800 ;
        RECT 194.800 375.600 195.600 375.800 ;
        RECT 196.400 375.600 198.000 376.400 ;
        RECT 201.000 375.600 202.000 376.400 ;
        RECT 204.400 375.800 206.800 376.600 ;
        RECT 193.200 373.600 194.000 375.200 ;
        RECT 194.800 374.800 195.600 375.000 ;
        RECT 194.800 374.200 199.200 374.800 ;
        RECT 198.400 374.000 199.200 374.200 ;
        RECT 180.400 367.400 181.200 373.000 ;
        RECT 189.800 372.600 191.800 373.400 ;
        RECT 195.600 372.600 198.800 373.400 ;
        RECT 201.200 372.800 202.000 375.600 ;
        RECT 206.000 375.200 206.800 375.800 ;
        RECT 206.000 374.600 207.800 375.200 ;
        RECT 207.000 373.400 207.800 374.600 ;
        RECT 210.800 374.600 211.600 379.800 ;
        RECT 212.400 376.000 213.200 379.800 ;
        RECT 212.400 375.200 213.400 376.000 ;
        RECT 215.600 375.800 216.400 379.800 ;
        RECT 217.200 376.000 218.000 379.800 ;
        RECT 220.400 376.000 221.200 379.800 ;
        RECT 217.200 375.800 221.200 376.000 ;
        RECT 210.800 374.000 212.000 374.600 ;
        RECT 207.000 372.600 210.800 373.400 ;
        RECT 181.800 372.000 182.600 372.200 ;
        RECT 183.600 372.000 184.400 372.400 ;
        RECT 186.800 372.000 187.600 372.400 ;
        RECT 204.400 372.000 205.200 372.600 ;
        RECT 211.400 372.000 212.000 374.000 ;
        RECT 181.800 371.400 205.200 372.000 ;
        RECT 211.200 371.400 212.000 372.000 ;
        RECT 211.200 369.600 211.800 371.400 ;
        RECT 212.600 370.800 213.400 375.200 ;
        RECT 215.800 374.400 216.400 375.800 ;
        RECT 217.400 375.400 221.000 375.800 ;
        RECT 222.000 375.200 222.800 379.800 ;
        RECT 226.800 375.200 227.600 379.800 ;
        RECT 230.000 376.400 230.800 379.800 ;
        RECT 233.800 376.400 234.600 379.800 ;
        RECT 230.000 375.800 231.000 376.400 ;
        RECT 233.800 375.800 235.600 376.400 ;
        RECT 219.600 374.400 220.400 374.800 ;
        RECT 222.000 374.600 224.200 375.200 ;
        RECT 226.800 374.600 229.400 375.200 ;
        RECT 214.000 374.300 214.800 374.400 ;
        RECT 215.600 374.300 218.200 374.400 ;
        RECT 214.000 373.700 218.200 374.300 ;
        RECT 219.600 373.800 221.200 374.400 ;
        RECT 214.000 373.600 214.800 373.700 ;
        RECT 215.600 373.600 218.200 373.700 ;
        RECT 220.400 373.600 221.200 373.800 ;
        RECT 190.000 369.400 190.800 369.600 ;
        RECT 185.400 369.000 190.800 369.400 ;
        RECT 184.600 368.800 190.800 369.000 ;
        RECT 191.800 369.000 200.400 369.600 ;
        RECT 182.000 368.000 183.600 368.800 ;
        RECT 184.600 368.200 186.000 368.800 ;
        RECT 191.800 368.200 192.400 369.000 ;
        RECT 199.600 368.800 200.400 369.000 ;
        RECT 202.800 369.000 211.800 369.600 ;
        RECT 202.800 368.800 203.600 369.000 ;
        RECT 183.000 367.600 183.600 368.000 ;
        RECT 186.600 367.600 192.400 368.200 ;
        RECT 193.000 367.600 195.600 368.400 ;
        RECT 180.400 366.800 182.400 367.400 ;
        RECT 183.000 366.800 187.200 367.600 ;
        RECT 181.800 366.200 182.400 366.800 ;
        RECT 181.800 365.600 182.800 366.200 ;
        RECT 182.000 362.200 182.800 365.600 ;
        RECT 185.200 362.200 186.000 366.800 ;
        RECT 188.400 362.200 189.200 365.000 ;
        RECT 190.000 362.200 190.800 365.000 ;
        RECT 191.600 362.200 192.400 367.000 ;
        RECT 194.800 362.200 195.600 367.000 ;
        RECT 198.000 362.200 198.800 368.400 ;
        RECT 206.000 367.600 208.600 368.400 ;
        RECT 201.200 366.800 205.400 367.600 ;
        RECT 199.600 362.200 200.400 365.000 ;
        RECT 201.200 362.200 202.000 365.000 ;
        RECT 202.800 362.200 203.600 365.000 ;
        RECT 206.000 362.200 206.800 367.600 ;
        RECT 211.200 367.400 211.800 369.000 ;
        RECT 209.200 366.800 211.800 367.400 ;
        RECT 212.400 370.300 213.400 370.800 ;
        RECT 215.600 370.300 216.400 370.400 ;
        RECT 212.400 370.200 216.400 370.300 ;
        RECT 217.600 370.200 218.200 373.600 ;
        RECT 218.800 372.300 219.600 373.200 ;
        RECT 220.400 372.300 221.200 372.400 ;
        RECT 218.800 371.700 221.200 372.300 ;
        RECT 218.800 371.600 219.600 371.700 ;
        RECT 220.400 371.600 221.200 371.700 ;
        RECT 222.000 371.600 222.800 373.200 ;
        RECT 223.600 371.600 224.200 374.600 ;
        RECT 227.000 372.400 227.800 373.200 ;
        RECT 226.800 371.600 227.800 372.400 ;
        RECT 228.800 373.000 229.400 374.600 ;
        RECT 230.400 374.400 231.000 375.800 ;
        RECT 230.000 373.600 231.000 374.400 ;
        RECT 228.800 372.200 229.800 373.000 ;
        RECT 223.600 370.800 224.800 371.600 ;
        RECT 223.600 370.200 224.200 370.800 ;
        RECT 228.800 370.200 229.400 372.200 ;
        RECT 230.400 370.200 231.000 373.600 ;
        RECT 212.400 369.700 217.000 370.200 ;
        RECT 209.200 362.200 210.000 366.800 ;
        RECT 212.400 362.200 213.200 369.700 ;
        RECT 215.600 369.600 217.000 369.700 ;
        RECT 217.600 369.600 218.600 370.200 ;
        RECT 216.400 368.400 217.000 369.600 ;
        RECT 216.400 367.600 217.200 368.400 ;
        RECT 217.800 362.200 218.600 369.600 ;
        RECT 222.000 369.600 224.200 370.200 ;
        RECT 226.800 369.600 229.400 370.200 ;
        RECT 222.000 362.200 222.800 369.600 ;
        RECT 226.800 362.200 227.600 369.600 ;
        RECT 230.000 369.200 231.000 370.200 ;
        RECT 230.000 362.200 230.800 369.200 ;
        RECT 233.200 368.800 234.000 370.400 ;
        RECT 234.800 362.200 235.600 375.800 ;
        RECT 236.400 373.600 237.200 375.200 ;
        RECT 238.000 373.800 238.800 379.800 ;
        RECT 244.400 376.600 245.200 379.800 ;
        RECT 246.000 377.000 246.800 379.800 ;
        RECT 247.600 377.000 248.400 379.800 ;
        RECT 249.200 377.000 250.000 379.800 ;
        RECT 252.400 377.000 253.200 379.800 ;
        RECT 255.600 377.000 256.400 379.800 ;
        RECT 257.200 377.000 258.000 379.800 ;
        RECT 258.800 377.000 259.600 379.800 ;
        RECT 260.400 377.000 261.200 379.800 ;
        RECT 242.600 375.800 245.200 376.600 ;
        RECT 262.000 376.600 262.800 379.800 ;
        RECT 248.600 375.800 253.200 376.400 ;
        RECT 242.600 375.200 243.400 375.800 ;
        RECT 240.400 374.400 243.400 375.200 ;
        RECT 238.000 373.000 246.800 373.800 ;
        RECT 248.600 373.400 249.400 375.800 ;
        RECT 252.400 375.600 253.200 375.800 ;
        RECT 254.000 375.600 255.600 376.400 ;
        RECT 258.600 375.600 259.600 376.400 ;
        RECT 262.000 375.800 264.400 376.600 ;
        RECT 250.800 373.600 251.600 375.200 ;
        RECT 252.400 374.800 253.200 375.000 ;
        RECT 252.400 374.200 256.800 374.800 ;
        RECT 256.000 374.000 256.800 374.200 ;
        RECT 238.000 367.400 238.800 373.000 ;
        RECT 247.400 372.600 249.400 373.400 ;
        RECT 253.200 372.600 256.400 373.400 ;
        RECT 258.800 372.800 259.600 375.600 ;
        RECT 263.600 375.200 264.400 375.800 ;
        RECT 263.600 374.600 265.400 375.200 ;
        RECT 264.600 373.400 265.400 374.600 ;
        RECT 268.400 374.600 269.200 379.800 ;
        RECT 270.000 376.000 270.800 379.800 ;
        RECT 270.000 375.200 271.000 376.000 ;
        RECT 278.000 375.800 278.800 379.800 ;
        RECT 279.600 376.000 280.400 379.800 ;
        RECT 282.800 376.000 283.600 379.800 ;
        RECT 279.600 375.800 283.600 376.000 ;
        RECT 268.400 374.000 269.600 374.600 ;
        RECT 264.600 372.600 268.400 373.400 ;
        RECT 239.400 372.000 240.200 372.200 ;
        RECT 241.200 372.000 242.000 372.400 ;
        RECT 244.400 372.000 245.200 372.400 ;
        RECT 262.000 372.000 262.800 372.600 ;
        RECT 269.000 372.000 269.600 374.000 ;
        RECT 239.400 371.400 262.800 372.000 ;
        RECT 268.800 371.400 269.600 372.000 ;
        RECT 268.800 369.600 269.400 371.400 ;
        RECT 270.200 370.800 271.000 375.200 ;
        RECT 278.200 374.400 278.800 375.800 ;
        RECT 279.800 375.400 283.400 375.800 ;
        RECT 284.400 375.200 285.200 379.800 ;
        RECT 287.600 376.400 288.400 379.800 ;
        RECT 287.600 375.600 288.600 376.400 ;
        RECT 282.000 374.400 282.800 374.800 ;
        RECT 284.400 374.600 287.000 375.200 ;
        RECT 271.600 374.300 272.400 374.400 ;
        RECT 278.000 374.300 280.600 374.400 ;
        RECT 271.600 373.700 280.600 374.300 ;
        RECT 282.000 373.800 283.600 374.400 ;
        RECT 271.600 373.600 272.400 373.700 ;
        RECT 278.000 373.600 280.600 373.700 ;
        RECT 282.800 373.600 283.600 373.800 ;
        RECT 247.600 369.400 248.400 369.600 ;
        RECT 243.000 369.000 248.400 369.400 ;
        RECT 242.200 368.800 248.400 369.000 ;
        RECT 249.400 369.000 258.000 369.600 ;
        RECT 239.600 368.000 241.200 368.800 ;
        RECT 242.200 368.200 243.600 368.800 ;
        RECT 249.400 368.200 250.000 369.000 ;
        RECT 257.200 368.800 258.000 369.000 ;
        RECT 260.400 369.000 269.400 369.600 ;
        RECT 260.400 368.800 261.200 369.000 ;
        RECT 240.600 367.600 241.200 368.000 ;
        RECT 244.200 367.600 250.000 368.200 ;
        RECT 250.600 367.600 253.200 368.400 ;
        RECT 238.000 366.800 240.000 367.400 ;
        RECT 240.600 366.800 244.800 367.600 ;
        RECT 239.400 366.200 240.000 366.800 ;
        RECT 239.400 365.600 240.400 366.200 ;
        RECT 239.600 362.200 240.400 365.600 ;
        RECT 242.800 362.200 243.600 366.800 ;
        RECT 246.000 362.200 246.800 365.000 ;
        RECT 247.600 362.200 248.400 365.000 ;
        RECT 249.200 362.200 250.000 367.000 ;
        RECT 252.400 362.200 253.200 367.000 ;
        RECT 255.600 362.200 256.400 368.400 ;
        RECT 263.600 367.600 266.200 368.400 ;
        RECT 258.800 366.800 263.000 367.600 ;
        RECT 257.200 362.200 258.000 365.000 ;
        RECT 258.800 362.200 259.600 365.000 ;
        RECT 260.400 362.200 261.200 365.000 ;
        RECT 263.600 362.200 264.400 367.600 ;
        RECT 268.800 367.400 269.400 369.000 ;
        RECT 266.800 366.800 269.400 367.400 ;
        RECT 270.000 370.300 271.000 370.800 ;
        RECT 278.000 370.300 278.800 370.400 ;
        RECT 270.000 370.200 278.800 370.300 ;
        RECT 280.000 370.200 280.600 373.600 ;
        RECT 281.200 371.600 282.000 373.200 ;
        RECT 284.600 372.400 285.400 373.200 ;
        RECT 284.400 371.600 285.400 372.400 ;
        RECT 286.400 373.000 287.000 374.600 ;
        RECT 288.000 374.400 288.600 375.600 ;
        RECT 292.400 375.200 293.200 379.800 ;
        RECT 295.600 375.200 296.400 379.800 ;
        RECT 298.800 375.200 299.600 379.800 ;
        RECT 302.000 375.200 302.800 379.800 ;
        RECT 305.200 375.600 306.000 377.200 ;
        RECT 292.400 374.400 294.200 375.200 ;
        RECT 295.600 374.400 297.800 375.200 ;
        RECT 298.800 374.400 301.000 375.200 ;
        RECT 302.000 374.400 304.400 375.200 ;
        RECT 287.600 373.600 288.600 374.400 ;
        RECT 286.400 372.200 287.400 373.000 ;
        RECT 286.400 370.200 287.000 372.200 ;
        RECT 288.000 370.200 288.600 373.600 ;
        RECT 290.800 373.800 291.600 374.400 ;
        RECT 293.400 373.800 294.200 374.400 ;
        RECT 297.000 373.800 297.800 374.400 ;
        RECT 300.200 373.800 301.000 374.400 ;
        RECT 290.800 373.000 292.600 373.800 ;
        RECT 293.400 373.000 296.000 373.800 ;
        RECT 297.000 373.000 299.400 373.800 ;
        RECT 300.200 373.000 302.800 373.800 ;
        RECT 293.400 371.600 294.200 373.000 ;
        RECT 297.000 371.600 297.800 373.000 ;
        RECT 300.200 371.600 301.000 373.000 ;
        RECT 303.600 371.600 304.400 374.400 ;
        RECT 270.000 369.700 279.400 370.200 ;
        RECT 266.800 362.200 267.600 366.800 ;
        RECT 270.000 362.200 270.800 369.700 ;
        RECT 278.000 369.600 279.400 369.700 ;
        RECT 280.000 369.600 281.000 370.200 ;
        RECT 278.800 368.400 279.400 369.600 ;
        RECT 278.000 367.600 279.600 368.400 ;
        RECT 280.200 362.200 281.000 369.600 ;
        RECT 284.400 369.600 287.000 370.200 ;
        RECT 284.400 362.200 285.200 369.600 ;
        RECT 287.600 369.200 288.600 370.200 ;
        RECT 292.400 370.800 294.200 371.600 ;
        RECT 295.600 370.800 297.800 371.600 ;
        RECT 298.800 370.800 301.000 371.600 ;
        RECT 302.000 370.800 304.400 371.600 ;
        RECT 306.800 372.300 307.600 379.800 ;
        RECT 308.400 376.000 309.200 379.800 ;
        RECT 311.600 376.000 312.400 379.800 ;
        RECT 308.400 375.800 312.400 376.000 ;
        RECT 313.200 375.800 314.000 379.800 ;
        RECT 317.400 376.400 319.000 379.800 ;
        RECT 316.400 375.800 319.000 376.400 ;
        RECT 308.600 375.400 312.200 375.800 ;
        RECT 309.200 374.400 310.000 374.800 ;
        RECT 313.200 374.400 313.800 375.800 ;
        RECT 316.400 375.600 318.600 375.800 ;
        RECT 308.400 373.800 310.000 374.400 ;
        RECT 308.400 373.600 309.200 373.800 ;
        RECT 311.400 373.600 314.000 374.400 ;
        RECT 316.400 373.600 317.200 374.400 ;
        RECT 308.400 372.300 309.200 372.400 ;
        RECT 306.800 371.700 309.200 372.300 ;
        RECT 287.600 362.200 288.400 369.200 ;
        RECT 292.400 362.200 293.200 370.800 ;
        RECT 295.600 362.200 296.400 370.800 ;
        RECT 298.800 362.200 299.600 370.800 ;
        RECT 302.000 362.200 302.800 370.800 ;
        RECT 306.800 362.200 307.600 371.700 ;
        RECT 308.400 371.600 309.200 371.700 ;
        RECT 310.000 371.600 310.800 373.200 ;
        RECT 311.400 370.200 312.000 373.600 ;
        RECT 316.600 373.200 317.200 373.600 ;
        RECT 316.600 372.400 317.400 373.200 ;
        RECT 318.000 372.400 318.600 375.600 ;
        RECT 319.600 372.800 320.400 374.400 ;
        RECT 314.800 370.800 315.600 372.400 ;
        RECT 318.000 371.600 318.800 372.400 ;
        RECT 321.200 372.300 322.000 372.400 ;
        RECT 322.800 372.300 323.600 379.800 ;
        RECT 324.400 375.600 325.200 377.200 ;
        RECT 326.000 375.600 326.800 377.200 ;
        RECT 324.400 374.300 325.200 374.400 ;
        RECT 327.600 374.300 328.400 379.800 ;
        RECT 332.200 375.800 333.800 379.800 ;
        RECT 340.800 376.400 341.600 379.800 ;
        RECT 330.800 374.300 331.600 374.400 ;
        RECT 324.400 373.700 331.600 374.300 ;
        RECT 324.400 373.600 325.200 373.700 ;
        RECT 326.000 372.300 326.800 372.400 ;
        RECT 321.200 372.200 326.800 372.300 ;
        RECT 320.400 371.700 326.800 372.200 ;
        RECT 320.400 371.600 322.000 371.700 ;
        RECT 318.000 371.400 318.600 371.600 ;
        RECT 316.600 370.800 318.600 371.400 ;
        RECT 320.400 371.200 321.200 371.600 ;
        RECT 313.200 370.200 314.000 370.400 ;
        RECT 316.600 370.200 317.200 370.800 ;
        RECT 311.000 369.600 312.000 370.200 ;
        RECT 312.600 369.600 314.000 370.200 ;
        RECT 311.000 362.200 311.800 369.600 ;
        RECT 312.600 368.400 313.200 369.600 ;
        RECT 312.400 367.600 313.200 368.400 ;
        RECT 314.800 362.800 315.600 370.200 ;
        RECT 316.400 363.400 317.200 370.200 ;
        RECT 318.000 369.600 322.000 370.200 ;
        RECT 318.000 362.800 318.800 369.600 ;
        RECT 314.800 362.200 318.800 362.800 ;
        RECT 321.200 362.200 322.000 369.600 ;
        RECT 322.800 362.200 323.600 371.700 ;
        RECT 326.000 371.600 326.800 371.700 ;
        RECT 327.600 362.200 328.400 373.700 ;
        RECT 330.800 372.800 331.600 373.700 ;
        RECT 332.600 372.400 333.200 375.800 ;
        RECT 340.800 375.600 342.800 376.400 ;
        RECT 334.000 373.600 334.800 374.400 ;
        RECT 340.800 374.200 341.600 375.600 ;
        RECT 347.200 374.200 348.000 379.800 ;
        RECT 351.200 374.200 352.000 379.800 ;
        RECT 356.400 375.600 357.200 377.200 ;
        RECT 340.800 373.800 342.600 374.200 ;
        RECT 347.200 373.800 349.000 374.200 ;
        RECT 341.000 373.600 342.600 373.800 ;
        RECT 347.400 373.600 349.000 373.800 ;
        RECT 334.000 373.200 334.600 373.600 ;
        RECT 333.800 372.400 334.600 373.200 ;
        RECT 329.200 372.200 330.000 372.400 ;
        RECT 329.200 371.600 330.800 372.200 ;
        RECT 332.400 371.600 333.200 372.400 ;
        RECT 330.000 371.200 330.800 371.600 ;
        RECT 332.600 371.400 333.200 371.600 ;
        RECT 332.600 370.800 334.600 371.400 ;
        RECT 335.600 370.800 336.400 372.400 ;
        RECT 338.800 371.600 340.400 372.400 ;
        RECT 334.000 370.200 334.600 370.800 ;
        RECT 329.200 369.600 333.200 370.200 ;
        RECT 329.200 362.200 330.000 369.600 ;
        RECT 332.400 362.800 333.200 369.600 ;
        RECT 334.000 363.400 334.800 370.200 ;
        RECT 335.600 362.800 336.400 370.200 ;
        RECT 337.200 369.600 338.000 371.200 ;
        RECT 342.000 370.400 342.600 373.600 ;
        RECT 345.200 371.600 347.600 372.400 ;
        RECT 342.000 369.600 342.800 370.400 ;
        RECT 343.600 369.600 344.400 371.200 ;
        RECT 348.400 370.400 349.000 373.600 ;
        RECT 350.200 373.800 352.000 374.200 ;
        RECT 350.200 373.600 351.800 373.800 ;
        RECT 350.200 370.400 350.800 373.600 ;
        RECT 352.400 371.600 354.000 372.400 ;
        RECT 348.400 369.600 349.200 370.400 ;
        RECT 350.000 369.600 350.800 370.400 ;
        RECT 354.800 369.600 355.600 371.200 ;
        RECT 340.400 367.600 341.200 369.200 ;
        RECT 342.000 367.000 342.600 369.600 ;
        RECT 345.200 368.300 346.000 368.400 ;
        RECT 346.800 368.300 347.600 369.200 ;
        RECT 345.200 367.700 347.600 368.300 ;
        RECT 345.200 367.600 346.000 367.700 ;
        RECT 346.800 367.600 347.600 367.700 ;
        RECT 348.400 367.000 349.000 369.600 ;
        RECT 339.000 366.400 342.600 367.000 ;
        RECT 339.000 366.200 339.600 366.400 ;
        RECT 332.400 362.200 336.400 362.800 ;
        RECT 338.800 362.200 339.600 366.200 ;
        RECT 342.000 366.200 342.600 366.400 ;
        RECT 345.400 366.400 349.000 367.000 ;
        RECT 350.200 367.000 350.800 369.600 ;
        RECT 351.600 368.300 352.400 369.200 ;
        RECT 356.400 368.300 357.200 368.400 ;
        RECT 351.600 367.700 357.200 368.300 ;
        RECT 351.600 367.600 352.400 367.700 ;
        RECT 356.400 367.600 357.200 367.700 ;
        RECT 350.200 366.400 353.800 367.000 ;
        RECT 345.400 366.200 346.000 366.400 ;
        RECT 342.000 362.200 342.800 366.200 ;
        RECT 345.200 362.200 346.000 366.200 ;
        RECT 348.400 362.200 349.200 366.400 ;
        RECT 350.200 366.200 350.800 366.400 ;
        RECT 350.000 362.200 350.800 366.200 ;
        RECT 353.200 366.200 353.800 366.400 ;
        RECT 353.200 362.200 354.000 366.200 ;
        RECT 358.000 362.200 358.800 379.800 ;
        RECT 362.200 375.800 363.800 379.800 ;
        RECT 361.200 373.600 362.000 374.400 ;
        RECT 361.400 373.200 362.000 373.600 ;
        RECT 361.400 372.400 362.200 373.200 ;
        RECT 362.800 372.400 363.400 375.800 ;
        RECT 367.600 375.600 368.400 377.200 ;
        RECT 364.400 374.300 365.200 374.400 ;
        RECT 369.200 374.300 370.000 379.800 ;
        RECT 373.800 375.800 375.400 379.800 ;
        RECT 372.400 374.300 373.200 374.400 ;
        RECT 364.400 373.700 373.200 374.300 ;
        RECT 364.400 372.800 365.200 373.700 ;
        RECT 359.600 370.800 360.400 372.400 ;
        RECT 362.800 371.600 363.600 372.400 ;
        RECT 366.000 372.200 366.800 372.400 ;
        RECT 365.200 371.600 366.800 372.200 ;
        RECT 362.800 371.400 363.400 371.600 ;
        RECT 361.400 370.800 363.400 371.400 ;
        RECT 365.200 371.200 366.000 371.600 ;
        RECT 361.400 370.200 362.000 370.800 ;
        RECT 359.600 362.800 360.400 370.200 ;
        RECT 361.200 363.400 362.000 370.200 ;
        RECT 362.800 369.600 366.800 370.200 ;
        RECT 362.800 362.800 363.600 369.600 ;
        RECT 359.600 362.200 363.600 362.800 ;
        RECT 366.000 362.200 366.800 369.600 ;
        RECT 369.200 362.200 370.000 373.700 ;
        RECT 372.400 372.800 373.200 373.700 ;
        RECT 374.200 372.400 374.800 375.800 ;
        RECT 375.600 373.600 376.400 374.400 ;
        RECT 380.000 374.200 380.800 379.800 ;
        RECT 379.000 373.800 380.800 374.200 ;
        RECT 388.800 374.200 389.600 379.800 ;
        RECT 395.200 374.200 396.000 379.800 ;
        RECT 399.600 377.600 400.400 379.800 ;
        RECT 398.000 375.600 398.800 377.200 ;
        RECT 399.800 374.400 400.400 377.600 ;
        RECT 404.400 375.200 405.200 379.800 ;
        RECT 407.600 375.200 408.400 379.800 ;
        RECT 417.200 376.000 418.000 379.800 ;
        RECT 404.400 374.400 408.400 375.200 ;
        RECT 388.800 373.800 390.600 374.200 ;
        RECT 395.200 373.800 397.000 374.200 ;
        RECT 379.000 373.600 380.600 373.800 ;
        RECT 389.000 373.600 390.600 373.800 ;
        RECT 395.400 373.600 397.000 373.800 ;
        RECT 399.600 373.600 400.400 374.400 ;
        RECT 375.600 373.200 376.200 373.600 ;
        RECT 375.400 372.400 376.200 373.200 ;
        RECT 370.800 372.200 371.600 372.400 ;
        RECT 370.800 371.600 372.400 372.200 ;
        RECT 374.000 371.600 374.800 372.400 ;
        RECT 371.600 371.200 372.400 371.600 ;
        RECT 374.200 371.400 374.800 371.600 ;
        RECT 374.200 370.800 376.200 371.400 ;
        RECT 377.200 370.800 378.000 372.400 ;
        RECT 375.600 370.200 376.200 370.800 ;
        RECT 379.000 370.400 379.600 373.600 ;
        RECT 381.200 371.600 382.800 372.400 ;
        RECT 386.800 371.600 388.400 372.400 ;
        RECT 370.800 369.600 374.800 370.200 ;
        RECT 370.800 362.200 371.600 369.600 ;
        RECT 374.000 362.800 374.800 369.600 ;
        RECT 375.600 363.400 376.400 370.200 ;
        RECT 377.200 362.800 378.000 370.200 ;
        RECT 378.800 369.600 379.600 370.400 ;
        RECT 383.600 369.600 384.400 371.200 ;
        RECT 385.200 369.600 386.000 371.200 ;
        RECT 390.000 370.400 390.600 373.600 ;
        RECT 393.200 371.600 394.800 372.400 ;
        RECT 390.000 369.600 390.800 370.400 ;
        RECT 391.600 369.600 392.400 371.200 ;
        RECT 396.400 370.400 397.000 373.600 ;
        RECT 396.400 369.600 397.200 370.400 ;
        RECT 399.800 370.200 400.400 373.600 ;
        RECT 401.200 372.300 402.000 372.400 ;
        RECT 402.800 372.300 403.600 372.400 ;
        RECT 401.200 371.700 403.600 372.300 ;
        RECT 401.200 370.800 402.000 371.700 ;
        RECT 402.800 371.600 403.600 371.700 ;
        RECT 407.600 371.600 408.400 374.400 ;
        RECT 404.400 370.800 408.400 371.600 ;
        RECT 379.000 367.000 379.600 369.600 ;
        RECT 380.400 367.600 381.200 369.200 ;
        RECT 383.700 368.300 384.300 369.600 ;
        RECT 383.700 367.700 387.500 368.300 ;
        RECT 386.900 367.000 387.500 367.700 ;
        RECT 388.400 367.600 389.200 369.200 ;
        RECT 390.000 367.000 390.600 369.600 ;
        RECT 394.800 367.600 395.600 369.200 ;
        RECT 396.400 367.000 397.000 369.600 ;
        RECT 399.600 369.400 401.400 370.200 ;
        RECT 379.000 366.400 382.600 367.000 ;
        RECT 379.000 366.200 379.600 366.400 ;
        RECT 374.000 362.200 378.000 362.800 ;
        RECT 378.800 362.200 379.600 366.200 ;
        RECT 382.000 366.200 382.600 366.400 ;
        RECT 386.900 366.400 390.600 367.000 ;
        RECT 393.400 366.400 397.000 367.000 ;
        RECT 386.900 366.200 387.600 366.400 ;
        RECT 382.000 362.200 382.800 366.200 ;
        RECT 386.800 362.200 387.600 366.200 ;
        RECT 390.000 366.200 390.600 366.400 ;
        RECT 390.000 362.200 390.800 366.200 ;
        RECT 393.200 362.200 394.000 366.400 ;
        RECT 396.400 366.200 397.000 366.400 ;
        RECT 396.400 362.200 397.200 366.200 ;
        RECT 400.600 364.400 401.400 369.400 ;
        RECT 400.600 363.600 402.000 364.400 ;
        RECT 400.600 362.200 401.400 363.600 ;
        RECT 404.400 362.200 405.200 370.800 ;
        RECT 407.600 362.200 408.400 370.800 ;
        RECT 417.000 375.200 418.000 376.000 ;
        RECT 417.000 370.800 417.800 375.200 ;
        RECT 418.800 374.600 419.600 379.800 ;
        RECT 425.200 376.600 426.000 379.800 ;
        RECT 426.800 377.000 427.600 379.800 ;
        RECT 428.400 377.000 429.200 379.800 ;
        RECT 430.000 377.000 430.800 379.800 ;
        RECT 431.600 377.000 432.400 379.800 ;
        RECT 434.800 377.000 435.600 379.800 ;
        RECT 438.000 377.000 438.800 379.800 ;
        RECT 439.600 377.000 440.400 379.800 ;
        RECT 441.200 377.000 442.000 379.800 ;
        RECT 423.600 375.800 426.000 376.600 ;
        RECT 442.800 376.600 443.600 379.800 ;
        RECT 423.600 375.200 424.400 375.800 ;
        RECT 418.400 374.000 419.600 374.600 ;
        RECT 422.600 374.600 424.400 375.200 ;
        RECT 428.400 375.600 429.400 376.400 ;
        RECT 432.400 375.600 434.000 376.400 ;
        RECT 434.800 375.800 439.400 376.400 ;
        RECT 442.800 375.800 445.400 376.600 ;
        RECT 434.800 375.600 435.600 375.800 ;
        RECT 418.400 372.000 419.000 374.000 ;
        RECT 422.600 373.400 423.400 374.600 ;
        RECT 419.600 372.600 423.400 373.400 ;
        RECT 428.400 372.800 429.200 375.600 ;
        RECT 434.800 374.800 435.600 375.000 ;
        RECT 431.200 374.200 435.600 374.800 ;
        RECT 431.200 374.000 432.000 374.200 ;
        RECT 436.400 373.600 437.200 375.200 ;
        RECT 438.600 373.400 439.400 375.800 ;
        RECT 444.600 375.200 445.400 375.800 ;
        RECT 444.600 374.400 447.600 375.200 ;
        RECT 449.200 373.800 450.000 379.800 ;
        RECT 431.600 372.600 434.800 373.400 ;
        RECT 438.600 372.600 440.600 373.400 ;
        RECT 441.200 373.000 450.000 373.800 ;
        RECT 425.200 372.000 426.000 372.600 ;
        RECT 442.800 372.000 443.600 372.400 ;
        RECT 446.000 372.000 446.800 372.400 ;
        RECT 447.800 372.000 448.600 372.200 ;
        RECT 418.400 371.400 419.200 372.000 ;
        RECT 425.200 371.400 448.600 372.000 ;
        RECT 417.000 370.000 418.000 370.800 ;
        RECT 417.200 362.200 418.000 370.000 ;
        RECT 418.600 369.600 419.200 371.400 ;
        RECT 418.600 369.000 427.600 369.600 ;
        RECT 418.600 367.400 419.200 369.000 ;
        RECT 426.800 368.800 427.600 369.000 ;
        RECT 430.000 369.000 438.600 369.600 ;
        RECT 430.000 368.800 430.800 369.000 ;
        RECT 421.800 367.600 424.400 368.400 ;
        RECT 418.600 366.800 421.200 367.400 ;
        RECT 420.400 362.200 421.200 366.800 ;
        RECT 423.600 362.200 424.400 367.600 ;
        RECT 425.000 366.800 429.200 367.600 ;
        RECT 426.800 362.200 427.600 365.000 ;
        RECT 428.400 362.200 429.200 365.000 ;
        RECT 430.000 362.200 430.800 365.000 ;
        RECT 431.600 362.200 432.400 368.400 ;
        RECT 434.800 367.600 437.400 368.400 ;
        RECT 438.000 368.200 438.600 369.000 ;
        RECT 439.600 369.400 440.400 369.600 ;
        RECT 439.600 369.000 445.000 369.400 ;
        RECT 439.600 368.800 445.800 369.000 ;
        RECT 444.400 368.200 445.800 368.800 ;
        RECT 438.000 367.600 443.800 368.200 ;
        RECT 446.800 368.000 448.400 368.800 ;
        RECT 446.800 367.600 447.400 368.000 ;
        RECT 434.800 362.200 435.600 367.000 ;
        RECT 438.000 362.200 438.800 367.000 ;
        RECT 443.200 366.800 447.400 367.600 ;
        RECT 449.200 367.400 450.000 373.000 ;
        RECT 448.000 366.800 450.000 367.400 ;
        RECT 450.800 373.800 451.600 379.800 ;
        RECT 457.200 376.600 458.000 379.800 ;
        RECT 458.800 377.000 459.600 379.800 ;
        RECT 460.400 377.000 461.200 379.800 ;
        RECT 462.000 377.000 462.800 379.800 ;
        RECT 465.200 377.000 466.000 379.800 ;
        RECT 468.400 377.000 469.200 379.800 ;
        RECT 470.000 377.000 470.800 379.800 ;
        RECT 471.600 377.000 472.400 379.800 ;
        RECT 473.200 377.000 474.000 379.800 ;
        RECT 455.400 375.800 458.000 376.600 ;
        RECT 474.800 376.600 475.600 379.800 ;
        RECT 461.400 375.800 466.000 376.400 ;
        RECT 455.400 375.200 456.200 375.800 ;
        RECT 453.200 374.400 456.200 375.200 ;
        RECT 450.800 373.000 459.600 373.800 ;
        RECT 461.400 373.400 462.200 375.800 ;
        RECT 465.200 375.600 466.000 375.800 ;
        RECT 466.800 375.600 468.400 376.400 ;
        RECT 471.400 375.600 472.400 376.400 ;
        RECT 474.800 375.800 477.200 376.600 ;
        RECT 463.600 373.600 464.400 375.200 ;
        RECT 465.200 374.800 466.000 375.000 ;
        RECT 465.200 374.200 469.600 374.800 ;
        RECT 468.800 374.000 469.600 374.200 ;
        RECT 450.800 367.400 451.600 373.000 ;
        RECT 460.200 372.600 462.200 373.400 ;
        RECT 466.000 372.600 469.200 373.400 ;
        RECT 471.600 372.800 472.400 375.600 ;
        RECT 476.400 375.200 477.200 375.800 ;
        RECT 476.400 374.600 478.200 375.200 ;
        RECT 477.400 373.400 478.200 374.600 ;
        RECT 481.200 374.600 482.000 379.800 ;
        RECT 482.800 376.000 483.600 379.800 ;
        RECT 482.800 375.200 483.800 376.000 ;
        RECT 481.200 374.000 482.400 374.600 ;
        RECT 477.400 372.600 481.200 373.400 ;
        RECT 452.200 372.000 453.000 372.200 ;
        RECT 455.600 372.000 456.400 372.400 ;
        RECT 457.200 372.000 458.000 372.400 ;
        RECT 474.800 372.000 475.600 372.600 ;
        RECT 481.800 372.000 482.400 374.000 ;
        RECT 452.200 371.400 475.600 372.000 ;
        RECT 481.600 371.400 482.400 372.000 ;
        RECT 481.600 369.600 482.200 371.400 ;
        RECT 483.000 370.800 483.800 375.200 ;
        RECT 487.600 375.200 488.400 379.800 ;
        RECT 490.800 375.200 491.600 379.800 ;
        RECT 494.000 375.200 494.800 379.800 ;
        RECT 497.200 375.200 498.000 379.800 ;
        RECT 503.000 376.400 503.800 379.800 ;
        RECT 502.000 375.800 503.800 376.400 ;
        RECT 505.200 375.800 506.000 379.800 ;
        RECT 506.800 376.000 507.600 379.800 ;
        RECT 510.000 376.000 510.800 379.800 ;
        RECT 515.400 378.400 516.200 379.000 ;
        RECT 515.400 377.600 517.200 378.400 ;
        RECT 515.400 376.000 516.200 377.600 ;
        RECT 519.600 377.000 520.400 379.000 ;
        RECT 506.800 375.800 510.800 376.000 ;
        RECT 487.600 374.400 489.400 375.200 ;
        RECT 490.800 374.400 493.000 375.200 ;
        RECT 494.000 374.400 496.200 375.200 ;
        RECT 497.200 374.400 499.600 375.200 ;
        RECT 486.000 373.800 486.800 374.400 ;
        RECT 488.600 373.800 489.400 374.400 ;
        RECT 492.200 373.800 493.000 374.400 ;
        RECT 495.400 373.800 496.200 374.400 ;
        RECT 486.000 373.000 487.800 373.800 ;
        RECT 488.600 373.000 491.200 373.800 ;
        RECT 492.200 373.000 494.600 373.800 ;
        RECT 495.400 373.000 498.000 373.800 ;
        RECT 488.600 371.600 489.400 373.000 ;
        RECT 492.200 371.600 493.000 373.000 ;
        RECT 495.400 371.600 496.200 373.000 ;
        RECT 498.800 371.600 499.600 374.400 ;
        RECT 500.400 373.600 501.200 375.200 ;
        RECT 460.400 369.400 461.200 369.600 ;
        RECT 455.800 369.000 461.200 369.400 ;
        RECT 455.000 368.800 461.200 369.000 ;
        RECT 462.200 369.000 470.800 369.600 ;
        RECT 452.400 368.000 454.000 368.800 ;
        RECT 455.000 368.200 456.400 368.800 ;
        RECT 462.200 368.200 462.800 369.000 ;
        RECT 470.000 368.800 470.800 369.000 ;
        RECT 473.200 369.000 482.200 369.600 ;
        RECT 473.200 368.800 474.000 369.000 ;
        RECT 453.400 367.600 454.000 368.000 ;
        RECT 457.000 367.600 462.800 368.200 ;
        RECT 463.400 367.600 466.000 368.400 ;
        RECT 450.800 366.800 452.800 367.400 ;
        RECT 453.400 366.800 457.600 367.600 ;
        RECT 439.600 362.200 440.400 365.000 ;
        RECT 441.200 362.200 442.000 365.000 ;
        RECT 444.400 362.200 445.200 366.800 ;
        RECT 448.000 366.200 448.600 366.800 ;
        RECT 447.600 365.600 448.600 366.200 ;
        RECT 452.200 366.200 452.800 366.800 ;
        RECT 452.200 365.600 453.200 366.200 ;
        RECT 447.600 362.200 448.400 365.600 ;
        RECT 452.400 362.200 453.200 365.600 ;
        RECT 455.600 362.200 456.400 366.800 ;
        RECT 458.800 362.200 459.600 365.000 ;
        RECT 460.400 362.200 461.200 365.000 ;
        RECT 462.000 362.200 462.800 367.000 ;
        RECT 465.200 362.200 466.000 367.000 ;
        RECT 468.400 362.200 469.200 368.400 ;
        RECT 476.400 367.600 479.000 368.400 ;
        RECT 471.600 366.800 475.800 367.600 ;
        RECT 470.000 362.200 470.800 365.000 ;
        RECT 471.600 362.200 472.400 365.000 ;
        RECT 473.200 362.200 474.000 365.000 ;
        RECT 476.400 362.200 477.200 367.600 ;
        RECT 481.600 367.400 482.200 369.000 ;
        RECT 479.600 366.800 482.200 367.400 ;
        RECT 482.800 370.000 483.800 370.800 ;
        RECT 487.600 370.800 489.400 371.600 ;
        RECT 490.800 370.800 493.000 371.600 ;
        RECT 494.000 370.800 496.200 371.600 ;
        RECT 497.200 370.800 499.600 371.600 ;
        RECT 502.000 372.300 502.800 375.800 ;
        RECT 505.400 374.400 506.000 375.800 ;
        RECT 507.000 375.400 510.600 375.800 ;
        RECT 514.600 375.400 516.200 376.000 ;
        RECT 514.600 375.000 515.400 375.400 ;
        RECT 509.200 374.400 510.000 374.800 ;
        RECT 514.600 374.400 515.200 375.000 ;
        RECT 519.800 374.800 520.400 377.000 ;
        RECT 521.200 376.000 522.000 379.800 ;
        RECT 524.400 376.000 525.200 379.800 ;
        RECT 521.200 375.800 525.200 376.000 ;
        RECT 526.000 375.800 526.800 379.800 ;
        RECT 527.600 375.800 528.400 379.800 ;
        RECT 529.200 376.000 530.000 379.800 ;
        RECT 532.400 376.000 533.200 379.800 ;
        RECT 529.200 375.800 533.200 376.000 ;
        RECT 521.400 375.400 525.000 375.800 ;
        RECT 505.200 373.600 507.800 374.400 ;
        RECT 509.200 374.300 510.800 374.400 ;
        RECT 511.600 374.300 512.400 374.400 ;
        RECT 509.200 373.800 512.400 374.300 ;
        RECT 510.000 373.700 512.400 373.800 ;
        RECT 510.000 373.600 510.800 373.700 ;
        RECT 511.600 373.600 512.400 373.700 ;
        RECT 513.200 373.600 515.200 374.400 ;
        RECT 516.200 374.200 520.400 374.800 ;
        RECT 522.000 374.400 522.800 374.800 ;
        RECT 526.000 374.400 526.600 375.800 ;
        RECT 527.800 374.400 528.400 375.800 ;
        RECT 529.400 375.400 533.000 375.800 ;
        RECT 531.600 374.400 532.400 374.800 ;
        RECT 516.200 373.800 517.200 374.200 ;
        RECT 502.000 371.700 505.900 372.300 ;
        RECT 479.600 362.200 480.400 366.800 ;
        RECT 482.800 362.200 483.600 370.000 ;
        RECT 487.600 362.200 488.400 370.800 ;
        RECT 490.800 362.200 491.600 370.800 ;
        RECT 494.000 362.200 494.800 370.800 ;
        RECT 497.200 362.200 498.000 370.800 ;
        RECT 502.000 362.200 502.800 371.700 ;
        RECT 505.300 370.400 505.900 371.700 ;
        RECT 507.200 370.400 507.800 373.600 ;
        RECT 508.400 371.600 509.200 373.200 ;
        RECT 510.000 372.300 510.800 372.400 ;
        RECT 513.200 372.300 514.000 372.400 ;
        RECT 510.000 371.700 514.000 372.300 ;
        RECT 510.000 371.600 510.800 371.700 ;
        RECT 513.200 370.800 514.000 371.700 ;
        RECT 503.600 368.800 504.400 370.400 ;
        RECT 505.200 370.200 506.000 370.400 ;
        RECT 505.200 369.600 506.600 370.200 ;
        RECT 507.200 369.600 509.200 370.400 ;
        RECT 514.600 369.800 515.200 373.600 ;
        RECT 515.800 373.000 517.200 373.800 ;
        RECT 521.200 373.800 522.800 374.400 ;
        RECT 521.200 373.600 522.000 373.800 ;
        RECT 524.200 373.600 526.800 374.400 ;
        RECT 527.600 373.600 530.200 374.400 ;
        RECT 531.600 373.800 533.200 374.400 ;
        RECT 537.600 374.200 538.400 379.800 ;
        RECT 544.200 378.400 545.000 379.000 ;
        RECT 543.600 377.600 545.000 378.400 ;
        RECT 544.200 376.000 545.000 377.600 ;
        RECT 548.400 377.000 549.200 379.000 ;
        RECT 543.400 375.400 545.000 376.000 ;
        RECT 543.400 375.000 544.200 375.400 ;
        RECT 543.400 374.400 544.000 375.000 ;
        RECT 548.600 374.800 549.200 377.000 ;
        RECT 537.600 373.800 539.400 374.200 ;
        RECT 532.400 373.600 533.200 373.800 ;
        RECT 537.800 373.600 539.400 373.800 ;
        RECT 542.000 373.600 544.000 374.400 ;
        RECT 545.000 374.200 549.200 374.800 ;
        RECT 550.000 375.400 550.800 379.800 ;
        RECT 554.200 378.400 555.400 379.800 ;
        RECT 554.200 377.800 555.600 378.400 ;
        RECT 558.800 377.800 559.600 379.800 ;
        RECT 563.200 378.400 564.000 379.800 ;
        RECT 563.200 377.800 565.200 378.400 ;
        RECT 554.800 377.000 555.600 377.800 ;
        RECT 559.000 377.200 559.600 377.800 ;
        RECT 559.000 376.600 561.800 377.200 ;
        RECT 561.000 376.400 561.800 376.600 ;
        RECT 562.800 376.400 563.600 377.200 ;
        RECT 564.400 377.000 565.200 377.800 ;
        RECT 553.000 375.400 553.800 375.600 ;
        RECT 550.000 374.800 553.800 375.400 ;
        RECT 545.000 373.800 546.000 374.200 ;
        RECT 516.600 371.000 517.200 373.000 ;
        RECT 518.000 371.600 518.800 373.200 ;
        RECT 519.600 371.600 520.400 373.200 ;
        RECT 522.800 371.600 523.600 373.200 ;
        RECT 524.200 372.300 524.800 373.600 ;
        RECT 524.200 371.700 528.300 372.300 ;
        RECT 516.600 370.400 520.400 371.000 ;
        RECT 506.000 368.400 506.600 369.600 ;
        RECT 506.000 367.600 506.800 368.400 ;
        RECT 507.400 362.200 508.200 369.600 ;
        RECT 514.600 369.200 516.200 369.800 ;
        RECT 515.400 362.200 516.200 369.200 ;
        RECT 519.800 367.000 520.400 370.400 ;
        RECT 524.200 370.200 524.800 371.700 ;
        RECT 527.700 370.400 528.300 371.700 ;
        RECT 526.000 370.200 526.800 370.400 ;
        RECT 519.600 363.000 520.400 367.000 ;
        RECT 523.800 369.600 524.800 370.200 ;
        RECT 525.400 369.600 526.800 370.200 ;
        RECT 527.600 370.200 528.400 370.400 ;
        RECT 529.600 370.200 530.200 373.600 ;
        RECT 530.800 371.600 531.600 373.200 ;
        RECT 535.600 371.600 537.200 372.400 ;
        RECT 527.600 369.600 529.000 370.200 ;
        RECT 529.600 369.600 530.600 370.200 ;
        RECT 534.000 369.600 534.800 371.200 ;
        RECT 538.800 370.400 539.400 373.600 ;
        RECT 540.400 372.300 541.200 372.400 ;
        RECT 542.000 372.300 542.800 372.400 ;
        RECT 540.400 371.700 542.800 372.300 ;
        RECT 540.400 371.600 541.200 371.700 ;
        RECT 542.000 370.800 542.800 371.700 ;
        RECT 538.800 369.600 539.600 370.400 ;
        RECT 543.400 369.800 544.000 373.600 ;
        RECT 544.600 373.000 546.000 373.800 ;
        RECT 545.400 371.000 546.000 373.000 ;
        RECT 546.800 371.600 547.600 373.200 ;
        RECT 548.400 371.600 549.200 373.200 ;
        RECT 550.000 371.400 550.800 374.800 ;
        RECT 557.000 374.200 557.800 374.400 ;
        RECT 562.800 374.200 563.400 376.400 ;
        RECT 567.600 375.000 568.400 379.800 ;
        RECT 571.800 378.300 572.600 379.800 ;
        RECT 577.200 378.300 578.000 378.400 ;
        RECT 571.800 377.700 578.000 378.300 ;
        RECT 571.800 376.400 572.600 377.700 ;
        RECT 577.200 377.600 578.000 377.700 ;
        RECT 570.800 375.800 572.600 376.400 ;
        RECT 578.800 376.000 579.600 379.800 ;
        RECT 582.000 376.000 582.800 379.800 ;
        RECT 578.800 375.800 582.800 376.000 ;
        RECT 583.600 375.800 584.400 379.800 ;
        RECT 585.200 375.800 586.000 379.800 ;
        RECT 586.800 376.000 587.600 379.800 ;
        RECT 590.000 376.000 590.800 379.800 ;
        RECT 593.200 376.400 594.000 379.800 ;
        RECT 586.800 375.800 590.800 376.000 ;
        RECT 593.000 375.800 594.000 376.400 ;
        RECT 566.000 374.200 567.600 374.400 ;
        RECT 556.600 373.600 567.600 374.200 ;
        RECT 569.200 373.600 570.000 375.200 ;
        RECT 554.800 372.800 555.600 373.000 ;
        RECT 551.800 372.200 555.600 372.800 ;
        RECT 556.600 372.400 557.200 373.600 ;
        RECT 563.800 373.400 564.600 373.600 ;
        RECT 562.800 372.400 563.600 372.600 ;
        RECT 565.400 372.400 566.200 372.600 ;
        RECT 551.800 372.000 552.600 372.200 ;
        RECT 556.400 371.600 557.200 372.400 ;
        RECT 561.200 371.800 566.200 372.400 ;
        RECT 561.200 371.600 562.000 371.800 ;
        RECT 553.400 371.400 554.200 371.600 ;
        RECT 545.400 370.400 549.200 371.000 ;
        RECT 523.800 362.200 524.600 369.600 ;
        RECT 525.400 368.400 526.000 369.600 ;
        RECT 525.200 367.600 526.000 368.400 ;
        RECT 528.400 368.400 529.000 369.600 ;
        RECT 528.400 367.600 529.200 368.400 ;
        RECT 529.800 362.200 530.600 369.600 ;
        RECT 537.200 367.600 538.000 369.200 ;
        RECT 538.800 367.000 539.400 369.600 ;
        RECT 543.400 369.200 545.000 369.800 ;
        RECT 535.800 366.400 539.400 367.000 ;
        RECT 535.800 366.200 536.400 366.400 ;
        RECT 535.600 362.200 536.400 366.200 ;
        RECT 538.800 366.200 539.400 366.400 ;
        RECT 538.800 362.200 539.600 366.200 ;
        RECT 544.200 362.200 545.000 369.200 ;
        RECT 548.600 367.000 549.200 370.400 ;
        RECT 548.400 363.000 549.200 367.000 ;
        RECT 550.000 370.800 554.200 371.400 ;
        RECT 550.000 362.200 550.800 370.800 ;
        RECT 556.600 370.400 557.200 371.600 ;
        RECT 562.800 371.000 568.400 371.200 ;
        RECT 562.600 370.800 568.400 371.000 ;
        RECT 554.800 369.800 557.200 370.400 ;
        RECT 558.600 370.600 568.400 370.800 ;
        RECT 558.600 370.200 563.400 370.600 ;
        RECT 554.800 368.800 555.400 369.800 ;
        RECT 554.000 368.000 555.400 368.800 ;
        RECT 557.000 369.000 557.800 369.200 ;
        RECT 558.600 369.000 559.200 370.200 ;
        RECT 557.000 368.400 559.200 369.000 ;
        RECT 559.800 369.000 565.200 369.600 ;
        RECT 559.800 368.800 560.600 369.000 ;
        RECT 564.400 368.800 565.200 369.000 ;
        RECT 558.200 367.400 559.000 367.600 ;
        RECT 561.000 367.400 561.800 367.600 ;
        RECT 554.800 366.200 555.600 367.000 ;
        RECT 558.200 366.800 561.800 367.400 ;
        RECT 559.000 366.200 559.600 366.800 ;
        RECT 564.400 366.200 565.200 367.000 ;
        RECT 554.200 362.200 555.400 366.200 ;
        RECT 558.800 362.200 559.600 366.200 ;
        RECT 563.200 365.600 565.200 366.200 ;
        RECT 563.200 362.200 564.000 365.600 ;
        RECT 567.600 362.200 568.400 370.600 ;
        RECT 570.800 362.200 571.600 375.800 ;
        RECT 579.000 375.400 582.600 375.800 ;
        RECT 579.600 374.400 580.400 374.800 ;
        RECT 583.600 374.400 584.200 375.800 ;
        RECT 585.400 374.400 586.000 375.800 ;
        RECT 587.000 375.400 590.600 375.800 ;
        RECT 589.200 374.400 590.000 374.800 ;
        RECT 593.000 374.400 593.600 375.800 ;
        RECT 596.400 375.200 597.200 379.800 ;
        RECT 599.600 376.400 600.400 379.800 ;
        RECT 594.600 374.600 597.200 375.200 ;
        RECT 599.400 375.600 600.400 376.400 ;
        RECT 578.800 373.800 580.400 374.400 ;
        RECT 578.800 373.600 579.600 373.800 ;
        RECT 581.800 373.600 584.400 374.400 ;
        RECT 585.200 373.600 587.800 374.400 ;
        RECT 589.200 373.800 590.800 374.400 ;
        RECT 590.000 373.600 590.800 373.800 ;
        RECT 591.600 374.300 592.400 374.400 ;
        RECT 593.000 374.300 594.000 374.400 ;
        RECT 591.600 373.700 594.000 374.300 ;
        RECT 591.600 373.600 592.400 373.700 ;
        RECT 593.000 373.600 594.000 373.700 ;
        RECT 577.200 372.300 578.000 372.400 ;
        RECT 580.400 372.300 581.200 373.200 ;
        RECT 577.200 371.700 581.200 372.300 ;
        RECT 577.200 371.600 578.000 371.700 ;
        RECT 580.400 371.600 581.200 371.700 ;
        RECT 572.400 368.800 573.200 370.400 ;
        RECT 581.800 370.200 582.400 373.600 ;
        RECT 587.200 372.300 587.800 373.600 ;
        RECT 583.700 371.700 587.800 372.300 ;
        RECT 583.700 370.400 584.300 371.700 ;
        RECT 583.600 370.200 584.400 370.400 ;
        RECT 581.400 369.600 582.400 370.200 ;
        RECT 583.000 369.600 584.400 370.200 ;
        RECT 585.200 370.200 586.000 370.400 ;
        RECT 587.200 370.200 587.800 371.700 ;
        RECT 588.400 371.600 589.200 373.200 ;
        RECT 593.000 370.200 593.600 373.600 ;
        RECT 594.600 373.000 595.200 374.600 ;
        RECT 599.400 374.400 600.000 375.600 ;
        RECT 602.800 375.200 603.600 379.800 ;
        RECT 601.000 374.600 603.600 375.200 ;
        RECT 599.400 373.600 600.400 374.400 ;
        RECT 594.200 372.200 595.200 373.000 ;
        RECT 594.600 370.200 595.200 372.200 ;
        RECT 596.200 372.400 597.000 373.200 ;
        RECT 596.200 372.300 597.200 372.400 ;
        RECT 598.000 372.300 598.800 372.400 ;
        RECT 596.200 371.700 598.800 372.300 ;
        RECT 596.200 371.600 597.200 371.700 ;
        RECT 598.000 371.600 598.800 371.700 ;
        RECT 599.400 370.200 600.000 373.600 ;
        RECT 601.000 373.000 601.600 374.600 ;
        RECT 600.600 372.200 601.600 373.000 ;
        RECT 601.000 370.200 601.600 372.200 ;
        RECT 602.600 372.400 603.400 373.200 ;
        RECT 602.600 371.600 603.600 372.400 ;
        RECT 585.200 369.600 586.600 370.200 ;
        RECT 587.200 369.600 588.200 370.200 ;
        RECT 581.400 362.200 582.200 369.600 ;
        RECT 583.000 368.400 583.600 369.600 ;
        RECT 582.800 367.600 583.600 368.400 ;
        RECT 586.000 368.400 586.600 369.600 ;
        RECT 586.000 367.600 586.800 368.400 ;
        RECT 587.400 362.200 588.200 369.600 ;
        RECT 593.000 369.200 594.000 370.200 ;
        RECT 594.600 369.600 597.200 370.200 ;
        RECT 593.200 362.200 594.000 369.200 ;
        RECT 596.400 362.200 597.200 369.600 ;
        RECT 599.400 369.200 600.400 370.200 ;
        RECT 601.000 369.600 603.600 370.200 ;
        RECT 599.600 362.200 600.400 369.200 ;
        RECT 602.800 362.200 603.600 369.600 ;
        RECT 604.400 362.200 605.200 379.800 ;
        RECT 609.200 377.800 610.000 379.800 ;
        RECT 606.000 375.600 606.800 377.200 ;
        RECT 609.200 374.400 609.800 377.800 ;
        RECT 610.800 376.300 611.600 377.200 ;
        RECT 612.400 376.300 613.200 377.200 ;
        RECT 610.800 375.700 613.200 376.300 ;
        RECT 610.800 375.600 611.600 375.700 ;
        RECT 612.400 375.600 613.200 375.700 ;
        RECT 609.200 373.600 610.000 374.400 ;
        RECT 607.600 370.800 608.400 372.400 ;
        RECT 609.200 370.400 609.800 373.600 ;
        RECT 609.200 370.200 610.000 370.400 ;
        RECT 608.200 369.400 610.000 370.200 ;
        RECT 614.000 370.300 614.800 379.800 ;
        RECT 616.200 378.400 617.000 379.800 ;
        RECT 615.600 377.600 617.000 378.400 ;
        RECT 616.200 376.400 617.000 377.600 ;
        RECT 616.200 375.800 618.000 376.400 ;
        RECT 620.400 376.000 621.200 379.800 ;
        RECT 623.600 376.000 624.400 379.800 ;
        RECT 620.400 375.800 624.400 376.000 ;
        RECT 625.200 375.800 626.000 379.800 ;
        RECT 626.800 377.000 627.600 379.000 ;
        RECT 615.600 370.300 616.400 370.400 ;
        RECT 614.000 369.700 616.400 370.300 ;
        RECT 608.200 362.200 609.000 369.400 ;
        RECT 614.000 362.200 614.800 369.700 ;
        RECT 615.600 368.800 616.400 369.700 ;
        RECT 617.200 362.200 618.000 375.800 ;
        RECT 620.600 375.400 624.200 375.800 ;
        RECT 618.800 373.600 619.600 375.200 ;
        RECT 621.200 374.400 622.000 374.800 ;
        RECT 625.200 374.400 625.800 375.800 ;
        RECT 626.800 374.800 627.400 377.000 ;
        RECT 631.000 376.000 631.800 379.000 ;
        RECT 631.000 375.400 632.600 376.000 ;
        RECT 636.400 375.800 637.200 379.800 ;
        RECT 638.000 376.000 638.800 379.800 ;
        RECT 641.200 376.000 642.000 379.800 ;
        RECT 645.400 376.400 646.200 379.800 ;
        RECT 649.200 377.800 650.000 379.800 ;
        RECT 638.000 375.800 642.000 376.000 ;
        RECT 644.400 375.800 646.200 376.400 ;
        RECT 631.800 375.000 632.600 375.400 ;
        RECT 620.400 373.800 622.000 374.400 ;
        RECT 620.400 373.600 621.200 373.800 ;
        RECT 623.400 373.600 626.000 374.400 ;
        RECT 626.800 374.200 631.000 374.800 ;
        RECT 630.000 373.800 631.000 374.200 ;
        RECT 632.000 374.400 632.600 375.000 ;
        RECT 636.600 374.400 637.200 375.800 ;
        RECT 638.200 375.400 641.800 375.800 ;
        RECT 640.400 374.400 641.200 374.800 ;
        RECT 632.000 374.300 634.000 374.400 ;
        RECT 634.800 374.300 635.600 374.400 ;
        RECT 620.400 372.300 621.200 372.400 ;
        RECT 622.000 372.300 622.800 373.200 ;
        RECT 620.400 371.700 622.800 372.300 ;
        RECT 620.400 371.600 621.200 371.700 ;
        RECT 622.000 371.600 622.800 371.700 ;
        RECT 623.400 370.200 624.000 373.600 ;
        RECT 626.800 371.600 627.600 373.200 ;
        RECT 628.400 371.600 629.200 373.200 ;
        RECT 630.000 373.000 631.400 373.800 ;
        RECT 632.000 373.700 635.600 374.300 ;
        RECT 632.000 373.600 634.000 373.700 ;
        RECT 634.800 373.600 635.600 373.700 ;
        RECT 636.400 373.600 639.000 374.400 ;
        RECT 640.400 373.800 642.000 374.400 ;
        RECT 641.200 373.600 642.000 373.800 ;
        RECT 642.800 373.600 643.600 375.200 ;
        RECT 630.000 371.000 630.600 373.000 ;
        RECT 626.800 370.400 630.600 371.000 ;
        RECT 625.200 370.200 626.000 370.400 ;
        RECT 623.000 369.600 624.000 370.200 ;
        RECT 624.600 369.600 626.000 370.200 ;
        RECT 623.000 368.400 623.800 369.600 ;
        RECT 624.600 368.400 625.200 369.600 ;
        RECT 622.000 367.600 623.800 368.400 ;
        RECT 624.400 367.600 625.200 368.400 ;
        RECT 623.000 362.200 623.800 367.600 ;
        RECT 626.800 367.000 627.400 370.400 ;
        RECT 632.000 369.800 632.600 373.600 ;
        RECT 633.200 370.800 634.000 372.400 ;
        RECT 631.000 369.200 632.600 369.800 ;
        RECT 636.400 370.200 637.200 370.400 ;
        RECT 638.400 370.200 639.000 373.600 ;
        RECT 639.600 371.600 640.400 373.200 ;
        RECT 636.400 369.600 637.800 370.200 ;
        RECT 638.400 369.600 639.400 370.200 ;
        RECT 626.800 363.000 627.600 367.000 ;
        RECT 631.000 362.200 631.800 369.200 ;
        RECT 637.200 368.400 637.800 369.600 ;
        RECT 637.200 367.600 638.000 368.400 ;
        RECT 638.600 362.200 639.400 369.600 ;
        RECT 644.400 362.200 645.200 375.800 ;
        RECT 647.600 375.600 648.400 377.200 ;
        RECT 649.400 374.400 650.000 377.800 ;
        RECT 654.000 376.000 654.800 379.800 ;
        RECT 649.200 373.600 650.000 374.400 ;
        RECT 646.000 368.800 646.800 370.400 ;
        RECT 649.400 370.200 650.000 373.600 ;
        RECT 653.800 375.200 654.800 376.000 ;
        RECT 650.800 370.800 651.600 372.400 ;
        RECT 653.800 370.800 654.600 375.200 ;
        RECT 655.600 374.600 656.400 379.800 ;
        RECT 662.000 376.600 662.800 379.800 ;
        RECT 663.600 377.000 664.400 379.800 ;
        RECT 665.200 377.000 666.000 379.800 ;
        RECT 666.800 377.000 667.600 379.800 ;
        RECT 668.400 377.000 669.200 379.800 ;
        RECT 671.600 377.000 672.400 379.800 ;
        RECT 674.800 377.000 675.600 379.800 ;
        RECT 676.400 377.000 677.200 379.800 ;
        RECT 678.000 377.000 678.800 379.800 ;
        RECT 660.400 375.800 662.800 376.600 ;
        RECT 679.600 376.600 680.400 379.800 ;
        RECT 660.400 375.200 661.200 375.800 ;
        RECT 655.200 374.000 656.400 374.600 ;
        RECT 659.400 374.600 661.200 375.200 ;
        RECT 665.200 375.600 666.200 376.400 ;
        RECT 669.200 375.600 670.800 376.400 ;
        RECT 671.600 375.800 676.200 376.400 ;
        RECT 679.600 375.800 682.200 376.600 ;
        RECT 671.600 375.600 672.400 375.800 ;
        RECT 655.200 372.000 655.800 374.000 ;
        RECT 659.400 373.400 660.200 374.600 ;
        RECT 656.400 372.600 660.200 373.400 ;
        RECT 665.200 372.800 666.000 375.600 ;
        RECT 671.600 374.800 672.400 375.000 ;
        RECT 668.000 374.200 672.400 374.800 ;
        RECT 668.000 374.000 668.800 374.200 ;
        RECT 673.200 373.600 674.000 375.200 ;
        RECT 675.400 373.400 676.200 375.800 ;
        RECT 681.400 375.200 682.200 375.800 ;
        RECT 681.400 374.400 684.400 375.200 ;
        RECT 686.000 373.800 686.800 379.800 ;
        RECT 668.400 372.600 671.600 373.400 ;
        RECT 675.400 372.600 677.400 373.400 ;
        RECT 678.000 373.000 686.800 373.800 ;
        RECT 662.000 372.000 662.800 372.600 ;
        RECT 679.600 372.000 680.400 372.400 ;
        RECT 681.200 372.000 682.000 372.400 ;
        RECT 684.600 372.000 685.400 372.200 ;
        RECT 655.200 371.400 656.000 372.000 ;
        RECT 662.000 371.400 685.400 372.000 ;
        RECT 649.200 369.400 651.000 370.200 ;
        RECT 653.800 370.000 654.800 370.800 ;
        RECT 650.200 364.400 651.000 369.400 ;
        RECT 650.200 363.600 651.600 364.400 ;
        RECT 650.200 362.200 651.000 363.600 ;
        RECT 654.000 362.200 654.800 370.000 ;
        RECT 655.400 369.600 656.000 371.400 ;
        RECT 655.400 369.000 664.400 369.600 ;
        RECT 655.400 367.400 656.000 369.000 ;
        RECT 663.600 368.800 664.400 369.000 ;
        RECT 666.800 369.000 675.400 369.600 ;
        RECT 666.800 368.800 667.600 369.000 ;
        RECT 658.600 367.600 661.200 368.400 ;
        RECT 655.400 366.800 658.000 367.400 ;
        RECT 657.200 362.200 658.000 366.800 ;
        RECT 660.400 362.200 661.200 367.600 ;
        RECT 661.800 366.800 666.000 367.600 ;
        RECT 663.600 362.200 664.400 365.000 ;
        RECT 665.200 362.200 666.000 365.000 ;
        RECT 666.800 362.200 667.600 365.000 ;
        RECT 668.400 362.200 669.200 368.400 ;
        RECT 671.600 367.600 674.200 368.400 ;
        RECT 674.800 368.200 675.400 369.000 ;
        RECT 676.400 369.400 677.200 369.600 ;
        RECT 676.400 369.000 681.800 369.400 ;
        RECT 676.400 368.800 682.600 369.000 ;
        RECT 681.200 368.200 682.600 368.800 ;
        RECT 674.800 367.600 680.600 368.200 ;
        RECT 683.600 368.000 685.200 368.800 ;
        RECT 683.600 367.600 684.200 368.000 ;
        RECT 671.600 362.200 672.400 367.000 ;
        RECT 674.800 362.200 675.600 367.000 ;
        RECT 680.000 366.800 684.200 367.600 ;
        RECT 686.000 367.400 686.800 373.000 ;
        RECT 684.800 366.800 686.800 367.400 ;
        RECT 676.400 362.200 677.200 365.000 ;
        RECT 678.000 362.200 678.800 365.000 ;
        RECT 681.200 362.200 682.000 366.800 ;
        RECT 684.800 366.200 685.400 366.800 ;
        RECT 684.400 365.600 685.400 366.200 ;
        RECT 684.400 362.200 685.200 365.600 ;
        RECT 1.200 351.400 2.000 359.800 ;
        RECT 5.600 356.400 6.400 359.800 ;
        RECT 4.400 355.800 6.400 356.400 ;
        RECT 10.000 355.800 10.800 359.800 ;
        RECT 14.200 355.800 15.400 359.800 ;
        RECT 4.400 355.000 5.200 355.800 ;
        RECT 10.000 355.200 10.600 355.800 ;
        RECT 7.800 354.600 11.400 355.200 ;
        RECT 14.000 355.000 14.800 355.800 ;
        RECT 7.800 354.400 8.600 354.600 ;
        RECT 10.600 354.400 11.400 354.600 ;
        RECT 4.400 353.000 5.200 353.200 ;
        RECT 9.000 353.000 9.800 353.200 ;
        RECT 4.400 352.400 9.800 353.000 ;
        RECT 10.400 353.000 12.600 353.600 ;
        RECT 10.400 351.800 11.000 353.000 ;
        RECT 11.800 352.800 12.600 353.000 ;
        RECT 14.200 353.200 15.600 354.000 ;
        RECT 14.200 352.200 14.800 353.200 ;
        RECT 6.200 351.400 11.000 351.800 ;
        RECT 1.200 351.200 11.000 351.400 ;
        RECT 12.400 351.600 14.800 352.200 ;
        RECT 18.800 352.300 19.600 359.800 ;
        RECT 21.200 353.600 22.000 354.400 ;
        RECT 21.200 352.400 21.800 353.600 ;
        RECT 22.600 352.400 23.400 359.800 ;
        RECT 27.600 353.600 28.400 354.400 ;
        RECT 27.600 352.400 28.200 353.600 ;
        RECT 29.000 352.400 29.800 359.800 ;
        RECT 20.400 352.300 21.800 352.400 ;
        RECT 18.800 351.800 21.800 352.300 ;
        RECT 18.800 351.700 21.200 351.800 ;
        RECT 1.200 351.000 7.000 351.200 ;
        RECT 1.200 350.800 6.800 351.000 ;
        RECT 12.400 350.400 13.000 351.600 ;
        RECT 18.800 351.200 19.600 351.700 ;
        RECT 20.400 351.600 21.200 351.700 ;
        RECT 22.400 351.600 24.400 352.400 ;
        RECT 26.800 351.800 28.200 352.400 ;
        RECT 28.800 351.800 29.800 352.400 ;
        RECT 35.800 352.400 36.600 359.800 ;
        RECT 37.200 353.600 38.000 354.400 ;
        RECT 37.400 352.400 38.000 353.600 ;
        RECT 40.400 353.600 41.200 354.400 ;
        RECT 40.400 352.400 41.000 353.600 ;
        RECT 41.800 352.400 42.600 359.800 ;
        RECT 49.800 352.800 50.600 359.800 ;
        RECT 54.000 355.000 54.800 359.000 ;
        RECT 35.800 351.800 36.800 352.400 ;
        RECT 37.400 351.800 38.800 352.400 ;
        RECT 26.800 351.600 27.600 351.800 ;
        RECT 15.400 350.600 19.600 351.200 ;
        RECT 15.400 350.400 16.200 350.600 ;
        RECT 7.600 350.200 8.400 350.400 ;
        RECT 3.400 349.600 8.400 350.200 ;
        RECT 12.400 349.600 13.200 350.400 ;
        RECT 17.000 349.800 17.800 350.000 ;
        RECT 3.400 349.400 4.200 349.600 ;
        RECT 5.000 348.400 5.800 348.600 ;
        RECT 12.400 348.400 13.000 349.600 ;
        RECT 14.000 349.200 17.800 349.800 ;
        RECT 14.000 349.000 14.800 349.200 ;
        RECT 2.000 347.800 13.000 348.400 ;
        RECT 2.000 347.600 3.600 347.800 ;
        RECT 1.200 342.200 2.000 347.000 ;
        RECT 6.200 345.600 6.800 347.800 ;
        RECT 11.800 347.600 12.600 347.800 ;
        RECT 18.800 347.200 19.600 350.600 ;
        RECT 22.400 348.400 23.000 351.600 ;
        RECT 23.600 348.800 24.400 350.400 ;
        RECT 28.800 348.400 29.400 351.800 ;
        RECT 30.000 348.800 30.800 350.400 ;
        RECT 34.800 348.800 35.600 350.400 ;
        RECT 36.200 350.300 36.800 351.800 ;
        RECT 38.000 351.600 38.800 351.800 ;
        RECT 39.600 351.800 41.000 352.400 ;
        RECT 41.600 351.800 42.600 352.400 ;
        RECT 49.000 352.200 50.600 352.800 ;
        RECT 39.600 351.600 40.400 351.800 ;
        RECT 39.700 350.300 40.300 351.600 ;
        RECT 36.200 349.700 40.300 350.300 ;
        RECT 36.200 348.400 36.800 349.700 ;
        RECT 41.600 348.400 42.200 351.800 ;
        RECT 42.800 348.800 43.600 350.400 ;
        RECT 46.000 350.300 46.800 350.400 ;
        RECT 47.600 350.300 48.400 351.200 ;
        RECT 46.000 349.700 48.400 350.300 ;
        RECT 46.000 349.600 46.800 349.700 ;
        RECT 47.600 349.600 48.400 349.700 ;
        RECT 49.000 348.400 49.600 352.200 ;
        RECT 54.200 351.600 54.800 355.000 ;
        RECT 51.000 351.000 54.800 351.600 ;
        RECT 51.000 349.000 51.600 351.000 ;
        RECT 20.400 347.600 23.000 348.400 ;
        RECT 25.200 348.200 26.000 348.400 ;
        RECT 24.400 347.600 26.000 348.200 ;
        RECT 26.800 347.600 29.400 348.400 ;
        RECT 31.600 348.200 32.400 348.400 ;
        RECT 30.800 347.600 32.400 348.200 ;
        RECT 33.200 348.200 34.000 348.400 ;
        RECT 33.200 347.600 34.800 348.200 ;
        RECT 36.200 347.600 38.800 348.400 ;
        RECT 39.600 347.600 42.200 348.400 ;
        RECT 44.400 348.200 45.200 348.400 ;
        RECT 43.600 347.600 45.200 348.200 ;
        RECT 47.600 347.600 49.600 348.400 ;
        RECT 50.200 348.200 51.600 349.000 ;
        RECT 52.400 348.800 53.200 350.400 ;
        RECT 54.000 348.800 54.800 350.400 ;
        RECT 15.800 346.600 19.600 347.200 ;
        RECT 15.800 346.400 16.600 346.600 ;
        RECT 4.400 344.200 5.200 345.000 ;
        RECT 6.000 344.800 6.800 345.600 ;
        RECT 7.800 345.400 8.600 345.600 ;
        RECT 7.800 344.800 10.600 345.400 ;
        RECT 10.000 344.200 10.600 344.800 ;
        RECT 14.000 344.200 14.800 345.000 ;
        RECT 4.400 343.600 6.400 344.200 ;
        RECT 5.600 342.200 6.400 343.600 ;
        RECT 10.000 342.200 10.800 344.200 ;
        RECT 14.000 343.600 15.400 344.200 ;
        RECT 14.200 342.200 15.400 343.600 ;
        RECT 18.800 342.200 19.600 346.600 ;
        RECT 20.600 346.200 21.200 347.600 ;
        RECT 24.400 347.200 25.200 347.600 ;
        RECT 22.200 346.200 25.800 346.600 ;
        RECT 27.000 346.200 27.600 347.600 ;
        RECT 30.800 347.200 31.600 347.600 ;
        RECT 34.000 347.200 34.800 347.600 ;
        RECT 28.600 346.200 32.200 346.600 ;
        RECT 33.400 346.200 37.000 346.600 ;
        RECT 38.000 346.200 38.600 347.600 ;
        RECT 39.800 346.200 40.400 347.600 ;
        RECT 43.600 347.200 44.400 347.600 ;
        RECT 49.000 347.000 49.600 347.600 ;
        RECT 50.600 347.800 51.600 348.200 ;
        RECT 50.600 347.200 54.800 347.800 ;
        RECT 49.000 346.600 49.800 347.000 ;
        RECT 41.400 346.200 45.000 346.600 ;
        RECT 20.400 342.200 21.200 346.200 ;
        RECT 22.000 346.000 26.000 346.200 ;
        RECT 22.000 342.200 22.800 346.000 ;
        RECT 25.200 342.200 26.000 346.000 ;
        RECT 26.800 342.200 27.600 346.200 ;
        RECT 28.400 346.000 32.400 346.200 ;
        RECT 28.400 342.200 29.200 346.000 ;
        RECT 31.600 342.200 32.400 346.000 ;
        RECT 33.200 346.000 37.200 346.200 ;
        RECT 33.200 342.200 34.000 346.000 ;
        RECT 36.400 342.200 37.200 346.000 ;
        RECT 38.000 342.200 38.800 346.200 ;
        RECT 39.600 342.200 40.400 346.200 ;
        RECT 41.200 346.000 45.200 346.200 ;
        RECT 49.000 346.000 50.600 346.600 ;
        RECT 41.200 342.200 42.000 346.000 ;
        RECT 44.400 342.200 45.200 346.000 ;
        RECT 49.800 343.000 50.600 346.000 ;
        RECT 54.200 345.000 54.800 347.200 ;
        RECT 55.600 346.800 56.400 348.400 ;
        RECT 57.200 346.200 58.000 359.800 ;
        RECT 58.800 351.600 59.600 353.200 ;
        RECT 64.200 352.800 65.000 359.800 ;
        RECT 68.400 355.000 69.200 359.000 ;
        RECT 63.400 352.200 65.000 352.800 ;
        RECT 62.000 349.600 62.800 351.200 ;
        RECT 63.400 350.400 64.000 352.200 ;
        RECT 68.600 351.600 69.200 355.000 ;
        RECT 70.800 353.600 71.600 354.400 ;
        RECT 70.800 352.400 71.400 353.600 ;
        RECT 72.200 352.400 73.000 359.800 ;
        RECT 70.000 351.800 71.400 352.400 ;
        RECT 72.000 351.800 73.000 352.400 ;
        RECT 79.000 352.400 79.800 359.800 ;
        RECT 80.400 353.600 81.200 354.400 ;
        RECT 80.600 352.400 81.200 353.600 ;
        RECT 83.600 353.600 84.400 354.400 ;
        RECT 83.600 352.400 84.200 353.600 ;
        RECT 85.000 352.400 85.800 359.800 ;
        RECT 91.400 358.400 92.200 359.800 ;
        RECT 91.400 357.600 93.200 358.400 ;
        RECT 90.000 353.600 90.800 354.400 ;
        RECT 90.000 352.400 90.600 353.600 ;
        RECT 91.400 352.400 92.200 357.600 ;
        RECT 97.200 352.800 98.000 359.800 ;
        RECT 79.000 351.800 80.000 352.400 ;
        RECT 80.600 351.800 82.000 352.400 ;
        RECT 70.000 351.600 70.800 351.800 ;
        RECT 65.400 351.000 69.200 351.600 ;
        RECT 63.400 349.600 64.400 350.400 ;
        RECT 63.400 348.400 64.000 349.600 ;
        RECT 65.400 349.000 66.000 351.000 ;
        RECT 62.000 347.600 64.000 348.400 ;
        RECT 64.600 348.200 66.000 349.000 ;
        RECT 66.800 348.800 67.600 350.400 ;
        RECT 68.400 348.800 69.200 350.400 ;
        RECT 72.000 348.400 72.600 351.800 ;
        RECT 73.200 348.800 74.000 350.400 ;
        RECT 78.000 348.800 78.800 350.400 ;
        RECT 79.400 348.400 80.000 351.800 ;
        RECT 81.200 351.600 82.000 351.800 ;
        RECT 82.800 351.800 84.200 352.400 ;
        RECT 84.800 351.800 85.800 352.400 ;
        RECT 89.200 351.800 90.600 352.400 ;
        RECT 91.200 351.800 92.200 352.400 ;
        RECT 97.000 351.800 98.000 352.800 ;
        RECT 100.400 352.400 101.200 359.800 ;
        RECT 98.600 351.800 101.200 352.400 ;
        RECT 104.600 352.400 105.400 359.800 ;
        RECT 115.800 354.400 116.600 359.800 ;
        RECT 119.600 355.000 120.400 359.000 ;
        RECT 106.000 353.600 106.800 354.400 ;
        RECT 114.800 353.600 116.600 354.400 ;
        RECT 117.200 353.600 118.000 354.400 ;
        RECT 106.200 352.400 106.800 353.600 ;
        RECT 115.800 352.400 116.600 353.600 ;
        RECT 117.400 352.400 118.000 353.600 ;
        RECT 104.600 351.800 105.600 352.400 ;
        RECT 106.200 351.800 107.600 352.400 ;
        RECT 115.800 351.800 116.800 352.400 ;
        RECT 117.400 351.800 118.800 352.400 ;
        RECT 82.800 351.600 83.600 351.800 ;
        RECT 81.300 350.300 81.900 351.600 ;
        RECT 84.800 350.300 85.400 351.800 ;
        RECT 89.200 351.600 90.000 351.800 ;
        RECT 81.300 349.700 85.400 350.300 ;
        RECT 84.800 348.400 85.400 349.700 ;
        RECT 86.000 348.800 86.800 350.400 ;
        RECT 91.200 348.400 91.800 351.800 ;
        RECT 92.400 348.800 93.200 350.400 ;
        RECT 97.000 348.400 97.600 351.800 ;
        RECT 98.600 349.800 99.200 351.800 ;
        RECT 98.200 349.000 99.200 349.800 ;
        RECT 63.400 347.000 64.000 347.600 ;
        RECT 65.000 347.800 66.000 348.200 ;
        RECT 65.000 347.200 69.200 347.800 ;
        RECT 70.000 347.600 72.600 348.400 ;
        RECT 74.800 348.200 75.600 348.400 ;
        RECT 74.000 347.600 75.600 348.200 ;
        RECT 76.400 348.200 77.200 348.400 ;
        RECT 76.400 347.600 78.000 348.200 ;
        RECT 79.400 347.600 82.000 348.400 ;
        RECT 82.800 347.600 85.400 348.400 ;
        RECT 87.600 348.200 88.400 348.400 ;
        RECT 86.800 347.600 88.400 348.200 ;
        RECT 89.200 347.600 91.800 348.400 ;
        RECT 94.000 348.300 94.800 348.400 ;
        RECT 95.600 348.300 96.400 348.400 ;
        RECT 94.000 348.200 96.400 348.300 ;
        RECT 93.200 347.700 96.400 348.200 ;
        RECT 93.200 347.600 94.800 347.700 ;
        RECT 95.600 347.600 96.400 347.700 ;
        RECT 97.000 347.600 98.000 348.400 ;
        RECT 63.400 346.600 64.200 347.000 ;
        RECT 57.200 345.600 59.000 346.200 ;
        RECT 63.400 346.000 65.000 346.600 ;
        RECT 54.000 343.000 54.800 345.000 ;
        RECT 58.200 342.200 59.000 345.600 ;
        RECT 64.200 343.000 65.000 346.000 ;
        RECT 68.600 345.000 69.200 347.200 ;
        RECT 70.200 346.200 70.800 347.600 ;
        RECT 74.000 347.200 74.800 347.600 ;
        RECT 77.200 347.200 78.000 347.600 ;
        RECT 71.800 346.200 75.400 346.600 ;
        RECT 76.600 346.200 80.200 346.600 ;
        RECT 81.200 346.200 81.800 347.600 ;
        RECT 83.000 346.200 83.600 347.600 ;
        RECT 86.800 347.200 87.600 347.600 ;
        RECT 84.600 346.200 88.200 346.600 ;
        RECT 89.400 346.200 90.000 347.600 ;
        RECT 93.200 347.200 94.000 347.600 ;
        RECT 91.000 346.200 94.600 346.600 ;
        RECT 97.000 346.200 97.600 347.600 ;
        RECT 98.600 347.400 99.200 349.000 ;
        RECT 100.200 349.600 101.200 350.400 ;
        RECT 100.200 348.800 101.000 349.600 ;
        RECT 103.600 348.800 104.400 350.400 ;
        RECT 105.000 348.400 105.600 351.800 ;
        RECT 106.800 351.600 107.600 351.800 ;
        RECT 114.800 348.800 115.600 350.400 ;
        RECT 116.200 348.400 116.800 351.800 ;
        RECT 118.000 351.600 118.800 351.800 ;
        RECT 119.600 351.600 120.200 355.000 ;
        RECT 123.800 352.800 124.600 359.800 ;
        RECT 123.800 352.200 125.400 352.800 ;
        RECT 119.600 351.000 123.400 351.600 ;
        RECT 119.600 348.800 120.400 350.400 ;
        RECT 121.200 348.800 122.000 350.400 ;
        RECT 122.800 349.000 123.400 351.000 ;
        RECT 102.000 348.200 102.800 348.400 ;
        RECT 102.000 347.600 103.600 348.200 ;
        RECT 105.000 347.600 107.600 348.400 ;
        RECT 113.200 348.200 114.000 348.400 ;
        RECT 113.200 347.600 114.800 348.200 ;
        RECT 116.200 347.600 118.800 348.400 ;
        RECT 122.800 348.200 124.200 349.000 ;
        RECT 124.800 348.400 125.400 352.200 ;
        RECT 130.800 352.300 131.600 359.800 ;
        RECT 133.200 353.600 134.000 354.400 ;
        RECT 133.200 352.400 133.800 353.600 ;
        RECT 134.600 352.400 135.400 359.800 ;
        RECT 139.600 353.600 140.400 354.400 ;
        RECT 139.600 352.400 140.200 353.600 ;
        RECT 141.000 352.400 141.800 359.800 ;
        RECT 132.400 352.300 133.800 352.400 ;
        RECT 130.800 351.800 133.800 352.300 ;
        RECT 134.400 351.800 135.400 352.400 ;
        RECT 138.800 351.800 140.200 352.400 ;
        RECT 140.800 351.800 141.800 352.400 ;
        RECT 147.800 352.400 148.600 359.800 ;
        RECT 149.200 353.600 150.000 354.400 ;
        RECT 149.400 352.400 150.000 353.600 ;
        RECT 152.400 353.600 153.200 354.400 ;
        RECT 152.400 352.400 153.000 353.600 ;
        RECT 153.800 352.400 154.600 359.800 ;
        RECT 158.800 353.600 159.600 354.400 ;
        RECT 158.800 352.400 159.400 353.600 ;
        RECT 160.200 352.400 161.000 359.800 ;
        RECT 165.200 353.600 166.000 354.400 ;
        RECT 165.200 352.400 165.800 353.600 ;
        RECT 166.600 352.400 167.400 359.800 ;
        RECT 172.400 356.400 173.200 359.800 ;
        RECT 172.200 355.800 173.200 356.400 ;
        RECT 172.200 355.200 172.800 355.800 ;
        RECT 175.600 355.200 176.400 359.800 ;
        RECT 178.800 357.000 179.600 359.800 ;
        RECT 180.400 357.000 181.200 359.800 ;
        RECT 147.800 351.800 148.800 352.400 ;
        RECT 149.400 351.800 150.800 352.400 ;
        RECT 130.800 351.700 133.200 351.800 ;
        RECT 126.000 350.300 126.800 351.200 ;
        RECT 127.600 350.300 128.400 350.400 ;
        RECT 126.000 349.700 128.400 350.300 ;
        RECT 126.000 349.600 126.800 349.700 ;
        RECT 127.600 349.600 128.400 349.700 ;
        RECT 122.800 347.800 123.800 348.200 ;
        RECT 98.600 346.800 101.200 347.400 ;
        RECT 102.800 347.200 103.600 347.600 ;
        RECT 68.400 343.000 69.200 345.000 ;
        RECT 70.000 342.200 70.800 346.200 ;
        RECT 71.600 346.000 75.600 346.200 ;
        RECT 71.600 342.200 72.400 346.000 ;
        RECT 74.800 342.200 75.600 346.000 ;
        RECT 76.400 346.000 80.400 346.200 ;
        RECT 76.400 342.200 77.200 346.000 ;
        RECT 79.600 342.200 80.400 346.000 ;
        RECT 81.200 342.200 82.000 346.200 ;
        RECT 82.800 342.200 83.600 346.200 ;
        RECT 84.400 346.000 88.400 346.200 ;
        RECT 84.400 342.200 85.200 346.000 ;
        RECT 87.600 342.200 88.400 346.000 ;
        RECT 89.200 342.200 90.000 346.200 ;
        RECT 90.800 346.000 94.800 346.200 ;
        RECT 90.800 342.200 91.600 346.000 ;
        RECT 94.000 342.200 94.800 346.000 ;
        RECT 97.000 345.600 98.000 346.200 ;
        RECT 97.200 342.200 98.000 345.600 ;
        RECT 100.400 342.200 101.200 346.800 ;
        RECT 102.200 346.200 105.800 346.600 ;
        RECT 106.800 346.200 107.400 347.600 ;
        RECT 114.000 347.200 114.800 347.600 ;
        RECT 113.400 346.200 117.000 346.600 ;
        RECT 118.000 346.200 118.600 347.600 ;
        RECT 119.600 347.200 123.800 347.800 ;
        RECT 124.800 347.600 126.800 348.400 ;
        RECT 102.000 346.000 106.000 346.200 ;
        RECT 102.000 342.200 102.800 346.000 ;
        RECT 105.200 342.200 106.000 346.000 ;
        RECT 106.800 344.300 107.600 346.200 ;
        RECT 113.200 346.000 117.200 346.200 ;
        RECT 111.600 344.300 112.400 344.400 ;
        RECT 106.800 343.700 112.400 344.300 ;
        RECT 106.800 342.200 107.600 343.700 ;
        RECT 111.600 343.600 112.400 343.700 ;
        RECT 113.200 342.200 114.000 346.000 ;
        RECT 116.400 342.200 117.200 346.000 ;
        RECT 118.000 342.200 118.800 346.200 ;
        RECT 119.600 345.000 120.200 347.200 ;
        RECT 124.800 347.000 125.400 347.600 ;
        RECT 124.600 346.600 125.400 347.000 ;
        RECT 123.800 346.000 125.400 346.600 ;
        RECT 119.600 343.000 120.400 345.000 ;
        RECT 123.800 344.400 124.600 346.000 ;
        RECT 129.200 344.800 130.000 346.400 ;
        RECT 122.800 343.600 124.600 344.400 ;
        RECT 123.800 343.000 124.600 343.600 ;
        RECT 130.800 342.200 131.600 351.700 ;
        RECT 132.400 351.600 133.200 351.700 ;
        RECT 132.400 350.300 133.200 350.400 ;
        RECT 134.400 350.300 135.000 351.800 ;
        RECT 138.800 351.600 139.600 351.800 ;
        RECT 132.400 349.700 135.000 350.300 ;
        RECT 132.400 349.600 133.200 349.700 ;
        RECT 134.400 348.400 135.000 349.700 ;
        RECT 135.600 348.800 136.400 350.400 ;
        RECT 140.800 348.400 141.400 351.800 ;
        RECT 142.000 348.800 142.800 350.400 ;
        RECT 146.800 348.800 147.600 350.400 ;
        RECT 148.200 348.400 148.800 351.800 ;
        RECT 150.000 351.600 150.800 351.800 ;
        RECT 151.600 351.800 153.000 352.400 ;
        RECT 151.600 351.600 152.400 351.800 ;
        RECT 153.600 351.600 155.600 352.400 ;
        RECT 158.000 351.800 159.400 352.400 ;
        RECT 160.000 351.800 161.000 352.400 ;
        RECT 164.400 351.800 165.800 352.400 ;
        RECT 166.400 351.800 167.400 352.400 ;
        RECT 170.800 354.600 172.800 355.200 ;
        RECT 158.000 351.600 158.800 351.800 ;
        RECT 153.600 348.400 154.200 351.600 ;
        RECT 154.800 350.300 155.600 350.400 ;
        RECT 156.400 350.300 157.200 350.400 ;
        RECT 154.800 349.700 157.200 350.300 ;
        RECT 154.800 348.800 155.600 349.700 ;
        RECT 156.400 349.600 157.200 349.700 ;
        RECT 160.000 348.400 160.600 351.800 ;
        RECT 164.400 351.600 165.200 351.800 ;
        RECT 166.400 350.400 167.000 351.800 ;
        RECT 161.200 348.800 162.000 350.400 ;
        RECT 166.000 349.600 167.000 350.400 ;
        RECT 166.400 348.400 167.000 349.600 ;
        RECT 167.600 348.800 168.400 350.400 ;
        RECT 170.800 349.000 171.600 354.600 ;
        RECT 173.400 354.400 177.600 355.200 ;
        RECT 182.000 355.000 182.800 359.800 ;
        RECT 185.200 355.000 186.000 359.800 ;
        RECT 173.400 354.000 174.000 354.400 ;
        RECT 172.400 353.200 174.000 354.000 ;
        RECT 177.000 353.800 182.800 354.400 ;
        RECT 175.000 353.200 176.400 353.800 ;
        RECT 175.000 353.000 181.200 353.200 ;
        RECT 175.800 352.600 181.200 353.000 ;
        RECT 180.400 352.400 181.200 352.600 ;
        RECT 182.200 353.000 182.800 353.800 ;
        RECT 183.400 353.600 186.000 354.400 ;
        RECT 188.400 353.600 189.200 359.800 ;
        RECT 190.000 357.000 190.800 359.800 ;
        RECT 191.600 357.000 192.400 359.800 ;
        RECT 193.200 357.000 194.000 359.800 ;
        RECT 191.600 354.400 195.800 355.200 ;
        RECT 196.400 354.400 197.200 359.800 ;
        RECT 199.600 355.200 200.400 359.800 ;
        RECT 199.600 354.600 202.200 355.200 ;
        RECT 196.400 353.600 199.000 354.400 ;
        RECT 190.000 353.000 190.800 353.200 ;
        RECT 182.200 352.400 190.800 353.000 ;
        RECT 193.200 353.000 194.000 353.200 ;
        RECT 201.600 353.000 202.200 354.600 ;
        RECT 193.200 352.400 202.200 353.000 ;
        RECT 201.600 350.600 202.200 352.400 ;
        RECT 202.800 352.000 203.600 359.800 ;
        RECT 206.000 352.400 206.800 359.800 ;
        RECT 207.600 352.400 208.400 352.600 ;
        RECT 202.800 351.200 203.800 352.000 ;
        RECT 206.000 351.800 208.400 352.400 ;
        RECT 210.400 351.800 212.000 359.800 ;
        RECT 213.800 352.400 214.600 352.600 ;
        RECT 215.600 352.400 216.400 359.800 ;
        RECT 218.000 353.600 218.800 354.400 ;
        RECT 218.000 352.400 218.600 353.600 ;
        RECT 219.400 352.400 220.200 359.800 ;
        RECT 213.800 351.800 216.400 352.400 ;
        RECT 217.200 351.800 218.600 352.400 ;
        RECT 219.200 351.800 220.200 352.400 ;
        RECT 172.200 350.000 195.600 350.600 ;
        RECT 201.600 350.000 202.400 350.600 ;
        RECT 172.200 349.800 173.000 350.000 ;
        RECT 175.600 349.600 176.400 350.000 ;
        RECT 177.200 349.600 178.000 350.000 ;
        RECT 194.800 349.400 195.600 350.000 ;
        RECT 132.400 347.600 135.000 348.400 ;
        RECT 137.200 348.200 138.000 348.400 ;
        RECT 136.400 347.600 138.000 348.200 ;
        RECT 138.800 347.600 141.400 348.400 ;
        RECT 143.600 348.200 144.400 348.400 ;
        RECT 142.800 347.600 144.400 348.200 ;
        RECT 145.200 348.200 146.000 348.400 ;
        RECT 145.200 347.600 146.800 348.200 ;
        RECT 148.200 347.600 150.800 348.400 ;
        RECT 151.600 347.600 154.200 348.400 ;
        RECT 156.400 348.200 157.200 348.400 ;
        RECT 155.600 347.600 157.200 348.200 ;
        RECT 158.000 347.600 160.600 348.400 ;
        RECT 162.800 348.200 163.600 348.400 ;
        RECT 162.000 347.600 163.600 348.200 ;
        RECT 164.400 347.600 167.000 348.400 ;
        RECT 169.200 348.200 170.000 348.400 ;
        RECT 168.400 347.600 170.000 348.200 ;
        RECT 170.800 348.200 179.600 349.000 ;
        RECT 180.200 348.600 182.200 349.400 ;
        RECT 186.000 348.600 189.200 349.400 ;
        RECT 132.600 346.200 133.200 347.600 ;
        RECT 136.400 347.200 137.200 347.600 ;
        RECT 134.200 346.200 137.800 346.600 ;
        RECT 139.000 346.200 139.600 347.600 ;
        RECT 142.800 347.200 143.600 347.600 ;
        RECT 146.000 347.200 146.800 347.600 ;
        RECT 140.600 346.200 144.200 346.600 ;
        RECT 145.400 346.200 149.000 346.600 ;
        RECT 150.000 346.200 150.600 347.600 ;
        RECT 151.800 346.200 152.400 347.600 ;
        RECT 155.600 347.200 156.400 347.600 ;
        RECT 153.400 346.200 157.000 346.600 ;
        RECT 158.200 346.200 158.800 347.600 ;
        RECT 162.000 347.200 162.800 347.600 ;
        RECT 159.800 346.200 163.400 346.600 ;
        RECT 164.600 346.200 165.200 347.600 ;
        RECT 168.400 347.200 169.200 347.600 ;
        RECT 166.200 346.200 169.800 346.600 ;
        RECT 132.400 342.200 133.200 346.200 ;
        RECT 134.000 346.000 138.000 346.200 ;
        RECT 134.000 342.200 134.800 346.000 ;
        RECT 137.200 342.200 138.000 346.000 ;
        RECT 138.800 342.200 139.600 346.200 ;
        RECT 140.400 346.000 144.400 346.200 ;
        RECT 140.400 342.200 141.200 346.000 ;
        RECT 143.600 342.200 144.400 346.000 ;
        RECT 145.200 346.000 149.200 346.200 ;
        RECT 145.200 342.200 146.000 346.000 ;
        RECT 148.400 342.200 149.200 346.000 ;
        RECT 150.000 342.200 150.800 346.200 ;
        RECT 151.600 342.200 152.400 346.200 ;
        RECT 153.200 346.000 157.200 346.200 ;
        RECT 153.200 342.200 154.000 346.000 ;
        RECT 156.400 342.200 157.200 346.000 ;
        RECT 158.000 342.200 158.800 346.200 ;
        RECT 159.600 346.000 163.600 346.200 ;
        RECT 159.600 342.200 160.400 346.000 ;
        RECT 162.800 342.200 163.600 346.000 ;
        RECT 164.400 342.200 165.200 346.200 ;
        RECT 166.000 346.000 170.000 346.200 ;
        RECT 166.000 342.200 166.800 346.000 ;
        RECT 169.200 342.200 170.000 346.000 ;
        RECT 170.800 342.200 171.600 348.200 ;
        RECT 173.200 346.800 176.200 347.600 ;
        RECT 175.400 346.200 176.200 346.800 ;
        RECT 181.400 346.200 182.200 348.600 ;
        RECT 183.600 346.800 184.400 348.400 ;
        RECT 188.800 347.800 189.600 348.000 ;
        RECT 185.200 347.200 189.600 347.800 ;
        RECT 185.200 347.000 186.000 347.200 ;
        RECT 191.600 346.400 192.400 349.200 ;
        RECT 197.400 348.600 201.200 349.400 ;
        RECT 197.400 347.400 198.200 348.600 ;
        RECT 201.800 348.000 202.400 350.000 ;
        RECT 185.200 346.200 186.000 346.400 ;
        RECT 175.400 345.400 178.000 346.200 ;
        RECT 181.400 345.600 186.000 346.200 ;
        RECT 186.800 345.600 188.400 346.400 ;
        RECT 191.400 345.600 192.400 346.400 ;
        RECT 196.400 346.800 198.200 347.400 ;
        RECT 201.200 347.400 202.400 348.000 ;
        RECT 203.000 348.300 203.800 351.200 ;
        RECT 210.800 350.400 211.400 351.800 ;
        RECT 217.200 351.600 218.000 351.800 ;
        RECT 212.600 350.400 213.400 350.600 ;
        RECT 210.800 349.600 211.600 350.400 ;
        RECT 212.600 349.800 214.200 350.400 ;
        RECT 213.400 349.600 214.200 349.800 ;
        RECT 210.800 348.400 211.400 349.600 ;
        RECT 206.000 348.300 207.600 348.400 ;
        RECT 203.000 347.700 207.600 348.300 ;
        RECT 196.400 346.200 197.200 346.800 ;
        RECT 177.200 342.200 178.000 345.400 ;
        RECT 194.800 345.400 197.200 346.200 ;
        RECT 178.800 342.200 179.600 345.000 ;
        RECT 180.400 342.200 181.200 345.000 ;
        RECT 182.000 342.200 182.800 345.000 ;
        RECT 185.200 342.200 186.000 345.000 ;
        RECT 188.400 342.200 189.200 345.000 ;
        RECT 190.000 342.200 190.800 345.000 ;
        RECT 191.600 342.200 192.400 345.000 ;
        RECT 193.200 342.200 194.000 345.000 ;
        RECT 194.800 342.200 195.600 345.400 ;
        RECT 201.200 342.200 202.000 347.400 ;
        RECT 203.000 346.800 203.800 347.700 ;
        RECT 206.000 347.600 207.600 347.700 ;
        RECT 208.800 347.600 209.600 348.400 ;
        RECT 209.000 347.200 209.600 347.600 ;
        RECT 210.400 347.800 211.400 348.400 ;
        RECT 212.000 348.600 212.800 348.800 ;
        RECT 212.000 348.400 214.800 348.600 ;
        RECT 219.200 348.400 219.800 351.800 ;
        RECT 223.600 351.200 224.400 359.800 ;
        RECT 227.800 358.400 228.600 359.800 ;
        RECT 227.800 357.600 229.200 358.400 ;
        RECT 227.800 352.400 228.600 357.600 ;
        RECT 232.600 352.400 233.400 359.800 ;
        RECT 234.000 354.300 234.800 354.400 ;
        RECT 236.400 354.300 237.200 354.400 ;
        RECT 234.000 353.700 237.200 354.300 ;
        RECT 234.000 353.600 234.800 353.700 ;
        RECT 236.400 353.600 237.200 353.700 ;
        RECT 234.200 352.400 234.800 353.600 ;
        RECT 227.800 351.800 229.200 352.400 ;
        RECT 232.600 351.800 233.600 352.400 ;
        RECT 234.200 351.800 235.600 352.400 ;
        RECT 223.600 350.800 227.600 351.200 ;
        RECT 223.600 350.600 227.800 350.800 ;
        RECT 220.400 348.800 221.200 350.400 ;
        RECT 227.000 350.000 227.800 350.600 ;
        RECT 228.600 350.400 229.200 351.800 ;
        RECT 225.600 348.400 226.400 349.200 ;
        RECT 212.000 348.300 216.400 348.400 ;
        RECT 217.200 348.300 219.800 348.400 ;
        RECT 212.000 348.000 219.800 348.300 ;
        RECT 222.000 348.300 222.800 348.400 ;
        RECT 225.200 348.300 226.200 348.400 ;
        RECT 222.000 348.200 226.200 348.300 ;
        RECT 214.200 347.800 219.800 348.000 ;
        RECT 207.600 346.800 208.400 347.000 ;
        RECT 202.800 346.000 203.800 346.800 ;
        RECT 206.000 346.200 208.400 346.800 ;
        RECT 209.000 346.400 209.800 347.200 ;
        RECT 202.800 342.200 203.600 346.000 ;
        RECT 206.000 342.200 206.800 346.200 ;
        RECT 210.400 345.800 211.000 347.800 ;
        RECT 214.800 347.700 219.800 347.800 ;
        RECT 214.800 347.600 216.400 347.700 ;
        RECT 217.200 347.600 219.800 347.700 ;
        RECT 221.200 347.700 226.200 348.200 ;
        RECT 221.200 347.600 222.800 347.700 ;
        RECT 225.200 347.600 226.200 347.700 ;
        RECT 211.600 346.400 213.200 347.200 ;
        RECT 213.800 346.800 214.600 347.000 ;
        RECT 213.800 346.200 216.400 346.800 ;
        RECT 217.400 346.200 218.000 347.600 ;
        RECT 221.200 347.200 222.000 347.600 ;
        RECT 227.200 347.000 227.800 350.000 ;
        RECT 228.400 349.600 229.200 350.400 ;
        RECT 219.000 346.200 222.600 346.600 ;
        RECT 225.400 346.400 227.800 347.000 ;
        RECT 210.400 344.400 212.000 345.800 ;
        RECT 209.200 343.600 212.000 344.400 ;
        RECT 210.400 342.200 212.000 343.600 ;
        RECT 215.600 342.200 216.400 346.200 ;
        RECT 217.200 342.200 218.000 346.200 ;
        RECT 218.800 346.000 222.800 346.200 ;
        RECT 218.800 342.200 219.600 346.000 ;
        RECT 222.000 342.200 222.800 346.000 ;
        RECT 223.600 344.800 224.400 346.400 ;
        RECT 225.400 344.200 226.000 346.400 ;
        RECT 228.600 346.200 229.200 349.600 ;
        RECT 231.600 348.800 232.400 350.400 ;
        RECT 233.000 348.400 233.600 351.800 ;
        RECT 234.800 351.600 235.600 351.800 ;
        RECT 230.000 348.200 230.800 348.400 ;
        RECT 233.000 348.300 235.600 348.400 ;
        RECT 236.400 348.300 237.200 348.400 ;
        RECT 230.000 347.600 231.600 348.200 ;
        RECT 233.000 347.700 237.200 348.300 ;
        RECT 233.000 347.600 235.600 347.700 ;
        RECT 230.800 347.200 231.600 347.600 ;
        RECT 230.200 346.200 233.800 346.600 ;
        RECT 234.800 346.200 235.400 347.600 ;
        RECT 236.400 346.800 237.200 347.700 ;
        RECT 238.000 346.200 238.800 359.800 ;
        RECT 242.800 356.400 243.600 359.800 ;
        RECT 242.600 355.800 243.600 356.400 ;
        RECT 242.600 355.200 243.200 355.800 ;
        RECT 246.000 355.200 246.800 359.800 ;
        RECT 249.200 357.000 250.000 359.800 ;
        RECT 250.800 357.000 251.600 359.800 ;
        RECT 241.200 354.600 243.200 355.200 ;
        RECT 239.600 351.600 240.400 353.200 ;
        RECT 241.200 349.000 242.000 354.600 ;
        RECT 243.800 354.400 248.000 355.200 ;
        RECT 252.400 355.000 253.200 359.800 ;
        RECT 255.600 355.000 256.400 359.800 ;
        RECT 243.800 354.000 244.400 354.400 ;
        RECT 242.800 353.200 244.400 354.000 ;
        RECT 247.400 353.800 253.200 354.400 ;
        RECT 245.400 353.200 246.800 353.800 ;
        RECT 245.400 353.000 251.600 353.200 ;
        RECT 246.200 352.600 251.600 353.000 ;
        RECT 250.800 352.400 251.600 352.600 ;
        RECT 252.600 353.000 253.200 353.800 ;
        RECT 253.800 353.600 256.400 354.400 ;
        RECT 258.800 353.600 259.600 359.800 ;
        RECT 260.400 357.000 261.200 359.800 ;
        RECT 262.000 357.000 262.800 359.800 ;
        RECT 263.600 357.000 264.400 359.800 ;
        RECT 262.000 354.400 266.200 355.200 ;
        RECT 266.800 354.400 267.600 359.800 ;
        RECT 270.000 355.200 270.800 359.800 ;
        RECT 270.000 354.600 272.600 355.200 ;
        RECT 266.800 353.600 269.400 354.400 ;
        RECT 260.400 353.000 261.200 353.200 ;
        RECT 252.600 352.400 261.200 353.000 ;
        RECT 263.600 353.000 264.400 353.200 ;
        RECT 272.000 353.000 272.600 354.600 ;
        RECT 263.600 352.400 272.600 353.000 ;
        RECT 272.000 350.600 272.600 352.400 ;
        RECT 273.200 352.000 274.000 359.800 ;
        RECT 273.200 351.200 274.200 352.000 ;
        RECT 242.600 350.000 266.000 350.600 ;
        RECT 272.000 350.000 272.800 350.600 ;
        RECT 242.600 349.800 243.400 350.000 ;
        RECT 244.400 349.600 245.200 350.000 ;
        RECT 247.600 349.600 248.400 350.000 ;
        RECT 265.200 349.400 266.000 350.000 ;
        RECT 241.200 348.200 250.000 349.000 ;
        RECT 250.600 348.600 252.600 349.400 ;
        RECT 256.400 348.600 259.600 349.400 ;
        RECT 225.200 342.200 226.000 344.200 ;
        RECT 228.400 342.200 229.200 346.200 ;
        RECT 230.000 346.000 234.000 346.200 ;
        RECT 230.000 342.200 230.800 346.000 ;
        RECT 233.200 342.200 234.000 346.000 ;
        RECT 234.800 342.200 235.600 346.200 ;
        RECT 238.000 345.600 239.800 346.200 ;
        RECT 239.000 342.200 239.800 345.600 ;
        RECT 241.200 342.200 242.000 348.200 ;
        RECT 243.600 346.800 246.600 347.600 ;
        RECT 245.800 346.200 246.600 346.800 ;
        RECT 251.800 346.200 252.600 348.600 ;
        RECT 254.000 346.800 254.800 348.400 ;
        RECT 259.200 347.800 260.000 348.000 ;
        RECT 255.600 347.200 260.000 347.800 ;
        RECT 255.600 347.000 256.400 347.200 ;
        RECT 262.000 346.400 262.800 349.200 ;
        RECT 267.800 348.600 271.600 349.400 ;
        RECT 267.800 347.400 268.600 348.600 ;
        RECT 272.200 348.000 272.800 350.000 ;
        RECT 255.600 346.200 256.400 346.400 ;
        RECT 245.800 345.400 248.400 346.200 ;
        RECT 251.800 345.600 256.400 346.200 ;
        RECT 257.200 345.600 258.800 346.400 ;
        RECT 261.800 345.600 262.800 346.400 ;
        RECT 266.800 346.800 268.600 347.400 ;
        RECT 271.600 347.400 272.800 348.000 ;
        RECT 266.800 346.200 267.600 346.800 ;
        RECT 247.600 342.200 248.400 345.400 ;
        RECT 265.200 345.400 267.600 346.200 ;
        RECT 249.200 342.200 250.000 345.000 ;
        RECT 250.800 342.200 251.600 345.000 ;
        RECT 252.400 342.200 253.200 345.000 ;
        RECT 255.600 342.200 256.400 345.000 ;
        RECT 258.800 342.200 259.600 345.000 ;
        RECT 260.400 342.200 261.200 345.000 ;
        RECT 262.000 342.200 262.800 345.000 ;
        RECT 263.600 342.200 264.400 345.000 ;
        RECT 265.200 342.200 266.000 345.400 ;
        RECT 271.600 342.200 272.400 347.400 ;
        RECT 273.400 346.800 274.200 351.200 ;
        RECT 282.800 351.200 283.600 359.800 ;
        RECT 286.000 351.200 286.800 359.800 ;
        RECT 289.200 351.200 290.000 359.800 ;
        RECT 292.400 351.200 293.200 359.800 ;
        RECT 295.600 352.300 296.400 359.800 ;
        RECT 297.200 352.300 298.000 352.400 ;
        RECT 295.600 351.700 298.000 352.300 ;
        RECT 282.800 350.400 284.600 351.200 ;
        RECT 286.000 350.400 288.200 351.200 ;
        RECT 289.200 350.400 291.400 351.200 ;
        RECT 292.400 350.400 294.800 351.200 ;
        RECT 283.800 349.000 284.600 350.400 ;
        RECT 287.400 349.000 288.200 350.400 ;
        RECT 290.600 349.000 291.400 350.400 ;
        RECT 281.200 348.200 283.000 349.000 ;
        RECT 283.800 348.200 286.400 349.000 ;
        RECT 287.400 348.200 289.800 349.000 ;
        RECT 290.600 348.200 293.200 349.000 ;
        RECT 281.200 347.600 282.000 348.200 ;
        RECT 283.800 347.600 284.600 348.200 ;
        RECT 287.400 347.600 288.200 348.200 ;
        RECT 290.600 347.600 291.400 348.200 ;
        RECT 294.000 347.600 294.800 350.400 ;
        RECT 273.200 346.000 274.200 346.800 ;
        RECT 282.800 346.800 284.600 347.600 ;
        RECT 286.000 346.800 288.200 347.600 ;
        RECT 289.200 346.800 291.400 347.600 ;
        RECT 292.400 346.800 294.800 347.600 ;
        RECT 273.200 342.200 274.000 346.000 ;
        RECT 282.800 342.200 283.600 346.800 ;
        RECT 286.000 342.200 286.800 346.800 ;
        RECT 289.200 342.200 290.000 346.800 ;
        RECT 292.400 342.200 293.200 346.800 ;
        RECT 295.600 342.200 296.400 351.700 ;
        RECT 297.200 351.600 298.000 351.700 ;
        RECT 298.800 346.800 299.600 348.400 ;
        RECT 297.200 344.800 298.000 346.400 ;
        RECT 300.400 346.200 301.200 359.800 ;
        RECT 305.800 358.400 306.600 359.800 ;
        RECT 305.800 357.600 307.600 358.400 ;
        RECT 304.400 353.600 305.200 354.400 ;
        RECT 302.000 351.600 302.800 353.200 ;
        RECT 304.400 352.400 305.000 353.600 ;
        RECT 305.800 352.400 306.600 357.600 ;
        RECT 310.000 355.800 310.800 359.800 ;
        RECT 310.200 355.600 310.800 355.800 ;
        RECT 313.200 355.800 314.000 359.800 ;
        RECT 313.200 355.600 313.800 355.800 ;
        RECT 310.200 355.000 313.800 355.600 ;
        RECT 310.200 352.400 310.800 355.000 ;
        RECT 311.600 352.800 312.400 354.400 ;
        RECT 316.400 352.400 317.200 359.800 ;
        RECT 319.600 359.200 323.600 359.800 ;
        RECT 319.600 352.400 320.400 359.200 ;
        RECT 303.600 351.800 305.000 352.400 ;
        RECT 305.600 351.800 306.600 352.400 ;
        RECT 303.600 351.600 304.400 351.800 ;
        RECT 305.600 348.400 306.200 351.800 ;
        RECT 310.000 351.600 310.800 352.400 ;
        RECT 306.800 348.800 307.600 350.400 ;
        RECT 310.200 348.400 310.800 351.600 ;
        RECT 314.800 350.800 315.600 352.400 ;
        RECT 316.400 351.800 320.400 352.400 ;
        RECT 321.200 351.600 322.000 358.600 ;
        RECT 322.800 351.800 323.600 359.200 ;
        RECT 324.400 352.400 325.200 359.800 ;
        RECT 327.600 359.200 331.600 359.800 ;
        RECT 327.600 352.400 328.400 359.200 ;
        RECT 324.400 351.800 328.400 352.400 ;
        RECT 329.200 351.800 330.000 358.600 ;
        RECT 330.800 351.800 331.600 359.200 ;
        RECT 332.400 352.400 333.200 359.800 ;
        RECT 335.600 359.200 339.600 359.800 ;
        RECT 335.600 352.400 336.400 359.200 ;
        RECT 332.400 351.800 336.400 352.400 ;
        RECT 337.200 351.800 338.000 358.600 ;
        RECT 338.800 351.800 339.600 359.200 ;
        RECT 342.000 355.800 342.800 359.800 ;
        RECT 342.200 355.600 342.800 355.800 ;
        RECT 345.200 355.800 346.000 359.800 ;
        RECT 346.800 359.200 350.800 359.800 ;
        RECT 345.200 355.600 345.800 355.800 ;
        RECT 342.200 355.000 345.800 355.600 ;
        RECT 343.600 352.800 344.400 354.400 ;
        RECT 345.200 352.400 345.800 355.000 ;
        RECT 321.200 351.200 321.800 351.600 ;
        RECT 329.200 351.200 329.800 351.800 ;
        RECT 337.200 351.200 337.800 351.800 ;
        RECT 317.200 350.400 318.000 350.800 ;
        RECT 319.800 350.600 321.800 351.200 ;
        RECT 319.800 350.400 320.400 350.600 ;
        RECT 312.400 349.600 314.000 350.400 ;
        RECT 316.400 349.800 318.000 350.400 ;
        RECT 316.400 349.600 317.200 349.800 ;
        RECT 319.600 349.600 320.400 350.400 ;
        RECT 322.800 349.600 323.600 351.200 ;
        RECT 325.200 350.400 326.000 350.800 ;
        RECT 327.800 350.600 329.800 351.200 ;
        RECT 327.800 350.400 328.400 350.600 ;
        RECT 324.400 349.800 326.000 350.400 ;
        RECT 324.400 349.600 325.200 349.800 ;
        RECT 327.600 349.600 328.400 350.400 ;
        RECT 330.800 349.600 331.600 351.200 ;
        RECT 333.200 350.400 334.000 350.800 ;
        RECT 335.800 350.600 337.800 351.200 ;
        RECT 335.800 350.400 336.400 350.600 ;
        RECT 332.400 349.800 334.000 350.400 ;
        RECT 332.400 349.600 333.200 349.800 ;
        RECT 335.600 349.600 336.400 350.400 ;
        RECT 338.800 349.600 339.600 351.200 ;
        RECT 340.400 350.800 341.200 352.400 ;
        RECT 345.200 351.600 346.000 352.400 ;
        RECT 346.800 351.800 347.600 359.200 ;
        RECT 348.400 351.800 349.200 358.600 ;
        RECT 350.000 352.400 350.800 359.200 ;
        RECT 353.200 352.400 354.000 359.800 ;
        RECT 354.800 355.800 355.600 359.800 ;
        RECT 355.000 355.600 355.600 355.800 ;
        RECT 358.000 355.800 358.800 359.800 ;
        RECT 358.000 355.600 358.600 355.800 ;
        RECT 355.000 355.000 358.600 355.600 ;
        RECT 355.000 352.400 355.600 355.000 ;
        RECT 356.400 352.800 357.200 354.400 ;
        RECT 350.000 351.800 354.000 352.400 ;
        RECT 342.000 349.600 343.600 350.400 ;
        RECT 303.600 347.600 306.200 348.400 ;
        RECT 308.400 348.200 309.200 348.400 ;
        RECT 307.600 347.600 309.200 348.200 ;
        RECT 310.200 348.200 311.800 348.400 ;
        RECT 310.200 347.800 312.000 348.200 ;
        RECT 303.800 346.200 304.400 347.600 ;
        RECT 307.600 347.200 308.400 347.600 ;
        RECT 305.400 346.200 309.000 346.600 ;
        RECT 300.400 345.600 302.200 346.200 ;
        RECT 301.400 344.400 302.200 345.600 ;
        RECT 301.400 343.600 302.800 344.400 ;
        RECT 301.400 342.200 302.200 343.600 ;
        RECT 303.600 342.200 304.400 346.200 ;
        RECT 305.200 346.000 309.200 346.200 ;
        RECT 305.200 342.200 306.000 346.000 ;
        RECT 308.400 342.200 309.200 346.000 ;
        RECT 311.200 342.200 312.000 347.800 ;
        RECT 318.000 347.600 318.800 349.200 ;
        RECT 319.800 346.200 320.400 349.600 ;
        RECT 321.000 348.800 321.800 349.600 ;
        RECT 321.200 348.400 321.800 348.800 ;
        RECT 321.200 347.600 322.000 348.400 ;
        RECT 326.000 347.600 326.800 349.200 ;
        RECT 327.800 346.200 328.400 349.600 ;
        RECT 329.000 348.800 329.800 349.600 ;
        RECT 329.200 348.400 329.800 348.800 ;
        RECT 329.200 347.600 330.000 348.400 ;
        RECT 334.000 347.600 334.800 349.200 ;
        RECT 335.800 346.200 336.400 349.600 ;
        RECT 337.000 348.800 337.800 349.600 ;
        RECT 337.200 348.400 337.800 348.800 ;
        RECT 345.200 348.400 345.800 351.600 ;
        RECT 348.600 351.200 349.200 351.800 ;
        RECT 354.800 351.600 355.600 352.400 ;
        RECT 346.800 349.600 347.600 351.200 ;
        RECT 348.600 350.600 350.600 351.200 ;
        RECT 350.000 350.400 350.600 350.600 ;
        RECT 352.400 350.400 353.200 350.800 ;
        RECT 350.000 349.600 350.800 350.400 ;
        RECT 352.400 349.800 354.000 350.400 ;
        RECT 353.200 349.600 354.000 349.800 ;
        RECT 348.600 348.800 349.400 349.600 ;
        RECT 348.600 348.400 349.200 348.800 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 344.200 348.200 345.800 348.400 ;
        RECT 344.000 347.800 345.800 348.200 ;
        RECT 346.800 348.300 347.600 348.400 ;
        RECT 348.400 348.300 349.200 348.400 ;
        RECT 319.400 342.200 321.000 346.200 ;
        RECT 327.400 342.200 329.000 346.200 ;
        RECT 335.400 342.200 337.000 346.200 ;
        RECT 344.000 342.200 344.800 347.800 ;
        RECT 346.800 347.700 349.200 348.300 ;
        RECT 346.800 347.600 347.600 347.700 ;
        RECT 348.400 347.600 349.200 347.700 ;
        RECT 350.000 346.200 350.600 349.600 ;
        RECT 351.600 347.600 352.400 349.200 ;
        RECT 355.000 348.400 355.600 351.600 ;
        RECT 359.600 350.800 360.400 352.400 ;
        RECT 361.200 351.600 362.000 353.200 ;
        RECT 357.200 349.600 358.800 350.400 ;
        RECT 361.200 350.300 362.000 350.400 ;
        RECT 362.800 350.300 363.600 359.800 ;
        RECT 366.000 351.600 366.800 353.200 ;
        RECT 361.200 349.700 363.600 350.300 ;
        RECT 361.200 349.600 362.000 349.700 ;
        RECT 355.000 348.200 356.600 348.400 ;
        RECT 355.000 347.800 356.800 348.200 ;
        RECT 349.400 342.200 351.000 346.200 ;
        RECT 356.000 342.200 356.800 347.800 ;
        RECT 362.800 346.200 363.600 349.700 ;
        RECT 364.400 346.800 365.200 348.400 ;
        RECT 367.600 346.200 368.400 359.800 ;
        RECT 370.800 352.400 371.600 359.800 ;
        RECT 374.000 359.200 378.000 359.800 ;
        RECT 374.000 352.400 374.800 359.200 ;
        RECT 370.800 351.800 374.800 352.400 ;
        RECT 375.600 351.800 376.400 358.600 ;
        RECT 377.200 351.800 378.000 359.200 ;
        RECT 380.400 355.800 381.200 359.800 ;
        RECT 380.600 355.600 381.200 355.800 ;
        RECT 383.600 355.800 384.400 359.800 ;
        RECT 383.600 355.600 384.200 355.800 ;
        RECT 380.600 355.000 384.200 355.600 ;
        RECT 382.000 352.800 382.800 354.400 ;
        RECT 383.600 352.400 384.200 355.000 ;
        RECT 375.600 351.200 376.200 351.800 ;
        RECT 371.600 350.400 372.400 350.800 ;
        RECT 374.200 350.600 376.200 351.200 ;
        RECT 374.200 350.400 374.800 350.600 ;
        RECT 370.800 349.800 372.400 350.400 ;
        RECT 370.800 349.600 371.600 349.800 ;
        RECT 374.000 349.600 374.800 350.400 ;
        RECT 377.200 349.600 378.000 351.200 ;
        RECT 378.800 350.800 379.600 352.400 ;
        RECT 383.600 351.600 384.400 352.400 ;
        RECT 386.800 352.000 387.600 359.800 ;
        RECT 390.000 355.200 390.800 359.800 ;
        RECT 380.400 349.600 382.000 350.400 ;
        RECT 369.200 346.800 370.000 348.400 ;
        RECT 372.400 347.600 373.200 349.200 ;
        RECT 374.200 346.200 374.800 349.600 ;
        RECT 375.400 348.800 376.200 349.600 ;
        RECT 375.600 348.400 376.200 348.800 ;
        RECT 383.600 348.400 384.200 351.600 ;
        RECT 375.600 347.600 376.400 348.400 ;
        RECT 382.600 348.200 384.200 348.400 ;
        RECT 382.400 347.800 384.200 348.200 ;
        RECT 386.600 351.200 387.600 352.000 ;
        RECT 388.200 354.600 390.800 355.200 ;
        RECT 388.200 353.000 388.800 354.600 ;
        RECT 393.200 354.400 394.000 359.800 ;
        RECT 396.400 357.000 397.200 359.800 ;
        RECT 398.000 357.000 398.800 359.800 ;
        RECT 399.600 357.000 400.400 359.800 ;
        RECT 394.600 354.400 398.800 355.200 ;
        RECT 391.400 353.600 394.000 354.400 ;
        RECT 401.200 353.600 402.000 359.800 ;
        RECT 404.400 355.000 405.200 359.800 ;
        RECT 407.600 355.000 408.400 359.800 ;
        RECT 409.200 357.000 410.000 359.800 ;
        RECT 410.800 357.000 411.600 359.800 ;
        RECT 414.000 355.200 414.800 359.800 ;
        RECT 417.200 356.400 418.000 359.800 ;
        RECT 417.200 355.800 418.200 356.400 ;
        RECT 417.600 355.200 418.200 355.800 ;
        RECT 412.800 354.400 417.000 355.200 ;
        RECT 417.600 354.600 419.600 355.200 ;
        RECT 404.400 353.600 407.000 354.400 ;
        RECT 407.600 353.800 413.400 354.400 ;
        RECT 416.400 354.000 417.000 354.400 ;
        RECT 396.400 353.000 397.200 353.200 ;
        RECT 388.200 352.400 397.200 353.000 ;
        RECT 399.600 353.000 400.400 353.200 ;
        RECT 407.600 353.000 408.200 353.800 ;
        RECT 414.000 353.200 415.400 353.800 ;
        RECT 416.400 353.200 418.000 354.000 ;
        RECT 399.600 352.400 408.200 353.000 ;
        RECT 409.200 353.000 415.400 353.200 ;
        RECT 409.200 352.600 414.600 353.000 ;
        RECT 409.200 352.400 410.000 352.600 ;
        RECT 361.800 345.600 363.600 346.200 ;
        RECT 366.600 345.600 368.400 346.200 ;
        RECT 361.800 342.200 362.600 345.600 ;
        RECT 366.600 344.400 367.400 345.600 ;
        RECT 366.000 343.600 367.400 344.400 ;
        RECT 366.600 342.200 367.400 343.600 ;
        RECT 373.800 342.200 375.400 346.200 ;
        RECT 382.400 342.200 383.200 347.800 ;
        RECT 386.600 346.800 387.400 351.200 ;
        RECT 388.200 350.600 388.800 352.400 ;
        RECT 388.000 350.000 388.800 350.600 ;
        RECT 394.800 350.000 418.200 350.600 ;
        RECT 388.000 348.000 388.600 350.000 ;
        RECT 394.800 349.400 395.600 350.000 ;
        RECT 412.400 349.600 413.200 350.000 ;
        RECT 415.600 349.600 416.400 350.000 ;
        RECT 417.400 349.800 418.200 350.000 ;
        RECT 389.200 348.600 393.000 349.400 ;
        RECT 388.000 347.400 389.200 348.000 ;
        RECT 385.200 346.300 386.000 346.400 ;
        RECT 386.600 346.300 387.600 346.800 ;
        RECT 385.200 345.700 387.600 346.300 ;
        RECT 385.200 345.600 386.000 345.700 ;
        RECT 386.800 342.200 387.600 345.700 ;
        RECT 388.400 342.200 389.200 347.400 ;
        RECT 392.200 347.400 393.000 348.600 ;
        RECT 392.200 346.800 394.000 347.400 ;
        RECT 393.200 346.200 394.000 346.800 ;
        RECT 398.000 346.400 398.800 349.200 ;
        RECT 401.200 348.600 404.400 349.400 ;
        RECT 408.200 348.600 410.200 349.400 ;
        RECT 418.800 349.000 419.600 354.600 ;
        RECT 422.000 354.300 422.800 354.400 ;
        RECT 426.000 354.300 426.800 354.400 ;
        RECT 422.000 353.700 426.800 354.300 ;
        RECT 422.000 353.600 422.800 353.700 ;
        RECT 426.000 353.600 426.800 353.700 ;
        RECT 426.000 352.400 426.600 353.600 ;
        RECT 427.400 352.400 428.200 359.800 ;
        RECT 425.200 351.800 426.600 352.400 ;
        RECT 427.200 351.800 428.200 352.400 ;
        RECT 425.200 351.600 426.000 351.800 ;
        RECT 400.800 347.800 401.600 348.000 ;
        RECT 400.800 347.200 405.200 347.800 ;
        RECT 404.400 347.000 405.200 347.200 ;
        RECT 406.000 346.800 406.800 348.400 ;
        RECT 393.200 345.400 395.600 346.200 ;
        RECT 398.000 345.600 399.000 346.400 ;
        RECT 402.000 345.600 403.600 346.400 ;
        RECT 404.400 346.200 405.200 346.400 ;
        RECT 408.200 346.200 409.000 348.600 ;
        RECT 410.800 348.200 419.600 349.000 ;
        RECT 427.200 348.400 427.800 351.800 ;
        RECT 428.400 348.800 429.200 350.400 ;
        RECT 414.200 346.800 417.200 347.600 ;
        RECT 414.200 346.200 415.000 346.800 ;
        RECT 404.400 345.600 409.000 346.200 ;
        RECT 394.800 342.200 395.600 345.400 ;
        RECT 412.400 345.400 415.000 346.200 ;
        RECT 396.400 342.200 397.200 345.000 ;
        RECT 398.000 342.200 398.800 345.000 ;
        RECT 399.600 342.200 400.400 345.000 ;
        RECT 401.200 342.200 402.000 345.000 ;
        RECT 404.400 342.200 405.200 345.000 ;
        RECT 407.600 342.200 408.400 345.000 ;
        RECT 409.200 342.200 410.000 345.000 ;
        RECT 410.800 342.200 411.600 345.000 ;
        RECT 412.400 342.200 413.200 345.400 ;
        RECT 418.800 342.200 419.600 348.200 ;
        RECT 425.200 347.600 427.800 348.400 ;
        RECT 430.000 348.200 430.800 348.400 ;
        RECT 429.200 347.600 430.800 348.200 ;
        RECT 425.400 346.200 426.000 347.600 ;
        RECT 429.200 347.200 430.000 347.600 ;
        RECT 431.600 346.800 432.400 348.400 ;
        RECT 427.000 346.200 430.600 346.600 ;
        RECT 433.200 346.200 434.000 359.800 ;
        RECT 434.800 351.600 435.600 353.200 ;
        RECT 438.000 352.000 438.800 359.800 ;
        RECT 441.200 355.200 442.000 359.800 ;
        RECT 437.800 351.200 438.800 352.000 ;
        RECT 439.400 354.600 442.000 355.200 ;
        RECT 439.400 353.000 440.000 354.600 ;
        RECT 444.400 354.400 445.200 359.800 ;
        RECT 447.600 357.000 448.400 359.800 ;
        RECT 449.200 357.000 450.000 359.800 ;
        RECT 450.800 357.000 451.600 359.800 ;
        RECT 445.800 354.400 450.000 355.200 ;
        RECT 442.600 353.600 445.200 354.400 ;
        RECT 452.400 353.600 453.200 359.800 ;
        RECT 455.600 355.000 456.400 359.800 ;
        RECT 458.800 355.000 459.600 359.800 ;
        RECT 460.400 357.000 461.200 359.800 ;
        RECT 462.000 357.000 462.800 359.800 ;
        RECT 465.200 355.200 466.000 359.800 ;
        RECT 468.400 356.400 469.200 359.800 ;
        RECT 468.400 355.800 469.400 356.400 ;
        RECT 468.800 355.200 469.400 355.800 ;
        RECT 464.000 354.400 468.200 355.200 ;
        RECT 468.800 354.600 470.800 355.200 ;
        RECT 455.600 353.600 458.200 354.400 ;
        RECT 458.800 353.800 464.600 354.400 ;
        RECT 467.600 354.000 468.200 354.400 ;
        RECT 447.600 353.000 448.400 353.200 ;
        RECT 439.400 352.400 448.400 353.000 ;
        RECT 450.800 353.000 451.600 353.200 ;
        RECT 458.800 353.000 459.400 353.800 ;
        RECT 465.200 353.200 466.600 353.800 ;
        RECT 467.600 353.200 469.200 354.000 ;
        RECT 450.800 352.400 459.400 353.000 ;
        RECT 460.400 353.000 466.600 353.200 ;
        RECT 460.400 352.600 465.800 353.000 ;
        RECT 460.400 352.400 461.200 352.600 ;
        RECT 437.800 346.800 438.600 351.200 ;
        RECT 439.400 350.600 440.000 352.400 ;
        RECT 439.200 350.000 440.000 350.600 ;
        RECT 446.000 350.000 469.400 350.600 ;
        RECT 439.200 348.000 439.800 350.000 ;
        RECT 446.000 349.400 446.800 350.000 ;
        RECT 457.200 349.600 458.000 350.000 ;
        RECT 463.600 349.600 464.400 350.000 ;
        RECT 468.600 349.800 469.400 350.000 ;
        RECT 440.400 348.600 444.200 349.400 ;
        RECT 439.200 347.400 440.400 348.000 ;
        RECT 425.200 342.200 426.000 346.200 ;
        RECT 426.800 346.000 430.800 346.200 ;
        RECT 426.800 342.200 427.600 346.000 ;
        RECT 430.000 342.200 430.800 346.000 ;
        RECT 433.200 345.600 435.000 346.200 ;
        RECT 437.800 346.000 438.800 346.800 ;
        RECT 434.200 342.200 435.000 345.600 ;
        RECT 438.000 342.200 438.800 346.000 ;
        RECT 439.600 342.200 440.400 347.400 ;
        RECT 443.400 347.400 444.200 348.600 ;
        RECT 443.400 346.800 445.200 347.400 ;
        RECT 444.400 346.200 445.200 346.800 ;
        RECT 449.200 346.400 450.000 349.200 ;
        RECT 452.400 348.600 455.600 349.400 ;
        RECT 459.400 348.600 461.400 349.400 ;
        RECT 470.000 349.000 470.800 354.600 ;
        RECT 452.000 347.800 452.800 348.000 ;
        RECT 452.000 347.200 456.400 347.800 ;
        RECT 455.600 347.000 456.400 347.200 ;
        RECT 457.200 346.800 458.000 348.400 ;
        RECT 444.400 345.400 446.800 346.200 ;
        RECT 449.200 345.600 450.200 346.400 ;
        RECT 453.200 345.600 454.800 346.400 ;
        RECT 455.600 346.200 456.400 346.400 ;
        RECT 459.400 346.200 460.200 348.600 ;
        RECT 462.000 348.200 470.800 349.000 ;
        RECT 465.400 346.800 468.400 347.600 ;
        RECT 465.400 346.200 466.200 346.800 ;
        RECT 455.600 345.600 460.200 346.200 ;
        RECT 446.000 342.200 446.800 345.400 ;
        RECT 463.600 345.400 466.200 346.200 ;
        RECT 447.600 342.200 448.400 345.000 ;
        RECT 449.200 342.200 450.000 345.000 ;
        RECT 450.800 342.200 451.600 345.000 ;
        RECT 452.400 342.200 453.200 345.000 ;
        RECT 455.600 342.200 456.400 345.000 ;
        RECT 458.800 342.200 459.600 345.000 ;
        RECT 460.400 342.200 461.200 345.000 ;
        RECT 462.000 342.200 462.800 345.000 ;
        RECT 463.600 342.200 464.400 345.400 ;
        RECT 470.000 342.200 470.800 348.200 ;
        RECT 471.600 346.800 472.400 348.400 ;
        RECT 473.200 346.200 474.000 359.800 ;
        RECT 474.800 351.600 475.600 354.400 ;
        RECT 479.000 352.400 479.800 359.800 ;
        RECT 480.400 353.600 481.200 354.400 ;
        RECT 480.600 352.400 481.200 353.600 ;
        RECT 479.000 351.800 480.000 352.400 ;
        RECT 480.600 351.800 482.000 352.400 ;
        RECT 478.000 348.800 478.800 350.400 ;
        RECT 479.400 348.400 480.000 351.800 ;
        RECT 481.200 351.600 482.000 351.800 ;
        RECT 482.800 351.200 483.600 359.800 ;
        RECT 487.000 355.800 488.200 359.800 ;
        RECT 491.600 355.800 492.400 359.800 ;
        RECT 496.000 356.400 496.800 359.800 ;
        RECT 496.000 355.800 498.000 356.400 ;
        RECT 487.600 355.000 488.400 355.800 ;
        RECT 491.800 355.200 492.400 355.800 ;
        RECT 491.000 354.600 494.600 355.200 ;
        RECT 497.200 355.000 498.000 355.800 ;
        RECT 491.000 354.400 491.800 354.600 ;
        RECT 493.800 354.400 494.600 354.600 ;
        RECT 486.800 353.200 488.200 354.000 ;
        RECT 487.600 352.200 488.200 353.200 ;
        RECT 489.800 353.000 492.000 353.600 ;
        RECT 489.800 352.800 490.600 353.000 ;
        RECT 487.600 351.600 490.000 352.200 ;
        RECT 482.800 350.600 487.000 351.200 ;
        RECT 476.400 348.200 477.200 348.400 ;
        RECT 476.400 347.600 478.000 348.200 ;
        RECT 479.400 347.600 482.000 348.400 ;
        RECT 477.200 347.200 478.000 347.600 ;
        RECT 476.600 346.200 480.200 346.600 ;
        RECT 481.200 346.200 481.800 347.600 ;
        RECT 482.800 347.200 483.600 350.600 ;
        RECT 486.200 350.400 487.000 350.600 ;
        RECT 484.600 349.800 485.400 350.000 ;
        RECT 484.600 349.200 488.400 349.800 ;
        RECT 487.600 349.000 488.400 349.200 ;
        RECT 489.400 348.400 490.000 351.600 ;
        RECT 491.400 351.800 492.000 353.000 ;
        RECT 492.600 353.000 493.400 353.200 ;
        RECT 497.200 353.000 498.000 353.200 ;
        RECT 492.600 352.400 498.000 353.000 ;
        RECT 491.400 351.400 496.200 351.800 ;
        RECT 500.400 351.400 501.200 359.800 ;
        RECT 491.400 351.200 501.200 351.400 ;
        RECT 495.400 351.000 501.200 351.200 ;
        RECT 495.600 350.800 501.200 351.000 ;
        RECT 502.000 351.400 502.800 359.800 ;
        RECT 506.400 356.400 507.200 359.800 ;
        RECT 505.200 355.800 507.200 356.400 ;
        RECT 510.800 355.800 511.600 359.800 ;
        RECT 515.000 355.800 516.200 359.800 ;
        RECT 505.200 355.000 506.000 355.800 ;
        RECT 510.800 355.200 511.400 355.800 ;
        RECT 508.600 354.600 512.200 355.200 ;
        RECT 514.800 355.000 515.600 355.800 ;
        RECT 508.600 354.400 509.400 354.600 ;
        RECT 511.400 354.400 512.200 354.600 ;
        RECT 515.800 354.000 517.200 354.400 ;
        RECT 515.000 353.600 517.200 354.000 ;
        RECT 505.200 353.000 506.000 353.200 ;
        RECT 509.800 353.000 510.600 353.200 ;
        RECT 505.200 352.400 510.600 353.000 ;
        RECT 511.200 353.000 513.400 353.600 ;
        RECT 511.200 351.800 511.800 353.000 ;
        RECT 512.600 352.800 513.400 353.000 ;
        RECT 515.000 353.200 516.400 353.600 ;
        RECT 515.000 352.200 515.600 353.200 ;
        RECT 507.000 351.400 511.800 351.800 ;
        RECT 502.000 351.200 511.800 351.400 ;
        RECT 513.200 351.600 515.600 352.200 ;
        RECT 502.000 351.000 507.800 351.200 ;
        RECT 502.000 350.800 507.600 351.000 ;
        RECT 494.000 350.200 494.800 350.400 ;
        RECT 508.400 350.300 509.200 350.400 ;
        RECT 510.000 350.300 510.800 350.400 ;
        RECT 508.400 350.200 510.800 350.300 ;
        RECT 494.000 349.600 499.000 350.200 ;
        RECT 498.200 349.400 499.000 349.600 ;
        RECT 504.200 349.700 510.800 350.200 ;
        RECT 504.200 349.600 509.200 349.700 ;
        RECT 510.000 349.600 510.800 349.700 ;
        RECT 504.200 349.400 505.000 349.600 ;
        RECT 496.600 348.400 497.400 348.600 ;
        RECT 505.800 348.400 506.600 348.600 ;
        RECT 513.200 348.400 513.800 351.600 ;
        RECT 519.600 351.200 520.400 359.800 ;
        RECT 516.200 350.600 520.400 351.200 ;
        RECT 516.200 350.400 517.000 350.600 ;
        RECT 517.800 349.800 518.600 350.000 ;
        RECT 514.800 349.200 518.600 349.800 ;
        RECT 514.800 349.000 515.600 349.200 ;
        RECT 489.400 347.800 500.400 348.400 ;
        RECT 489.800 347.600 490.600 347.800 ;
        RECT 495.600 347.600 496.400 347.800 ;
        RECT 498.800 347.600 500.400 347.800 ;
        RECT 502.800 347.800 513.800 348.400 ;
        RECT 502.800 347.600 504.400 347.800 ;
        RECT 482.800 346.600 486.600 347.200 ;
        RECT 473.200 345.600 475.000 346.200 ;
        RECT 474.200 344.400 475.000 345.600 ;
        RECT 473.200 343.600 475.000 344.400 ;
        RECT 474.200 342.200 475.000 343.600 ;
        RECT 476.400 346.000 480.400 346.200 ;
        RECT 476.400 342.200 477.200 346.000 ;
        RECT 479.600 342.200 480.400 346.000 ;
        RECT 481.200 342.200 482.000 346.200 ;
        RECT 482.800 342.200 483.600 346.600 ;
        RECT 485.800 346.400 486.600 346.600 ;
        RECT 495.600 345.600 496.200 347.600 ;
        RECT 493.800 345.400 494.600 345.600 ;
        RECT 487.600 344.200 488.400 345.000 ;
        RECT 491.800 344.800 494.600 345.400 ;
        RECT 495.600 344.800 496.400 345.600 ;
        RECT 491.800 344.200 492.400 344.800 ;
        RECT 497.200 344.200 498.000 345.000 ;
        RECT 487.000 343.600 488.400 344.200 ;
        RECT 487.000 342.200 488.200 343.600 ;
        RECT 491.600 342.200 492.400 344.200 ;
        RECT 496.000 343.600 498.000 344.200 ;
        RECT 496.000 342.200 496.800 343.600 ;
        RECT 500.400 342.200 501.200 347.000 ;
        RECT 502.000 342.200 502.800 347.000 ;
        RECT 507.000 345.600 507.600 347.800 ;
        RECT 512.600 347.600 513.400 347.800 ;
        RECT 519.600 347.200 520.400 350.600 ;
        RECT 516.600 346.600 520.400 347.200 ;
        RECT 516.600 346.400 517.400 346.600 ;
        RECT 505.200 344.200 506.000 345.000 ;
        RECT 506.800 344.800 507.600 345.600 ;
        RECT 508.600 345.400 509.400 345.600 ;
        RECT 508.600 344.800 511.400 345.400 ;
        RECT 510.800 344.200 511.400 344.800 ;
        RECT 514.800 344.200 515.600 345.000 ;
        RECT 505.200 343.600 507.200 344.200 ;
        RECT 506.400 342.200 507.200 343.600 ;
        RECT 510.800 342.200 511.600 344.200 ;
        RECT 514.800 343.600 516.200 344.200 ;
        RECT 515.000 342.200 516.200 343.600 ;
        RECT 519.600 342.200 520.400 346.600 ;
        RECT 521.200 344.800 522.000 346.400 ;
        RECT 522.800 342.200 523.600 359.800 ;
        RECT 525.200 353.600 526.000 354.400 ;
        RECT 525.200 352.400 525.800 353.600 ;
        RECT 526.600 352.400 527.400 359.800 ;
        RECT 524.400 351.800 525.800 352.400 ;
        RECT 526.400 351.800 527.400 352.400 ;
        RECT 530.800 355.000 531.600 359.000 ;
        RECT 524.400 351.600 525.200 351.800 ;
        RECT 526.400 350.400 527.000 351.800 ;
        RECT 530.800 351.600 531.400 355.000 ;
        RECT 535.000 352.800 535.800 359.800 ;
        RECT 535.000 352.200 536.600 352.800 ;
        RECT 530.800 351.000 534.600 351.600 ;
        RECT 526.000 349.600 527.000 350.400 ;
        RECT 526.400 348.400 527.000 349.600 ;
        RECT 527.600 348.800 528.400 350.400 ;
        RECT 530.800 348.800 531.600 350.400 ;
        RECT 532.400 348.800 533.200 350.400 ;
        RECT 534.000 349.000 534.600 351.000 ;
        RECT 524.400 347.600 527.000 348.400 ;
        RECT 529.200 348.200 530.000 348.400 ;
        RECT 528.400 347.600 530.000 348.200 ;
        RECT 534.000 348.200 535.400 349.000 ;
        RECT 536.000 348.400 536.600 352.200 ;
        RECT 543.000 352.400 543.800 359.800 ;
        RECT 544.400 353.600 545.200 354.400 ;
        RECT 544.600 352.400 545.200 353.600 ;
        RECT 549.400 352.400 550.200 359.800 ;
        RECT 550.800 353.600 551.600 354.400 ;
        RECT 551.000 352.400 551.600 353.600 ;
        RECT 554.000 353.600 554.800 354.400 ;
        RECT 554.000 352.400 554.600 353.600 ;
        RECT 555.400 352.400 556.200 359.800 ;
        RECT 543.000 351.800 544.000 352.400 ;
        RECT 544.600 351.800 546.000 352.400 ;
        RECT 537.200 350.300 538.000 351.200 ;
        RECT 538.800 350.300 539.600 350.400 ;
        RECT 537.200 349.700 539.600 350.300 ;
        RECT 537.200 349.600 538.000 349.700 ;
        RECT 538.800 349.600 539.600 349.700 ;
        RECT 542.000 348.800 542.800 350.400 ;
        RECT 543.400 348.400 544.000 351.800 ;
        RECT 545.200 351.600 546.000 351.800 ;
        RECT 548.400 351.600 550.400 352.400 ;
        RECT 551.000 351.800 552.400 352.400 ;
        RECT 551.600 351.600 552.400 351.800 ;
        RECT 553.200 351.800 554.600 352.400 ;
        RECT 555.200 351.800 556.200 352.400 ;
        RECT 553.200 351.600 554.000 351.800 ;
        RECT 548.400 348.800 549.200 350.400 ;
        RECT 549.800 348.400 550.400 351.600 ;
        RECT 551.600 350.300 552.400 350.400 ;
        RECT 555.200 350.300 555.800 351.800 ;
        RECT 551.600 349.700 555.800 350.300 ;
        RECT 551.600 349.600 552.400 349.700 ;
        RECT 555.200 348.400 555.800 349.700 ;
        RECT 556.400 348.800 557.200 350.400 ;
        RECT 534.000 347.800 535.000 348.200 ;
        RECT 524.600 346.200 525.200 347.600 ;
        RECT 528.400 347.200 529.200 347.600 ;
        RECT 530.800 347.200 535.000 347.800 ;
        RECT 536.000 347.600 538.000 348.400 ;
        RECT 540.400 348.200 541.200 348.400 ;
        RECT 543.400 348.300 546.000 348.400 ;
        RECT 546.800 348.300 547.600 348.400 ;
        RECT 543.400 348.200 547.600 348.300 ;
        RECT 540.400 347.600 542.000 348.200 ;
        RECT 543.400 347.700 548.400 348.200 ;
        RECT 543.400 347.600 546.000 347.700 ;
        RECT 546.800 347.600 548.400 347.700 ;
        RECT 549.800 347.600 552.400 348.400 ;
        RECT 553.200 347.600 555.800 348.400 ;
        RECT 558.000 348.300 558.800 348.400 ;
        RECT 559.600 348.300 560.400 359.800 ;
        RECT 562.800 351.600 563.600 353.200 ;
        RECT 558.000 348.200 560.400 348.300 ;
        RECT 557.200 347.700 560.400 348.200 ;
        RECT 557.200 347.600 558.800 347.700 ;
        RECT 526.200 346.200 529.800 346.600 ;
        RECT 524.400 342.200 525.200 346.200 ;
        RECT 526.000 346.000 530.000 346.200 ;
        RECT 526.000 342.200 526.800 346.000 ;
        RECT 529.200 342.200 530.000 346.000 ;
        RECT 530.800 345.000 531.400 347.200 ;
        RECT 536.000 347.000 536.600 347.600 ;
        RECT 541.200 347.200 542.000 347.600 ;
        RECT 535.800 346.600 536.600 347.000 ;
        RECT 535.000 346.400 536.600 346.600 ;
        RECT 534.000 346.000 536.600 346.400 ;
        RECT 540.600 346.200 544.200 346.600 ;
        RECT 545.200 346.200 545.800 347.600 ;
        RECT 547.600 347.200 548.400 347.600 ;
        RECT 547.000 346.200 550.600 346.600 ;
        RECT 551.600 346.200 552.200 347.600 ;
        RECT 553.400 346.200 554.000 347.600 ;
        RECT 557.200 347.200 558.000 347.600 ;
        RECT 555.000 346.200 558.600 346.600 ;
        RECT 540.400 346.000 544.400 346.200 ;
        RECT 534.000 345.600 535.800 346.000 ;
        RECT 530.800 343.000 531.600 345.000 ;
        RECT 535.000 343.000 535.800 345.600 ;
        RECT 540.400 342.200 541.200 346.000 ;
        RECT 543.600 342.200 544.400 346.000 ;
        RECT 545.200 342.200 546.000 346.200 ;
        RECT 546.800 346.000 550.800 346.200 ;
        RECT 546.800 342.200 547.600 346.000 ;
        RECT 550.000 342.200 550.800 346.000 ;
        RECT 551.600 342.200 552.400 346.200 ;
        RECT 553.200 342.200 554.000 346.200 ;
        RECT 554.800 346.000 558.800 346.200 ;
        RECT 554.800 342.200 555.600 346.000 ;
        RECT 558.000 342.200 558.800 346.000 ;
        RECT 559.600 342.200 560.400 347.700 ;
        RECT 562.800 348.300 563.600 348.400 ;
        RECT 564.400 348.300 565.200 359.800 ;
        RECT 576.200 358.400 577.000 359.800 ;
        RECT 576.200 357.600 578.000 358.400 ;
        RECT 576.200 352.800 577.000 357.600 ;
        RECT 580.400 355.000 581.200 359.000 ;
        RECT 575.400 352.200 577.000 352.800 ;
        RECT 574.000 349.600 574.800 351.200 ;
        RECT 575.400 348.400 576.000 352.200 ;
        RECT 580.600 351.600 581.200 355.000 ;
        RECT 585.800 352.800 586.600 359.800 ;
        RECT 590.000 355.000 590.800 359.000 ;
        RECT 577.400 351.000 581.200 351.600 ;
        RECT 585.000 352.200 586.600 352.800 ;
        RECT 577.400 349.000 578.000 351.000 ;
        RECT 562.800 347.700 565.200 348.300 ;
        RECT 562.800 347.600 563.600 347.700 ;
        RECT 561.200 344.800 562.000 346.400 ;
        RECT 564.400 346.200 565.200 347.700 ;
        RECT 566.000 346.800 566.800 348.400 ;
        RECT 574.000 347.600 576.000 348.400 ;
        RECT 576.600 348.200 578.000 349.000 ;
        RECT 578.800 348.800 579.600 350.400 ;
        RECT 580.400 348.800 581.200 350.400 ;
        RECT 583.600 349.600 584.400 351.200 ;
        RECT 585.000 348.400 585.600 352.200 ;
        RECT 590.200 351.600 590.800 355.000 ;
        RECT 587.000 351.000 590.800 351.600 ;
        RECT 591.600 351.400 592.400 359.800 ;
        RECT 596.000 356.400 596.800 359.800 ;
        RECT 594.800 355.800 596.800 356.400 ;
        RECT 600.400 355.800 601.200 359.800 ;
        RECT 604.600 355.800 605.800 359.800 ;
        RECT 594.800 355.000 595.600 355.800 ;
        RECT 600.400 355.200 601.000 355.800 ;
        RECT 598.200 354.600 601.800 355.200 ;
        RECT 604.400 355.000 605.200 355.800 ;
        RECT 598.200 354.400 599.000 354.600 ;
        RECT 601.000 354.400 601.800 354.600 ;
        RECT 594.800 353.000 595.600 353.200 ;
        RECT 599.400 353.000 600.200 353.200 ;
        RECT 594.800 352.400 600.200 353.000 ;
        RECT 600.800 353.000 603.000 353.600 ;
        RECT 600.800 351.800 601.400 353.000 ;
        RECT 602.200 352.800 603.000 353.000 ;
        RECT 604.600 353.200 606.000 354.000 ;
        RECT 604.600 352.200 605.200 353.200 ;
        RECT 596.600 351.400 601.400 351.800 ;
        RECT 591.600 351.200 601.400 351.400 ;
        RECT 602.800 351.600 605.200 352.200 ;
        RECT 591.600 351.000 597.400 351.200 ;
        RECT 587.000 349.000 587.600 351.000 ;
        RECT 591.600 350.800 597.200 351.000 ;
        RECT 575.400 347.000 576.000 347.600 ;
        RECT 577.000 347.800 578.000 348.200 ;
        RECT 577.000 347.200 581.200 347.800 ;
        RECT 583.600 347.600 585.600 348.400 ;
        RECT 586.200 348.200 587.600 349.000 ;
        RECT 588.400 348.800 589.200 350.400 ;
        RECT 590.000 348.800 590.800 350.400 ;
        RECT 598.000 350.300 598.800 350.400 ;
        RECT 599.600 350.300 600.400 350.400 ;
        RECT 598.000 350.200 600.400 350.300 ;
        RECT 593.800 349.700 600.400 350.200 ;
        RECT 593.800 349.600 598.800 349.700 ;
        RECT 599.600 349.600 600.400 349.700 ;
        RECT 593.800 349.400 594.600 349.600 ;
        RECT 595.400 348.400 596.200 348.600 ;
        RECT 602.800 348.400 603.400 351.600 ;
        RECT 606.000 351.200 606.800 352.400 ;
        RECT 609.200 351.200 610.000 359.800 ;
        RECT 613.400 352.400 614.200 359.800 ;
        RECT 614.800 353.600 615.600 354.400 ;
        RECT 615.000 352.400 615.600 353.600 ;
        RECT 618.000 353.600 618.800 354.400 ;
        RECT 618.000 352.400 618.600 353.600 ;
        RECT 619.400 352.400 620.200 359.800 ;
        RECT 613.400 351.800 614.400 352.400 ;
        RECT 615.000 351.800 616.400 352.400 ;
        RECT 605.800 350.600 610.000 351.200 ;
        RECT 605.800 350.400 606.600 350.600 ;
        RECT 607.400 349.800 608.200 350.000 ;
        RECT 604.400 349.200 608.200 349.800 ;
        RECT 604.400 349.000 605.200 349.200 ;
        RECT 563.400 345.600 565.200 346.200 ;
        RECT 575.400 346.600 576.200 347.000 ;
        RECT 575.400 346.000 577.000 346.600 ;
        RECT 563.400 342.200 564.200 345.600 ;
        RECT 576.200 343.000 577.000 346.000 ;
        RECT 580.600 345.000 581.200 347.200 ;
        RECT 585.000 347.000 585.600 347.600 ;
        RECT 586.600 347.800 587.600 348.200 ;
        RECT 592.400 347.800 603.400 348.400 ;
        RECT 586.600 347.200 590.800 347.800 ;
        RECT 592.400 347.600 594.000 347.800 ;
        RECT 596.400 347.600 597.200 347.800 ;
        RECT 602.200 347.600 603.000 347.800 ;
        RECT 585.000 346.600 585.800 347.000 ;
        RECT 585.000 346.000 586.600 346.600 ;
        RECT 580.400 343.000 581.200 345.000 ;
        RECT 585.800 344.400 586.600 346.000 ;
        RECT 590.200 345.000 590.800 347.200 ;
        RECT 585.200 343.600 586.600 344.400 ;
        RECT 585.800 343.000 586.600 343.600 ;
        RECT 590.000 343.000 590.800 345.000 ;
        RECT 591.600 342.200 592.400 347.000 ;
        RECT 596.600 345.600 597.200 347.600 ;
        RECT 609.200 347.200 610.000 350.600 ;
        RECT 613.800 350.400 614.400 351.800 ;
        RECT 615.600 351.600 616.400 351.800 ;
        RECT 617.200 351.800 618.600 352.400 ;
        RECT 619.200 351.800 620.200 352.400 ;
        RECT 623.600 355.000 624.400 359.000 ;
        RECT 617.200 351.600 618.000 351.800 ;
        RECT 612.400 348.800 613.200 350.400 ;
        RECT 613.800 349.600 614.800 350.400 ;
        RECT 615.700 350.300 616.300 351.600 ;
        RECT 619.200 350.300 619.800 351.800 ;
        RECT 623.600 351.600 624.200 355.000 ;
        RECT 627.800 352.800 628.600 359.800 ;
        RECT 627.800 352.200 629.400 352.800 ;
        RECT 623.600 351.000 627.400 351.600 ;
        RECT 615.700 349.700 619.800 350.300 ;
        RECT 613.800 348.400 614.400 349.600 ;
        RECT 619.200 348.400 619.800 349.700 ;
        RECT 620.400 348.800 621.200 350.400 ;
        RECT 623.600 348.800 624.400 350.400 ;
        RECT 625.200 348.800 626.000 350.400 ;
        RECT 626.800 349.000 627.400 351.000 ;
        RECT 610.800 348.200 611.600 348.400 ;
        RECT 610.800 347.600 612.400 348.200 ;
        RECT 613.800 347.600 616.400 348.400 ;
        RECT 617.200 347.600 619.800 348.400 ;
        RECT 622.000 348.200 622.800 348.400 ;
        RECT 621.200 347.600 622.800 348.200 ;
        RECT 626.800 348.200 628.200 349.000 ;
        RECT 628.800 348.400 629.400 352.200 ;
        RECT 635.800 352.400 636.600 359.800 ;
        RECT 637.200 353.600 638.000 354.400 ;
        RECT 637.400 352.400 638.000 353.600 ;
        RECT 640.400 353.600 641.200 354.400 ;
        RECT 640.400 352.400 641.000 353.600 ;
        RECT 641.800 352.400 642.600 359.800 ;
        RECT 635.800 351.800 636.800 352.400 ;
        RECT 637.400 351.800 638.800 352.400 ;
        RECT 630.000 350.300 630.800 351.200 ;
        RECT 633.200 350.300 634.000 350.400 ;
        RECT 630.000 349.700 634.000 350.300 ;
        RECT 630.000 349.600 630.800 349.700 ;
        RECT 633.200 349.600 634.000 349.700 ;
        RECT 634.800 348.800 635.600 350.400 ;
        RECT 636.200 350.300 636.800 351.800 ;
        RECT 638.000 351.600 638.800 351.800 ;
        RECT 639.600 351.800 641.000 352.400 ;
        RECT 641.600 351.800 642.600 352.400 ;
        RECT 646.600 352.600 647.400 359.800 ;
        RECT 646.600 351.800 648.400 352.600 ;
        RECT 639.600 351.600 640.400 351.800 ;
        RECT 639.700 350.300 640.300 351.600 ;
        RECT 636.200 349.700 640.300 350.300 ;
        RECT 636.200 348.400 636.800 349.700 ;
        RECT 641.600 348.400 642.200 351.800 ;
        RECT 642.800 348.800 643.600 350.400 ;
        RECT 646.000 349.600 646.800 351.200 ;
        RECT 647.600 350.400 648.200 351.800 ;
        RECT 650.800 351.200 651.600 359.800 ;
        RECT 655.000 355.800 656.200 359.800 ;
        RECT 659.600 355.800 660.400 359.800 ;
        RECT 664.000 356.400 664.800 359.800 ;
        RECT 664.000 355.800 666.000 356.400 ;
        RECT 655.600 355.000 656.400 355.800 ;
        RECT 659.800 355.200 660.400 355.800 ;
        RECT 659.000 354.600 662.600 355.200 ;
        RECT 665.200 355.000 666.000 355.800 ;
        RECT 659.000 354.400 659.800 354.600 ;
        RECT 661.800 354.400 662.600 354.600 ;
        RECT 654.800 353.200 656.200 354.000 ;
        RECT 655.600 352.200 656.200 353.200 ;
        RECT 657.800 353.000 660.000 353.600 ;
        RECT 657.800 352.800 658.600 353.000 ;
        RECT 655.600 351.600 658.000 352.200 ;
        RECT 650.800 350.600 655.000 351.200 ;
        RECT 647.600 349.600 648.400 350.400 ;
        RECT 647.600 348.400 648.200 349.600 ;
        RECT 626.800 347.800 627.800 348.200 ;
        RECT 611.600 347.200 612.400 347.600 ;
        RECT 606.200 346.600 610.000 347.200 ;
        RECT 606.200 346.400 607.000 346.600 ;
        RECT 594.800 344.200 595.600 345.000 ;
        RECT 596.400 344.800 597.200 345.600 ;
        RECT 598.200 345.400 599.000 345.600 ;
        RECT 598.200 344.800 601.000 345.400 ;
        RECT 600.400 344.200 601.000 344.800 ;
        RECT 604.400 344.200 605.200 345.000 ;
        RECT 594.800 343.600 596.800 344.200 ;
        RECT 596.000 342.200 596.800 343.600 ;
        RECT 600.400 342.200 601.200 344.200 ;
        RECT 604.400 343.600 605.800 344.200 ;
        RECT 604.600 342.200 605.800 343.600 ;
        RECT 609.200 342.200 610.000 346.600 ;
        RECT 611.000 346.200 614.600 346.600 ;
        RECT 615.600 346.200 616.200 347.600 ;
        RECT 617.400 346.200 618.000 347.600 ;
        RECT 621.200 347.200 622.000 347.600 ;
        RECT 623.600 347.200 627.800 347.800 ;
        RECT 628.800 347.600 630.800 348.400 ;
        RECT 633.200 348.200 634.000 348.400 ;
        RECT 633.200 347.600 634.800 348.200 ;
        RECT 636.200 347.600 638.800 348.400 ;
        RECT 639.600 347.600 642.200 348.400 ;
        RECT 644.400 348.300 645.200 348.400 ;
        RECT 646.000 348.300 646.800 348.400 ;
        RECT 644.400 348.200 646.800 348.300 ;
        RECT 643.600 347.700 646.800 348.200 ;
        RECT 643.600 347.600 645.200 347.700 ;
        RECT 646.000 347.600 646.800 347.700 ;
        RECT 647.600 347.600 648.400 348.400 ;
        RECT 619.000 346.200 622.600 346.600 ;
        RECT 610.800 346.000 614.800 346.200 ;
        RECT 610.800 342.200 611.600 346.000 ;
        RECT 614.000 342.200 614.800 346.000 ;
        RECT 615.600 342.200 616.400 346.200 ;
        RECT 617.200 342.200 618.000 346.200 ;
        RECT 618.800 346.000 622.800 346.200 ;
        RECT 618.800 342.200 619.600 346.000 ;
        RECT 622.000 342.200 622.800 346.000 ;
        RECT 623.600 345.000 624.200 347.200 ;
        RECT 628.800 347.000 629.400 347.600 ;
        RECT 634.000 347.200 634.800 347.600 ;
        RECT 628.600 346.600 629.400 347.000 ;
        RECT 627.800 346.000 629.400 346.600 ;
        RECT 633.400 346.200 637.000 346.600 ;
        RECT 638.000 346.200 638.600 347.600 ;
        RECT 639.800 346.200 640.400 347.600 ;
        RECT 643.600 347.200 644.400 347.600 ;
        RECT 641.400 346.200 645.000 346.600 ;
        RECT 633.200 346.000 637.200 346.200 ;
        RECT 623.600 343.000 624.400 345.000 ;
        RECT 627.800 344.400 628.600 346.000 ;
        RECT 626.800 343.600 628.600 344.400 ;
        RECT 627.800 343.000 628.600 343.600 ;
        RECT 633.200 342.200 634.000 346.000 ;
        RECT 636.400 342.200 637.200 346.000 ;
        RECT 638.000 342.200 638.800 346.200 ;
        RECT 639.600 342.200 640.400 346.200 ;
        RECT 641.200 346.000 645.200 346.200 ;
        RECT 641.200 342.200 642.000 346.000 ;
        RECT 644.400 342.200 645.200 346.000 ;
        RECT 647.600 344.200 648.200 347.600 ;
        RECT 650.800 347.200 651.600 350.600 ;
        RECT 654.200 350.400 655.000 350.600 ;
        RECT 652.600 349.800 653.400 350.000 ;
        RECT 652.600 349.200 656.400 349.800 ;
        RECT 655.600 349.000 656.400 349.200 ;
        RECT 657.400 348.400 658.000 351.600 ;
        RECT 659.400 351.800 660.000 353.000 ;
        RECT 660.600 353.000 661.400 353.200 ;
        RECT 665.200 353.000 666.000 353.200 ;
        RECT 660.600 352.400 666.000 353.000 ;
        RECT 659.400 351.400 664.200 351.800 ;
        RECT 668.400 351.400 669.200 359.800 ;
        RECT 670.600 352.600 671.400 359.800 ;
        RECT 675.400 352.600 676.200 359.800 ;
        RECT 670.600 351.800 672.400 352.600 ;
        RECT 675.400 351.800 677.200 352.600 ;
        RECT 659.400 351.200 669.200 351.400 ;
        RECT 663.400 351.000 669.200 351.200 ;
        RECT 663.600 350.800 669.200 351.000 ;
        RECT 662.000 350.200 662.800 350.400 ;
        RECT 662.000 349.600 667.000 350.200 ;
        RECT 670.000 349.600 670.800 351.200 ;
        RECT 666.200 349.400 667.000 349.600 ;
        RECT 664.600 348.400 665.400 348.600 ;
        RECT 671.600 348.400 672.200 351.800 ;
        RECT 673.200 350.300 674.000 350.400 ;
        RECT 674.800 350.300 675.600 351.200 ;
        RECT 673.200 349.700 675.600 350.300 ;
        RECT 673.200 349.600 674.000 349.700 ;
        RECT 674.800 349.600 675.600 349.700 ;
        RECT 676.400 348.400 677.000 351.800 ;
        RECT 657.400 347.800 668.400 348.400 ;
        RECT 657.800 347.600 658.600 347.800 ;
        RECT 650.800 346.600 654.600 347.200 ;
        RECT 649.200 344.800 650.000 346.400 ;
        RECT 647.600 342.200 648.400 344.200 ;
        RECT 650.800 342.200 651.600 346.600 ;
        RECT 653.800 346.400 654.600 346.600 ;
        RECT 663.600 345.600 664.200 347.800 ;
        RECT 666.800 347.600 668.400 347.800 ;
        RECT 671.600 347.600 672.400 348.400 ;
        RECT 676.400 347.600 677.200 348.400 ;
        RECT 681.200 348.300 682.000 359.800 ;
        RECT 678.100 347.700 682.000 348.300 ;
        RECT 661.800 345.400 662.600 345.600 ;
        RECT 655.600 344.200 656.400 345.000 ;
        RECT 659.800 344.800 662.600 345.400 ;
        RECT 663.600 344.800 664.400 345.600 ;
        RECT 659.800 344.200 660.400 344.800 ;
        RECT 665.200 344.200 666.000 345.000 ;
        RECT 655.000 343.600 656.400 344.200 ;
        RECT 655.000 342.200 656.200 343.600 ;
        RECT 659.600 342.200 660.400 344.200 ;
        RECT 664.000 343.600 666.000 344.200 ;
        RECT 664.000 342.200 664.800 343.600 ;
        RECT 668.400 342.200 669.200 347.000 ;
        RECT 671.600 344.400 672.200 347.600 ;
        RECT 673.200 344.800 674.000 346.400 ;
        RECT 676.400 344.400 677.000 347.600 ;
        RECT 678.100 346.400 678.700 347.700 ;
        RECT 678.000 344.800 678.800 346.400 ;
        RECT 679.600 344.800 680.400 346.400 ;
        RECT 671.600 342.200 672.400 344.400 ;
        RECT 676.400 342.200 677.200 344.400 ;
        RECT 681.200 342.200 682.000 347.700 ;
        RECT 1.200 335.000 2.000 339.800 ;
        RECT 5.600 338.400 6.400 339.800 ;
        RECT 4.400 337.800 6.400 338.400 ;
        RECT 10.000 337.800 10.800 339.800 ;
        RECT 14.200 338.400 15.400 339.800 ;
        RECT 14.000 337.800 15.400 338.400 ;
        RECT 4.400 337.000 5.200 337.800 ;
        RECT 10.000 337.200 10.600 337.800 ;
        RECT 6.000 336.400 6.800 337.200 ;
        RECT 7.800 336.600 10.600 337.200 ;
        RECT 14.000 337.000 14.800 337.800 ;
        RECT 7.800 336.400 8.600 336.600 ;
        RECT 2.000 334.200 3.600 334.400 ;
        RECT 6.200 334.200 6.800 336.400 ;
        RECT 15.800 335.400 16.600 335.600 ;
        RECT 18.800 335.400 19.600 339.800 ;
        RECT 20.400 335.800 21.200 339.800 ;
        RECT 22.000 336.000 22.800 339.800 ;
        RECT 25.200 336.000 26.000 339.800 ;
        RECT 22.000 335.800 26.000 336.000 ;
        RECT 26.800 335.800 27.600 339.800 ;
        RECT 28.400 336.000 29.200 339.800 ;
        RECT 31.600 336.000 32.400 339.800 ;
        RECT 37.000 336.000 37.800 339.000 ;
        RECT 41.200 337.000 42.000 339.000 ;
        RECT 28.400 335.800 32.400 336.000 ;
        RECT 15.800 334.800 19.600 335.400 ;
        RECT 11.800 334.200 12.600 334.400 ;
        RECT 2.000 333.600 13.000 334.200 ;
        RECT 5.000 333.400 5.800 333.600 ;
        RECT 3.400 332.400 4.200 332.600 ;
        RECT 12.400 332.400 13.000 333.600 ;
        RECT 14.000 332.800 14.800 333.000 ;
        RECT 3.400 331.800 8.400 332.400 ;
        RECT 7.600 331.600 8.400 331.800 ;
        RECT 12.400 331.600 13.200 332.400 ;
        RECT 14.000 332.200 17.800 332.800 ;
        RECT 17.000 332.000 17.800 332.200 ;
        RECT 1.200 331.000 6.800 331.200 ;
        RECT 1.200 330.800 7.000 331.000 ;
        RECT 1.200 330.600 11.000 330.800 ;
        RECT 1.200 322.200 2.000 330.600 ;
        RECT 6.200 330.200 11.000 330.600 ;
        RECT 4.400 329.000 9.800 329.600 ;
        RECT 4.400 328.800 5.200 329.000 ;
        RECT 9.000 328.800 9.800 329.000 ;
        RECT 10.400 329.000 11.000 330.200 ;
        RECT 12.400 330.400 13.000 331.600 ;
        RECT 15.400 331.400 16.200 331.600 ;
        RECT 18.800 331.400 19.600 334.800 ;
        RECT 20.600 334.400 21.200 335.800 ;
        RECT 22.200 335.400 25.800 335.800 ;
        RECT 24.400 334.400 25.200 334.800 ;
        RECT 27.000 334.400 27.600 335.800 ;
        RECT 28.600 335.400 32.200 335.800 ;
        RECT 36.200 335.400 37.800 336.000 ;
        RECT 36.200 335.000 37.000 335.400 ;
        RECT 30.800 334.400 31.600 334.800 ;
        RECT 36.200 334.400 36.800 335.000 ;
        RECT 41.400 334.800 42.000 337.000 ;
        RECT 42.800 335.000 43.600 339.800 ;
        RECT 47.200 338.400 48.000 339.800 ;
        RECT 46.000 337.800 48.000 338.400 ;
        RECT 51.600 337.800 52.400 339.800 ;
        RECT 55.800 338.400 57.000 339.800 ;
        RECT 55.600 337.800 57.000 338.400 ;
        RECT 46.000 337.000 46.800 337.800 ;
        RECT 51.600 337.200 52.200 337.800 ;
        RECT 47.600 336.400 48.400 337.200 ;
        RECT 49.400 336.600 52.200 337.200 ;
        RECT 55.600 337.000 56.400 337.800 ;
        RECT 49.400 336.400 50.200 336.600 ;
        RECT 20.400 333.600 23.000 334.400 ;
        RECT 24.400 333.800 26.000 334.400 ;
        RECT 25.200 333.600 26.000 333.800 ;
        RECT 26.800 333.600 29.400 334.400 ;
        RECT 30.800 333.800 32.400 334.400 ;
        RECT 31.600 333.600 32.400 333.800 ;
        RECT 33.200 334.300 34.000 334.400 ;
        RECT 34.800 334.300 36.800 334.400 ;
        RECT 33.200 333.700 36.800 334.300 ;
        RECT 37.800 334.200 42.000 334.800 ;
        RECT 43.600 334.200 45.200 334.400 ;
        RECT 47.800 334.200 48.400 336.400 ;
        RECT 57.400 335.400 58.200 335.600 ;
        RECT 60.400 335.400 61.200 339.800 ;
        RECT 64.600 338.400 65.400 339.800 ;
        RECT 64.600 337.600 66.000 338.400 ;
        RECT 64.600 336.400 65.400 337.600 ;
        RECT 57.400 334.800 61.200 335.400 ;
        RECT 63.600 335.800 65.400 336.400 ;
        RECT 66.800 335.800 67.600 339.800 ;
        RECT 70.000 337.800 70.800 339.800 ;
        RECT 53.400 334.200 54.200 334.400 ;
        RECT 37.800 333.800 38.800 334.200 ;
        RECT 33.200 333.600 34.000 333.700 ;
        RECT 34.800 333.600 36.800 333.700 ;
        RECT 15.400 330.800 19.600 331.400 ;
        RECT 12.400 329.800 14.800 330.400 ;
        RECT 11.800 329.000 12.600 329.200 ;
        RECT 10.400 328.400 12.600 329.000 ;
        RECT 14.200 328.800 14.800 329.800 ;
        RECT 14.200 328.000 15.600 328.800 ;
        RECT 18.800 328.300 19.600 330.800 ;
        RECT 20.400 330.200 21.200 330.400 ;
        RECT 22.400 330.200 23.000 333.600 ;
        RECT 23.600 331.600 24.400 333.200 ;
        RECT 25.200 332.300 26.000 332.400 ;
        RECT 28.800 332.300 29.400 333.600 ;
        RECT 25.200 331.700 29.400 332.300 ;
        RECT 25.200 331.600 26.000 331.700 ;
        RECT 26.800 330.200 27.600 330.400 ;
        RECT 28.800 330.200 29.400 331.700 ;
        RECT 30.000 331.600 30.800 333.200 ;
        RECT 31.600 332.300 32.400 332.400 ;
        RECT 34.800 332.300 35.600 332.400 ;
        RECT 31.600 331.700 35.600 332.300 ;
        RECT 31.600 331.600 32.400 331.700 ;
        RECT 34.800 330.800 35.600 331.700 ;
        RECT 20.400 329.600 21.800 330.200 ;
        RECT 22.400 329.600 23.400 330.200 ;
        RECT 26.800 329.600 28.200 330.200 ;
        RECT 28.800 329.600 29.800 330.200 ;
        RECT 21.200 328.400 21.800 329.600 ;
        RECT 22.600 328.400 23.400 329.600 ;
        RECT 27.600 328.400 28.200 329.600 ;
        RECT 21.200 328.300 22.000 328.400 ;
        RECT 18.800 327.700 22.000 328.300 ;
        RECT 7.800 327.400 8.600 327.600 ;
        RECT 10.600 327.400 11.400 327.600 ;
        RECT 4.400 326.200 5.200 327.000 ;
        RECT 7.800 326.800 11.400 327.400 ;
        RECT 10.000 326.200 10.600 326.800 ;
        RECT 14.000 326.200 14.800 327.000 ;
        RECT 4.400 325.600 6.400 326.200 ;
        RECT 5.600 322.200 6.400 325.600 ;
        RECT 10.000 322.200 10.800 326.200 ;
        RECT 14.200 322.200 15.400 326.200 ;
        RECT 18.800 322.200 19.600 327.700 ;
        RECT 21.200 327.600 22.000 327.700 ;
        RECT 22.600 327.600 24.400 328.400 ;
        RECT 27.600 327.600 28.400 328.400 ;
        RECT 22.600 322.200 23.400 327.600 ;
        RECT 29.000 322.200 29.800 329.600 ;
        RECT 36.200 329.800 36.800 333.600 ;
        RECT 37.400 333.000 38.800 333.800 ;
        RECT 43.600 333.600 54.600 334.200 ;
        RECT 46.600 333.400 47.400 333.600 ;
        RECT 38.200 331.000 38.800 333.000 ;
        RECT 39.600 331.600 40.400 333.200 ;
        RECT 41.200 331.600 42.000 333.200 ;
        RECT 45.000 332.400 45.800 332.600 ;
        RECT 47.600 332.400 48.400 332.600 ;
        RECT 54.000 332.400 54.600 333.600 ;
        RECT 55.600 332.800 56.400 333.000 ;
        RECT 45.000 331.800 50.000 332.400 ;
        RECT 49.200 331.600 50.000 331.800 ;
        RECT 54.000 331.600 54.800 332.400 ;
        RECT 55.600 332.200 59.400 332.800 ;
        RECT 58.600 332.000 59.400 332.200 ;
        RECT 42.800 331.000 48.400 331.200 ;
        RECT 38.200 330.400 42.000 331.000 ;
        RECT 36.200 329.200 37.800 329.800 ;
        RECT 37.000 322.200 37.800 329.200 ;
        RECT 41.400 327.000 42.000 330.400 ;
        RECT 41.200 323.000 42.000 327.000 ;
        RECT 42.800 330.800 48.600 331.000 ;
        RECT 42.800 330.600 52.600 330.800 ;
        RECT 42.800 322.200 43.600 330.600 ;
        RECT 47.800 330.200 52.600 330.600 ;
        RECT 46.000 329.000 51.400 329.600 ;
        RECT 46.000 328.800 46.800 329.000 ;
        RECT 50.600 328.800 51.400 329.000 ;
        RECT 52.000 329.000 52.600 330.200 ;
        RECT 54.000 330.400 54.600 331.600 ;
        RECT 57.000 331.400 57.800 331.600 ;
        RECT 60.400 331.400 61.200 334.800 ;
        RECT 62.000 333.600 62.800 335.200 ;
        RECT 57.000 330.800 61.200 331.400 ;
        RECT 54.000 329.800 56.400 330.400 ;
        RECT 53.400 329.000 54.200 329.200 ;
        RECT 52.000 328.400 54.200 329.000 ;
        RECT 55.800 328.800 56.400 329.800 ;
        RECT 55.800 328.000 57.200 328.800 ;
        RECT 49.400 327.400 50.200 327.600 ;
        RECT 52.200 327.400 53.000 327.600 ;
        RECT 46.000 326.200 46.800 327.000 ;
        RECT 49.400 326.800 53.000 327.400 ;
        RECT 51.600 326.200 52.200 326.800 ;
        RECT 55.600 326.200 56.400 327.000 ;
        RECT 46.000 325.600 48.000 326.200 ;
        RECT 47.200 322.200 48.000 325.600 ;
        RECT 51.600 322.200 52.400 326.200 ;
        RECT 55.800 322.200 57.000 326.200 ;
        RECT 60.400 322.200 61.200 330.800 ;
        RECT 63.600 322.200 64.400 335.800 ;
        RECT 66.800 332.400 67.400 335.800 ;
        RECT 70.000 335.600 70.600 337.800 ;
        RECT 71.600 335.600 72.400 337.200 ;
        RECT 68.200 335.000 70.600 335.600 ;
        RECT 73.200 335.000 74.000 339.800 ;
        RECT 77.600 338.400 78.400 339.800 ;
        RECT 76.400 337.800 78.400 338.400 ;
        RECT 82.000 337.800 82.800 339.800 ;
        RECT 86.200 338.400 87.400 339.800 ;
        RECT 86.000 337.800 87.400 338.400 ;
        RECT 76.400 337.000 77.200 337.800 ;
        RECT 82.000 337.200 82.600 337.800 ;
        RECT 78.000 336.400 78.800 337.200 ;
        RECT 79.800 336.600 82.600 337.200 ;
        RECT 86.000 337.000 86.800 337.800 ;
        RECT 79.800 336.400 80.600 336.600 ;
        RECT 66.800 331.600 67.600 332.400 ;
        RECT 68.200 332.000 68.800 335.000 ;
        RECT 69.800 333.600 70.800 334.400 ;
        RECT 71.600 334.300 72.400 334.400 ;
        RECT 74.000 334.300 75.600 334.400 ;
        RECT 71.600 334.200 75.600 334.300 ;
        RECT 78.200 334.200 78.800 336.400 ;
        RECT 87.800 335.400 88.600 335.600 ;
        RECT 90.800 335.400 91.600 339.800 ;
        RECT 92.400 336.000 93.200 339.800 ;
        RECT 95.600 336.000 96.400 339.800 ;
        RECT 92.400 335.800 96.400 336.000 ;
        RECT 97.200 335.800 98.000 339.800 ;
        RECT 98.800 336.000 99.600 339.800 ;
        RECT 102.000 336.000 102.800 339.800 ;
        RECT 98.800 335.800 102.800 336.000 ;
        RECT 103.600 335.800 104.400 339.800 ;
        RECT 92.600 335.400 96.200 335.800 ;
        RECT 87.800 334.800 91.600 335.400 ;
        RECT 83.800 334.200 84.600 334.400 ;
        RECT 71.600 333.700 85.000 334.200 ;
        RECT 71.600 333.600 72.400 333.700 ;
        RECT 74.000 333.600 85.000 333.700 ;
        RECT 69.600 332.800 70.400 333.600 ;
        RECT 77.000 333.400 77.800 333.600 ;
        RECT 75.400 332.400 76.200 332.600 ;
        RECT 84.400 332.400 85.000 333.600 ;
        RECT 86.000 332.800 86.800 333.000 ;
        RECT 75.400 332.300 80.400 332.400 ;
        RECT 81.200 332.300 82.000 332.400 ;
        RECT 65.200 328.800 66.000 330.400 ;
        RECT 66.800 330.200 67.400 331.600 ;
        RECT 68.200 331.400 69.000 332.000 ;
        RECT 75.400 331.800 82.000 332.300 ;
        RECT 79.600 331.700 82.000 331.800 ;
        RECT 79.600 331.600 80.400 331.700 ;
        RECT 81.200 331.600 82.000 331.700 ;
        RECT 84.400 331.600 85.200 332.400 ;
        RECT 86.000 332.200 89.800 332.800 ;
        RECT 89.000 332.000 89.800 332.200 ;
        RECT 68.200 331.200 72.400 331.400 ;
        RECT 68.400 330.800 72.400 331.200 ;
        RECT 66.800 329.600 68.200 330.200 ;
        RECT 67.400 324.400 68.200 329.600 ;
        RECT 66.800 323.600 68.200 324.400 ;
        RECT 67.400 322.200 68.200 323.600 ;
        RECT 71.600 322.200 72.400 330.800 ;
        RECT 73.200 331.000 78.800 331.200 ;
        RECT 73.200 330.800 79.000 331.000 ;
        RECT 73.200 330.600 83.000 330.800 ;
        RECT 73.200 322.200 74.000 330.600 ;
        RECT 78.200 330.200 83.000 330.600 ;
        RECT 76.400 329.000 81.800 329.600 ;
        RECT 76.400 328.800 77.200 329.000 ;
        RECT 81.000 328.800 81.800 329.000 ;
        RECT 82.400 329.000 83.000 330.200 ;
        RECT 84.400 330.400 85.000 331.600 ;
        RECT 87.400 331.400 88.200 331.600 ;
        RECT 90.800 331.400 91.600 334.800 ;
        RECT 93.200 334.400 94.000 334.800 ;
        RECT 97.200 334.400 97.800 335.800 ;
        RECT 99.000 335.400 102.600 335.800 ;
        RECT 99.600 334.400 100.400 334.800 ;
        RECT 103.600 334.400 104.200 335.800 ;
        RECT 110.000 335.000 110.800 339.800 ;
        RECT 114.400 338.400 115.200 339.800 ;
        RECT 113.200 337.800 115.200 338.400 ;
        RECT 118.800 337.800 119.600 339.800 ;
        RECT 123.000 338.400 124.200 339.800 ;
        RECT 122.800 337.800 124.200 338.400 ;
        RECT 113.200 337.000 114.000 337.800 ;
        RECT 118.800 337.200 119.400 337.800 ;
        RECT 114.800 336.400 115.600 337.200 ;
        RECT 116.600 336.600 119.400 337.200 ;
        RECT 122.800 337.000 123.600 337.800 ;
        RECT 116.600 336.400 117.400 336.600 ;
        RECT 92.400 333.800 94.000 334.400 ;
        RECT 95.400 334.300 98.000 334.400 ;
        RECT 98.800 334.300 100.400 334.400 ;
        RECT 95.400 333.800 100.400 334.300 ;
        RECT 92.400 333.600 93.200 333.800 ;
        RECT 95.400 333.700 99.600 333.800 ;
        RECT 95.400 333.600 98.000 333.700 ;
        RECT 98.800 333.600 99.600 333.700 ;
        RECT 101.800 333.600 104.400 334.400 ;
        RECT 110.800 334.200 112.400 334.400 ;
        RECT 115.000 334.200 115.600 336.400 ;
        RECT 124.600 335.400 125.400 335.600 ;
        RECT 127.600 335.400 128.400 339.800 ;
        RECT 131.800 338.400 132.600 339.800 ;
        RECT 136.600 338.400 137.400 339.800 ;
        RECT 130.800 337.600 132.600 338.400 ;
        RECT 135.600 337.600 137.400 338.400 ;
        RECT 131.800 336.400 132.600 337.600 ;
        RECT 136.600 336.400 137.400 337.600 ;
        RECT 124.600 334.800 128.400 335.400 ;
        RECT 130.800 335.800 132.600 336.400 ;
        RECT 135.600 335.800 137.400 336.400 ;
        RECT 118.000 334.200 118.800 334.400 ;
        RECT 120.600 334.200 121.400 334.400 ;
        RECT 127.600 334.300 128.400 334.800 ;
        RECT 129.200 334.300 130.000 335.200 ;
        RECT 110.800 333.600 121.800 334.200 ;
        RECT 94.000 331.600 94.800 333.200 ;
        RECT 87.400 330.800 91.600 331.400 ;
        RECT 84.400 329.800 86.800 330.400 ;
        RECT 83.800 329.000 84.600 329.200 ;
        RECT 82.400 328.400 84.600 329.000 ;
        RECT 86.200 328.800 86.800 329.800 ;
        RECT 86.200 328.000 87.600 328.800 ;
        RECT 79.800 327.400 80.600 327.600 ;
        RECT 82.600 327.400 83.400 327.600 ;
        RECT 76.400 326.200 77.200 327.000 ;
        RECT 79.800 326.800 83.400 327.400 ;
        RECT 82.000 326.200 82.600 326.800 ;
        RECT 86.000 326.200 86.800 327.000 ;
        RECT 76.400 325.600 78.400 326.200 ;
        RECT 77.600 322.200 78.400 325.600 ;
        RECT 82.000 322.200 82.800 326.200 ;
        RECT 86.200 322.200 87.400 326.200 ;
        RECT 90.800 322.200 91.600 330.800 ;
        RECT 95.400 330.200 96.000 333.600 ;
        RECT 98.800 332.300 99.600 332.400 ;
        RECT 100.400 332.300 101.200 333.200 ;
        RECT 98.800 331.700 101.200 332.300 ;
        RECT 98.800 331.600 99.600 331.700 ;
        RECT 100.400 331.600 101.200 331.700 ;
        RECT 101.800 332.300 102.400 333.600 ;
        RECT 113.800 333.400 114.600 333.600 ;
        RECT 112.200 332.400 113.000 332.600 ;
        RECT 114.800 332.400 115.600 332.600 ;
        RECT 108.400 332.300 109.200 332.400 ;
        RECT 101.800 331.700 109.200 332.300 ;
        RECT 112.200 331.800 117.200 332.400 ;
        RECT 97.200 330.200 98.000 330.400 ;
        RECT 101.800 330.200 102.400 331.700 ;
        RECT 108.400 331.600 109.200 331.700 ;
        RECT 116.400 331.600 117.200 331.800 ;
        RECT 110.000 331.000 115.600 331.200 ;
        RECT 110.000 330.800 115.800 331.000 ;
        RECT 110.000 330.600 119.800 330.800 ;
        RECT 103.600 330.200 104.400 330.400 ;
        RECT 95.000 329.600 96.000 330.200 ;
        RECT 96.600 329.600 98.000 330.200 ;
        RECT 101.400 329.600 102.400 330.200 ;
        RECT 103.000 329.600 104.400 330.200 ;
        RECT 95.000 322.200 95.800 329.600 ;
        RECT 96.600 328.400 97.200 329.600 ;
        RECT 96.400 327.600 97.200 328.400 ;
        RECT 101.400 322.200 102.200 329.600 ;
        RECT 103.000 328.400 103.600 329.600 ;
        RECT 102.800 327.600 103.600 328.400 ;
        RECT 110.000 322.200 110.800 330.600 ;
        RECT 115.000 330.200 119.800 330.600 ;
        RECT 113.200 329.000 118.600 329.600 ;
        RECT 113.200 328.800 114.000 329.000 ;
        RECT 117.800 328.800 118.600 329.000 ;
        RECT 119.200 329.000 119.800 330.200 ;
        RECT 121.200 330.400 121.800 333.600 ;
        RECT 127.600 333.700 130.000 334.300 ;
        RECT 122.800 332.800 123.600 333.000 ;
        RECT 122.800 332.200 126.600 332.800 ;
        RECT 125.800 332.000 126.600 332.200 ;
        RECT 124.200 331.400 125.000 331.600 ;
        RECT 127.600 331.400 128.400 333.700 ;
        RECT 129.200 333.600 130.000 333.700 ;
        RECT 124.200 330.800 128.400 331.400 ;
        RECT 121.200 329.800 123.600 330.400 ;
        RECT 120.600 329.000 121.400 329.200 ;
        RECT 119.200 328.400 121.400 329.000 ;
        RECT 123.000 328.800 123.600 329.800 ;
        RECT 123.000 328.000 124.400 328.800 ;
        RECT 116.600 327.400 117.400 327.600 ;
        RECT 119.400 327.400 120.200 327.600 ;
        RECT 113.200 326.200 114.000 327.000 ;
        RECT 116.600 326.800 120.200 327.400 ;
        RECT 118.800 326.200 119.400 326.800 ;
        RECT 122.800 326.200 123.600 327.000 ;
        RECT 113.200 325.600 115.200 326.200 ;
        RECT 114.400 322.200 115.200 325.600 ;
        RECT 118.800 322.200 119.600 326.200 ;
        RECT 123.000 322.200 124.200 326.200 ;
        RECT 127.600 322.200 128.400 330.800 ;
        RECT 130.800 322.200 131.600 335.800 ;
        RECT 134.000 333.600 134.800 335.200 ;
        RECT 132.400 328.800 133.200 330.400 ;
        RECT 135.600 322.200 136.400 335.800 ;
        RECT 137.200 330.300 138.000 330.400 ;
        RECT 138.800 330.300 139.600 339.800 ;
        RECT 140.400 335.600 141.200 337.200 ;
        RECT 142.000 335.800 142.800 339.800 ;
        RECT 146.400 336.200 148.000 339.800 ;
        RECT 142.000 335.200 144.200 335.800 ;
        RECT 145.200 335.400 146.800 335.600 ;
        RECT 143.400 335.000 144.200 335.200 ;
        RECT 144.800 334.800 146.800 335.400 ;
        RECT 144.800 334.400 145.400 334.800 ;
        RECT 142.000 333.800 145.400 334.400 ;
        RECT 142.000 333.600 143.600 333.800 ;
        RECT 146.000 333.400 146.800 334.200 ;
        RECT 146.000 332.800 146.600 333.400 ;
        RECT 144.000 332.200 146.600 332.800 ;
        RECT 147.400 332.800 148.000 336.200 ;
        RECT 151.600 335.800 152.400 339.800 ;
        RECT 148.600 334.800 149.400 335.600 ;
        RECT 150.000 335.200 152.400 335.800 ;
        RECT 150.000 335.000 150.800 335.200 ;
        RECT 148.800 334.400 149.400 334.800 ;
        RECT 148.800 333.600 149.600 334.400 ;
        RECT 150.800 333.600 152.400 334.400 ;
        RECT 153.200 333.600 154.000 335.200 ;
        RECT 154.800 334.300 155.600 339.800 ;
        RECT 157.000 338.400 157.800 339.800 ;
        RECT 157.000 337.600 158.800 338.400 ;
        RECT 157.000 336.400 157.800 337.600 ;
        RECT 157.000 335.800 158.800 336.400 ;
        RECT 161.200 336.000 162.000 339.800 ;
        RECT 164.400 336.000 165.200 339.800 ;
        RECT 161.200 335.800 165.200 336.000 ;
        RECT 166.000 335.800 166.800 339.800 ;
        RECT 169.200 336.000 170.000 339.800 ;
        RECT 156.400 334.300 157.200 334.400 ;
        RECT 154.800 333.700 157.200 334.300 ;
        RECT 147.400 332.400 148.400 332.800 ;
        RECT 147.400 332.200 149.200 332.400 ;
        RECT 144.000 332.000 144.800 332.200 ;
        RECT 147.800 331.600 149.200 332.200 ;
        RECT 151.700 332.300 152.300 333.600 ;
        RECT 154.800 332.300 155.600 333.700 ;
        RECT 156.400 333.600 157.200 333.700 ;
        RECT 151.700 331.700 155.600 332.300 ;
        RECT 146.200 331.400 147.000 331.600 ;
        RECT 137.200 329.700 139.600 330.300 ;
        RECT 143.600 330.800 147.000 331.400 ;
        RECT 143.600 330.200 144.200 330.800 ;
        RECT 147.800 330.200 148.400 331.600 ;
        RECT 154.800 330.300 155.600 331.700 ;
        RECT 156.400 330.300 157.200 330.400 ;
        RECT 137.200 328.800 138.000 329.700 ;
        RECT 138.800 322.200 139.600 329.700 ;
        RECT 142.000 329.600 144.200 330.200 ;
        RECT 142.000 322.200 142.800 329.600 ;
        RECT 143.400 329.400 144.200 329.600 ;
        RECT 146.400 329.600 148.400 330.200 ;
        RECT 150.000 329.600 152.400 330.200 ;
        RECT 146.400 324.400 148.000 329.600 ;
        RECT 150.000 329.400 150.800 329.600 ;
        RECT 145.200 323.600 148.000 324.400 ;
        RECT 146.400 322.200 148.000 323.600 ;
        RECT 151.600 322.200 152.400 329.600 ;
        RECT 154.800 329.700 157.200 330.300 ;
        RECT 154.800 322.200 155.600 329.700 ;
        RECT 156.400 328.800 157.200 329.700 ;
        RECT 158.000 322.200 158.800 335.800 ;
        RECT 161.400 335.400 165.000 335.800 ;
        RECT 159.600 333.600 160.400 335.200 ;
        RECT 162.000 334.400 162.800 334.800 ;
        RECT 166.000 334.400 166.600 335.800 ;
        RECT 169.000 335.200 170.000 336.000 ;
        RECT 161.200 333.800 162.800 334.400 ;
        RECT 161.200 333.600 162.000 333.800 ;
        RECT 164.200 333.600 166.800 334.400 ;
        RECT 162.800 331.600 163.600 333.200 ;
        RECT 164.200 330.200 164.800 333.600 ;
        RECT 166.000 332.300 166.800 332.400 ;
        RECT 169.000 332.300 169.800 335.200 ;
        RECT 170.800 334.600 171.600 339.800 ;
        RECT 177.200 336.600 178.000 339.800 ;
        RECT 178.800 337.000 179.600 339.800 ;
        RECT 180.400 337.000 181.200 339.800 ;
        RECT 182.000 337.000 182.800 339.800 ;
        RECT 183.600 337.000 184.400 339.800 ;
        RECT 186.800 337.000 187.600 339.800 ;
        RECT 190.000 337.000 190.800 339.800 ;
        RECT 191.600 337.000 192.400 339.800 ;
        RECT 193.200 337.000 194.000 339.800 ;
        RECT 175.600 335.800 178.000 336.600 ;
        RECT 194.800 336.600 195.600 339.800 ;
        RECT 175.600 335.200 176.400 335.800 ;
        RECT 166.000 331.700 169.800 332.300 ;
        RECT 166.000 331.600 166.800 331.700 ;
        RECT 169.000 330.800 169.800 331.700 ;
        RECT 170.400 334.000 171.600 334.600 ;
        RECT 174.600 334.600 176.400 335.200 ;
        RECT 180.400 335.600 181.400 336.400 ;
        RECT 184.400 335.600 186.000 336.400 ;
        RECT 186.800 335.800 191.400 336.400 ;
        RECT 194.800 335.800 197.400 336.600 ;
        RECT 186.800 335.600 187.600 335.800 ;
        RECT 170.400 332.000 171.000 334.000 ;
        RECT 174.600 333.400 175.400 334.600 ;
        RECT 171.600 332.600 175.400 333.400 ;
        RECT 180.400 332.800 181.200 335.600 ;
        RECT 186.800 334.800 187.600 335.000 ;
        RECT 183.200 334.200 187.600 334.800 ;
        RECT 183.200 334.000 184.000 334.200 ;
        RECT 188.400 333.600 189.200 335.200 ;
        RECT 190.600 333.400 191.400 335.800 ;
        RECT 196.600 335.200 197.400 335.800 ;
        RECT 196.600 334.400 199.600 335.200 ;
        RECT 201.200 333.800 202.000 339.800 ;
        RECT 204.400 336.400 205.200 339.800 ;
        RECT 183.600 332.600 186.800 333.400 ;
        RECT 190.600 332.600 192.600 333.400 ;
        RECT 193.200 333.000 202.000 333.800 ;
        RECT 177.200 332.000 178.000 332.600 ;
        RECT 194.800 332.000 195.600 332.400 ;
        RECT 198.000 332.000 198.800 332.400 ;
        RECT 199.800 332.000 200.600 332.200 ;
        RECT 170.400 331.400 171.200 332.000 ;
        RECT 177.200 331.400 200.600 332.000 ;
        RECT 166.000 330.300 166.800 330.400 ;
        RECT 167.600 330.300 168.400 330.400 ;
        RECT 166.000 330.200 168.400 330.300 ;
        RECT 163.800 329.600 164.800 330.200 ;
        RECT 165.400 329.700 168.400 330.200 ;
        RECT 169.000 330.000 170.000 330.800 ;
        RECT 165.400 329.600 166.800 329.700 ;
        RECT 167.600 329.600 168.400 329.700 ;
        RECT 163.800 324.400 164.600 329.600 ;
        RECT 165.400 328.400 166.000 329.600 ;
        RECT 165.200 327.600 166.000 328.400 ;
        RECT 162.800 323.600 164.600 324.400 ;
        RECT 163.800 322.200 164.600 323.600 ;
        RECT 169.200 322.200 170.000 330.000 ;
        RECT 170.600 329.600 171.200 331.400 ;
        RECT 170.600 329.000 179.600 329.600 ;
        RECT 170.600 327.400 171.200 329.000 ;
        RECT 178.800 328.800 179.600 329.000 ;
        RECT 182.000 329.000 190.600 329.600 ;
        RECT 182.000 328.800 182.800 329.000 ;
        RECT 173.800 327.600 176.400 328.400 ;
        RECT 170.600 326.800 173.200 327.400 ;
        RECT 172.400 322.200 173.200 326.800 ;
        RECT 175.600 322.200 176.400 327.600 ;
        RECT 177.000 326.800 181.200 327.600 ;
        RECT 178.800 322.200 179.600 325.000 ;
        RECT 180.400 322.200 181.200 325.000 ;
        RECT 182.000 322.200 182.800 325.000 ;
        RECT 183.600 322.200 184.400 328.400 ;
        RECT 186.800 327.600 189.400 328.400 ;
        RECT 190.000 328.200 190.600 329.000 ;
        RECT 191.600 329.400 192.400 329.600 ;
        RECT 191.600 329.000 197.000 329.400 ;
        RECT 191.600 328.800 197.800 329.000 ;
        RECT 196.400 328.200 197.800 328.800 ;
        RECT 190.000 327.600 195.800 328.200 ;
        RECT 198.800 328.000 200.400 328.800 ;
        RECT 198.800 327.600 199.400 328.000 ;
        RECT 186.800 322.200 187.600 327.000 ;
        RECT 190.000 322.200 190.800 327.000 ;
        RECT 195.200 326.800 199.400 327.600 ;
        RECT 201.200 327.400 202.000 333.000 ;
        RECT 204.200 335.800 205.200 336.400 ;
        RECT 204.200 334.400 204.800 335.800 ;
        RECT 207.600 335.200 208.400 339.800 ;
        RECT 205.800 334.600 208.400 335.200 ;
        RECT 209.200 335.200 210.000 339.800 ;
        RECT 212.400 336.400 213.200 339.800 ;
        RECT 212.400 335.800 213.400 336.400 ;
        RECT 215.600 335.800 216.400 339.800 ;
        RECT 217.200 336.000 218.000 339.800 ;
        RECT 220.400 336.000 221.200 339.800 ;
        RECT 217.200 335.800 221.200 336.000 ;
        RECT 209.200 334.600 211.800 335.200 ;
        RECT 204.200 333.600 205.200 334.400 ;
        RECT 204.200 330.200 204.800 333.600 ;
        RECT 205.800 333.000 206.400 334.600 ;
        RECT 205.400 332.200 206.400 333.000 ;
        RECT 209.400 332.400 210.200 333.200 ;
        RECT 205.800 330.200 206.400 332.200 ;
        RECT 209.200 331.600 210.200 332.400 ;
        RECT 211.200 333.000 211.800 334.600 ;
        RECT 212.800 334.400 213.400 335.800 ;
        RECT 215.800 334.400 216.400 335.800 ;
        RECT 217.400 335.400 221.000 335.800 ;
        RECT 219.600 334.400 220.400 334.800 ;
        RECT 212.400 333.600 213.400 334.400 ;
        RECT 215.600 333.600 218.200 334.400 ;
        RECT 219.600 333.800 221.200 334.400 ;
        RECT 220.400 333.600 221.200 333.800 ;
        RECT 211.200 332.200 212.200 333.000 ;
        RECT 211.200 330.200 211.800 332.200 ;
        RECT 212.800 330.400 213.400 333.600 ;
        RECT 204.200 329.200 205.200 330.200 ;
        RECT 205.800 329.600 208.400 330.200 ;
        RECT 200.000 326.800 202.000 327.400 ;
        RECT 191.600 322.200 192.400 325.000 ;
        RECT 193.200 322.200 194.000 325.000 ;
        RECT 196.400 322.200 197.200 326.800 ;
        RECT 200.000 326.200 200.600 326.800 ;
        RECT 199.600 325.600 200.600 326.200 ;
        RECT 199.600 322.200 200.400 325.600 ;
        RECT 204.400 322.200 205.200 329.200 ;
        RECT 207.600 322.200 208.400 329.600 ;
        RECT 209.200 329.600 211.800 330.200 ;
        RECT 209.200 322.200 210.000 329.600 ;
        RECT 212.400 329.200 213.400 330.400 ;
        RECT 215.600 330.200 216.400 330.400 ;
        RECT 217.600 330.200 218.200 333.600 ;
        RECT 218.800 332.300 219.600 333.200 ;
        RECT 222.000 332.300 222.800 339.800 ;
        RECT 226.800 337.600 227.600 339.800 ;
        RECT 223.600 335.600 224.400 337.200 ;
        RECT 226.800 334.400 227.400 337.600 ;
        RECT 228.400 336.300 229.200 337.200 ;
        RECT 230.000 336.300 230.800 336.400 ;
        RECT 228.400 335.700 230.800 336.300 ;
        RECT 231.600 336.000 232.400 339.800 ;
        RECT 228.400 335.600 229.200 335.700 ;
        RECT 230.000 335.600 230.800 335.700 ;
        RECT 231.400 335.200 232.400 336.000 ;
        RECT 226.800 333.600 227.600 334.400 ;
        RECT 228.400 334.300 229.200 334.400 ;
        RECT 231.400 334.300 232.200 335.200 ;
        RECT 233.200 334.600 234.000 339.800 ;
        RECT 239.600 336.600 240.400 339.800 ;
        RECT 241.200 337.000 242.000 339.800 ;
        RECT 242.800 337.000 243.600 339.800 ;
        RECT 244.400 337.000 245.200 339.800 ;
        RECT 246.000 337.000 246.800 339.800 ;
        RECT 249.200 337.000 250.000 339.800 ;
        RECT 252.400 337.000 253.200 339.800 ;
        RECT 254.000 337.000 254.800 339.800 ;
        RECT 255.600 337.000 256.400 339.800 ;
        RECT 238.000 335.800 240.400 336.600 ;
        RECT 257.200 336.600 258.000 339.800 ;
        RECT 238.000 335.200 238.800 335.800 ;
        RECT 228.400 333.700 232.200 334.300 ;
        RECT 228.400 333.600 229.200 333.700 ;
        RECT 218.800 331.700 222.800 332.300 ;
        RECT 218.800 331.600 219.600 331.700 ;
        RECT 215.600 329.600 217.000 330.200 ;
        RECT 217.600 329.600 218.600 330.200 ;
        RECT 212.400 322.200 213.200 329.200 ;
        RECT 216.400 328.400 217.000 329.600 ;
        RECT 216.400 327.600 217.200 328.400 ;
        RECT 217.800 322.200 218.600 329.600 ;
        RECT 222.000 322.200 222.800 331.700 ;
        RECT 225.200 330.800 226.000 332.400 ;
        RECT 226.800 330.200 227.400 333.600 ;
        RECT 231.400 330.800 232.200 333.700 ;
        RECT 232.800 334.000 234.000 334.600 ;
        RECT 237.000 334.600 238.800 335.200 ;
        RECT 242.800 335.600 243.800 336.400 ;
        RECT 246.800 335.600 248.400 336.400 ;
        RECT 249.200 335.800 253.800 336.400 ;
        RECT 257.200 335.800 259.800 336.600 ;
        RECT 249.200 335.600 250.000 335.800 ;
        RECT 232.800 332.000 233.400 334.000 ;
        RECT 237.000 333.400 237.800 334.600 ;
        RECT 234.000 332.600 237.800 333.400 ;
        RECT 242.800 332.800 243.600 335.600 ;
        RECT 249.200 334.800 250.000 335.000 ;
        RECT 245.600 334.200 250.000 334.800 ;
        RECT 245.600 334.000 246.400 334.200 ;
        RECT 250.800 333.600 251.600 335.200 ;
        RECT 253.000 333.400 253.800 335.800 ;
        RECT 259.000 335.200 259.800 335.800 ;
        RECT 259.000 334.400 262.000 335.200 ;
        RECT 263.600 333.800 264.400 339.800 ;
        RECT 246.000 332.600 249.200 333.400 ;
        RECT 253.000 332.600 255.000 333.400 ;
        RECT 255.600 333.000 264.400 333.800 ;
        RECT 239.600 332.000 240.400 332.600 ;
        RECT 257.200 332.000 258.000 332.400 ;
        RECT 262.200 332.000 263.000 332.200 ;
        RECT 232.800 331.400 233.600 332.000 ;
        RECT 239.600 331.400 263.000 332.000 ;
        RECT 225.800 329.400 227.600 330.200 ;
        RECT 231.400 330.000 232.400 330.800 ;
        RECT 225.800 322.200 226.600 329.400 ;
        RECT 231.600 322.200 232.400 330.000 ;
        RECT 233.000 329.600 233.600 331.400 ;
        RECT 233.000 329.000 242.000 329.600 ;
        RECT 233.000 327.400 233.600 329.000 ;
        RECT 241.200 328.800 242.000 329.000 ;
        RECT 244.400 329.000 253.000 329.600 ;
        RECT 244.400 328.800 245.200 329.000 ;
        RECT 236.200 327.600 238.800 328.400 ;
        RECT 233.000 326.800 235.600 327.400 ;
        RECT 234.800 322.200 235.600 326.800 ;
        RECT 238.000 322.200 238.800 327.600 ;
        RECT 239.400 326.800 243.600 327.600 ;
        RECT 241.200 322.200 242.000 325.000 ;
        RECT 242.800 322.200 243.600 325.000 ;
        RECT 244.400 322.200 245.200 325.000 ;
        RECT 246.000 322.200 246.800 328.400 ;
        RECT 249.200 327.600 251.800 328.400 ;
        RECT 252.400 328.200 253.000 329.000 ;
        RECT 254.000 329.400 254.800 329.600 ;
        RECT 254.000 329.000 259.400 329.400 ;
        RECT 254.000 328.800 260.200 329.000 ;
        RECT 258.800 328.200 260.200 328.800 ;
        RECT 252.400 327.600 258.200 328.200 ;
        RECT 261.200 328.000 262.800 328.800 ;
        RECT 261.200 327.600 261.800 328.000 ;
        RECT 249.200 322.200 250.000 327.000 ;
        RECT 252.400 322.200 253.200 327.000 ;
        RECT 257.600 326.800 261.800 327.600 ;
        RECT 263.600 327.400 264.400 333.000 ;
        RECT 262.400 326.800 264.400 327.400 ;
        RECT 270.000 333.800 270.800 339.800 ;
        RECT 276.400 336.600 277.200 339.800 ;
        RECT 278.000 337.000 278.800 339.800 ;
        RECT 279.600 337.000 280.400 339.800 ;
        RECT 281.200 337.000 282.000 339.800 ;
        RECT 284.400 337.000 285.200 339.800 ;
        RECT 287.600 337.000 288.400 339.800 ;
        RECT 289.200 337.000 290.000 339.800 ;
        RECT 290.800 337.000 291.600 339.800 ;
        RECT 292.400 337.000 293.200 339.800 ;
        RECT 274.600 335.800 277.200 336.600 ;
        RECT 294.000 336.600 294.800 339.800 ;
        RECT 280.600 335.800 285.200 336.400 ;
        RECT 274.600 335.200 275.400 335.800 ;
        RECT 272.400 334.400 275.400 335.200 ;
        RECT 270.000 333.000 278.800 333.800 ;
        RECT 280.600 333.400 281.400 335.800 ;
        RECT 284.400 335.600 285.200 335.800 ;
        RECT 286.000 335.600 287.600 336.400 ;
        RECT 290.600 335.600 291.600 336.400 ;
        RECT 294.000 335.800 296.400 336.600 ;
        RECT 282.800 333.600 283.600 335.200 ;
        RECT 284.400 334.800 285.200 335.000 ;
        RECT 284.400 334.200 288.800 334.800 ;
        RECT 288.000 334.000 288.800 334.200 ;
        RECT 270.000 327.400 270.800 333.000 ;
        RECT 279.400 332.600 281.400 333.400 ;
        RECT 285.200 332.600 288.400 333.400 ;
        RECT 290.800 332.800 291.600 335.600 ;
        RECT 295.600 335.200 296.400 335.800 ;
        RECT 295.600 334.600 297.400 335.200 ;
        RECT 296.600 333.400 297.400 334.600 ;
        RECT 300.400 334.600 301.200 339.800 ;
        RECT 302.000 336.000 302.800 339.800 ;
        RECT 302.000 335.200 303.000 336.000 ;
        RECT 305.200 335.800 306.000 339.800 ;
        RECT 306.800 336.000 307.600 339.800 ;
        RECT 310.000 336.000 310.800 339.800 ;
        RECT 306.800 335.800 310.800 336.000 ;
        RECT 311.600 335.800 312.400 339.800 ;
        RECT 313.200 336.000 314.000 339.800 ;
        RECT 316.400 336.000 317.200 339.800 ;
        RECT 313.200 335.800 317.200 336.000 ;
        RECT 318.600 338.400 319.400 339.800 ;
        RECT 318.600 337.600 320.400 338.400 ;
        RECT 318.600 336.400 319.400 337.600 ;
        RECT 318.600 335.800 320.400 336.400 ;
        RECT 325.400 335.800 327.000 339.800 ;
        RECT 333.400 338.400 335.000 339.800 ;
        RECT 332.400 337.600 335.000 338.400 ;
        RECT 333.400 335.800 335.000 337.600 ;
        RECT 341.400 335.800 343.000 339.800 ;
        RECT 349.400 338.400 351.000 339.800 ;
        RECT 348.400 337.600 351.000 338.400 ;
        RECT 349.400 335.800 351.000 337.600 ;
        RECT 357.800 336.400 359.400 339.800 ;
        RECT 365.400 338.400 366.200 339.800 ;
        RECT 364.400 337.600 366.200 338.400 ;
        RECT 365.400 336.400 366.200 337.600 ;
        RECT 357.800 335.800 360.400 336.400 ;
        RECT 300.400 334.000 301.600 334.600 ;
        RECT 296.600 332.600 300.400 333.400 ;
        RECT 271.400 332.000 272.200 332.200 ;
        RECT 276.400 332.000 277.200 332.400 ;
        RECT 294.000 332.000 294.800 332.600 ;
        RECT 301.000 332.000 301.600 334.000 ;
        RECT 271.400 331.400 294.800 332.000 ;
        RECT 300.800 331.400 301.600 332.000 ;
        RECT 300.800 329.600 301.400 331.400 ;
        RECT 302.200 330.800 303.000 335.200 ;
        RECT 305.400 334.400 306.000 335.800 ;
        RECT 307.000 335.400 310.600 335.800 ;
        RECT 309.200 334.400 310.000 334.800 ;
        RECT 311.800 334.400 312.400 335.800 ;
        RECT 313.400 335.400 317.000 335.800 ;
        RECT 315.600 334.400 316.400 334.800 ;
        RECT 303.600 334.300 304.400 334.400 ;
        RECT 305.200 334.300 307.800 334.400 ;
        RECT 303.600 333.700 307.800 334.300 ;
        RECT 309.200 334.300 310.800 334.400 ;
        RECT 311.600 334.300 314.200 334.400 ;
        RECT 309.200 333.800 314.200 334.300 ;
        RECT 315.600 333.800 317.200 334.400 ;
        RECT 303.600 333.600 304.400 333.700 ;
        RECT 305.200 333.600 307.800 333.700 ;
        RECT 310.000 333.700 314.200 333.800 ;
        RECT 310.000 333.600 310.800 333.700 ;
        RECT 311.600 333.600 314.200 333.700 ;
        RECT 316.400 333.600 317.200 333.800 ;
        RECT 279.600 329.400 280.400 329.600 ;
        RECT 275.000 329.000 280.400 329.400 ;
        RECT 274.200 328.800 280.400 329.000 ;
        RECT 281.400 329.000 290.000 329.600 ;
        RECT 271.600 328.000 273.200 328.800 ;
        RECT 274.200 328.200 275.600 328.800 ;
        RECT 281.400 328.200 282.000 329.000 ;
        RECT 289.200 328.800 290.000 329.000 ;
        RECT 292.400 329.000 301.400 329.600 ;
        RECT 292.400 328.800 293.200 329.000 ;
        RECT 272.600 327.600 273.200 328.000 ;
        RECT 276.200 327.600 282.000 328.200 ;
        RECT 282.600 327.600 285.200 328.400 ;
        RECT 270.000 326.800 272.000 327.400 ;
        RECT 272.600 326.800 276.800 327.600 ;
        RECT 254.000 322.200 254.800 325.000 ;
        RECT 255.600 322.200 256.400 325.000 ;
        RECT 258.800 322.200 259.600 326.800 ;
        RECT 262.400 326.200 263.000 326.800 ;
        RECT 262.000 325.600 263.000 326.200 ;
        RECT 271.400 326.200 272.000 326.800 ;
        RECT 271.400 325.600 272.400 326.200 ;
        RECT 262.000 322.200 262.800 325.600 ;
        RECT 271.600 322.200 272.400 325.600 ;
        RECT 274.800 322.200 275.600 326.800 ;
        RECT 278.000 322.200 278.800 325.000 ;
        RECT 279.600 322.200 280.400 325.000 ;
        RECT 281.200 322.200 282.000 327.000 ;
        RECT 284.400 322.200 285.200 327.000 ;
        RECT 287.600 322.200 288.400 328.400 ;
        RECT 295.600 327.600 298.200 328.400 ;
        RECT 290.800 326.800 295.000 327.600 ;
        RECT 289.200 322.200 290.000 325.000 ;
        RECT 290.800 322.200 291.600 325.000 ;
        RECT 292.400 322.200 293.200 325.000 ;
        RECT 295.600 322.200 296.400 327.600 ;
        RECT 300.800 327.400 301.400 329.000 ;
        RECT 298.800 326.800 301.400 327.400 ;
        RECT 302.000 330.000 303.000 330.800 ;
        RECT 303.600 330.300 304.400 330.400 ;
        RECT 305.200 330.300 306.000 330.400 ;
        RECT 303.600 330.200 306.000 330.300 ;
        RECT 307.200 330.200 307.800 333.600 ;
        RECT 308.400 331.600 309.200 333.200 ;
        RECT 311.600 330.200 312.400 330.400 ;
        RECT 313.600 330.200 314.200 333.600 ;
        RECT 314.800 331.600 315.600 333.200 ;
        RECT 298.800 322.200 299.600 326.800 ;
        RECT 302.000 322.200 302.800 330.000 ;
        RECT 303.600 329.700 306.600 330.200 ;
        RECT 303.600 329.600 304.400 329.700 ;
        RECT 305.200 329.600 306.600 329.700 ;
        RECT 307.200 329.600 308.200 330.200 ;
        RECT 311.600 329.600 313.000 330.200 ;
        RECT 313.600 329.600 314.600 330.200 ;
        RECT 306.000 328.400 306.600 329.600 ;
        RECT 306.000 327.600 306.800 328.400 ;
        RECT 307.400 322.200 308.200 329.600 ;
        RECT 312.400 328.400 313.000 329.600 ;
        RECT 312.400 327.600 313.200 328.400 ;
        RECT 313.800 322.200 314.600 329.600 ;
        RECT 318.000 328.800 318.800 330.400 ;
        RECT 319.600 322.200 320.400 335.800 ;
        RECT 321.200 333.600 322.000 335.200 ;
        RECT 324.400 333.600 325.200 334.400 ;
        RECT 324.600 333.200 325.200 333.600 ;
        RECT 324.600 332.400 325.400 333.200 ;
        RECT 326.000 332.400 326.600 335.800 ;
        RECT 327.600 332.800 328.400 334.400 ;
        RECT 332.400 333.600 333.200 334.400 ;
        RECT 332.600 333.200 333.200 333.600 ;
        RECT 332.600 332.400 333.400 333.200 ;
        RECT 334.000 332.400 334.600 335.800 ;
        RECT 335.600 334.300 336.400 334.400 ;
        RECT 340.400 334.300 341.200 334.400 ;
        RECT 335.600 333.700 341.200 334.300 ;
        RECT 335.600 332.800 336.400 333.700 ;
        RECT 340.400 333.600 341.200 333.700 ;
        RECT 340.600 333.200 341.200 333.600 ;
        RECT 340.600 332.400 341.400 333.200 ;
        RECT 342.000 332.400 342.600 335.800 ;
        RECT 343.600 332.800 344.400 334.400 ;
        RECT 348.400 333.600 349.200 334.400 ;
        RECT 348.600 333.200 349.200 333.600 ;
        RECT 348.600 332.400 349.400 333.200 ;
        RECT 350.000 332.400 350.600 335.800 ;
        RECT 358.200 335.600 360.400 335.800 ;
        RECT 364.400 335.800 366.200 336.400 ;
        RECT 370.200 335.800 371.800 339.800 ;
        RECT 378.200 338.400 379.000 339.800 ;
        RECT 381.000 338.400 381.800 339.800 ;
        RECT 378.200 337.600 379.600 338.400 ;
        RECT 380.400 337.600 381.800 338.400 ;
        RECT 378.200 336.400 379.000 337.600 ;
        RECT 377.200 335.800 379.000 336.400 ;
        RECT 381.000 336.400 381.800 337.600 ;
        RECT 381.000 335.800 382.800 336.400 ;
        RECT 387.800 335.800 389.400 339.800 ;
        RECT 393.800 336.400 394.600 339.800 ;
        RECT 393.800 335.800 395.600 336.400 ;
        RECT 401.000 335.800 402.600 339.800 ;
        RECT 406.000 335.800 406.800 339.800 ;
        RECT 407.600 336.000 408.400 339.800 ;
        RECT 410.800 336.000 411.600 339.800 ;
        RECT 415.000 338.400 415.800 339.800 ;
        RECT 414.000 337.600 415.800 338.400 ;
        RECT 415.000 336.400 415.800 337.600 ;
        RECT 407.600 335.800 411.600 336.000 ;
        RECT 414.000 335.800 415.800 336.400 ;
        RECT 422.000 336.000 422.800 339.800 ;
        RECT 425.200 336.000 426.000 339.800 ;
        RECT 422.000 335.800 426.000 336.000 ;
        RECT 351.600 332.800 352.400 334.400 ;
        RECT 356.400 332.800 357.200 334.400 ;
        RECT 358.200 332.400 358.800 335.600 ;
        RECT 359.600 333.600 360.400 334.400 ;
        RECT 361.200 334.300 362.000 334.400 ;
        RECT 362.800 334.300 363.600 335.200 ;
        RECT 361.200 333.700 363.600 334.300 ;
        RECT 361.200 333.600 362.000 333.700 ;
        RECT 362.800 333.600 363.600 333.700 ;
        RECT 359.600 333.200 360.200 333.600 ;
        RECT 359.400 332.400 360.200 333.200 ;
        RECT 322.800 330.800 323.600 332.400 ;
        RECT 326.000 331.600 326.800 332.400 ;
        RECT 329.200 332.200 330.000 332.400 ;
        RECT 328.400 331.600 330.000 332.200 ;
        RECT 326.000 331.400 326.600 331.600 ;
        RECT 324.600 330.800 326.600 331.400 ;
        RECT 328.400 331.200 329.200 331.600 ;
        RECT 330.800 330.800 331.600 332.400 ;
        RECT 334.000 331.600 334.800 332.400 ;
        RECT 337.200 332.200 338.000 332.400 ;
        RECT 336.400 331.600 338.000 332.200 ;
        RECT 334.000 331.400 334.600 331.600 ;
        RECT 332.600 330.800 334.600 331.400 ;
        RECT 336.400 331.200 337.200 331.600 ;
        RECT 338.800 330.800 339.600 332.400 ;
        RECT 342.000 331.600 342.800 332.400 ;
        RECT 345.200 332.200 346.000 332.400 ;
        RECT 344.400 331.600 346.000 332.200 ;
        RECT 342.000 331.400 342.600 331.600 ;
        RECT 340.600 330.800 342.600 331.400 ;
        RECT 344.400 331.200 345.200 331.600 ;
        RECT 346.800 330.800 347.600 332.400 ;
        RECT 350.000 331.600 350.800 332.400 ;
        RECT 353.200 332.200 354.000 332.400 ;
        RECT 352.400 331.600 354.000 332.200 ;
        RECT 354.800 332.200 355.600 332.400 ;
        RECT 354.800 331.600 356.400 332.200 ;
        RECT 358.000 331.600 358.800 332.400 ;
        RECT 350.000 331.400 350.600 331.600 ;
        RECT 348.600 330.800 350.600 331.400 ;
        RECT 352.400 331.200 353.200 331.600 ;
        RECT 355.600 331.200 356.400 331.600 ;
        RECT 358.200 331.400 358.800 331.600 ;
        RECT 358.200 330.800 360.200 331.400 ;
        RECT 361.200 330.800 362.000 332.400 ;
        RECT 324.600 330.200 325.200 330.800 ;
        RECT 332.600 330.200 333.200 330.800 ;
        RECT 340.600 330.200 341.200 330.800 ;
        RECT 348.600 330.200 349.200 330.800 ;
        RECT 359.600 330.200 360.200 330.800 ;
        RECT 322.800 322.800 323.600 330.200 ;
        RECT 324.400 323.400 325.200 330.200 ;
        RECT 326.000 329.600 330.000 330.200 ;
        RECT 326.000 322.800 326.800 329.600 ;
        RECT 322.800 322.200 326.800 322.800 ;
        RECT 329.200 322.200 330.000 329.600 ;
        RECT 330.800 322.800 331.600 330.200 ;
        RECT 332.400 323.400 333.200 330.200 ;
        RECT 334.000 329.600 338.000 330.200 ;
        RECT 334.000 322.800 334.800 329.600 ;
        RECT 330.800 322.200 334.800 322.800 ;
        RECT 337.200 322.200 338.000 329.600 ;
        RECT 338.800 322.800 339.600 330.200 ;
        RECT 340.400 323.400 341.200 330.200 ;
        RECT 342.000 329.600 346.000 330.200 ;
        RECT 342.000 322.800 342.800 329.600 ;
        RECT 338.800 322.200 342.800 322.800 ;
        RECT 345.200 322.200 346.000 329.600 ;
        RECT 346.800 322.800 347.600 330.200 ;
        RECT 348.400 323.400 349.200 330.200 ;
        RECT 350.000 329.600 354.000 330.200 ;
        RECT 350.000 322.800 350.800 329.600 ;
        RECT 346.800 322.200 350.800 322.800 ;
        RECT 353.200 322.200 354.000 329.600 ;
        RECT 354.800 329.600 358.800 330.200 ;
        RECT 354.800 322.200 355.600 329.600 ;
        RECT 358.000 322.800 358.800 329.600 ;
        RECT 359.600 323.400 360.400 330.200 ;
        RECT 361.200 322.800 362.000 330.200 ;
        RECT 358.000 322.200 362.000 322.800 ;
        RECT 364.400 322.200 365.200 335.800 ;
        RECT 367.600 334.300 368.400 334.400 ;
        RECT 369.200 334.300 370.000 334.400 ;
        RECT 367.600 333.700 370.000 334.300 ;
        RECT 367.600 333.600 368.400 333.700 ;
        RECT 369.200 333.600 370.000 333.700 ;
        RECT 369.400 333.200 370.000 333.600 ;
        RECT 369.400 332.400 370.200 333.200 ;
        RECT 370.800 332.400 371.400 335.800 ;
        RECT 372.400 332.800 373.200 334.400 ;
        RECT 375.600 333.600 376.400 335.200 ;
        RECT 367.600 330.800 368.400 332.400 ;
        RECT 370.800 331.600 371.600 332.400 ;
        RECT 374.000 332.200 374.800 332.400 ;
        RECT 373.200 331.600 374.800 332.200 ;
        RECT 370.800 331.400 371.400 331.600 ;
        RECT 369.400 330.800 371.400 331.400 ;
        RECT 373.200 331.200 374.000 331.600 ;
        RECT 366.000 328.800 366.800 330.400 ;
        RECT 369.400 330.200 370.000 330.800 ;
        RECT 367.600 322.800 368.400 330.200 ;
        RECT 369.200 323.400 370.000 330.200 ;
        RECT 370.800 329.600 374.800 330.200 ;
        RECT 370.800 322.800 371.600 329.600 ;
        RECT 367.600 322.200 371.600 322.800 ;
        RECT 374.000 322.200 374.800 329.600 ;
        RECT 377.200 322.200 378.000 335.800 ;
        RECT 378.800 328.800 379.600 330.400 ;
        RECT 380.400 328.800 381.200 330.400 ;
        RECT 382.000 322.200 382.800 335.800 ;
        RECT 383.600 333.600 384.400 335.200 ;
        RECT 386.800 333.600 387.600 334.400 ;
        RECT 383.700 332.300 384.300 333.600 ;
        RECT 387.000 333.200 387.600 333.600 ;
        RECT 387.000 332.400 387.800 333.200 ;
        RECT 388.400 332.400 389.000 335.800 ;
        RECT 390.000 332.800 390.800 334.400 ;
        RECT 391.600 334.300 392.400 334.400 ;
        RECT 394.800 334.300 395.600 335.800 ;
        RECT 391.600 333.700 395.600 334.300 ;
        RECT 391.600 333.600 392.400 333.700 ;
        RECT 385.200 332.300 386.000 332.400 ;
        RECT 383.700 331.700 386.000 332.300 ;
        RECT 385.200 330.800 386.000 331.700 ;
        RECT 388.400 331.600 389.200 332.400 ;
        RECT 391.600 332.200 392.400 332.400 ;
        RECT 390.800 331.600 392.400 332.200 ;
        RECT 388.400 331.400 389.000 331.600 ;
        RECT 387.000 330.800 389.000 331.400 ;
        RECT 390.800 331.200 391.600 331.600 ;
        RECT 387.000 330.200 387.600 330.800 ;
        RECT 385.200 322.800 386.000 330.200 ;
        RECT 386.800 323.400 387.600 330.200 ;
        RECT 388.400 329.600 392.400 330.200 ;
        RECT 388.400 322.800 389.200 329.600 ;
        RECT 385.200 322.200 389.200 322.800 ;
        RECT 391.600 322.200 392.400 329.600 ;
        RECT 393.200 328.800 394.000 330.400 ;
        RECT 394.800 322.200 395.600 333.700 ;
        RECT 396.400 333.600 397.200 335.200 ;
        RECT 401.400 334.400 402.000 335.800 ;
        RECT 406.200 334.400 406.800 335.800 ;
        RECT 407.800 335.400 411.400 335.800 ;
        RECT 410.000 334.400 410.800 334.800 ;
        RECT 399.600 332.800 400.400 334.400 ;
        RECT 401.200 333.600 402.000 334.400 ;
        RECT 401.400 332.400 402.000 333.600 ;
        RECT 402.800 333.600 403.600 334.400 ;
        RECT 406.000 333.600 408.600 334.400 ;
        RECT 410.000 333.800 411.600 334.400 ;
        RECT 410.800 333.600 411.600 333.800 ;
        RECT 412.400 333.600 413.200 335.200 ;
        RECT 402.800 333.200 403.400 333.600 ;
        RECT 402.600 332.400 403.400 333.200 ;
        RECT 398.000 332.200 398.800 332.400 ;
        RECT 398.000 331.600 399.600 332.200 ;
        RECT 401.200 331.600 402.000 332.400 ;
        RECT 398.800 331.200 399.600 331.600 ;
        RECT 401.400 331.400 402.000 331.600 ;
        RECT 401.400 330.800 403.400 331.400 ;
        RECT 404.400 330.800 405.200 332.400 ;
        RECT 402.800 330.200 403.400 330.800 ;
        RECT 406.000 330.200 406.800 330.400 ;
        RECT 408.000 330.200 408.600 333.600 ;
        RECT 409.200 331.600 410.000 333.200 ;
        RECT 398.000 329.600 402.000 330.200 ;
        RECT 398.000 322.200 398.800 329.600 ;
        RECT 401.200 322.800 402.000 329.600 ;
        RECT 402.800 323.400 403.600 330.200 ;
        RECT 404.400 322.800 405.200 330.200 ;
        RECT 406.000 329.600 407.400 330.200 ;
        RECT 408.000 329.600 409.000 330.200 ;
        RECT 406.800 328.400 407.400 329.600 ;
        RECT 406.800 327.600 407.600 328.400 ;
        RECT 401.200 322.200 405.200 322.800 ;
        RECT 408.200 322.200 409.000 329.600 ;
        RECT 414.000 322.200 414.800 335.800 ;
        RECT 422.200 335.400 425.800 335.800 ;
        RECT 426.800 335.600 427.600 339.800 ;
        RECT 428.400 336.000 429.200 339.800 ;
        RECT 431.600 336.000 432.400 339.800 ;
        RECT 428.400 335.800 432.400 336.000 ;
        RECT 433.200 335.800 434.000 339.800 ;
        RECT 436.400 336.000 437.200 339.800 ;
        RECT 422.800 334.400 423.600 334.800 ;
        RECT 426.800 334.400 427.400 335.600 ;
        RECT 428.600 335.400 432.200 335.800 ;
        RECT 429.200 334.400 430.000 334.800 ;
        RECT 433.200 334.400 433.800 335.800 ;
        RECT 436.200 335.200 437.200 336.000 ;
        RECT 422.000 333.800 423.600 334.400 ;
        RECT 422.000 333.600 422.800 333.800 ;
        RECT 425.000 333.600 427.600 334.400 ;
        RECT 428.400 333.800 430.000 334.400 ;
        RECT 431.400 334.300 434.000 334.400 ;
        RECT 434.800 334.300 435.600 334.400 ;
        RECT 428.400 333.600 429.200 333.800 ;
        RECT 431.400 333.700 435.600 334.300 ;
        RECT 431.400 333.600 434.000 333.700 ;
        RECT 434.800 333.600 435.600 333.700 ;
        RECT 423.600 331.600 424.400 333.200 ;
        RECT 415.600 328.800 416.400 330.400 ;
        RECT 425.000 330.200 425.600 333.600 ;
        RECT 430.000 331.600 430.800 333.200 ;
        RECT 426.800 330.200 427.600 330.400 ;
        RECT 431.400 330.200 432.000 333.600 ;
        RECT 436.200 330.800 437.000 335.200 ;
        RECT 438.000 334.600 438.800 339.800 ;
        RECT 444.400 336.600 445.200 339.800 ;
        RECT 446.000 337.000 446.800 339.800 ;
        RECT 447.600 337.000 448.400 339.800 ;
        RECT 449.200 337.000 450.000 339.800 ;
        RECT 450.800 337.000 451.600 339.800 ;
        RECT 454.000 337.000 454.800 339.800 ;
        RECT 457.200 337.000 458.000 339.800 ;
        RECT 458.800 337.000 459.600 339.800 ;
        RECT 460.400 337.000 461.200 339.800 ;
        RECT 442.800 335.800 445.200 336.600 ;
        RECT 462.000 336.600 462.800 339.800 ;
        RECT 442.800 335.200 443.600 335.800 ;
        RECT 437.600 334.000 438.800 334.600 ;
        RECT 441.800 334.600 443.600 335.200 ;
        RECT 447.600 335.600 448.600 336.400 ;
        RECT 451.600 335.600 453.200 336.400 ;
        RECT 454.000 335.800 458.600 336.400 ;
        RECT 462.000 335.800 464.600 336.600 ;
        RECT 454.000 335.600 454.800 335.800 ;
        RECT 437.600 332.000 438.200 334.000 ;
        RECT 441.800 333.400 442.600 334.600 ;
        RECT 438.800 332.600 442.600 333.400 ;
        RECT 447.600 332.800 448.400 335.600 ;
        RECT 454.000 334.800 454.800 335.000 ;
        RECT 450.400 334.200 454.800 334.800 ;
        RECT 450.400 334.000 451.200 334.200 ;
        RECT 455.600 333.600 456.400 335.200 ;
        RECT 457.800 333.400 458.600 335.800 ;
        RECT 463.800 335.200 464.600 335.800 ;
        RECT 463.800 334.400 466.800 335.200 ;
        RECT 468.400 333.800 469.200 339.800 ;
        RECT 472.600 338.400 473.400 339.800 ;
        RECT 477.400 338.400 478.200 339.800 ;
        RECT 471.600 337.600 473.400 338.400 ;
        RECT 476.400 337.600 478.200 338.400 ;
        RECT 472.600 336.400 473.400 337.600 ;
        RECT 477.400 336.400 478.200 337.600 ;
        RECT 471.600 335.800 473.400 336.400 ;
        RECT 476.400 335.800 478.200 336.400 ;
        RECT 450.800 332.600 454.000 333.400 ;
        RECT 457.800 332.600 459.800 333.400 ;
        RECT 460.400 333.000 469.200 333.800 ;
        RECT 470.000 333.600 470.800 335.200 ;
        RECT 444.400 332.000 445.200 332.600 ;
        RECT 462.000 332.000 462.800 332.400 ;
        RECT 463.600 332.000 464.400 332.400 ;
        RECT 467.000 332.000 467.800 332.200 ;
        RECT 437.600 331.400 438.400 332.000 ;
        RECT 444.400 331.400 467.800 332.000 ;
        RECT 433.200 330.200 434.000 330.400 ;
        RECT 424.600 329.600 425.600 330.200 ;
        RECT 426.200 329.600 427.600 330.200 ;
        RECT 431.000 329.600 432.000 330.200 ;
        RECT 432.600 329.600 434.000 330.200 ;
        RECT 436.200 330.000 437.200 330.800 ;
        RECT 424.600 322.200 425.400 329.600 ;
        RECT 426.200 328.400 426.800 329.600 ;
        RECT 426.000 327.600 426.800 328.400 ;
        RECT 431.000 322.200 431.800 329.600 ;
        RECT 432.600 328.400 433.200 329.600 ;
        RECT 432.400 327.600 433.200 328.400 ;
        RECT 436.400 322.200 437.200 330.000 ;
        RECT 437.800 329.600 438.400 331.400 ;
        RECT 437.800 329.000 446.800 329.600 ;
        RECT 437.800 327.400 438.400 329.000 ;
        RECT 446.000 328.800 446.800 329.000 ;
        RECT 449.200 329.000 457.800 329.600 ;
        RECT 449.200 328.800 450.000 329.000 ;
        RECT 441.000 327.600 443.600 328.400 ;
        RECT 437.800 326.800 440.400 327.400 ;
        RECT 439.600 322.200 440.400 326.800 ;
        RECT 442.800 322.200 443.600 327.600 ;
        RECT 444.200 326.800 448.400 327.600 ;
        RECT 446.000 322.200 446.800 325.000 ;
        RECT 447.600 322.200 448.400 325.000 ;
        RECT 449.200 322.200 450.000 325.000 ;
        RECT 450.800 322.200 451.600 328.400 ;
        RECT 454.000 327.600 456.600 328.400 ;
        RECT 457.200 328.200 457.800 329.000 ;
        RECT 458.800 329.400 459.600 329.600 ;
        RECT 458.800 329.000 464.200 329.400 ;
        RECT 458.800 328.800 465.000 329.000 ;
        RECT 463.600 328.200 465.000 328.800 ;
        RECT 457.200 327.600 463.000 328.200 ;
        RECT 466.000 328.000 467.600 328.800 ;
        RECT 466.000 327.600 466.600 328.000 ;
        RECT 454.000 322.200 454.800 327.000 ;
        RECT 457.200 322.200 458.000 327.000 ;
        RECT 462.400 326.800 466.600 327.600 ;
        RECT 468.400 327.400 469.200 333.000 ;
        RECT 467.200 326.800 469.200 327.400 ;
        RECT 458.800 322.200 459.600 325.000 ;
        RECT 460.400 322.200 461.200 325.000 ;
        RECT 463.600 322.200 464.400 326.800 ;
        RECT 467.200 326.200 467.800 326.800 ;
        RECT 466.800 325.600 467.800 326.200 ;
        RECT 466.800 322.200 467.600 325.600 ;
        RECT 471.600 322.200 472.400 335.800 ;
        RECT 474.800 333.600 475.600 335.200 ;
        RECT 473.200 330.300 474.000 330.400 ;
        RECT 474.800 330.300 475.600 330.400 ;
        RECT 473.200 329.700 475.600 330.300 ;
        RECT 473.200 328.800 474.000 329.700 ;
        RECT 474.800 329.600 475.600 329.700 ;
        RECT 476.400 322.200 477.200 335.800 ;
        RECT 479.600 335.600 480.400 337.200 ;
        RECT 481.200 332.300 482.000 339.800 ;
        RECT 482.800 336.000 483.600 339.800 ;
        RECT 486.000 336.000 486.800 339.800 ;
        RECT 482.800 335.800 486.800 336.000 ;
        RECT 487.600 335.800 488.400 339.800 ;
        RECT 490.800 336.400 491.600 339.800 ;
        RECT 490.600 335.800 491.600 336.400 ;
        RECT 483.000 335.400 486.600 335.800 ;
        RECT 483.600 334.400 484.400 334.800 ;
        RECT 487.600 334.400 488.200 335.800 ;
        RECT 490.600 334.400 491.200 335.800 ;
        RECT 494.000 335.200 494.800 339.800 ;
        RECT 492.200 334.600 494.800 335.200 ;
        RECT 495.600 337.000 496.400 339.000 ;
        RECT 495.600 334.800 496.200 337.000 ;
        RECT 499.800 336.000 500.600 339.000 ;
        RECT 505.200 336.000 506.000 339.800 ;
        RECT 508.400 336.000 509.200 339.800 ;
        RECT 499.800 335.400 501.400 336.000 ;
        RECT 505.200 335.800 509.200 336.000 ;
        RECT 510.000 335.800 510.800 339.800 ;
        RECT 511.600 335.800 512.400 339.800 ;
        RECT 513.200 336.000 514.000 339.800 ;
        RECT 516.400 336.000 517.200 339.800 ;
        RECT 513.200 335.800 517.200 336.000 ;
        RECT 505.400 335.400 509.000 335.800 ;
        RECT 500.600 335.000 501.400 335.400 ;
        RECT 482.800 333.800 484.400 334.400 ;
        RECT 482.800 333.600 483.600 333.800 ;
        RECT 485.800 333.600 488.400 334.400 ;
        RECT 489.200 334.300 490.000 334.400 ;
        RECT 490.600 334.300 491.600 334.400 ;
        RECT 489.200 333.700 491.600 334.300 ;
        RECT 489.200 333.600 490.000 333.700 ;
        RECT 490.600 333.600 491.600 333.700 ;
        RECT 484.400 332.300 485.200 333.200 ;
        RECT 481.200 331.700 485.200 332.300 ;
        RECT 478.000 328.800 478.800 330.400 ;
        RECT 481.200 322.200 482.000 331.700 ;
        RECT 484.400 331.600 485.200 331.700 ;
        RECT 485.800 330.200 486.400 333.600 ;
        RECT 487.600 330.200 488.400 330.400 ;
        RECT 485.400 329.600 486.400 330.200 ;
        RECT 487.000 329.600 488.400 330.200 ;
        RECT 490.600 330.200 491.200 333.600 ;
        RECT 492.200 333.000 492.800 334.600 ;
        RECT 495.600 334.200 499.800 334.800 ;
        RECT 498.800 333.800 499.800 334.200 ;
        RECT 500.800 334.400 501.400 335.000 ;
        RECT 506.000 334.400 506.800 334.800 ;
        RECT 510.000 334.400 510.600 335.800 ;
        RECT 511.800 334.400 512.400 335.800 ;
        RECT 513.400 335.400 517.000 335.800 ;
        RECT 518.000 335.600 518.800 337.200 ;
        RECT 515.600 334.400 516.400 334.800 ;
        RECT 491.800 332.200 492.800 333.000 ;
        RECT 492.200 330.200 492.800 332.200 ;
        RECT 495.600 331.600 496.400 333.200 ;
        RECT 497.200 331.600 498.000 333.200 ;
        RECT 498.800 333.000 500.200 333.800 ;
        RECT 500.800 333.600 502.800 334.400 ;
        RECT 505.200 333.800 506.800 334.400 ;
        RECT 505.200 333.600 506.000 333.800 ;
        RECT 508.200 333.600 510.800 334.400 ;
        RECT 511.600 333.600 514.200 334.400 ;
        RECT 515.600 333.800 517.200 334.400 ;
        RECT 516.400 333.600 517.200 333.800 ;
        RECT 498.800 331.000 499.400 333.000 ;
        RECT 495.600 330.400 499.400 331.000 ;
        RECT 485.400 324.400 486.200 329.600 ;
        RECT 487.000 328.400 487.600 329.600 ;
        RECT 490.600 329.200 491.600 330.200 ;
        RECT 492.200 329.600 494.800 330.200 ;
        RECT 486.800 327.600 487.600 328.400 ;
        RECT 484.400 323.600 486.200 324.400 ;
        RECT 485.400 322.200 486.200 323.600 ;
        RECT 490.800 322.200 491.600 329.200 ;
        RECT 494.000 322.200 494.800 329.600 ;
        RECT 495.600 327.000 496.200 330.400 ;
        RECT 500.800 329.800 501.400 333.600 ;
        RECT 502.000 332.300 502.800 332.400 ;
        RECT 503.600 332.300 504.400 332.400 ;
        RECT 502.000 331.700 504.400 332.300 ;
        RECT 502.000 330.800 502.800 331.700 ;
        RECT 503.600 331.600 504.400 331.700 ;
        RECT 506.800 331.600 507.600 333.200 ;
        RECT 508.200 330.200 508.800 333.600 ;
        RECT 513.600 332.300 514.200 333.600 ;
        RECT 510.100 331.700 514.200 332.300 ;
        RECT 510.100 330.400 510.700 331.700 ;
        RECT 510.000 330.200 510.800 330.400 ;
        RECT 499.800 329.200 501.400 329.800 ;
        RECT 507.800 329.600 508.800 330.200 ;
        RECT 509.400 329.600 510.800 330.200 ;
        RECT 511.600 330.200 512.400 330.400 ;
        RECT 513.600 330.200 514.200 331.700 ;
        RECT 514.800 331.600 515.600 333.200 ;
        RECT 511.600 329.600 513.000 330.200 ;
        RECT 513.600 329.600 514.600 330.200 ;
        RECT 495.600 323.000 496.400 327.000 ;
        RECT 499.800 322.200 500.600 329.200 ;
        RECT 507.800 322.200 508.600 329.600 ;
        RECT 509.400 328.400 510.000 329.600 ;
        RECT 509.200 327.600 510.000 328.400 ;
        RECT 512.400 328.400 513.000 329.600 ;
        RECT 512.400 327.600 513.200 328.400 ;
        RECT 513.800 322.200 514.600 329.600 ;
        RECT 519.600 322.200 520.400 339.800 ;
        RECT 521.200 336.000 522.000 339.800 ;
        RECT 524.400 336.000 525.200 339.800 ;
        RECT 521.200 335.800 525.200 336.000 ;
        RECT 526.000 335.800 526.800 339.800 ;
        RECT 521.400 335.400 525.000 335.800 ;
        RECT 522.000 334.400 522.800 334.800 ;
        RECT 526.000 334.400 526.600 335.800 ;
        RECT 527.600 335.200 528.400 339.800 ;
        RECT 530.800 336.400 531.600 339.800 ;
        RECT 530.800 335.800 531.800 336.400 ;
        RECT 527.600 334.600 530.200 335.200 ;
        RECT 521.200 333.800 522.800 334.400 ;
        RECT 521.200 333.600 522.000 333.800 ;
        RECT 524.200 333.600 526.800 334.400 ;
        RECT 522.800 331.600 523.600 333.200 ;
        RECT 524.200 330.200 524.800 333.600 ;
        RECT 527.800 332.400 528.600 333.200 ;
        RECT 527.600 331.600 528.600 332.400 ;
        RECT 529.600 333.000 530.200 334.600 ;
        RECT 531.200 334.400 531.800 335.800 ;
        RECT 530.800 333.600 531.800 334.400 ;
        RECT 537.600 334.200 538.400 339.800 ;
        RECT 540.400 336.000 541.200 339.800 ;
        RECT 543.600 336.000 544.400 339.800 ;
        RECT 540.400 335.800 544.400 336.000 ;
        RECT 545.200 335.800 546.000 339.800 ;
        RECT 540.600 335.400 544.200 335.800 ;
        RECT 541.200 334.400 542.000 334.800 ;
        RECT 545.200 334.400 545.800 335.800 ;
        RECT 537.600 333.800 539.400 334.200 ;
        RECT 537.800 333.600 539.400 333.800 ;
        RECT 540.400 333.800 542.000 334.400 ;
        RECT 540.400 333.600 541.200 333.800 ;
        RECT 543.400 333.600 546.000 334.400 ;
        RECT 550.400 334.200 551.200 339.800 ;
        RECT 553.200 336.000 554.000 339.800 ;
        RECT 556.400 336.000 557.200 339.800 ;
        RECT 553.200 335.800 557.200 336.000 ;
        RECT 558.000 335.800 558.800 339.800 ;
        RECT 553.400 335.400 557.000 335.800 ;
        RECT 554.000 334.400 554.800 334.800 ;
        RECT 558.000 334.400 558.600 335.800 ;
        RECT 559.600 335.400 560.400 339.800 ;
        RECT 563.800 338.400 565.000 339.800 ;
        RECT 563.800 337.800 565.200 338.400 ;
        RECT 568.400 337.800 569.200 339.800 ;
        RECT 572.800 338.400 573.600 339.800 ;
        RECT 572.800 337.800 574.800 338.400 ;
        RECT 564.400 337.000 565.200 337.800 ;
        RECT 568.600 337.200 569.200 337.800 ;
        RECT 568.600 336.600 571.400 337.200 ;
        RECT 570.600 336.400 571.400 336.600 ;
        RECT 572.400 336.400 573.200 337.200 ;
        RECT 574.000 337.000 574.800 337.800 ;
        RECT 562.600 335.400 563.400 335.600 ;
        RECT 559.600 334.800 563.400 335.400 ;
        RECT 550.400 333.800 552.200 334.200 ;
        RECT 550.600 333.600 552.200 333.800 ;
        RECT 553.200 333.800 554.800 334.400 ;
        RECT 553.200 333.600 554.000 333.800 ;
        RECT 556.200 333.600 558.800 334.400 ;
        RECT 529.600 332.200 530.600 333.000 ;
        RECT 526.000 330.200 526.800 330.400 ;
        RECT 529.600 330.200 530.200 332.200 ;
        RECT 531.200 330.200 531.800 333.600 ;
        RECT 535.600 331.600 537.200 332.400 ;
        RECT 523.800 329.600 524.800 330.200 ;
        RECT 525.400 329.600 526.800 330.200 ;
        RECT 527.600 329.600 530.200 330.200 ;
        RECT 523.800 322.200 524.600 329.600 ;
        RECT 525.400 328.400 526.000 329.600 ;
        RECT 525.200 327.600 526.000 328.400 ;
        RECT 527.600 322.200 528.400 329.600 ;
        RECT 530.800 329.200 531.800 330.200 ;
        RECT 534.000 329.600 534.800 331.200 ;
        RECT 538.800 330.400 539.400 333.600 ;
        RECT 542.000 331.600 542.800 333.200 ;
        RECT 538.800 329.600 539.600 330.400 ;
        RECT 543.400 330.200 544.000 333.600 ;
        RECT 548.400 331.600 550.000 332.400 ;
        RECT 545.200 330.200 546.000 330.400 ;
        RECT 543.000 329.600 544.000 330.200 ;
        RECT 544.600 329.600 546.000 330.200 ;
        RECT 546.800 330.300 547.600 331.200 ;
        RECT 551.600 330.400 552.200 333.600 ;
        RECT 554.800 331.600 555.600 333.200 ;
        RECT 548.400 330.300 549.200 330.400 ;
        RECT 546.800 329.700 549.200 330.300 ;
        RECT 546.800 329.600 547.600 329.700 ;
        RECT 548.400 329.600 549.200 329.700 ;
        RECT 551.600 329.600 552.400 330.400 ;
        RECT 556.200 330.200 556.800 333.600 ;
        RECT 559.600 331.400 560.400 334.800 ;
        RECT 566.600 334.200 567.400 334.400 ;
        RECT 569.200 334.200 570.000 334.400 ;
        RECT 572.400 334.200 573.000 336.400 ;
        RECT 577.200 335.000 578.000 339.800 ;
        RECT 583.600 336.000 584.400 339.800 ;
        RECT 586.800 336.000 587.600 339.800 ;
        RECT 583.600 335.800 587.600 336.000 ;
        RECT 588.400 335.800 589.200 339.800 ;
        RECT 590.000 335.800 590.800 339.800 ;
        RECT 591.600 336.000 592.400 339.800 ;
        RECT 594.800 336.000 595.600 339.800 ;
        RECT 591.600 335.800 595.600 336.000 ;
        RECT 583.800 335.400 587.400 335.800 ;
        RECT 584.400 334.400 585.200 334.800 ;
        RECT 588.400 334.400 589.000 335.800 ;
        RECT 590.200 334.400 590.800 335.800 ;
        RECT 591.800 335.400 595.400 335.800 ;
        RECT 594.000 334.400 594.800 334.800 ;
        RECT 575.600 334.200 577.200 334.400 ;
        RECT 566.200 333.600 577.200 334.200 ;
        RECT 582.000 334.300 582.800 334.400 ;
        RECT 583.600 334.300 585.200 334.400 ;
        RECT 582.000 333.800 585.200 334.300 ;
        RECT 582.000 333.700 584.400 333.800 ;
        RECT 582.000 333.600 582.800 333.700 ;
        RECT 583.600 333.600 584.400 333.700 ;
        RECT 586.600 333.600 589.200 334.400 ;
        RECT 590.000 333.600 592.600 334.400 ;
        RECT 594.000 333.800 595.600 334.400 ;
        RECT 600.000 334.200 600.800 339.800 ;
        RECT 602.800 335.200 603.600 339.800 ;
        RECT 606.000 336.400 606.800 339.800 ;
        RECT 606.000 335.800 607.000 336.400 ;
        RECT 609.200 335.800 610.000 339.800 ;
        RECT 610.800 336.000 611.600 339.800 ;
        RECT 614.000 336.000 614.800 339.800 ;
        RECT 610.800 335.800 614.800 336.000 ;
        RECT 602.800 334.600 605.400 335.200 ;
        RECT 600.000 333.800 601.800 334.200 ;
        RECT 594.800 333.600 595.600 333.800 ;
        RECT 600.200 333.600 601.800 333.800 ;
        RECT 564.400 332.800 565.200 333.000 ;
        RECT 561.400 332.200 565.200 332.800 ;
        RECT 561.400 332.000 562.200 332.200 ;
        RECT 563.000 331.400 563.800 331.600 ;
        RECT 559.600 330.800 563.800 331.400 ;
        RECT 558.000 330.200 558.800 330.400 ;
        RECT 555.800 329.600 556.800 330.200 ;
        RECT 557.400 329.600 558.800 330.200 ;
        RECT 530.800 322.200 531.600 329.200 ;
        RECT 537.200 327.600 538.000 329.200 ;
        RECT 538.800 327.000 539.400 329.600 ;
        RECT 535.800 326.400 539.400 327.000 ;
        RECT 535.800 326.200 536.400 326.400 ;
        RECT 535.600 322.200 536.400 326.200 ;
        RECT 538.800 326.200 539.400 326.400 ;
        RECT 538.800 322.200 539.600 326.200 ;
        RECT 543.000 322.200 543.800 329.600 ;
        RECT 544.600 328.400 545.200 329.600 ;
        RECT 544.400 327.600 545.200 328.400 ;
        RECT 550.000 327.600 550.800 329.200 ;
        RECT 551.600 327.000 552.200 329.600 ;
        RECT 548.600 326.400 552.200 327.000 ;
        RECT 548.600 326.200 549.200 326.400 ;
        RECT 548.400 322.200 549.200 326.200 ;
        RECT 551.600 326.200 552.200 326.400 ;
        RECT 551.600 322.200 552.400 326.200 ;
        RECT 555.800 322.200 556.600 329.600 ;
        RECT 557.400 328.400 558.000 329.600 ;
        RECT 557.200 327.600 558.000 328.400 ;
        RECT 559.600 322.200 560.400 330.800 ;
        RECT 566.200 330.400 566.800 333.600 ;
        RECT 573.400 333.400 574.200 333.600 ;
        RECT 572.400 332.400 573.200 332.600 ;
        RECT 575.000 332.400 575.800 332.600 ;
        RECT 570.800 331.800 575.800 332.400 ;
        RECT 570.800 331.600 571.600 331.800 ;
        RECT 585.200 331.600 586.000 333.200 ;
        RECT 586.600 332.400 587.200 333.600 ;
        RECT 586.600 331.600 587.600 332.400 ;
        RECT 588.400 332.300 589.200 332.400 ;
        RECT 588.400 331.700 590.700 332.300 ;
        RECT 588.400 331.600 589.200 331.700 ;
        RECT 572.400 331.000 578.000 331.200 ;
        RECT 572.200 330.800 578.000 331.000 ;
        RECT 564.400 329.800 566.800 330.400 ;
        RECT 568.200 330.600 578.000 330.800 ;
        RECT 568.200 330.200 573.000 330.600 ;
        RECT 564.400 328.800 565.000 329.800 ;
        RECT 563.600 328.000 565.000 328.800 ;
        RECT 566.600 329.000 567.400 329.200 ;
        RECT 568.200 329.000 568.800 330.200 ;
        RECT 566.600 328.400 568.800 329.000 ;
        RECT 569.400 329.000 574.800 329.600 ;
        RECT 569.400 328.800 570.200 329.000 ;
        RECT 574.000 328.800 574.800 329.000 ;
        RECT 567.800 327.400 568.600 327.600 ;
        RECT 570.600 327.400 571.400 327.600 ;
        RECT 564.400 326.200 565.200 327.000 ;
        RECT 567.800 326.800 571.400 327.400 ;
        RECT 568.600 326.200 569.200 326.800 ;
        RECT 574.000 326.200 574.800 327.000 ;
        RECT 563.800 322.200 565.000 326.200 ;
        RECT 568.400 322.200 569.200 326.200 ;
        RECT 572.800 325.600 574.800 326.200 ;
        RECT 572.800 322.200 573.600 325.600 ;
        RECT 577.200 322.200 578.000 330.600 ;
        RECT 586.600 330.200 587.200 331.600 ;
        RECT 590.100 330.400 590.700 331.700 ;
        RECT 588.400 330.200 589.200 330.400 ;
        RECT 586.200 329.600 587.200 330.200 ;
        RECT 587.800 329.600 589.200 330.200 ;
        RECT 590.000 330.200 590.800 330.400 ;
        RECT 592.000 330.200 592.600 333.600 ;
        RECT 593.200 331.600 594.000 333.200 ;
        RECT 598.000 331.600 599.600 332.400 ;
        RECT 596.400 330.300 597.200 331.200 ;
        RECT 601.200 330.400 601.800 333.600 ;
        RECT 603.000 332.400 603.800 333.200 ;
        RECT 602.800 331.600 603.800 332.400 ;
        RECT 604.800 333.000 605.400 334.600 ;
        RECT 606.400 334.400 607.000 335.800 ;
        RECT 609.400 334.400 610.000 335.800 ;
        RECT 611.000 335.400 614.600 335.800 ;
        RECT 615.600 335.200 616.400 339.800 ;
        RECT 618.800 336.400 619.600 339.800 ;
        RECT 618.800 335.800 619.800 336.400 ;
        RECT 622.000 336.000 622.800 339.800 ;
        RECT 625.200 336.000 626.000 339.800 ;
        RECT 622.000 335.800 626.000 336.000 ;
        RECT 626.800 335.800 627.600 339.800 ;
        RECT 613.200 334.400 614.000 334.800 ;
        RECT 615.600 334.600 618.200 335.200 ;
        RECT 606.000 334.300 607.000 334.400 ;
        RECT 607.600 334.300 608.400 334.400 ;
        RECT 606.000 333.700 608.400 334.300 ;
        RECT 606.000 333.600 607.000 333.700 ;
        RECT 607.600 333.600 608.400 333.700 ;
        RECT 609.200 333.600 611.800 334.400 ;
        RECT 613.200 333.800 614.800 334.400 ;
        RECT 614.000 333.600 614.800 333.800 ;
        RECT 604.800 332.200 605.800 333.000 ;
        RECT 598.000 330.300 598.800 330.400 ;
        RECT 590.000 329.600 591.400 330.200 ;
        RECT 592.000 329.600 593.000 330.200 ;
        RECT 596.400 329.700 598.800 330.300 ;
        RECT 596.400 329.600 597.200 329.700 ;
        RECT 598.000 329.600 598.800 329.700 ;
        RECT 601.200 329.600 602.000 330.400 ;
        RECT 604.800 330.200 605.400 332.200 ;
        RECT 606.400 330.200 607.000 333.600 ;
        RECT 602.800 329.600 605.400 330.200 ;
        RECT 586.200 322.200 587.000 329.600 ;
        RECT 587.800 328.400 588.400 329.600 ;
        RECT 587.600 327.600 588.400 328.400 ;
        RECT 590.800 328.400 591.400 329.600 ;
        RECT 590.800 327.600 591.600 328.400 ;
        RECT 592.200 322.200 593.000 329.600 ;
        RECT 596.400 328.300 597.200 328.400 ;
        RECT 596.400 327.700 598.700 328.300 ;
        RECT 596.400 327.600 597.200 327.700 ;
        RECT 598.100 327.000 598.700 327.700 ;
        RECT 599.600 327.600 600.400 329.200 ;
        RECT 601.200 327.000 601.800 329.600 ;
        RECT 598.100 326.400 601.800 327.000 ;
        RECT 598.100 326.200 598.800 326.400 ;
        RECT 598.000 322.200 598.800 326.200 ;
        RECT 601.200 326.200 601.800 326.400 ;
        RECT 601.200 322.200 602.000 326.200 ;
        RECT 602.800 322.200 603.600 329.600 ;
        RECT 606.000 329.200 607.000 330.200 ;
        RECT 609.200 330.200 610.000 330.400 ;
        RECT 611.200 330.200 611.800 333.600 ;
        RECT 612.400 332.300 613.200 333.200 ;
        RECT 615.800 332.400 616.600 333.200 ;
        RECT 614.000 332.300 614.800 332.400 ;
        RECT 612.400 331.700 614.800 332.300 ;
        RECT 612.400 331.600 613.200 331.700 ;
        RECT 614.000 331.600 614.800 331.700 ;
        RECT 615.600 331.600 616.600 332.400 ;
        RECT 617.600 333.000 618.200 334.600 ;
        RECT 619.200 334.400 619.800 335.800 ;
        RECT 622.200 335.400 625.800 335.800 ;
        RECT 622.800 334.400 623.600 334.800 ;
        RECT 626.800 334.400 627.400 335.800 ;
        RECT 618.800 334.300 619.800 334.400 ;
        RECT 620.400 334.300 621.200 334.400 ;
        RECT 618.800 333.700 621.200 334.300 ;
        RECT 618.800 333.600 619.800 333.700 ;
        RECT 620.400 333.600 621.200 333.700 ;
        RECT 622.000 333.800 623.600 334.400 ;
        RECT 622.000 333.600 622.800 333.800 ;
        RECT 625.000 333.600 627.600 334.400 ;
        RECT 629.600 334.200 630.400 339.800 ;
        RECT 628.600 333.800 630.400 334.200 ;
        RECT 628.600 333.600 630.200 333.800 ;
        RECT 617.600 332.200 618.600 333.000 ;
        RECT 617.600 330.200 618.200 332.200 ;
        RECT 619.200 330.200 619.800 333.600 ;
        RECT 623.600 331.600 624.400 333.200 ;
        RECT 625.000 330.200 625.600 333.600 ;
        RECT 628.600 330.400 629.200 333.600 ;
        RECT 630.800 331.600 632.400 332.400 ;
        RECT 626.800 330.300 627.600 330.400 ;
        RECT 628.400 330.300 629.200 330.400 ;
        RECT 626.800 330.200 629.200 330.300 ;
        RECT 609.200 329.600 610.600 330.200 ;
        RECT 611.200 329.600 612.200 330.200 ;
        RECT 606.000 322.200 606.800 329.200 ;
        RECT 610.000 328.400 610.600 329.600 ;
        RECT 610.000 327.600 610.800 328.400 ;
        RECT 611.400 322.200 612.200 329.600 ;
        RECT 615.600 329.600 618.200 330.200 ;
        RECT 615.600 322.200 616.400 329.600 ;
        RECT 618.800 329.200 619.800 330.200 ;
        RECT 624.600 329.600 625.600 330.200 ;
        RECT 626.200 329.700 629.200 330.200 ;
        RECT 626.200 329.600 627.600 329.700 ;
        RECT 628.400 329.600 629.200 329.700 ;
        RECT 633.200 329.600 634.000 331.200 ;
        RECT 618.800 322.200 619.600 329.200 ;
        RECT 624.600 322.200 625.400 329.600 ;
        RECT 626.200 328.400 626.800 329.600 ;
        RECT 626.000 327.600 626.800 328.400 ;
        RECT 628.600 327.000 629.200 329.600 ;
        RECT 630.000 327.600 630.800 329.200 ;
        RECT 628.600 326.400 632.200 327.000 ;
        RECT 628.600 326.200 629.200 326.400 ;
        RECT 628.400 322.200 629.200 326.200 ;
        RECT 631.600 326.200 632.200 326.400 ;
        RECT 631.600 322.200 632.400 326.200 ;
        RECT 634.800 322.200 635.600 339.800 ;
        RECT 636.400 335.600 637.200 337.200 ;
        RECT 638.000 337.000 638.800 339.000 ;
        RECT 642.200 338.400 643.000 339.000 ;
        RECT 642.200 337.600 643.600 338.400 ;
        RECT 638.000 334.800 638.600 337.000 ;
        RECT 642.200 336.000 643.000 337.600 ;
        RECT 647.600 336.000 648.400 339.800 ;
        RECT 650.800 336.000 651.600 339.800 ;
        RECT 642.200 335.400 643.800 336.000 ;
        RECT 647.600 335.800 651.600 336.000 ;
        RECT 652.400 335.800 653.200 339.800 ;
        RECT 654.000 337.000 654.800 339.000 ;
        RECT 647.800 335.400 651.400 335.800 ;
        RECT 643.000 335.000 643.800 335.400 ;
        RECT 638.000 334.200 642.200 334.800 ;
        RECT 641.200 333.800 642.200 334.200 ;
        RECT 643.200 334.400 643.800 335.000 ;
        RECT 648.400 334.400 649.200 334.800 ;
        RECT 652.400 334.400 653.000 335.800 ;
        RECT 654.000 334.800 654.600 337.000 ;
        RECT 658.200 336.000 659.000 339.000 ;
        RECT 658.200 335.400 659.800 336.000 ;
        RECT 663.600 335.800 664.400 339.800 ;
        RECT 665.200 336.000 666.000 339.800 ;
        RECT 668.400 336.000 669.200 339.800 ;
        RECT 665.200 335.800 669.200 336.000 ;
        RECT 659.000 335.000 659.800 335.400 ;
        RECT 638.000 331.600 638.800 333.200 ;
        RECT 639.600 331.600 640.400 333.200 ;
        RECT 641.200 333.000 642.600 333.800 ;
        RECT 643.200 333.600 645.200 334.400 ;
        RECT 647.600 333.800 649.200 334.400 ;
        RECT 647.600 333.600 648.400 333.800 ;
        RECT 650.600 333.600 653.200 334.400 ;
        RECT 654.000 334.200 658.200 334.800 ;
        RECT 657.200 333.800 658.200 334.200 ;
        RECT 659.200 334.400 659.800 335.000 ;
        RECT 663.800 334.400 664.400 335.800 ;
        RECT 665.400 335.400 669.000 335.800 ;
        RECT 670.000 335.000 670.800 339.800 ;
        RECT 674.400 338.400 675.200 339.800 ;
        RECT 673.200 337.800 675.200 338.400 ;
        RECT 678.800 337.800 679.600 339.800 ;
        RECT 683.000 338.400 684.200 339.800 ;
        RECT 682.800 337.800 684.200 338.400 ;
        RECT 673.200 337.000 674.000 337.800 ;
        RECT 678.800 337.200 679.400 337.800 ;
        RECT 674.800 336.400 675.600 337.200 ;
        RECT 676.600 336.600 679.400 337.200 ;
        RECT 682.800 337.000 683.600 337.800 ;
        RECT 676.600 336.400 677.400 336.600 ;
        RECT 667.600 334.400 668.400 334.800 ;
        RECT 641.200 331.000 641.800 333.000 ;
        RECT 638.000 330.400 641.800 331.000 ;
        RECT 638.000 327.000 638.600 330.400 ;
        RECT 643.200 329.800 643.800 333.600 ;
        RECT 644.400 330.800 645.200 332.400 ;
        RECT 649.200 331.600 650.000 333.200 ;
        RECT 650.600 330.200 651.200 333.600 ;
        RECT 654.000 331.600 654.800 333.200 ;
        RECT 655.600 331.600 656.400 333.200 ;
        RECT 657.200 333.000 658.600 333.800 ;
        RECT 659.200 333.600 661.200 334.400 ;
        RECT 663.600 333.600 666.200 334.400 ;
        RECT 667.600 333.800 669.200 334.400 ;
        RECT 668.400 333.600 669.200 333.800 ;
        RECT 670.800 334.200 672.400 334.400 ;
        RECT 675.000 334.200 675.600 336.400 ;
        RECT 684.600 335.400 685.400 335.600 ;
        RECT 687.600 335.400 688.400 339.800 ;
        RECT 684.600 334.800 688.400 335.400 ;
        RECT 680.600 334.200 681.400 334.400 ;
        RECT 670.800 333.600 681.800 334.200 ;
        RECT 657.200 331.000 657.800 333.000 ;
        RECT 654.000 330.400 657.800 331.000 ;
        RECT 652.400 330.200 653.200 330.400 ;
        RECT 642.200 329.200 643.800 329.800 ;
        RECT 650.200 329.600 651.200 330.200 ;
        RECT 651.800 329.600 653.200 330.200 ;
        RECT 638.000 323.000 638.800 327.000 ;
        RECT 642.200 322.200 643.000 329.200 ;
        RECT 650.200 328.400 651.000 329.600 ;
        RECT 651.800 328.400 652.400 329.600 ;
        RECT 649.200 327.600 651.000 328.400 ;
        RECT 651.600 327.600 652.400 328.400 ;
        RECT 650.200 322.200 651.000 327.600 ;
        RECT 654.000 327.000 654.600 330.400 ;
        RECT 659.200 329.800 659.800 333.600 ;
        RECT 660.400 332.300 661.200 332.400 ;
        RECT 662.000 332.300 662.800 332.400 ;
        RECT 660.400 331.700 662.800 332.300 ;
        RECT 660.400 330.800 661.200 331.700 ;
        RECT 662.000 331.600 662.800 331.700 ;
        RECT 658.200 329.200 659.800 329.800 ;
        RECT 663.600 330.200 664.400 330.400 ;
        RECT 665.600 330.200 666.200 333.600 ;
        RECT 673.800 333.400 674.600 333.600 ;
        RECT 666.800 331.600 667.600 333.200 ;
        RECT 672.200 332.400 673.000 332.600 ;
        RECT 674.800 332.400 675.600 332.600 ;
        RECT 681.200 332.400 681.800 333.600 ;
        RECT 682.800 332.800 683.600 333.000 ;
        RECT 672.200 331.800 677.200 332.400 ;
        RECT 676.400 331.600 677.200 331.800 ;
        RECT 681.200 331.600 682.000 332.400 ;
        RECT 682.800 332.200 686.600 332.800 ;
        RECT 685.800 332.000 686.600 332.200 ;
        RECT 670.000 331.000 675.600 331.200 ;
        RECT 670.000 330.800 675.800 331.000 ;
        RECT 670.000 330.600 679.800 330.800 ;
        RECT 663.600 329.600 665.000 330.200 ;
        RECT 665.600 329.600 666.600 330.200 ;
        RECT 658.200 328.400 659.000 329.200 ;
        RECT 657.200 327.600 659.000 328.400 ;
        RECT 664.400 328.400 665.000 329.600 ;
        RECT 665.800 328.400 666.600 329.600 ;
        RECT 664.400 327.600 665.200 328.400 ;
        RECT 665.800 327.600 667.600 328.400 ;
        RECT 654.000 323.000 654.800 327.000 ;
        RECT 658.200 322.200 659.000 327.600 ;
        RECT 665.800 322.200 666.600 327.600 ;
        RECT 670.000 322.200 670.800 330.600 ;
        RECT 675.000 330.200 679.800 330.600 ;
        RECT 673.200 329.000 678.600 329.600 ;
        RECT 673.200 328.800 674.000 329.000 ;
        RECT 677.800 328.800 678.600 329.000 ;
        RECT 679.200 329.000 679.800 330.200 ;
        RECT 681.200 330.400 681.800 331.600 ;
        RECT 684.200 331.400 685.000 331.600 ;
        RECT 687.600 331.400 688.400 334.800 ;
        RECT 684.200 330.800 688.400 331.400 ;
        RECT 681.200 329.800 683.600 330.400 ;
        RECT 680.600 329.000 681.400 329.200 ;
        RECT 679.200 328.400 681.400 329.000 ;
        RECT 683.000 328.800 683.600 329.800 ;
        RECT 683.000 328.000 684.400 328.800 ;
        RECT 676.600 327.400 677.400 327.600 ;
        RECT 679.400 327.400 680.200 327.600 ;
        RECT 673.200 326.200 674.000 327.000 ;
        RECT 676.600 326.800 680.200 327.400 ;
        RECT 678.800 326.200 679.400 326.800 ;
        RECT 682.800 326.200 683.600 327.000 ;
        RECT 673.200 325.600 675.200 326.200 ;
        RECT 674.400 322.200 675.200 325.600 ;
        RECT 678.800 322.200 679.600 326.200 ;
        RECT 683.000 322.200 684.200 326.200 ;
        RECT 687.600 322.200 688.400 330.800 ;
        RECT 2.800 316.400 3.600 319.800 ;
        RECT 2.600 315.800 3.600 316.400 ;
        RECT 2.600 315.200 3.200 315.800 ;
        RECT 6.000 315.200 6.800 319.800 ;
        RECT 9.200 317.000 10.000 319.800 ;
        RECT 10.800 317.000 11.600 319.800 ;
        RECT 1.200 314.600 3.200 315.200 ;
        RECT 1.200 309.000 2.000 314.600 ;
        RECT 3.800 314.400 8.000 315.200 ;
        RECT 12.400 315.000 13.200 319.800 ;
        RECT 15.600 315.000 16.400 319.800 ;
        RECT 3.800 314.000 4.400 314.400 ;
        RECT 2.800 313.200 4.400 314.000 ;
        RECT 7.400 313.800 13.200 314.400 ;
        RECT 5.400 313.200 6.800 313.800 ;
        RECT 5.400 313.000 11.600 313.200 ;
        RECT 6.200 312.600 11.600 313.000 ;
        RECT 10.800 312.400 11.600 312.600 ;
        RECT 12.600 313.000 13.200 313.800 ;
        RECT 13.800 313.600 16.400 314.400 ;
        RECT 18.800 313.600 19.600 319.800 ;
        RECT 20.400 317.000 21.200 319.800 ;
        RECT 22.000 317.000 22.800 319.800 ;
        RECT 23.600 317.000 24.400 319.800 ;
        RECT 22.000 314.400 26.200 315.200 ;
        RECT 26.800 314.400 27.600 319.800 ;
        RECT 30.000 315.200 30.800 319.800 ;
        RECT 30.000 314.600 32.600 315.200 ;
        RECT 26.800 313.600 29.400 314.400 ;
        RECT 20.400 313.000 21.200 313.200 ;
        RECT 12.600 312.400 21.200 313.000 ;
        RECT 23.600 313.000 24.400 313.200 ;
        RECT 32.000 313.000 32.600 314.600 ;
        RECT 23.600 312.400 32.600 313.000 ;
        RECT 32.000 310.600 32.600 312.400 ;
        RECT 33.200 312.000 34.000 319.800 ;
        RECT 39.000 312.400 39.800 319.800 ;
        RECT 40.400 313.600 41.200 314.400 ;
        RECT 40.600 312.400 41.200 313.600 ;
        RECT 43.600 313.600 44.400 314.400 ;
        RECT 43.600 312.400 44.200 313.600 ;
        RECT 45.000 312.400 45.800 319.800 ;
        RECT 33.200 311.200 34.200 312.000 ;
        RECT 39.000 311.800 40.000 312.400 ;
        RECT 40.600 311.800 42.000 312.400 ;
        RECT 2.600 310.000 26.000 310.600 ;
        RECT 32.000 310.000 32.800 310.600 ;
        RECT 2.600 309.800 3.400 310.000 ;
        RECT 7.600 309.600 8.400 310.000 ;
        RECT 25.200 309.400 26.000 310.000 ;
        RECT 1.200 308.200 10.000 309.000 ;
        RECT 10.600 308.600 12.600 309.400 ;
        RECT 16.400 308.600 19.600 309.400 ;
        RECT 1.200 302.200 2.000 308.200 ;
        RECT 3.600 306.800 6.600 307.600 ;
        RECT 5.800 306.200 6.600 306.800 ;
        RECT 11.800 306.200 12.600 308.600 ;
        RECT 14.000 306.800 14.800 308.400 ;
        RECT 19.200 307.800 20.000 308.000 ;
        RECT 15.600 307.200 20.000 307.800 ;
        RECT 15.600 307.000 16.400 307.200 ;
        RECT 22.000 306.400 22.800 309.200 ;
        RECT 27.800 308.600 31.600 309.400 ;
        RECT 27.800 307.400 28.600 308.600 ;
        RECT 32.200 308.000 32.800 310.000 ;
        RECT 15.600 306.200 16.400 306.400 ;
        RECT 5.800 305.400 8.400 306.200 ;
        RECT 11.800 305.600 16.400 306.200 ;
        RECT 17.200 305.600 18.800 306.400 ;
        RECT 21.800 305.600 22.800 306.400 ;
        RECT 26.800 306.800 28.600 307.400 ;
        RECT 31.600 307.400 32.800 308.000 ;
        RECT 26.800 306.200 27.600 306.800 ;
        RECT 7.600 302.200 8.400 305.400 ;
        RECT 25.200 305.400 27.600 306.200 ;
        RECT 9.200 302.200 10.000 305.000 ;
        RECT 10.800 302.200 11.600 305.000 ;
        RECT 12.400 302.200 13.200 305.000 ;
        RECT 15.600 302.200 16.400 305.000 ;
        RECT 18.800 302.200 19.600 305.000 ;
        RECT 20.400 302.200 21.200 305.000 ;
        RECT 22.000 302.200 22.800 305.000 ;
        RECT 23.600 302.200 24.400 305.000 ;
        RECT 25.200 302.200 26.000 305.400 ;
        RECT 31.600 302.200 32.400 307.400 ;
        RECT 33.400 306.800 34.200 311.200 ;
        RECT 34.800 310.300 35.600 310.400 ;
        RECT 38.000 310.300 38.800 310.400 ;
        RECT 34.800 309.700 38.800 310.300 ;
        RECT 34.800 309.600 35.600 309.700 ;
        RECT 38.000 308.800 38.800 309.700 ;
        RECT 39.400 310.300 40.000 311.800 ;
        RECT 41.200 311.600 42.000 311.800 ;
        RECT 42.800 311.800 44.200 312.400 ;
        RECT 44.800 311.800 45.800 312.400 ;
        RECT 42.800 311.600 43.600 311.800 ;
        RECT 42.900 310.300 43.500 311.600 ;
        RECT 39.400 309.700 43.500 310.300 ;
        RECT 39.400 308.400 40.000 309.700 ;
        RECT 44.800 308.400 45.400 311.800 ;
        RECT 46.000 308.800 46.800 310.400 ;
        RECT 36.400 308.200 37.200 308.400 ;
        RECT 36.400 307.600 38.000 308.200 ;
        RECT 39.400 307.600 42.000 308.400 ;
        RECT 42.800 307.600 45.400 308.400 ;
        RECT 47.600 308.300 48.400 308.400 ;
        RECT 49.200 308.300 50.000 319.800 ;
        RECT 50.800 312.300 51.600 312.400 ;
        RECT 52.400 312.300 53.200 313.200 ;
        RECT 50.800 311.700 53.200 312.300 ;
        RECT 50.800 311.600 51.600 311.700 ;
        RECT 52.400 311.600 53.200 311.700 ;
        RECT 47.600 308.200 50.000 308.300 ;
        RECT 46.800 307.700 50.000 308.200 ;
        RECT 46.800 307.600 48.400 307.700 ;
        RECT 37.200 307.200 38.000 307.600 ;
        RECT 33.200 306.000 34.200 306.800 ;
        RECT 36.600 306.200 40.200 306.600 ;
        RECT 41.200 306.200 41.800 307.600 ;
        RECT 43.000 306.200 43.600 307.600 ;
        RECT 46.800 307.200 47.600 307.600 ;
        RECT 44.600 306.200 48.200 306.600 ;
        RECT 36.400 306.000 40.400 306.200 ;
        RECT 33.200 302.200 34.000 306.000 ;
        RECT 36.400 302.200 37.200 306.000 ;
        RECT 39.600 302.200 40.400 306.000 ;
        RECT 41.200 302.200 42.000 306.200 ;
        RECT 42.800 302.200 43.600 306.200 ;
        RECT 44.400 306.000 48.400 306.200 ;
        RECT 44.400 302.200 45.200 306.000 ;
        RECT 47.600 302.200 48.400 306.000 ;
        RECT 49.200 302.200 50.000 307.700 ;
        RECT 50.800 304.800 51.600 306.400 ;
        RECT 54.000 306.200 54.800 319.800 ;
        RECT 55.600 306.800 56.400 308.400 ;
        RECT 57.200 306.800 58.000 308.400 ;
        RECT 53.000 305.600 54.800 306.200 ;
        RECT 58.800 306.200 59.600 319.800 ;
        RECT 63.600 316.400 64.400 319.800 ;
        RECT 63.400 315.800 64.400 316.400 ;
        RECT 63.400 315.200 64.000 315.800 ;
        RECT 66.800 315.200 67.600 319.800 ;
        RECT 70.000 317.000 70.800 319.800 ;
        RECT 71.600 317.000 72.400 319.800 ;
        RECT 62.000 314.600 64.000 315.200 ;
        RECT 60.400 311.600 61.200 313.200 ;
        RECT 62.000 309.000 62.800 314.600 ;
        RECT 64.600 314.400 68.800 315.200 ;
        RECT 73.200 315.000 74.000 319.800 ;
        RECT 76.400 315.000 77.200 319.800 ;
        RECT 64.600 314.000 65.200 314.400 ;
        RECT 63.600 313.200 65.200 314.000 ;
        RECT 68.200 313.800 74.000 314.400 ;
        RECT 66.200 313.200 67.600 313.800 ;
        RECT 66.200 313.000 72.400 313.200 ;
        RECT 67.000 312.600 72.400 313.000 ;
        RECT 71.600 312.400 72.400 312.600 ;
        RECT 73.400 313.000 74.000 313.800 ;
        RECT 74.600 313.600 77.200 314.400 ;
        RECT 79.600 313.600 80.400 319.800 ;
        RECT 81.200 317.000 82.000 319.800 ;
        RECT 82.800 317.000 83.600 319.800 ;
        RECT 84.400 317.000 85.200 319.800 ;
        RECT 82.800 314.400 87.000 315.200 ;
        RECT 87.600 314.400 88.400 319.800 ;
        RECT 90.800 315.200 91.600 319.800 ;
        RECT 90.800 314.600 93.400 315.200 ;
        RECT 87.600 313.600 90.200 314.400 ;
        RECT 81.200 313.000 82.000 313.200 ;
        RECT 73.400 312.400 82.000 313.000 ;
        RECT 84.400 313.000 85.200 313.200 ;
        RECT 92.800 313.000 93.400 314.600 ;
        RECT 84.400 312.400 93.400 313.000 ;
        RECT 92.800 310.600 93.400 312.400 ;
        RECT 94.000 312.000 94.800 319.800 ;
        RECT 94.000 311.200 95.000 312.000 ;
        RECT 63.400 310.000 86.800 310.600 ;
        RECT 92.800 310.000 93.600 310.600 ;
        RECT 63.400 309.800 64.200 310.000 ;
        RECT 68.400 309.600 69.200 310.000 ;
        RECT 86.000 309.400 86.800 310.000 ;
        RECT 62.000 308.200 70.800 309.000 ;
        RECT 71.400 308.600 73.400 309.400 ;
        RECT 77.200 308.600 80.400 309.400 ;
        RECT 58.800 305.600 60.600 306.200 ;
        RECT 53.000 304.400 53.800 305.600 ;
        RECT 59.800 304.400 60.600 305.600 ;
        RECT 53.000 303.600 54.800 304.400 ;
        RECT 58.800 303.600 60.600 304.400 ;
        RECT 53.000 302.200 53.800 303.600 ;
        RECT 59.800 302.200 60.600 303.600 ;
        RECT 62.000 302.200 62.800 308.200 ;
        RECT 64.400 306.800 67.400 307.600 ;
        RECT 66.600 306.200 67.400 306.800 ;
        RECT 72.600 306.200 73.400 308.600 ;
        RECT 74.800 306.800 75.600 308.400 ;
        RECT 80.000 307.800 80.800 308.000 ;
        RECT 76.400 307.200 80.800 307.800 ;
        RECT 76.400 307.000 77.200 307.200 ;
        RECT 82.800 306.400 83.600 309.200 ;
        RECT 88.600 308.600 92.400 309.400 ;
        RECT 88.600 307.400 89.400 308.600 ;
        RECT 93.000 308.000 93.600 310.000 ;
        RECT 76.400 306.200 77.200 306.400 ;
        RECT 66.600 305.400 69.200 306.200 ;
        RECT 72.600 305.600 77.200 306.200 ;
        RECT 78.000 305.600 79.600 306.400 ;
        RECT 82.600 305.600 83.600 306.400 ;
        RECT 87.600 306.800 89.400 307.400 ;
        RECT 92.400 307.400 93.600 308.000 ;
        RECT 87.600 306.200 88.400 306.800 ;
        RECT 68.400 302.200 69.200 305.400 ;
        RECT 86.000 305.400 88.400 306.200 ;
        RECT 70.000 302.200 70.800 305.000 ;
        RECT 71.600 302.200 72.400 305.000 ;
        RECT 73.200 302.200 74.000 305.000 ;
        RECT 76.400 302.200 77.200 305.000 ;
        RECT 79.600 302.200 80.400 305.000 ;
        RECT 81.200 302.200 82.000 305.000 ;
        RECT 82.800 302.200 83.600 305.000 ;
        RECT 84.400 302.200 85.200 305.000 ;
        RECT 86.000 302.200 86.800 305.400 ;
        RECT 92.400 302.200 93.200 307.400 ;
        RECT 94.200 306.800 95.000 311.200 ;
        RECT 94.000 306.000 95.000 306.800 ;
        RECT 94.000 302.200 94.800 306.000 ;
        RECT 97.200 302.200 98.000 319.800 ;
        RECT 102.000 315.800 102.800 319.800 ;
        RECT 102.200 315.600 102.800 315.800 ;
        RECT 105.200 315.800 106.000 319.800 ;
        RECT 113.200 316.400 114.000 319.800 ;
        RECT 113.000 315.800 114.000 316.400 ;
        RECT 105.200 315.600 105.800 315.800 ;
        RECT 102.200 315.000 105.800 315.600 ;
        RECT 113.000 315.200 113.600 315.800 ;
        RECT 116.400 315.200 117.200 319.800 ;
        RECT 119.600 317.000 120.400 319.800 ;
        RECT 121.200 317.000 122.000 319.800 ;
        RECT 103.600 312.800 104.400 314.400 ;
        RECT 105.200 312.400 105.800 315.000 ;
        RECT 111.600 314.600 113.600 315.200 ;
        RECT 100.400 310.800 101.200 312.400 ;
        RECT 105.200 311.600 106.000 312.400 ;
        RECT 102.000 309.600 103.600 310.400 ;
        RECT 105.200 308.400 105.800 311.600 ;
        RECT 104.200 308.200 105.800 308.400 ;
        RECT 104.000 307.800 105.800 308.200 ;
        RECT 111.600 309.000 112.400 314.600 ;
        RECT 114.200 314.400 118.400 315.200 ;
        RECT 122.800 315.000 123.600 319.800 ;
        RECT 126.000 315.000 126.800 319.800 ;
        RECT 114.200 314.000 114.800 314.400 ;
        RECT 113.200 313.200 114.800 314.000 ;
        RECT 117.800 313.800 123.600 314.400 ;
        RECT 115.800 313.200 117.200 313.800 ;
        RECT 115.800 313.000 122.000 313.200 ;
        RECT 116.600 312.600 122.000 313.000 ;
        RECT 121.200 312.400 122.000 312.600 ;
        RECT 123.000 313.000 123.600 313.800 ;
        RECT 124.200 313.600 126.800 314.400 ;
        RECT 129.200 313.600 130.000 319.800 ;
        RECT 130.800 317.000 131.600 319.800 ;
        RECT 132.400 317.000 133.200 319.800 ;
        RECT 134.000 317.000 134.800 319.800 ;
        RECT 132.400 314.400 136.600 315.200 ;
        RECT 137.200 314.400 138.000 319.800 ;
        RECT 140.400 315.200 141.200 319.800 ;
        RECT 140.400 314.600 143.000 315.200 ;
        RECT 137.200 313.600 139.800 314.400 ;
        RECT 130.800 313.000 131.600 313.200 ;
        RECT 123.000 312.400 131.600 313.000 ;
        RECT 134.000 313.000 134.800 313.200 ;
        RECT 142.400 313.000 143.000 314.600 ;
        RECT 134.000 312.400 143.000 313.000 ;
        RECT 142.400 310.600 143.000 312.400 ;
        RECT 143.600 314.300 144.400 319.800 ;
        RECT 147.600 314.300 148.400 314.400 ;
        RECT 143.600 313.700 148.400 314.300 ;
        RECT 143.600 312.000 144.400 313.700 ;
        RECT 147.600 313.600 148.400 313.700 ;
        RECT 147.600 312.400 148.200 313.600 ;
        RECT 149.000 312.400 149.800 319.800 ;
        RECT 143.600 311.200 144.600 312.000 ;
        RECT 146.800 311.800 148.200 312.400 ;
        RECT 148.800 311.800 149.800 312.400 ;
        RECT 146.800 311.600 147.600 311.800 ;
        RECT 113.000 310.000 136.400 310.600 ;
        RECT 142.400 310.000 143.200 310.600 ;
        RECT 113.000 309.800 114.000 310.000 ;
        RECT 113.200 309.600 114.000 309.800 ;
        RECT 118.000 309.600 118.800 310.000 ;
        RECT 135.600 309.400 136.400 310.000 ;
        RECT 111.600 308.200 120.400 309.000 ;
        RECT 121.000 308.600 123.000 309.400 ;
        RECT 126.800 308.600 130.000 309.400 ;
        RECT 98.800 304.800 99.600 306.400 ;
        RECT 104.000 302.200 104.800 307.800 ;
        RECT 111.600 302.200 112.400 308.200 ;
        RECT 114.000 306.800 117.000 307.600 ;
        RECT 116.200 306.200 117.000 306.800 ;
        RECT 122.200 306.200 123.000 308.600 ;
        RECT 124.400 306.800 125.200 308.400 ;
        RECT 129.600 307.800 130.400 308.000 ;
        RECT 126.000 307.200 130.400 307.800 ;
        RECT 126.000 307.000 126.800 307.200 ;
        RECT 132.400 306.400 133.200 309.200 ;
        RECT 138.200 308.600 142.000 309.400 ;
        RECT 138.200 307.400 139.000 308.600 ;
        RECT 142.600 308.000 143.200 310.000 ;
        RECT 126.000 306.200 126.800 306.400 ;
        RECT 116.200 305.400 118.800 306.200 ;
        RECT 122.200 305.600 126.800 306.200 ;
        RECT 127.600 305.600 129.200 306.400 ;
        RECT 132.200 305.600 133.200 306.400 ;
        RECT 137.200 306.800 139.000 307.400 ;
        RECT 142.000 307.400 143.200 308.000 ;
        RECT 137.200 306.200 138.000 306.800 ;
        RECT 118.000 302.200 118.800 305.400 ;
        RECT 135.600 305.400 138.000 306.200 ;
        RECT 119.600 302.200 120.400 305.000 ;
        RECT 121.200 302.200 122.000 305.000 ;
        RECT 122.800 302.200 123.600 305.000 ;
        RECT 126.000 302.200 126.800 305.000 ;
        RECT 129.200 302.200 130.000 305.000 ;
        RECT 130.800 302.200 131.600 305.000 ;
        RECT 132.400 302.200 133.200 305.000 ;
        RECT 134.000 302.200 134.800 305.000 ;
        RECT 135.600 302.200 136.400 305.400 ;
        RECT 142.000 302.200 142.800 307.400 ;
        RECT 143.800 306.800 144.600 311.200 ;
        RECT 148.800 308.400 149.400 311.800 ;
        RECT 153.200 311.600 154.000 313.200 ;
        RECT 150.000 308.800 150.800 310.400 ;
        RECT 146.800 307.600 149.400 308.400 ;
        RECT 151.600 308.200 152.400 308.400 ;
        RECT 150.800 307.600 152.400 308.200 ;
        RECT 143.600 306.000 144.600 306.800 ;
        RECT 147.000 306.200 147.600 307.600 ;
        RECT 150.800 307.200 151.600 307.600 ;
        RECT 148.600 306.200 152.200 306.600 ;
        RECT 154.800 306.200 155.600 319.800 ;
        RECT 156.400 306.800 157.200 308.400 ;
        RECT 143.600 302.200 144.400 306.000 ;
        RECT 146.800 302.200 147.600 306.200 ;
        RECT 148.400 306.000 152.400 306.200 ;
        RECT 148.400 302.200 149.200 306.000 ;
        RECT 151.600 302.200 152.400 306.000 ;
        RECT 153.800 305.600 155.600 306.200 ;
        RECT 153.800 302.200 154.600 305.600 ;
        RECT 158.000 304.800 158.800 306.400 ;
        RECT 159.600 302.200 160.400 319.800 ;
        RECT 162.800 312.800 163.600 319.800 ;
        RECT 162.600 311.800 163.600 312.800 ;
        RECT 166.000 312.400 166.800 319.800 ;
        RECT 164.200 311.800 166.800 312.400 ;
        RECT 169.200 312.000 170.000 319.800 ;
        RECT 172.400 315.200 173.200 319.800 ;
        RECT 162.600 308.400 163.200 311.800 ;
        RECT 164.200 309.800 164.800 311.800 ;
        RECT 169.000 311.200 170.000 312.000 ;
        RECT 170.600 314.600 173.200 315.200 ;
        RECT 170.600 313.000 171.200 314.600 ;
        RECT 175.600 314.400 176.400 319.800 ;
        RECT 178.800 317.000 179.600 319.800 ;
        RECT 180.400 317.000 181.200 319.800 ;
        RECT 182.000 317.000 182.800 319.800 ;
        RECT 177.000 314.400 181.200 315.200 ;
        RECT 173.800 313.600 176.400 314.400 ;
        RECT 183.600 313.600 184.400 319.800 ;
        RECT 186.800 315.000 187.600 319.800 ;
        RECT 190.000 315.000 190.800 319.800 ;
        RECT 191.600 317.000 192.400 319.800 ;
        RECT 193.200 317.000 194.000 319.800 ;
        RECT 196.400 315.200 197.200 319.800 ;
        RECT 199.600 316.400 200.400 319.800 ;
        RECT 199.600 315.800 200.600 316.400 ;
        RECT 200.000 315.200 200.600 315.800 ;
        RECT 195.200 314.400 199.400 315.200 ;
        RECT 200.000 314.600 202.000 315.200 ;
        RECT 186.800 313.600 189.400 314.400 ;
        RECT 190.000 313.800 195.800 314.400 ;
        RECT 198.800 314.000 199.400 314.400 ;
        RECT 178.800 313.000 179.600 313.200 ;
        RECT 170.600 312.400 179.600 313.000 ;
        RECT 182.000 313.000 182.800 313.200 ;
        RECT 190.000 313.000 190.600 313.800 ;
        RECT 196.400 313.200 197.800 313.800 ;
        RECT 198.800 313.200 200.400 314.000 ;
        RECT 182.000 312.400 190.600 313.000 ;
        RECT 191.600 313.000 197.800 313.200 ;
        RECT 191.600 312.600 197.000 313.000 ;
        RECT 191.600 312.400 192.400 312.600 ;
        RECT 163.800 309.000 164.800 309.800 ;
        RECT 162.600 307.600 163.600 308.400 ;
        RECT 162.600 306.200 163.200 307.600 ;
        RECT 164.200 307.400 164.800 309.000 ;
        RECT 165.800 309.600 166.800 310.400 ;
        RECT 165.800 308.800 166.600 309.600 ;
        RECT 164.200 306.800 166.800 307.400 ;
        RECT 162.600 305.600 163.600 306.200 ;
        RECT 162.800 302.200 163.600 305.600 ;
        RECT 166.000 302.200 166.800 306.800 ;
        RECT 169.000 306.800 169.800 311.200 ;
        RECT 170.600 310.600 171.200 312.400 ;
        RECT 170.400 310.000 171.200 310.600 ;
        RECT 177.200 310.000 200.600 310.600 ;
        RECT 170.400 308.000 171.000 310.000 ;
        RECT 177.200 309.400 178.000 310.000 ;
        RECT 194.800 309.600 195.600 310.000 ;
        RECT 198.000 309.600 198.800 310.000 ;
        RECT 199.800 309.800 200.600 310.000 ;
        RECT 171.600 308.600 175.400 309.400 ;
        RECT 170.400 307.400 171.600 308.000 ;
        RECT 169.000 306.000 170.000 306.800 ;
        RECT 169.200 302.200 170.000 306.000 ;
        RECT 170.800 302.200 171.600 307.400 ;
        RECT 174.600 307.400 175.400 308.600 ;
        RECT 174.600 306.800 176.400 307.400 ;
        RECT 175.600 306.200 176.400 306.800 ;
        RECT 180.400 306.400 181.200 309.200 ;
        RECT 183.600 308.600 186.800 309.400 ;
        RECT 190.600 308.600 192.600 309.400 ;
        RECT 201.200 309.000 202.000 314.600 ;
        RECT 183.200 307.800 184.000 308.000 ;
        RECT 183.200 307.200 187.600 307.800 ;
        RECT 186.800 307.000 187.600 307.200 ;
        RECT 188.400 306.800 189.200 308.400 ;
        RECT 175.600 305.400 178.000 306.200 ;
        RECT 180.400 305.600 181.400 306.400 ;
        RECT 184.400 305.600 186.000 306.400 ;
        RECT 186.800 306.200 187.600 306.400 ;
        RECT 190.600 306.200 191.400 308.600 ;
        RECT 193.200 308.200 202.000 309.000 ;
        RECT 196.600 306.800 199.600 307.600 ;
        RECT 196.600 306.200 197.400 306.800 ;
        RECT 186.800 305.600 191.400 306.200 ;
        RECT 177.200 302.200 178.000 305.400 ;
        RECT 194.800 305.400 197.400 306.200 ;
        RECT 178.800 302.200 179.600 305.000 ;
        RECT 180.400 302.200 181.200 305.000 ;
        RECT 182.000 302.200 182.800 305.000 ;
        RECT 183.600 302.200 184.400 305.000 ;
        RECT 186.800 302.200 187.600 305.000 ;
        RECT 190.000 302.200 190.800 305.000 ;
        RECT 191.600 302.200 192.400 305.000 ;
        RECT 193.200 302.200 194.000 305.000 ;
        RECT 194.800 302.200 195.600 305.400 ;
        RECT 201.200 302.200 202.000 308.200 ;
        RECT 202.800 306.800 203.600 308.400 ;
        RECT 204.400 306.200 205.200 319.800 ;
        RECT 206.000 312.300 206.800 313.200 ;
        RECT 207.600 312.300 208.400 313.200 ;
        RECT 206.000 311.700 208.400 312.300 ;
        RECT 206.000 311.600 206.800 311.700 ;
        RECT 207.600 311.600 208.400 311.700 ;
        RECT 206.000 308.300 206.800 308.400 ;
        RECT 209.200 308.300 210.000 319.800 ;
        RECT 210.800 314.300 211.600 314.400 ;
        RECT 213.200 314.300 214.000 314.400 ;
        RECT 210.800 313.700 214.000 314.300 ;
        RECT 210.800 313.600 211.600 313.700 ;
        RECT 213.200 313.600 214.000 313.700 ;
        RECT 213.200 312.400 213.800 313.600 ;
        RECT 214.600 312.400 215.400 319.800 ;
        RECT 212.400 311.800 213.800 312.400 ;
        RECT 214.400 311.800 215.400 312.400 ;
        RECT 218.800 311.800 219.600 319.800 ;
        RECT 222.000 312.400 222.800 319.800 ;
        RECT 220.600 311.800 222.800 312.400 ;
        RECT 223.600 312.400 224.400 319.800 ;
        RECT 226.800 312.800 227.600 319.800 ;
        RECT 223.600 311.800 226.200 312.400 ;
        RECT 226.800 311.800 227.800 312.800 ;
        RECT 212.400 311.600 213.200 311.800 ;
        RECT 214.400 308.400 215.000 311.800 ;
        RECT 215.600 308.800 216.400 310.400 ;
        RECT 218.800 309.600 219.400 311.800 ;
        RECT 220.600 311.200 221.200 311.800 ;
        RECT 220.000 310.400 221.200 311.200 ;
        RECT 206.000 307.700 210.000 308.300 ;
        RECT 206.000 307.600 206.800 307.700 ;
        RECT 209.200 306.200 210.000 307.700 ;
        RECT 210.800 308.300 211.600 308.400 ;
        RECT 212.400 308.300 215.000 308.400 ;
        RECT 210.800 307.700 215.000 308.300 ;
        RECT 217.200 308.200 218.000 308.400 ;
        RECT 210.800 306.800 211.600 307.700 ;
        RECT 212.400 307.600 215.000 307.700 ;
        RECT 216.400 307.600 218.000 308.200 ;
        RECT 212.600 306.200 213.200 307.600 ;
        RECT 216.400 307.200 217.200 307.600 ;
        RECT 214.200 306.200 217.800 306.600 ;
        RECT 204.400 305.600 206.200 306.200 ;
        RECT 205.400 304.400 206.200 305.600 ;
        RECT 204.400 303.600 206.200 304.400 ;
        RECT 205.400 302.200 206.200 303.600 ;
        RECT 208.200 305.600 210.000 306.200 ;
        RECT 208.200 302.200 209.000 305.600 ;
        RECT 212.400 302.200 213.200 306.200 ;
        RECT 214.000 306.000 218.000 306.200 ;
        RECT 214.000 302.200 214.800 306.000 ;
        RECT 217.200 302.200 218.000 306.000 ;
        RECT 218.800 302.200 219.600 309.600 ;
        RECT 220.600 307.400 221.200 310.400 ;
        RECT 222.000 310.300 222.800 310.400 ;
        RECT 223.600 310.300 224.600 310.400 ;
        RECT 222.000 309.700 224.600 310.300 ;
        RECT 222.000 308.800 222.800 309.700 ;
        RECT 223.600 309.600 224.600 309.700 ;
        RECT 223.800 308.800 224.600 309.600 ;
        RECT 225.600 309.800 226.200 311.800 ;
        RECT 225.600 309.000 226.600 309.800 ;
        RECT 225.600 307.400 226.200 309.000 ;
        RECT 227.200 308.400 227.800 311.800 ;
        RECT 226.800 307.600 227.800 308.400 ;
        RECT 220.600 306.800 222.800 307.400 ;
        RECT 222.000 302.200 222.800 306.800 ;
        RECT 223.600 306.800 226.200 307.400 ;
        RECT 223.600 302.200 224.400 306.800 ;
        RECT 227.200 306.200 227.800 307.600 ;
        RECT 226.800 305.600 227.800 306.200 ;
        RECT 231.600 311.200 232.400 319.800 ;
        RECT 234.800 311.200 235.600 319.800 ;
        RECT 238.000 311.600 238.800 313.200 ;
        RECT 231.600 310.400 235.600 311.200 ;
        RECT 231.600 307.600 232.400 310.400 ;
        RECT 239.600 310.300 240.400 319.800 ;
        RECT 245.400 312.400 246.200 319.800 ;
        RECT 255.600 316.400 256.400 319.800 ;
        RECT 255.400 315.800 256.400 316.400 ;
        RECT 255.400 315.200 256.000 315.800 ;
        RECT 258.800 315.200 259.600 319.800 ;
        RECT 262.000 317.000 262.800 319.800 ;
        RECT 263.600 317.000 264.400 319.800 ;
        RECT 254.000 314.600 256.000 315.200 ;
        RECT 246.800 314.300 247.600 314.400 ;
        RECT 252.400 314.300 253.200 314.400 ;
        RECT 246.800 313.700 253.200 314.300 ;
        RECT 246.800 313.600 247.600 313.700 ;
        RECT 252.400 313.600 253.200 313.700 ;
        RECT 247.000 312.400 247.600 313.600 ;
        RECT 245.400 311.800 246.400 312.400 ;
        RECT 247.000 311.800 248.400 312.400 ;
        RECT 242.800 310.300 243.600 310.400 ;
        RECT 239.600 309.700 243.600 310.300 ;
        RECT 231.600 306.800 235.600 307.600 ;
        RECT 226.800 302.200 227.600 305.600 ;
        RECT 231.600 302.200 232.400 306.800 ;
        RECT 234.800 302.200 235.600 306.800 ;
        RECT 239.600 306.200 240.400 309.700 ;
        RECT 242.800 309.600 243.600 309.700 ;
        RECT 244.400 308.800 245.200 310.400 ;
        RECT 245.800 308.400 246.400 311.800 ;
        RECT 247.600 311.600 248.400 311.800 ;
        RECT 254.000 309.000 254.800 314.600 ;
        RECT 256.600 314.400 260.800 315.200 ;
        RECT 265.200 315.000 266.000 319.800 ;
        RECT 268.400 315.000 269.200 319.800 ;
        RECT 256.600 314.000 257.200 314.400 ;
        RECT 255.600 313.200 257.200 314.000 ;
        RECT 260.200 313.800 266.000 314.400 ;
        RECT 258.200 313.200 259.600 313.800 ;
        RECT 258.200 313.000 264.400 313.200 ;
        RECT 259.000 312.600 264.400 313.000 ;
        RECT 263.600 312.400 264.400 312.600 ;
        RECT 265.400 313.000 266.000 313.800 ;
        RECT 266.600 313.600 269.200 314.400 ;
        RECT 271.600 313.600 272.400 319.800 ;
        RECT 273.200 317.000 274.000 319.800 ;
        RECT 274.800 317.000 275.600 319.800 ;
        RECT 276.400 317.000 277.200 319.800 ;
        RECT 274.800 314.400 279.000 315.200 ;
        RECT 279.600 314.400 280.400 319.800 ;
        RECT 282.800 315.200 283.600 319.800 ;
        RECT 282.800 314.600 285.400 315.200 ;
        RECT 279.600 313.600 282.200 314.400 ;
        RECT 273.200 313.000 274.000 313.200 ;
        RECT 265.400 312.400 274.000 313.000 ;
        RECT 276.400 313.000 277.200 313.200 ;
        RECT 284.800 313.000 285.400 314.600 ;
        RECT 276.400 312.400 285.400 313.000 ;
        RECT 284.800 310.600 285.400 312.400 ;
        RECT 286.000 312.000 286.800 319.800 ;
        RECT 286.000 311.200 287.000 312.000 ;
        RECT 255.400 310.000 278.800 310.600 ;
        RECT 284.800 310.000 285.600 310.600 ;
        RECT 255.400 309.800 256.200 310.000 ;
        RECT 257.200 309.600 258.000 310.000 ;
        RECT 260.400 309.600 261.200 310.000 ;
        RECT 278.000 309.400 278.800 310.000 ;
        RECT 241.200 306.800 242.000 308.400 ;
        RECT 242.800 308.200 243.600 308.400 ;
        RECT 242.800 307.600 244.400 308.200 ;
        RECT 245.800 307.600 248.400 308.400 ;
        RECT 254.000 308.200 262.800 309.000 ;
        RECT 263.400 308.600 265.400 309.400 ;
        RECT 269.200 308.600 272.400 309.400 ;
        RECT 243.600 307.200 244.400 307.600 ;
        RECT 243.000 306.200 246.600 306.600 ;
        RECT 247.600 306.200 248.200 307.600 ;
        RECT 238.600 305.600 240.400 306.200 ;
        RECT 242.800 306.000 246.800 306.200 ;
        RECT 238.600 302.200 239.400 305.600 ;
        RECT 242.800 302.200 243.600 306.000 ;
        RECT 246.000 302.200 246.800 306.000 ;
        RECT 247.600 302.200 248.400 306.200 ;
        RECT 254.000 302.200 254.800 308.200 ;
        RECT 256.400 306.800 259.400 307.600 ;
        RECT 258.600 306.200 259.400 306.800 ;
        RECT 264.600 306.200 265.400 308.600 ;
        RECT 266.800 306.800 267.600 308.400 ;
        RECT 272.000 307.800 272.800 308.000 ;
        RECT 268.400 307.200 272.800 307.800 ;
        RECT 268.400 307.000 269.200 307.200 ;
        RECT 274.800 306.400 275.600 309.200 ;
        RECT 280.600 308.600 284.400 309.400 ;
        RECT 280.600 307.400 281.400 308.600 ;
        RECT 285.000 308.000 285.600 310.000 ;
        RECT 268.400 306.200 269.200 306.400 ;
        RECT 258.600 305.400 261.200 306.200 ;
        RECT 264.600 305.600 269.200 306.200 ;
        RECT 270.000 305.600 271.600 306.400 ;
        RECT 274.600 305.600 275.600 306.400 ;
        RECT 279.600 306.800 281.400 307.400 ;
        RECT 284.400 307.400 285.600 308.000 ;
        RECT 279.600 306.200 280.400 306.800 ;
        RECT 260.400 302.200 261.200 305.400 ;
        RECT 278.000 305.400 280.400 306.200 ;
        RECT 262.000 302.200 262.800 305.000 ;
        RECT 263.600 302.200 264.400 305.000 ;
        RECT 265.200 302.200 266.000 305.000 ;
        RECT 268.400 302.200 269.200 305.000 ;
        RECT 271.600 302.200 272.400 305.000 ;
        RECT 273.200 302.200 274.000 305.000 ;
        RECT 274.800 302.200 275.600 305.000 ;
        RECT 276.400 302.200 277.200 305.000 ;
        RECT 278.000 302.200 278.800 305.400 ;
        RECT 284.400 302.200 285.200 307.400 ;
        RECT 286.200 306.800 287.000 311.200 ;
        RECT 286.000 306.000 287.000 306.800 ;
        RECT 286.000 302.200 286.800 306.000 ;
        RECT 290.800 302.200 291.600 319.800 ;
        RECT 294.000 311.600 294.800 313.200 ;
        RECT 295.600 306.200 296.400 319.800 ;
        RECT 301.400 312.400 302.200 319.800 ;
        RECT 302.800 313.600 303.600 314.400 ;
        RECT 303.000 312.400 303.600 313.600 ;
        RECT 300.400 311.600 302.400 312.400 ;
        RECT 303.000 311.800 304.400 312.400 ;
        RECT 303.600 311.600 304.400 311.800 ;
        RECT 300.400 308.800 301.200 310.400 ;
        RECT 301.800 308.400 302.400 311.600 ;
        RECT 303.600 310.300 304.400 310.400 ;
        RECT 305.200 310.300 306.000 319.800 ;
        RECT 303.600 309.700 306.000 310.300 ;
        RECT 303.600 309.600 304.400 309.700 ;
        RECT 297.200 306.800 298.000 308.400 ;
        RECT 298.800 308.200 299.600 308.400 ;
        RECT 298.800 307.600 300.400 308.200 ;
        RECT 301.800 307.600 304.400 308.400 ;
        RECT 299.600 307.200 300.400 307.600 ;
        RECT 299.000 306.200 302.600 306.600 ;
        RECT 303.600 306.200 304.200 307.600 ;
        RECT 294.600 305.600 296.400 306.200 ;
        RECT 298.800 306.000 302.800 306.200 ;
        RECT 294.600 302.200 295.400 305.600 ;
        RECT 298.800 302.200 299.600 306.000 ;
        RECT 302.000 302.200 302.800 306.000 ;
        RECT 303.600 302.200 304.400 306.200 ;
        RECT 305.200 302.200 306.000 309.700 ;
        RECT 310.000 310.300 310.800 319.800 ;
        RECT 313.200 315.800 314.000 319.800 ;
        RECT 313.400 315.600 314.000 315.800 ;
        RECT 316.400 315.800 317.200 319.800 ;
        RECT 316.400 315.600 317.000 315.800 ;
        RECT 313.400 315.000 317.000 315.600 ;
        RECT 311.600 311.600 312.400 313.200 ;
        RECT 313.400 312.400 314.000 315.000 ;
        RECT 314.800 312.800 315.600 314.400 ;
        RECT 313.200 311.600 314.000 312.400 ;
        RECT 311.600 310.300 312.400 310.400 ;
        RECT 310.000 309.700 312.400 310.300 ;
        RECT 308.400 306.800 309.200 308.400 ;
        RECT 306.800 304.800 307.600 306.400 ;
        RECT 310.000 306.200 310.800 309.700 ;
        RECT 311.600 309.600 312.400 309.700 ;
        RECT 313.400 308.400 314.000 311.600 ;
        RECT 318.000 310.800 318.800 312.400 ;
        RECT 319.600 311.600 320.400 313.200 ;
        RECT 315.600 309.600 317.200 310.400 ;
        RECT 313.400 308.200 315.000 308.400 ;
        RECT 313.400 307.800 315.200 308.200 ;
        RECT 310.000 305.600 311.800 306.200 ;
        RECT 311.000 302.200 311.800 305.600 ;
        RECT 314.400 302.200 315.200 307.800 ;
        RECT 321.200 306.200 322.000 319.800 ;
        RECT 324.400 312.400 325.200 319.800 ;
        RECT 327.600 312.800 328.400 319.800 ;
        RECT 332.400 315.800 333.200 319.800 ;
        RECT 332.600 315.600 333.200 315.800 ;
        RECT 335.600 315.800 336.400 319.800 ;
        RECT 335.600 315.600 336.200 315.800 ;
        RECT 332.600 315.000 336.200 315.600 ;
        RECT 334.000 312.800 334.800 314.400 ;
        RECT 324.400 311.800 327.000 312.400 ;
        RECT 324.400 309.600 325.400 310.400 ;
        RECT 324.600 308.800 325.400 309.600 ;
        RECT 326.400 309.800 327.000 311.800 ;
        RECT 327.600 311.600 328.600 312.800 ;
        RECT 335.600 312.400 336.200 315.000 ;
        RECT 338.800 312.800 339.600 319.800 ;
        RECT 326.400 309.000 327.400 309.800 ;
        RECT 322.800 306.800 323.600 308.400 ;
        RECT 326.400 307.400 327.000 309.000 ;
        RECT 328.000 308.400 328.600 311.600 ;
        RECT 330.800 310.800 331.600 312.400 ;
        RECT 335.600 311.600 336.400 312.400 ;
        RECT 338.600 311.800 339.600 312.800 ;
        RECT 342.000 312.400 342.800 319.800 ;
        RECT 340.200 311.800 342.800 312.400 ;
        RECT 335.600 308.400 336.200 311.600 ;
        RECT 338.600 308.400 339.200 311.800 ;
        RECT 340.200 309.800 340.800 311.800 ;
        RECT 339.800 309.000 340.800 309.800 ;
        RECT 327.600 307.600 328.600 308.400 ;
        RECT 334.600 308.200 336.200 308.400 ;
        RECT 324.400 306.800 327.000 307.400 ;
        RECT 320.200 305.600 322.000 306.200 ;
        RECT 320.200 302.200 321.000 305.600 ;
        RECT 324.400 302.200 325.200 306.800 ;
        RECT 328.000 306.200 328.600 307.600 ;
        RECT 327.600 305.600 328.600 306.200 ;
        RECT 334.400 307.800 336.200 308.200 ;
        RECT 337.200 308.300 338.000 308.400 ;
        RECT 338.600 308.300 339.600 308.400 ;
        RECT 327.600 302.200 328.400 305.600 ;
        RECT 332.400 304.300 333.200 304.400 ;
        RECT 334.400 304.300 335.200 307.800 ;
        RECT 337.200 307.700 339.600 308.300 ;
        RECT 337.200 307.600 338.000 307.700 ;
        RECT 338.600 307.600 339.600 307.700 ;
        RECT 338.600 306.200 339.200 307.600 ;
        RECT 340.200 307.400 340.800 309.000 ;
        RECT 341.800 309.600 342.800 310.400 ;
        RECT 345.200 310.300 346.000 319.800 ;
        RECT 348.400 310.300 349.200 310.400 ;
        RECT 345.200 309.700 349.200 310.300 ;
        RECT 341.800 308.800 342.600 309.600 ;
        RECT 340.200 306.800 342.800 307.400 ;
        RECT 343.600 306.800 344.400 308.400 ;
        RECT 338.600 305.600 339.600 306.200 ;
        RECT 332.400 303.700 335.200 304.300 ;
        RECT 332.400 303.600 333.200 303.700 ;
        RECT 334.400 302.200 335.200 303.700 ;
        RECT 338.800 302.200 339.600 305.600 ;
        RECT 342.000 302.200 342.800 306.800 ;
        RECT 345.200 302.200 346.000 309.700 ;
        RECT 348.400 309.600 349.200 309.700 ;
        RECT 350.000 310.300 350.800 319.800 ;
        RECT 355.800 311.800 357.800 319.800 ;
        RECT 363.800 312.400 364.600 319.800 ;
        RECT 365.200 313.600 366.000 314.400 ;
        RECT 365.400 312.400 366.000 313.600 ;
        RECT 354.800 310.300 355.600 310.400 ;
        RECT 350.000 309.700 355.600 310.300 ;
        RECT 346.800 308.300 347.600 308.400 ;
        RECT 348.400 308.300 349.200 308.400 ;
        RECT 346.800 307.700 349.200 308.300 ;
        RECT 346.800 307.600 347.600 307.700 ;
        RECT 348.400 306.800 349.200 307.700 ;
        RECT 350.000 306.200 350.800 309.700 ;
        RECT 354.800 308.800 355.600 309.700 ;
        RECT 356.400 308.400 357.000 311.800 ;
        RECT 362.800 311.600 364.800 312.400 ;
        RECT 365.400 312.300 366.800 312.400 ;
        RECT 369.200 312.300 370.000 319.800 ;
        RECT 372.400 315.200 373.200 319.800 ;
        RECT 365.400 311.800 370.000 312.300 ;
        RECT 366.000 311.700 370.000 311.800 ;
        RECT 366.000 311.600 366.800 311.700 ;
        RECT 358.000 308.800 358.800 310.400 ;
        RECT 353.200 308.200 354.000 308.400 ;
        RECT 356.400 308.200 357.200 308.400 ;
        RECT 353.200 307.600 354.800 308.200 ;
        RECT 356.400 307.600 358.800 308.200 ;
        RECT 359.600 307.600 360.400 309.200 ;
        RECT 362.800 308.800 363.600 310.400 ;
        RECT 364.200 308.400 364.800 311.600 ;
        RECT 369.000 311.200 370.000 311.700 ;
        RECT 370.600 314.600 373.200 315.200 ;
        RECT 370.600 313.000 371.200 314.600 ;
        RECT 375.600 314.400 376.400 319.800 ;
        RECT 378.800 317.000 379.600 319.800 ;
        RECT 380.400 317.000 381.200 319.800 ;
        RECT 382.000 317.000 382.800 319.800 ;
        RECT 377.000 314.400 381.200 315.200 ;
        RECT 373.800 313.600 376.400 314.400 ;
        RECT 383.600 313.600 384.400 319.800 ;
        RECT 386.800 315.000 387.600 319.800 ;
        RECT 390.000 315.000 390.800 319.800 ;
        RECT 391.600 317.000 392.400 319.800 ;
        RECT 393.200 317.000 394.000 319.800 ;
        RECT 396.400 315.200 397.200 319.800 ;
        RECT 399.600 316.400 400.400 319.800 ;
        RECT 409.200 316.400 410.000 319.800 ;
        RECT 399.600 315.800 400.600 316.400 ;
        RECT 400.000 315.200 400.600 315.800 ;
        RECT 409.000 315.800 410.000 316.400 ;
        RECT 409.000 315.200 409.600 315.800 ;
        RECT 412.400 315.200 413.200 319.800 ;
        RECT 415.600 317.000 416.400 319.800 ;
        RECT 417.200 317.000 418.000 319.800 ;
        RECT 395.200 314.400 399.400 315.200 ;
        RECT 400.000 314.600 402.000 315.200 ;
        RECT 386.800 313.600 389.400 314.400 ;
        RECT 390.000 313.800 395.800 314.400 ;
        RECT 398.800 314.000 399.400 314.400 ;
        RECT 378.800 313.000 379.600 313.200 ;
        RECT 370.600 312.400 379.600 313.000 ;
        RECT 382.000 313.000 382.800 313.200 ;
        RECT 390.000 313.000 390.600 313.800 ;
        RECT 396.400 313.200 397.800 313.800 ;
        RECT 398.800 313.200 400.400 314.000 ;
        RECT 382.000 312.400 390.600 313.000 ;
        RECT 391.600 313.000 397.800 313.200 ;
        RECT 391.600 312.600 397.000 313.000 ;
        RECT 391.600 312.400 392.400 312.600 ;
        RECT 361.200 308.200 362.000 308.400 ;
        RECT 361.200 307.600 362.800 308.200 ;
        RECT 364.200 307.600 366.800 308.400 ;
        RECT 354.000 307.200 354.800 307.600 ;
        RECT 353.400 306.200 357.000 306.600 ;
        RECT 358.200 306.400 358.800 307.600 ;
        RECT 362.000 307.200 362.800 307.600 ;
        RECT 350.000 305.600 351.800 306.200 ;
        RECT 351.000 302.200 351.800 305.600 ;
        RECT 353.200 306.000 357.200 306.200 ;
        RECT 353.200 302.200 354.000 306.000 ;
        RECT 356.400 302.800 357.200 306.000 ;
        RECT 358.000 303.400 358.800 306.400 ;
        RECT 361.400 306.200 365.000 306.600 ;
        RECT 366.000 306.200 366.600 307.600 ;
        RECT 369.000 306.800 369.800 311.200 ;
        RECT 370.600 310.600 371.200 312.400 ;
        RECT 370.400 310.000 371.200 310.600 ;
        RECT 377.200 310.000 400.600 310.600 ;
        RECT 370.400 308.000 371.000 310.000 ;
        RECT 377.200 309.400 378.000 310.000 ;
        RECT 394.800 309.600 395.600 310.000 ;
        RECT 399.800 309.800 400.600 310.000 ;
        RECT 371.600 308.600 375.400 309.400 ;
        RECT 370.400 307.400 371.600 308.000 ;
        RECT 359.600 302.800 360.400 306.200 ;
        RECT 356.400 302.200 360.400 302.800 ;
        RECT 361.200 306.000 365.200 306.200 ;
        RECT 361.200 302.200 362.000 306.000 ;
        RECT 364.400 302.200 365.200 306.000 ;
        RECT 366.000 302.200 366.800 306.200 ;
        RECT 369.000 306.000 370.000 306.800 ;
        RECT 369.200 302.200 370.000 306.000 ;
        RECT 370.800 302.200 371.600 307.400 ;
        RECT 374.600 307.400 375.400 308.600 ;
        RECT 374.600 306.800 376.400 307.400 ;
        RECT 375.600 306.200 376.400 306.800 ;
        RECT 380.400 306.400 381.200 309.200 ;
        RECT 383.600 308.600 386.800 309.400 ;
        RECT 390.600 308.600 392.600 309.400 ;
        RECT 401.200 309.000 402.000 314.600 ;
        RECT 383.200 307.800 384.000 308.000 ;
        RECT 383.200 307.200 387.600 307.800 ;
        RECT 386.800 307.000 387.600 307.200 ;
        RECT 388.400 306.800 389.200 308.400 ;
        RECT 375.600 305.400 378.000 306.200 ;
        RECT 380.400 305.600 381.400 306.400 ;
        RECT 384.400 305.600 386.000 306.400 ;
        RECT 386.800 306.200 387.600 306.400 ;
        RECT 390.600 306.200 391.400 308.600 ;
        RECT 393.200 308.200 402.000 309.000 ;
        RECT 396.600 306.800 399.600 307.600 ;
        RECT 396.600 306.200 397.400 306.800 ;
        RECT 386.800 305.600 391.400 306.200 ;
        RECT 377.200 302.200 378.000 305.400 ;
        RECT 394.800 305.400 397.400 306.200 ;
        RECT 378.800 302.200 379.600 305.000 ;
        RECT 380.400 302.200 381.200 305.000 ;
        RECT 382.000 302.200 382.800 305.000 ;
        RECT 383.600 302.200 384.400 305.000 ;
        RECT 386.800 302.200 387.600 305.000 ;
        RECT 390.000 302.200 390.800 305.000 ;
        RECT 391.600 302.200 392.400 305.000 ;
        RECT 393.200 302.200 394.000 305.000 ;
        RECT 394.800 302.200 395.600 305.400 ;
        RECT 401.200 302.200 402.000 308.200 ;
        RECT 407.600 314.600 409.600 315.200 ;
        RECT 407.600 309.000 408.400 314.600 ;
        RECT 410.200 314.400 414.400 315.200 ;
        RECT 418.800 315.000 419.600 319.800 ;
        RECT 422.000 315.000 422.800 319.800 ;
        RECT 410.200 314.000 410.800 314.400 ;
        RECT 409.200 313.200 410.800 314.000 ;
        RECT 413.800 313.800 419.600 314.400 ;
        RECT 411.800 313.200 413.200 313.800 ;
        RECT 411.800 313.000 418.000 313.200 ;
        RECT 412.600 312.600 418.000 313.000 ;
        RECT 417.200 312.400 418.000 312.600 ;
        RECT 419.000 313.000 419.600 313.800 ;
        RECT 420.200 313.600 422.800 314.400 ;
        RECT 425.200 313.600 426.000 319.800 ;
        RECT 426.800 317.000 427.600 319.800 ;
        RECT 428.400 317.000 429.200 319.800 ;
        RECT 430.000 317.000 430.800 319.800 ;
        RECT 428.400 314.400 432.600 315.200 ;
        RECT 433.200 314.400 434.000 319.800 ;
        RECT 436.400 315.200 437.200 319.800 ;
        RECT 436.400 314.600 439.000 315.200 ;
        RECT 433.200 313.600 435.800 314.400 ;
        RECT 426.800 313.000 427.600 313.200 ;
        RECT 419.000 312.400 427.600 313.000 ;
        RECT 430.000 313.000 430.800 313.200 ;
        RECT 438.400 313.000 439.000 314.600 ;
        RECT 430.000 312.400 439.000 313.000 ;
        RECT 438.400 310.600 439.000 312.400 ;
        RECT 439.600 312.000 440.400 319.800 ;
        RECT 439.600 311.200 440.600 312.000 ;
        RECT 409.000 310.000 432.400 310.600 ;
        RECT 438.400 310.000 439.200 310.600 ;
        RECT 409.000 309.800 409.800 310.000 ;
        RECT 410.800 309.600 411.600 310.000 ;
        RECT 414.000 309.600 414.800 310.000 ;
        RECT 431.600 309.400 432.400 310.000 ;
        RECT 407.600 308.200 416.400 309.000 ;
        RECT 417.000 308.600 419.000 309.400 ;
        RECT 422.800 308.600 426.000 309.400 ;
        RECT 407.600 302.200 408.400 308.200 ;
        RECT 410.000 306.800 413.000 307.600 ;
        RECT 412.200 306.200 413.000 306.800 ;
        RECT 418.200 306.200 419.000 308.600 ;
        RECT 420.400 306.800 421.200 308.400 ;
        RECT 425.600 307.800 426.400 308.000 ;
        RECT 422.000 307.200 426.400 307.800 ;
        RECT 422.000 307.000 422.800 307.200 ;
        RECT 428.400 306.400 429.200 309.200 ;
        RECT 434.200 308.600 438.000 309.400 ;
        RECT 434.200 307.400 435.000 308.600 ;
        RECT 438.600 308.000 439.200 310.000 ;
        RECT 422.000 306.200 422.800 306.400 ;
        RECT 412.200 305.400 414.800 306.200 ;
        RECT 418.200 305.600 422.800 306.200 ;
        RECT 423.600 305.600 425.200 306.400 ;
        RECT 428.200 305.600 429.200 306.400 ;
        RECT 433.200 306.800 435.000 307.400 ;
        RECT 438.000 307.400 439.200 308.000 ;
        RECT 433.200 306.200 434.000 306.800 ;
        RECT 414.000 302.200 414.800 305.400 ;
        RECT 431.600 305.400 434.000 306.200 ;
        RECT 415.600 302.200 416.400 305.000 ;
        RECT 417.200 302.200 418.000 305.000 ;
        RECT 418.800 302.200 419.600 305.000 ;
        RECT 422.000 302.200 422.800 305.000 ;
        RECT 425.200 302.200 426.000 305.000 ;
        RECT 426.800 302.200 427.600 305.000 ;
        RECT 428.400 302.200 429.200 305.000 ;
        RECT 430.000 302.200 430.800 305.000 ;
        RECT 431.600 302.200 432.400 305.400 ;
        RECT 438.000 302.200 438.800 307.400 ;
        RECT 439.800 306.800 440.600 311.200 ;
        RECT 439.600 306.000 440.600 306.800 ;
        RECT 441.200 306.300 442.000 306.400 ;
        RECT 442.800 306.300 443.600 306.400 ;
        RECT 439.600 302.200 440.400 306.000 ;
        RECT 441.200 305.700 443.600 306.300 ;
        RECT 441.200 305.600 442.000 305.700 ;
        RECT 442.800 304.800 443.600 305.700 ;
        RECT 444.400 302.200 445.200 319.800 ;
        RECT 446.000 311.400 446.800 319.800 ;
        RECT 450.400 316.400 451.200 319.800 ;
        RECT 449.200 315.800 451.200 316.400 ;
        RECT 454.800 315.800 455.600 319.800 ;
        RECT 459.000 315.800 460.200 319.800 ;
        RECT 449.200 315.000 450.000 315.800 ;
        RECT 454.800 315.200 455.400 315.800 ;
        RECT 452.600 314.600 456.200 315.200 ;
        RECT 458.800 315.000 459.600 315.800 ;
        RECT 452.600 314.400 453.400 314.600 ;
        RECT 455.400 314.400 456.200 314.600 ;
        RECT 463.600 314.300 464.400 319.800 ;
        RECT 465.200 314.300 466.000 314.400 ;
        RECT 449.200 313.000 450.000 313.200 ;
        RECT 453.800 313.000 454.600 313.200 ;
        RECT 449.200 312.400 454.600 313.000 ;
        RECT 455.200 313.000 457.400 313.600 ;
        RECT 455.200 311.800 455.800 313.000 ;
        RECT 456.600 312.800 457.400 313.000 ;
        RECT 459.000 313.200 460.400 314.000 ;
        RECT 463.600 313.700 466.000 314.300 ;
        RECT 459.000 312.200 459.600 313.200 ;
        RECT 451.000 311.400 455.800 311.800 ;
        RECT 446.000 311.200 455.800 311.400 ;
        RECT 457.200 311.600 459.600 312.200 ;
        RECT 446.000 311.000 451.800 311.200 ;
        RECT 446.000 310.800 451.600 311.000 ;
        RECT 452.400 310.200 453.200 310.400 ;
        RECT 448.200 309.600 453.200 310.200 ;
        RECT 448.200 309.400 449.000 309.600 ;
        RECT 449.800 308.400 450.600 308.600 ;
        RECT 457.200 308.400 457.800 311.600 ;
        RECT 463.600 311.200 464.400 313.700 ;
        RECT 465.200 313.600 466.000 313.700 ;
        RECT 460.200 310.600 464.400 311.200 ;
        RECT 460.200 310.400 461.000 310.600 ;
        RECT 461.800 309.800 462.600 310.000 ;
        RECT 458.800 309.200 462.600 309.800 ;
        RECT 458.800 309.000 459.600 309.200 ;
        RECT 446.800 307.800 457.800 308.400 ;
        RECT 446.800 307.600 448.400 307.800 ;
        RECT 446.000 302.200 446.800 307.000 ;
        RECT 451.000 305.600 451.600 307.800 ;
        RECT 456.600 307.600 457.400 307.800 ;
        RECT 463.600 307.200 464.400 310.600 ;
        RECT 460.600 306.600 464.400 307.200 ;
        RECT 460.600 306.400 461.400 306.600 ;
        RECT 449.200 304.200 450.000 305.000 ;
        RECT 450.800 304.800 451.600 305.600 ;
        RECT 452.600 305.400 453.400 305.600 ;
        RECT 452.600 304.800 455.400 305.400 ;
        RECT 454.800 304.200 455.400 304.800 ;
        RECT 458.800 304.200 459.600 305.000 ;
        RECT 449.200 303.600 451.200 304.200 ;
        RECT 450.400 302.200 451.200 303.600 ;
        RECT 454.800 302.200 455.600 304.200 ;
        RECT 458.800 303.600 460.200 304.200 ;
        RECT 459.000 302.200 460.200 303.600 ;
        RECT 463.600 302.200 464.400 306.600 ;
        RECT 465.200 304.800 466.000 306.400 ;
        RECT 466.800 302.200 467.600 319.800 ;
        RECT 471.000 312.400 471.800 319.800 ;
        RECT 472.400 313.600 473.200 314.400 ;
        RECT 472.600 312.400 473.200 313.600 ;
        RECT 478.600 312.800 479.400 319.800 ;
        RECT 482.800 315.000 483.600 319.000 ;
        RECT 487.000 318.400 487.800 319.800 ;
        RECT 486.000 317.600 487.800 318.400 ;
        RECT 471.000 311.800 472.000 312.400 ;
        RECT 472.600 311.800 474.000 312.400 ;
        RECT 470.000 308.800 470.800 310.400 ;
        RECT 471.400 308.400 472.000 311.800 ;
        RECT 473.200 311.600 474.000 311.800 ;
        RECT 477.800 312.200 479.400 312.800 ;
        RECT 474.800 310.300 475.600 310.400 ;
        RECT 476.400 310.300 477.200 311.200 ;
        RECT 474.800 309.700 477.200 310.300 ;
        RECT 474.800 309.600 475.600 309.700 ;
        RECT 476.400 309.600 477.200 309.700 ;
        RECT 477.800 308.400 478.400 312.200 ;
        RECT 483.000 311.600 483.600 315.000 ;
        RECT 487.000 312.400 487.800 317.600 ;
        RECT 488.400 313.600 489.200 314.400 ;
        RECT 488.600 312.400 489.200 313.600 ;
        RECT 491.600 313.600 492.400 314.400 ;
        RECT 491.600 312.400 492.200 313.600 ;
        RECT 493.000 312.400 493.800 319.800 ;
        RECT 498.000 313.600 498.800 314.400 ;
        RECT 498.000 312.400 498.600 313.600 ;
        RECT 499.400 312.400 500.200 319.800 ;
        RECT 487.000 311.800 488.000 312.400 ;
        RECT 488.600 311.800 490.000 312.400 ;
        RECT 479.800 311.000 483.600 311.600 ;
        RECT 479.800 309.000 480.400 311.000 ;
        RECT 468.400 308.200 469.200 308.400 ;
        RECT 471.400 308.300 474.000 308.400 ;
        RECT 474.800 308.300 475.600 308.400 ;
        RECT 468.400 307.600 470.000 308.200 ;
        RECT 471.400 307.700 475.600 308.300 ;
        RECT 471.400 307.600 474.000 307.700 ;
        RECT 474.800 307.600 475.600 307.700 ;
        RECT 476.400 307.600 478.400 308.400 ;
        RECT 479.000 308.200 480.400 309.000 ;
        RECT 481.200 308.800 482.000 310.400 ;
        RECT 482.800 308.800 483.600 310.400 ;
        RECT 486.000 308.800 486.800 310.400 ;
        RECT 487.400 308.400 488.000 311.800 ;
        RECT 489.200 311.600 490.000 311.800 ;
        RECT 490.800 311.800 492.200 312.400 ;
        RECT 492.800 311.800 493.800 312.400 ;
        RECT 497.200 311.800 498.600 312.400 ;
        RECT 499.200 311.800 500.200 312.400 ;
        RECT 490.800 311.600 491.600 311.800 ;
        RECT 489.300 310.300 489.900 311.600 ;
        RECT 492.800 310.300 493.400 311.800 ;
        RECT 497.200 311.600 498.000 311.800 ;
        RECT 489.300 309.700 493.400 310.300 ;
        RECT 492.800 308.400 493.400 309.700 ;
        RECT 494.000 308.800 494.800 310.400 ;
        RECT 499.200 308.400 499.800 311.800 ;
        RECT 500.400 308.800 501.200 310.400 ;
        RECT 469.200 307.200 470.000 307.600 ;
        RECT 468.600 306.200 472.200 306.600 ;
        RECT 473.200 306.200 473.800 307.600 ;
        RECT 477.800 307.000 478.400 307.600 ;
        RECT 479.400 307.800 480.400 308.200 ;
        RECT 484.400 308.200 485.200 308.400 ;
        RECT 479.400 307.200 483.600 307.800 ;
        RECT 484.400 307.600 486.000 308.200 ;
        RECT 487.400 307.600 490.000 308.400 ;
        RECT 490.800 307.600 493.400 308.400 ;
        RECT 495.600 308.200 496.400 308.400 ;
        RECT 494.800 307.600 496.400 308.200 ;
        RECT 497.200 307.600 499.800 308.400 ;
        RECT 502.000 308.200 502.800 308.400 ;
        RECT 501.200 307.600 502.800 308.200 ;
        RECT 485.200 307.200 486.000 307.600 ;
        RECT 477.800 306.600 478.600 307.000 ;
        RECT 477.800 306.400 479.400 306.600 ;
        RECT 468.400 306.000 472.400 306.200 ;
        RECT 468.400 302.200 469.200 306.000 ;
        RECT 471.600 302.200 472.400 306.000 ;
        RECT 473.200 302.200 474.000 306.200 ;
        RECT 477.800 306.000 480.400 306.400 ;
        RECT 478.600 305.600 480.400 306.000 ;
        RECT 478.600 303.000 479.400 305.600 ;
        RECT 483.000 305.000 483.600 307.200 ;
        RECT 484.600 306.200 488.200 306.600 ;
        RECT 489.200 306.200 489.800 307.600 ;
        RECT 491.000 306.200 491.600 307.600 ;
        RECT 494.800 307.200 495.600 307.600 ;
        RECT 492.600 306.200 496.200 306.600 ;
        RECT 497.400 306.200 498.000 307.600 ;
        RECT 501.200 307.200 502.000 307.600 ;
        RECT 499.000 306.200 502.600 306.600 ;
        RECT 482.800 303.000 483.600 305.000 ;
        RECT 484.400 306.000 488.400 306.200 ;
        RECT 484.400 302.200 485.200 306.000 ;
        RECT 487.600 302.200 488.400 306.000 ;
        RECT 489.200 302.200 490.000 306.200 ;
        RECT 490.800 302.200 491.600 306.200 ;
        RECT 492.400 306.000 496.400 306.200 ;
        RECT 492.400 302.200 493.200 306.000 ;
        RECT 495.600 302.200 496.400 306.000 ;
        RECT 497.200 302.200 498.000 306.200 ;
        RECT 498.800 306.000 502.800 306.200 ;
        RECT 498.800 302.200 499.600 306.000 ;
        RECT 502.000 302.200 502.800 306.000 ;
        RECT 503.600 304.800 504.400 306.400 ;
        RECT 505.200 302.200 506.000 319.800 ;
        RECT 507.600 313.600 508.400 314.400 ;
        RECT 507.600 312.400 508.200 313.600 ;
        RECT 509.000 312.400 509.800 319.800 ;
        RECT 515.800 314.400 516.600 319.800 ;
        RECT 515.800 313.600 517.200 314.400 ;
        RECT 515.800 312.600 516.600 313.600 ;
        RECT 506.800 311.800 508.200 312.400 ;
        RECT 508.800 311.800 509.800 312.400 ;
        RECT 514.800 311.800 516.600 312.600 ;
        RECT 518.000 312.400 518.800 319.800 ;
        RECT 521.200 312.800 522.000 319.800 ;
        RECT 526.000 312.800 526.800 319.800 ;
        RECT 518.000 311.800 520.600 312.400 ;
        RECT 521.200 311.800 522.200 312.800 ;
        RECT 506.800 311.600 507.600 311.800 ;
        RECT 508.800 310.400 509.400 311.800 ;
        RECT 508.400 309.600 509.400 310.400 ;
        RECT 508.800 308.400 509.400 309.600 ;
        RECT 510.000 310.300 510.800 310.400 ;
        RECT 513.200 310.300 514.000 310.400 ;
        RECT 510.000 309.700 514.000 310.300 ;
        RECT 510.000 308.800 510.800 309.700 ;
        RECT 513.200 309.600 514.000 309.700 ;
        RECT 515.000 308.400 515.600 311.800 ;
        RECT 516.400 309.600 517.200 311.200 ;
        RECT 518.000 309.600 519.000 310.400 ;
        RECT 518.200 308.800 519.000 309.600 ;
        RECT 520.000 309.800 520.600 311.800 ;
        RECT 520.000 309.000 521.000 309.800 ;
        RECT 506.800 307.600 509.400 308.400 ;
        RECT 511.600 308.300 512.400 308.400 ;
        RECT 511.600 308.200 513.900 308.300 ;
        RECT 510.800 307.700 513.900 308.200 ;
        RECT 510.800 307.600 512.400 307.700 ;
        RECT 507.000 306.200 507.600 307.600 ;
        RECT 510.800 307.200 511.600 307.600 ;
        RECT 508.600 306.200 512.200 306.600 ;
        RECT 513.300 306.400 513.900 307.700 ;
        RECT 514.800 307.600 515.600 308.400 ;
        RECT 506.800 302.200 507.600 306.200 ;
        RECT 508.400 306.000 512.400 306.200 ;
        RECT 508.400 302.200 509.200 306.000 ;
        RECT 511.600 302.200 512.400 306.000 ;
        RECT 513.200 304.800 514.000 306.400 ;
        RECT 515.000 304.200 515.600 307.600 ;
        RECT 520.000 307.400 520.600 309.000 ;
        RECT 521.600 308.400 522.200 311.800 ;
        RECT 525.800 311.800 526.800 312.800 ;
        RECT 529.200 312.400 530.000 319.800 ;
        RECT 527.400 311.800 530.000 312.400 ;
        RECT 533.400 312.400 534.200 319.800 ;
        RECT 539.800 318.400 540.600 319.800 ;
        RECT 538.800 317.600 540.600 318.400 ;
        RECT 534.800 313.600 535.600 314.400 ;
        RECT 535.000 312.400 535.600 313.600 ;
        RECT 539.800 312.400 540.600 317.600 ;
        RECT 541.200 313.600 542.000 314.400 ;
        RECT 541.400 312.400 542.000 313.600 ;
        RECT 543.600 312.400 544.400 319.800 ;
        RECT 546.800 312.800 547.600 319.800 ;
        RECT 552.200 318.400 553.000 319.800 ;
        RECT 552.200 317.600 554.000 318.400 ;
        RECT 550.800 313.600 551.600 314.400 ;
        RECT 533.400 311.800 534.400 312.400 ;
        RECT 535.000 311.800 536.400 312.400 ;
        RECT 539.800 311.800 540.800 312.400 ;
        RECT 541.400 311.800 542.800 312.400 ;
        RECT 543.600 311.800 546.200 312.400 ;
        RECT 546.800 311.800 547.800 312.800 ;
        RECT 550.800 312.400 551.400 313.600 ;
        RECT 552.200 312.400 553.000 317.600 ;
        RECT 525.800 308.400 526.400 311.800 ;
        RECT 527.400 309.800 528.000 311.800 ;
        RECT 527.000 309.000 528.000 309.800 ;
        RECT 521.200 308.300 522.200 308.400 ;
        RECT 522.800 308.300 523.600 308.400 ;
        RECT 521.200 307.700 523.600 308.300 ;
        RECT 521.200 307.600 522.200 307.700 ;
        RECT 522.800 307.600 523.600 307.700 ;
        RECT 525.800 307.600 526.800 308.400 ;
        RECT 514.800 302.200 515.600 304.200 ;
        RECT 518.000 306.800 520.600 307.400 ;
        RECT 518.000 302.200 518.800 306.800 ;
        RECT 521.600 306.200 522.200 307.600 ;
        RECT 521.200 305.600 522.200 306.200 ;
        RECT 525.800 306.200 526.400 307.600 ;
        RECT 527.400 307.400 528.000 309.000 ;
        RECT 529.000 309.600 530.000 310.400 ;
        RECT 529.000 308.800 529.800 309.600 ;
        RECT 532.400 308.800 533.200 310.400 ;
        RECT 533.800 308.400 534.400 311.800 ;
        RECT 535.600 311.600 536.400 311.800 ;
        RECT 538.800 308.800 539.600 310.400 ;
        RECT 540.200 308.400 540.800 311.800 ;
        RECT 542.000 311.600 542.800 311.800 ;
        RECT 543.600 309.600 544.600 310.400 ;
        RECT 543.800 308.800 544.600 309.600 ;
        RECT 545.600 309.800 546.200 311.800 ;
        RECT 545.600 309.000 546.600 309.800 ;
        RECT 530.800 308.200 531.600 308.400 ;
        RECT 533.800 308.300 536.400 308.400 ;
        RECT 537.200 308.300 538.000 308.400 ;
        RECT 533.800 308.200 538.000 308.300 ;
        RECT 530.800 307.600 532.400 308.200 ;
        RECT 533.800 307.700 538.800 308.200 ;
        RECT 533.800 307.600 536.400 307.700 ;
        RECT 537.200 307.600 538.800 307.700 ;
        RECT 540.200 307.600 542.800 308.400 ;
        RECT 527.400 306.800 530.000 307.400 ;
        RECT 531.600 307.200 532.400 307.600 ;
        RECT 525.800 305.600 526.800 306.200 ;
        RECT 521.200 302.200 522.000 305.600 ;
        RECT 526.000 302.200 526.800 305.600 ;
        RECT 529.200 302.200 530.000 306.800 ;
        RECT 531.000 306.200 534.600 306.600 ;
        RECT 535.600 306.200 536.200 307.600 ;
        RECT 538.000 307.200 538.800 307.600 ;
        RECT 537.400 306.200 541.000 306.600 ;
        RECT 542.000 306.200 542.600 307.600 ;
        RECT 545.600 307.400 546.200 309.000 ;
        RECT 547.200 308.400 547.800 311.800 ;
        RECT 550.000 311.800 551.400 312.400 ;
        RECT 552.000 311.800 553.000 312.400 ;
        RECT 559.000 312.400 559.800 319.800 ;
        RECT 560.400 313.600 561.200 314.400 ;
        RECT 560.600 312.400 561.200 313.600 ;
        RECT 563.600 313.600 564.400 314.400 ;
        RECT 563.600 312.400 564.200 313.600 ;
        RECT 565.000 312.400 565.800 319.800 ;
        RECT 559.000 311.800 560.000 312.400 ;
        RECT 560.600 311.800 562.000 312.400 ;
        RECT 550.000 311.600 550.800 311.800 ;
        RECT 552.000 308.400 552.600 311.800 ;
        RECT 553.200 308.800 554.000 310.400 ;
        RECT 558.000 308.800 558.800 310.400 ;
        RECT 559.400 308.400 560.000 311.800 ;
        RECT 561.200 311.600 562.000 311.800 ;
        RECT 562.800 311.800 564.200 312.400 ;
        RECT 564.800 311.800 565.800 312.400 ;
        RECT 562.800 311.600 563.600 311.800 ;
        RECT 564.800 308.400 565.400 311.800 ;
        RECT 566.000 310.300 566.800 310.400 ;
        RECT 567.600 310.300 568.400 310.400 ;
        RECT 566.000 309.700 568.400 310.300 ;
        RECT 566.000 308.800 566.800 309.700 ;
        RECT 567.600 309.600 568.400 309.700 ;
        RECT 546.800 307.600 547.800 308.400 ;
        RECT 550.000 307.600 552.600 308.400 ;
        RECT 554.800 308.200 555.600 308.400 ;
        RECT 554.000 307.600 555.600 308.200 ;
        RECT 556.400 308.200 557.200 308.400 ;
        RECT 556.400 307.600 558.000 308.200 ;
        RECT 559.400 307.600 562.000 308.400 ;
        RECT 562.800 307.600 565.400 308.400 ;
        RECT 567.600 308.300 568.400 308.400 ;
        RECT 569.200 308.300 570.000 319.800 ;
        RECT 577.200 311.400 578.000 319.800 ;
        RECT 581.600 316.400 582.400 319.800 ;
        RECT 580.400 315.800 582.400 316.400 ;
        RECT 586.000 315.800 586.800 319.800 ;
        RECT 590.200 315.800 591.400 319.800 ;
        RECT 580.400 315.000 581.200 315.800 ;
        RECT 586.000 315.200 586.600 315.800 ;
        RECT 583.800 314.600 587.400 315.200 ;
        RECT 590.000 315.000 590.800 315.800 ;
        RECT 583.800 314.400 584.600 314.600 ;
        RECT 586.600 314.400 587.400 314.600 ;
        RECT 580.400 313.000 581.200 313.200 ;
        RECT 585.000 313.000 585.800 313.200 ;
        RECT 580.400 312.400 585.800 313.000 ;
        RECT 586.400 313.000 588.600 313.600 ;
        RECT 586.400 311.800 587.000 313.000 ;
        RECT 587.800 312.800 588.600 313.000 ;
        RECT 590.200 313.200 591.600 314.000 ;
        RECT 590.200 312.200 590.800 313.200 ;
        RECT 582.200 311.400 587.000 311.800 ;
        RECT 577.200 311.200 587.000 311.400 ;
        RECT 588.400 311.600 590.800 312.200 ;
        RECT 577.200 311.000 583.000 311.200 ;
        RECT 577.200 310.800 582.800 311.000 ;
        RECT 583.600 310.200 584.400 310.400 ;
        RECT 579.400 309.600 584.400 310.200 ;
        RECT 579.400 309.400 580.200 309.600 ;
        RECT 581.000 308.400 581.800 308.600 ;
        RECT 588.400 308.400 589.000 311.600 ;
        RECT 594.800 311.200 595.600 319.800 ;
        RECT 599.000 312.400 599.800 319.800 ;
        RECT 600.400 313.600 601.200 314.400 ;
        RECT 600.600 312.400 601.200 313.600 ;
        RECT 603.600 313.600 604.400 314.400 ;
        RECT 603.600 312.400 604.200 313.600 ;
        RECT 605.000 312.400 605.800 319.800 ;
        RECT 599.000 311.800 600.000 312.400 ;
        RECT 600.600 311.800 602.000 312.400 ;
        RECT 591.400 310.600 595.600 311.200 ;
        RECT 591.400 310.400 592.200 310.600 ;
        RECT 593.000 309.800 593.800 310.000 ;
        RECT 590.000 309.200 593.800 309.800 ;
        RECT 590.000 309.000 590.800 309.200 ;
        RECT 567.600 308.200 570.000 308.300 ;
        RECT 566.800 307.700 570.000 308.200 ;
        RECT 566.800 307.600 568.400 307.700 ;
        RECT 543.600 306.800 546.200 307.400 ;
        RECT 530.800 306.000 534.800 306.200 ;
        RECT 530.800 302.200 531.600 306.000 ;
        RECT 534.000 302.200 534.800 306.000 ;
        RECT 535.600 302.200 536.400 306.200 ;
        RECT 537.200 306.000 541.200 306.200 ;
        RECT 537.200 302.200 538.000 306.000 ;
        RECT 540.400 302.200 541.200 306.000 ;
        RECT 542.000 302.200 542.800 306.200 ;
        RECT 543.600 302.200 544.400 306.800 ;
        RECT 547.200 306.200 547.800 307.600 ;
        RECT 550.200 306.200 550.800 307.600 ;
        RECT 554.000 307.200 554.800 307.600 ;
        RECT 557.200 307.200 558.000 307.600 ;
        RECT 551.800 306.200 555.400 306.600 ;
        RECT 556.600 306.200 560.200 306.600 ;
        RECT 561.200 306.200 561.800 307.600 ;
        RECT 563.000 306.200 563.600 307.600 ;
        RECT 566.800 307.200 567.600 307.600 ;
        RECT 564.600 306.200 568.200 306.600 ;
        RECT 546.800 305.600 547.800 306.200 ;
        RECT 546.800 302.200 547.600 305.600 ;
        RECT 550.000 302.200 550.800 306.200 ;
        RECT 551.600 306.000 555.600 306.200 ;
        RECT 551.600 302.200 552.400 306.000 ;
        RECT 554.800 302.200 555.600 306.000 ;
        RECT 556.400 306.000 560.400 306.200 ;
        RECT 556.400 302.200 557.200 306.000 ;
        RECT 559.600 302.200 560.400 306.000 ;
        RECT 561.200 302.200 562.000 306.200 ;
        RECT 562.800 302.200 563.600 306.200 ;
        RECT 564.400 306.000 568.400 306.200 ;
        RECT 564.400 302.200 565.200 306.000 ;
        RECT 567.600 302.200 568.400 306.000 ;
        RECT 569.200 302.200 570.000 307.700 ;
        RECT 578.000 307.800 589.000 308.400 ;
        RECT 578.000 307.600 579.600 307.800 ;
        RECT 570.800 304.800 571.600 306.400 ;
        RECT 577.200 302.200 578.000 307.000 ;
        RECT 582.200 305.600 582.800 307.800 ;
        RECT 587.800 307.600 588.600 307.800 ;
        RECT 594.800 307.200 595.600 310.600 ;
        RECT 598.000 308.800 598.800 310.400 ;
        RECT 599.400 310.300 600.000 311.800 ;
        RECT 601.200 311.600 602.000 311.800 ;
        RECT 602.800 311.800 604.200 312.400 ;
        RECT 604.800 311.800 605.800 312.400 ;
        RECT 609.200 315.000 610.000 319.000 ;
        RECT 602.800 311.600 603.600 311.800 ;
        RECT 602.900 310.300 603.500 311.600 ;
        RECT 599.400 309.700 603.500 310.300 ;
        RECT 599.400 308.400 600.000 309.700 ;
        RECT 604.800 308.400 605.400 311.800 ;
        RECT 609.200 311.600 609.800 315.000 ;
        RECT 613.400 312.800 614.200 319.800 ;
        RECT 613.400 312.200 615.000 312.800 ;
        RECT 609.200 311.000 613.000 311.600 ;
        RECT 606.000 308.800 606.800 310.400 ;
        RECT 609.200 308.800 610.000 310.400 ;
        RECT 610.800 308.800 611.600 310.400 ;
        RECT 612.400 309.000 613.000 311.000 ;
        RECT 596.400 308.200 597.200 308.400 ;
        RECT 596.400 307.600 598.000 308.200 ;
        RECT 599.400 307.600 602.000 308.400 ;
        RECT 602.800 307.600 605.400 308.400 ;
        RECT 607.600 308.200 608.400 308.400 ;
        RECT 606.800 307.600 608.400 308.200 ;
        RECT 612.400 308.200 613.800 309.000 ;
        RECT 614.400 308.400 615.000 312.200 ;
        RECT 618.800 312.400 619.600 319.800 ;
        RECT 622.000 312.800 622.800 319.800 ;
        RECT 618.800 311.800 621.400 312.400 ;
        RECT 622.000 311.800 623.000 312.800 ;
        RECT 615.600 309.600 616.400 311.200 ;
        RECT 618.800 309.600 619.800 310.400 ;
        RECT 619.000 308.800 619.800 309.600 ;
        RECT 620.800 309.800 621.400 311.800 ;
        RECT 620.800 309.000 621.800 309.800 ;
        RECT 612.400 307.800 613.400 308.200 ;
        RECT 597.200 307.200 598.000 307.600 ;
        RECT 591.800 306.600 595.600 307.200 ;
        RECT 591.800 306.400 592.600 306.600 ;
        RECT 580.400 304.200 581.200 305.000 ;
        RECT 582.000 304.800 582.800 305.600 ;
        RECT 583.800 305.400 584.600 305.600 ;
        RECT 583.800 304.800 586.600 305.400 ;
        RECT 586.000 304.200 586.600 304.800 ;
        RECT 590.000 304.200 590.800 305.000 ;
        RECT 580.400 303.600 582.400 304.200 ;
        RECT 581.600 302.200 582.400 303.600 ;
        RECT 586.000 302.200 586.800 304.200 ;
        RECT 590.000 303.600 591.400 304.200 ;
        RECT 590.200 302.200 591.400 303.600 ;
        RECT 594.800 302.200 595.600 306.600 ;
        RECT 596.600 306.200 600.200 306.600 ;
        RECT 601.200 306.200 601.800 307.600 ;
        RECT 603.000 306.200 603.600 307.600 ;
        RECT 606.800 307.200 607.600 307.600 ;
        RECT 609.200 307.200 613.400 307.800 ;
        RECT 614.400 307.600 616.400 308.400 ;
        RECT 604.600 306.200 608.200 306.600 ;
        RECT 596.400 306.000 600.400 306.200 ;
        RECT 596.400 302.200 597.200 306.000 ;
        RECT 599.600 302.200 600.400 306.000 ;
        RECT 601.200 302.200 602.000 306.200 ;
        RECT 602.800 302.200 603.600 306.200 ;
        RECT 604.400 306.000 608.400 306.200 ;
        RECT 604.400 302.200 605.200 306.000 ;
        RECT 607.600 302.200 608.400 306.000 ;
        RECT 609.200 305.000 609.800 307.200 ;
        RECT 614.400 307.000 615.000 307.600 ;
        RECT 620.800 307.400 621.400 309.000 ;
        RECT 622.400 308.400 623.000 311.800 ;
        RECT 626.800 310.300 627.600 319.800 ;
        RECT 632.200 318.400 633.000 319.800 ;
        RECT 637.000 318.400 637.800 319.800 ;
        RECT 632.200 317.600 634.000 318.400 ;
        RECT 636.400 317.600 637.800 318.400 ;
        RECT 630.800 313.600 631.600 314.400 ;
        RECT 628.400 311.600 629.200 313.200 ;
        RECT 630.800 312.400 631.400 313.600 ;
        RECT 632.200 312.400 633.000 317.600 ;
        RECT 637.000 312.400 637.800 317.600 ;
        RECT 630.000 311.800 631.400 312.400 ;
        RECT 632.000 311.800 633.000 312.400 ;
        RECT 636.400 311.800 637.800 312.400 ;
        RECT 630.000 311.600 630.800 311.800 ;
        RECT 630.100 310.300 630.700 311.600 ;
        RECT 626.800 309.700 630.700 310.300 ;
        RECT 622.000 307.600 623.000 308.400 ;
        RECT 614.200 306.600 615.000 307.000 ;
        RECT 613.400 306.400 615.000 306.600 ;
        RECT 612.400 306.000 615.000 306.400 ;
        RECT 618.800 306.800 621.400 307.400 ;
        RECT 612.400 305.600 614.200 306.000 ;
        RECT 609.200 303.000 610.000 305.000 ;
        RECT 613.400 303.000 614.200 305.600 ;
        RECT 618.800 302.200 619.600 306.800 ;
        RECT 622.400 306.200 623.000 307.600 ;
        RECT 625.200 306.800 626.000 308.400 ;
        RECT 622.000 305.600 623.000 306.200 ;
        RECT 626.800 306.200 627.600 309.700 ;
        RECT 632.000 308.400 632.600 311.800 ;
        RECT 636.400 310.400 637.000 311.800 ;
        RECT 641.200 311.200 642.000 319.800 ;
        RECT 638.000 310.800 642.000 311.200 ;
        RECT 637.800 310.600 642.000 310.800 ;
        RECT 633.200 308.800 634.000 310.400 ;
        RECT 636.400 309.600 637.200 310.400 ;
        RECT 637.800 310.000 638.600 310.600 ;
        RECT 630.000 307.600 632.600 308.400 ;
        RECT 634.800 308.200 635.600 308.400 ;
        RECT 634.000 307.600 635.600 308.200 ;
        RECT 630.200 306.200 630.800 307.600 ;
        RECT 634.000 307.200 634.800 307.600 ;
        RECT 631.800 306.200 635.400 306.600 ;
        RECT 636.400 306.200 637.000 309.600 ;
        RECT 637.800 307.000 638.400 310.000 ;
        RECT 639.200 308.400 640.000 309.200 ;
        RECT 639.400 307.600 640.400 308.400 ;
        RECT 637.800 306.400 640.200 307.000 ;
        RECT 626.800 305.600 628.600 306.200 ;
        RECT 622.000 302.200 622.800 305.600 ;
        RECT 627.800 302.200 628.600 305.600 ;
        RECT 630.000 302.200 630.800 306.200 ;
        RECT 631.600 306.000 635.600 306.200 ;
        RECT 631.600 302.200 632.400 306.000 ;
        RECT 634.800 302.200 635.600 306.000 ;
        RECT 636.400 302.200 637.200 306.200 ;
        RECT 639.600 304.200 640.200 306.400 ;
        RECT 641.200 304.800 642.000 306.400 ;
        RECT 639.600 302.200 640.400 304.200 ;
        RECT 642.800 302.200 643.600 319.800 ;
        RECT 649.800 312.800 650.600 319.800 ;
        RECT 654.000 315.000 654.800 319.000 ;
        RECT 649.000 312.200 650.600 312.800 ;
        RECT 646.000 310.300 646.800 310.400 ;
        RECT 647.600 310.300 648.400 311.200 ;
        RECT 646.000 309.700 648.400 310.300 ;
        RECT 646.000 309.600 646.800 309.700 ;
        RECT 647.600 309.600 648.400 309.700 ;
        RECT 649.000 308.400 649.600 312.200 ;
        RECT 654.200 311.600 654.800 315.000 ;
        RECT 658.200 312.400 659.000 319.800 ;
        RECT 659.600 313.600 660.400 314.400 ;
        RECT 659.800 312.400 660.400 313.600 ;
        RECT 662.800 313.600 663.600 314.400 ;
        RECT 662.800 312.400 663.400 313.600 ;
        RECT 664.200 312.400 665.000 319.800 ;
        RECT 658.200 311.800 659.200 312.400 ;
        RECT 659.800 311.800 661.200 312.400 ;
        RECT 651.000 311.000 654.800 311.600 ;
        RECT 651.000 309.000 651.600 311.000 ;
        RECT 647.600 307.600 649.600 308.400 ;
        RECT 650.200 308.200 651.600 309.000 ;
        RECT 652.400 308.800 653.200 310.400 ;
        RECT 654.000 308.800 654.800 310.400 ;
        RECT 657.200 308.800 658.000 310.400 ;
        RECT 658.600 310.300 659.200 311.800 ;
        RECT 660.400 311.600 661.200 311.800 ;
        RECT 662.000 311.800 663.400 312.400 ;
        RECT 664.000 311.800 665.000 312.400 ;
        RECT 662.000 311.600 662.800 311.800 ;
        RECT 662.100 310.300 662.700 311.600 ;
        RECT 664.000 310.400 664.600 311.800 ;
        RECT 668.400 311.400 669.200 319.800 ;
        RECT 672.800 316.400 673.600 319.800 ;
        RECT 671.600 315.800 673.600 316.400 ;
        RECT 677.200 315.800 678.000 319.800 ;
        RECT 681.400 315.800 682.600 319.800 ;
        RECT 671.600 315.000 672.400 315.800 ;
        RECT 677.200 315.200 677.800 315.800 ;
        RECT 675.000 314.600 678.600 315.200 ;
        RECT 681.200 315.000 682.000 315.800 ;
        RECT 675.000 314.400 675.800 314.600 ;
        RECT 677.800 314.400 678.600 314.600 ;
        RECT 671.600 313.000 672.400 313.200 ;
        RECT 676.200 313.000 677.000 313.200 ;
        RECT 671.600 312.400 677.000 313.000 ;
        RECT 677.600 313.000 679.800 313.600 ;
        RECT 677.600 311.800 678.200 313.000 ;
        RECT 679.000 312.800 679.800 313.000 ;
        RECT 681.400 313.200 682.800 314.000 ;
        RECT 681.400 312.200 682.000 313.200 ;
        RECT 673.400 311.400 678.200 311.800 ;
        RECT 668.400 311.200 678.200 311.400 ;
        RECT 679.600 311.600 682.000 312.200 ;
        RECT 668.400 311.000 674.200 311.200 ;
        RECT 668.400 310.800 674.000 311.000 ;
        RECT 658.600 309.700 662.700 310.300 ;
        RECT 658.600 308.400 659.200 309.700 ;
        RECT 663.600 309.600 664.600 310.400 ;
        RECT 664.000 308.400 664.600 309.600 ;
        RECT 665.200 308.800 666.000 310.400 ;
        RECT 674.800 310.200 675.600 310.400 ;
        RECT 670.600 309.600 675.600 310.200 ;
        RECT 670.600 309.400 671.400 309.600 ;
        RECT 673.200 309.400 674.000 309.600 ;
        RECT 672.200 308.400 673.000 308.600 ;
        RECT 679.600 308.400 680.200 311.600 ;
        RECT 686.000 311.200 686.800 319.800 ;
        RECT 682.600 310.600 686.800 311.200 ;
        RECT 682.600 310.400 683.400 310.600 ;
        RECT 684.200 309.800 685.000 310.000 ;
        RECT 681.200 309.200 685.000 309.800 ;
        RECT 681.200 309.000 682.000 309.200 ;
        RECT 649.000 307.000 649.600 307.600 ;
        RECT 650.600 307.800 651.600 308.200 ;
        RECT 655.600 308.200 656.400 308.400 ;
        RECT 650.600 307.200 654.800 307.800 ;
        RECT 655.600 307.600 657.200 308.200 ;
        RECT 658.600 307.600 661.200 308.400 ;
        RECT 662.000 307.600 664.600 308.400 ;
        RECT 666.800 308.200 667.600 308.400 ;
        RECT 666.000 307.600 667.600 308.200 ;
        RECT 669.200 307.800 680.200 308.400 ;
        RECT 669.200 307.600 670.800 307.800 ;
        RECT 656.400 307.200 657.200 307.600 ;
        RECT 649.000 306.600 649.800 307.000 ;
        RECT 649.000 306.400 650.600 306.600 ;
        RECT 644.400 304.800 645.200 306.400 ;
        RECT 649.000 306.000 651.600 306.400 ;
        RECT 649.800 305.600 651.600 306.000 ;
        RECT 649.800 303.000 650.600 305.600 ;
        RECT 654.200 305.000 654.800 307.200 ;
        RECT 655.800 306.200 659.400 306.600 ;
        RECT 660.400 306.200 661.000 307.600 ;
        RECT 662.200 306.200 662.800 307.600 ;
        RECT 666.000 307.200 666.800 307.600 ;
        RECT 663.800 306.200 667.400 306.600 ;
        RECT 654.000 303.000 654.800 305.000 ;
        RECT 655.600 306.000 659.600 306.200 ;
        RECT 655.600 302.200 656.400 306.000 ;
        RECT 658.800 302.200 659.600 306.000 ;
        RECT 660.400 302.200 661.200 306.200 ;
        RECT 662.000 302.200 662.800 306.200 ;
        RECT 663.600 306.000 667.600 306.200 ;
        RECT 663.600 302.200 664.400 306.000 ;
        RECT 666.800 302.200 667.600 306.000 ;
        RECT 668.400 302.200 669.200 307.000 ;
        RECT 673.400 305.600 674.000 307.800 ;
        RECT 676.400 307.600 677.200 307.800 ;
        RECT 679.000 307.600 679.800 307.800 ;
        RECT 686.000 307.200 686.800 310.600 ;
        RECT 683.000 306.600 686.800 307.200 ;
        RECT 683.000 306.400 683.800 306.600 ;
        RECT 671.600 304.200 672.400 305.000 ;
        RECT 673.200 304.800 674.000 305.600 ;
        RECT 675.000 305.400 675.800 305.600 ;
        RECT 675.000 304.800 677.800 305.400 ;
        RECT 677.200 304.200 677.800 304.800 ;
        RECT 681.200 304.200 682.000 305.000 ;
        RECT 671.600 303.600 673.600 304.200 ;
        RECT 672.800 302.200 673.600 303.600 ;
        RECT 677.200 302.200 678.000 304.200 ;
        RECT 681.200 303.600 682.600 304.200 ;
        RECT 681.400 302.200 682.600 303.600 ;
        RECT 686.000 302.200 686.800 306.600 ;
        RECT 2.800 294.300 3.600 299.800 ;
        RECT 4.400 296.000 5.200 299.800 ;
        RECT 7.600 296.000 8.400 299.800 ;
        RECT 4.400 295.800 8.400 296.000 ;
        RECT 9.200 295.800 10.000 299.800 ;
        RECT 10.800 295.800 11.600 299.800 ;
        RECT 12.400 296.000 13.200 299.800 ;
        RECT 15.600 296.000 16.400 299.800 ;
        RECT 12.400 295.800 16.400 296.000 ;
        RECT 17.800 296.400 18.600 299.800 ;
        RECT 17.800 295.800 19.600 296.400 ;
        RECT 22.000 295.800 22.800 299.800 ;
        RECT 23.600 296.000 24.400 299.800 ;
        RECT 26.800 296.000 27.600 299.800 ;
        RECT 23.600 295.800 27.600 296.000 ;
        RECT 28.400 296.000 29.200 299.800 ;
        RECT 31.600 296.000 32.400 299.800 ;
        RECT 28.400 295.800 32.400 296.000 ;
        RECT 33.200 295.800 34.000 299.800 ;
        RECT 34.800 295.800 35.600 299.800 ;
        RECT 36.400 296.000 37.200 299.800 ;
        RECT 39.600 296.000 40.400 299.800 ;
        RECT 36.400 295.800 40.400 296.000 ;
        RECT 4.600 295.400 8.200 295.800 ;
        RECT 5.200 294.400 6.000 294.800 ;
        RECT 9.200 294.400 9.800 295.800 ;
        RECT 11.000 294.400 11.600 295.800 ;
        RECT 12.600 295.400 16.200 295.800 ;
        RECT 14.800 294.400 15.600 294.800 ;
        RECT 4.400 294.300 6.000 294.400 ;
        RECT 2.800 293.800 6.000 294.300 ;
        RECT 2.800 293.700 5.200 293.800 ;
        RECT 2.800 282.200 3.600 293.700 ;
        RECT 4.400 293.600 5.200 293.700 ;
        RECT 7.400 293.600 10.000 294.400 ;
        RECT 10.800 293.600 13.400 294.400 ;
        RECT 14.800 293.800 16.400 294.400 ;
        RECT 15.600 293.600 16.400 293.800 ;
        RECT 6.000 291.600 6.800 293.200 ;
        RECT 7.400 290.200 8.000 293.600 ;
        RECT 12.800 292.300 13.400 293.600 ;
        RECT 9.300 291.700 13.400 292.300 ;
        RECT 9.300 290.400 9.900 291.700 ;
        RECT 9.200 290.200 10.000 290.400 ;
        RECT 7.000 289.600 8.000 290.200 ;
        RECT 8.600 289.600 10.000 290.200 ;
        RECT 10.800 290.200 11.600 290.400 ;
        RECT 12.800 290.200 13.400 291.700 ;
        RECT 14.000 291.600 14.800 293.200 ;
        RECT 10.800 289.600 12.200 290.200 ;
        RECT 12.800 289.600 13.800 290.200 ;
        RECT 7.000 284.400 7.800 289.600 ;
        RECT 8.600 288.400 9.200 289.600 ;
        RECT 8.400 287.600 9.200 288.400 ;
        RECT 11.600 288.400 12.200 289.600 ;
        RECT 11.600 287.600 12.400 288.400 ;
        RECT 6.000 283.600 7.800 284.400 ;
        RECT 7.000 282.200 7.800 283.600 ;
        RECT 13.000 282.200 13.800 289.600 ;
        RECT 17.200 287.600 18.000 290.400 ;
        RECT 18.800 290.300 19.600 295.800 ;
        RECT 20.400 293.600 21.200 295.200 ;
        RECT 22.200 294.400 22.800 295.800 ;
        RECT 23.800 295.400 27.400 295.800 ;
        RECT 28.600 295.400 32.200 295.800 ;
        RECT 26.000 294.400 26.800 294.800 ;
        RECT 29.200 294.400 30.000 294.800 ;
        RECT 33.200 294.400 33.800 295.800 ;
        RECT 35.000 294.400 35.600 295.800 ;
        RECT 36.600 295.400 40.200 295.800 ;
        RECT 38.800 294.400 39.600 294.800 ;
        RECT 22.000 293.600 24.600 294.400 ;
        RECT 26.000 293.800 27.600 294.400 ;
        RECT 26.800 293.600 27.600 293.800 ;
        RECT 28.400 293.800 30.000 294.400 ;
        RECT 28.400 293.600 29.200 293.800 ;
        RECT 31.400 293.600 34.000 294.400 ;
        RECT 34.800 293.600 37.400 294.400 ;
        RECT 38.800 294.300 40.400 294.400 ;
        RECT 41.200 294.300 42.000 299.800 ;
        RECT 42.800 295.600 43.600 297.200 ;
        RECT 47.000 296.400 47.800 299.800 ;
        RECT 46.000 295.800 47.800 296.400 ;
        RECT 49.200 295.800 50.000 299.800 ;
        RECT 50.800 296.000 51.600 299.800 ;
        RECT 54.000 296.000 54.800 299.800 ;
        RECT 50.800 295.800 54.800 296.000 ;
        RECT 55.600 295.800 56.400 299.800 ;
        RECT 57.200 296.000 58.000 299.800 ;
        RECT 60.400 296.000 61.200 299.800 ;
        RECT 57.200 295.800 61.200 296.000 ;
        RECT 38.800 293.800 42.000 294.300 ;
        RECT 39.600 293.700 42.000 293.800 ;
        RECT 39.600 293.600 40.400 293.700 ;
        RECT 22.000 290.300 22.800 290.400 ;
        RECT 18.800 290.200 22.800 290.300 ;
        RECT 24.000 290.200 24.600 293.600 ;
        RECT 25.200 292.300 26.000 293.200 ;
        RECT 26.800 292.300 27.600 292.400 ;
        RECT 25.200 291.700 27.600 292.300 ;
        RECT 25.200 291.600 26.000 291.700 ;
        RECT 26.800 291.600 27.600 291.700 ;
        RECT 30.000 291.600 30.800 293.200 ;
        RECT 31.400 292.300 32.000 293.600 ;
        RECT 31.400 291.700 35.500 292.300 ;
        RECT 31.400 290.200 32.000 291.700 ;
        RECT 34.900 290.400 35.500 291.700 ;
        RECT 33.200 290.200 34.000 290.400 ;
        RECT 18.800 289.700 23.400 290.200 ;
        RECT 18.800 282.200 19.600 289.700 ;
        RECT 22.000 289.600 23.400 289.700 ;
        RECT 24.000 289.600 25.000 290.200 ;
        RECT 22.800 288.400 23.400 289.600 ;
        RECT 22.800 287.600 23.600 288.400 ;
        RECT 24.200 282.200 25.000 289.600 ;
        RECT 31.000 289.600 32.000 290.200 ;
        RECT 32.600 289.600 34.000 290.200 ;
        RECT 34.800 290.200 35.600 290.400 ;
        RECT 36.800 290.200 37.400 293.600 ;
        RECT 38.000 291.600 38.800 293.200 ;
        RECT 34.800 289.600 36.200 290.200 ;
        RECT 36.800 289.600 37.800 290.200 ;
        RECT 31.000 282.200 31.800 289.600 ;
        RECT 32.600 288.400 33.200 289.600 ;
        RECT 32.400 287.600 33.200 288.400 ;
        RECT 35.600 288.400 36.200 289.600 ;
        RECT 35.600 287.600 36.400 288.400 ;
        RECT 37.000 284.400 37.800 289.600 ;
        RECT 37.000 283.600 38.800 284.400 ;
        RECT 37.000 282.200 37.800 283.600 ;
        RECT 41.200 282.200 42.000 293.700 ;
        RECT 44.400 293.600 45.200 295.200 ;
        RECT 46.000 292.300 46.800 295.800 ;
        RECT 49.400 294.400 50.000 295.800 ;
        RECT 51.000 295.400 54.600 295.800 ;
        RECT 53.200 294.400 54.000 294.800 ;
        RECT 55.800 294.400 56.400 295.800 ;
        RECT 57.400 295.400 61.000 295.800 ;
        RECT 59.600 294.400 60.400 294.800 ;
        RECT 49.200 293.600 51.800 294.400 ;
        RECT 53.200 293.800 54.800 294.400 ;
        RECT 54.000 293.600 54.800 293.800 ;
        RECT 55.600 293.600 58.200 294.400 ;
        RECT 59.600 293.800 61.200 294.400 ;
        RECT 60.400 293.600 61.200 293.800 ;
        RECT 62.000 293.800 62.800 299.800 ;
        RECT 68.400 296.600 69.200 299.800 ;
        RECT 70.000 297.000 70.800 299.800 ;
        RECT 71.600 297.000 72.400 299.800 ;
        RECT 73.200 297.000 74.000 299.800 ;
        RECT 76.400 297.000 77.200 299.800 ;
        RECT 79.600 297.000 80.400 299.800 ;
        RECT 81.200 297.000 82.000 299.800 ;
        RECT 82.800 297.000 83.600 299.800 ;
        RECT 84.400 297.000 85.200 299.800 ;
        RECT 66.600 295.800 69.200 296.600 ;
        RECT 86.000 296.600 86.800 299.800 ;
        RECT 72.600 295.800 77.200 296.400 ;
        RECT 66.600 295.200 67.400 295.800 ;
        RECT 64.400 294.400 67.400 295.200 ;
        RECT 46.000 291.700 49.900 292.300 ;
        RECT 46.000 282.200 46.800 291.700 ;
        RECT 49.300 290.400 49.900 291.700 ;
        RECT 47.600 288.800 48.400 290.400 ;
        RECT 49.200 290.200 50.000 290.400 ;
        RECT 51.200 290.200 51.800 293.600 ;
        RECT 52.400 291.600 53.200 293.200 ;
        RECT 55.600 290.200 56.400 290.400 ;
        RECT 57.600 290.200 58.200 293.600 ;
        RECT 58.800 292.300 59.600 293.200 ;
        RECT 62.000 293.000 70.800 293.800 ;
        RECT 72.600 293.400 73.400 295.800 ;
        RECT 76.400 295.600 77.200 295.800 ;
        RECT 78.000 295.600 79.600 296.400 ;
        RECT 82.600 295.600 83.600 296.400 ;
        RECT 86.000 295.800 88.400 296.600 ;
        RECT 74.800 293.600 75.600 295.200 ;
        RECT 76.400 294.800 77.200 295.000 ;
        RECT 76.400 294.200 80.800 294.800 ;
        RECT 80.000 294.000 80.800 294.200 ;
        RECT 60.400 292.300 61.200 292.400 ;
        RECT 58.800 291.700 61.200 292.300 ;
        RECT 58.800 291.600 59.600 291.700 ;
        RECT 60.400 291.600 61.200 291.700 ;
        RECT 49.200 289.600 50.600 290.200 ;
        RECT 51.200 289.600 52.200 290.200 ;
        RECT 55.600 289.600 57.000 290.200 ;
        RECT 57.600 289.600 58.600 290.200 ;
        RECT 50.000 288.400 50.600 289.600 ;
        RECT 50.000 287.600 50.800 288.400 ;
        RECT 51.400 282.200 52.200 289.600 ;
        RECT 56.400 288.400 57.000 289.600 ;
        RECT 56.400 287.600 57.200 288.400 ;
        RECT 57.800 282.200 58.600 289.600 ;
        RECT 62.000 287.400 62.800 293.000 ;
        RECT 71.400 292.600 73.400 293.400 ;
        RECT 77.200 292.600 80.400 293.400 ;
        RECT 82.800 292.800 83.600 295.600 ;
        RECT 87.600 295.200 88.400 295.800 ;
        RECT 87.600 294.600 89.400 295.200 ;
        RECT 88.600 293.400 89.400 294.600 ;
        RECT 92.400 294.600 93.200 299.800 ;
        RECT 94.000 296.000 94.800 299.800 ;
        RECT 97.800 296.400 98.600 299.800 ;
        RECT 94.000 295.200 95.000 296.000 ;
        RECT 97.800 295.800 99.600 296.400 ;
        RECT 102.000 295.800 102.800 299.800 ;
        RECT 103.600 296.000 104.400 299.800 ;
        RECT 106.800 296.000 107.600 299.800 ;
        RECT 103.600 295.800 107.600 296.000 ;
        RECT 109.000 298.400 109.800 299.800 ;
        RECT 109.000 297.600 110.800 298.400 ;
        RECT 109.000 296.400 109.800 297.600 ;
        RECT 109.000 295.800 110.800 296.400 ;
        RECT 92.400 294.000 93.600 294.600 ;
        RECT 88.600 292.600 92.400 293.400 ;
        RECT 63.400 292.000 64.200 292.200 ;
        RECT 68.400 292.000 69.200 292.400 ;
        RECT 86.000 292.000 86.800 292.600 ;
        RECT 93.000 292.000 93.600 294.000 ;
        RECT 63.400 291.400 86.800 292.000 ;
        RECT 92.800 291.400 93.600 292.000 ;
        RECT 92.800 289.600 93.400 291.400 ;
        RECT 94.200 290.800 95.000 295.200 ;
        RECT 95.600 294.300 96.400 294.400 ;
        RECT 98.800 294.300 99.600 295.800 ;
        RECT 95.600 293.700 99.600 294.300 ;
        RECT 95.600 293.600 96.400 293.700 ;
        RECT 71.600 289.400 72.400 289.600 ;
        RECT 67.000 289.000 72.400 289.400 ;
        RECT 66.200 288.800 72.400 289.000 ;
        RECT 73.400 289.000 82.000 289.600 ;
        RECT 63.600 288.000 65.200 288.800 ;
        RECT 66.200 288.200 67.600 288.800 ;
        RECT 73.400 288.200 74.000 289.000 ;
        RECT 81.200 288.800 82.000 289.000 ;
        RECT 84.400 289.000 93.400 289.600 ;
        RECT 84.400 288.800 85.200 289.000 ;
        RECT 64.600 287.600 65.200 288.000 ;
        RECT 68.200 287.600 74.000 288.200 ;
        RECT 74.600 287.600 77.200 288.400 ;
        RECT 62.000 286.800 64.000 287.400 ;
        RECT 64.600 286.800 68.800 287.600 ;
        RECT 63.400 286.200 64.000 286.800 ;
        RECT 63.400 285.600 64.400 286.200 ;
        RECT 63.600 282.200 64.400 285.600 ;
        RECT 66.800 282.200 67.600 286.800 ;
        RECT 70.000 282.200 70.800 285.000 ;
        RECT 71.600 282.200 72.400 285.000 ;
        RECT 73.200 282.200 74.000 287.000 ;
        RECT 76.400 282.200 77.200 287.000 ;
        RECT 79.600 282.200 80.400 288.400 ;
        RECT 87.600 287.600 90.200 288.400 ;
        RECT 82.800 286.800 87.000 287.600 ;
        RECT 81.200 282.200 82.000 285.000 ;
        RECT 82.800 282.200 83.600 285.000 ;
        RECT 84.400 282.200 85.200 285.000 ;
        RECT 87.600 282.200 88.400 287.600 ;
        RECT 92.800 287.400 93.400 289.000 ;
        RECT 90.800 286.800 93.400 287.400 ;
        RECT 94.000 290.000 95.000 290.800 ;
        RECT 90.800 282.200 91.600 286.800 ;
        RECT 94.000 282.200 94.800 290.000 ;
        RECT 97.200 288.800 98.000 290.400 ;
        RECT 98.800 282.200 99.600 293.700 ;
        RECT 100.400 294.300 101.200 295.200 ;
        RECT 102.200 294.400 102.800 295.800 ;
        RECT 103.800 295.400 107.400 295.800 ;
        RECT 106.000 294.400 106.800 294.800 ;
        RECT 102.000 294.300 104.600 294.400 ;
        RECT 100.400 293.700 104.600 294.300 ;
        RECT 106.000 293.800 107.600 294.400 ;
        RECT 100.400 293.600 101.200 293.700 ;
        RECT 102.000 293.600 104.600 293.700 ;
        RECT 106.800 293.600 107.600 293.800 ;
        RECT 100.400 290.300 101.200 290.400 ;
        RECT 102.000 290.300 102.800 290.400 ;
        RECT 100.400 290.200 102.800 290.300 ;
        RECT 104.000 290.200 104.600 293.600 ;
        RECT 105.200 291.600 106.000 293.200 ;
        RECT 100.400 289.700 103.400 290.200 ;
        RECT 100.400 289.600 101.200 289.700 ;
        RECT 102.000 289.600 103.400 289.700 ;
        RECT 104.000 289.600 105.000 290.200 ;
        RECT 102.800 288.400 103.400 289.600 ;
        RECT 102.800 287.600 103.600 288.400 ;
        RECT 104.200 282.200 105.000 289.600 ;
        RECT 108.400 288.800 109.200 290.400 ;
        RECT 110.000 282.200 110.800 295.800 ;
        RECT 111.600 293.600 112.400 295.200 ;
        RECT 118.000 293.800 118.800 299.800 ;
        RECT 124.400 296.600 125.200 299.800 ;
        RECT 126.000 297.000 126.800 299.800 ;
        RECT 127.600 297.000 128.400 299.800 ;
        RECT 129.200 297.000 130.000 299.800 ;
        RECT 132.400 297.000 133.200 299.800 ;
        RECT 135.600 297.000 136.400 299.800 ;
        RECT 137.200 297.000 138.000 299.800 ;
        RECT 138.800 297.000 139.600 299.800 ;
        RECT 140.400 297.000 141.200 299.800 ;
        RECT 122.600 295.800 125.200 296.600 ;
        RECT 142.000 296.600 142.800 299.800 ;
        RECT 128.600 295.800 133.200 296.400 ;
        RECT 122.600 295.200 123.400 295.800 ;
        RECT 120.400 294.400 123.400 295.200 ;
        RECT 118.000 293.000 126.800 293.800 ;
        RECT 128.600 293.400 129.400 295.800 ;
        RECT 132.400 295.600 133.200 295.800 ;
        RECT 134.000 295.600 135.600 296.400 ;
        RECT 138.600 295.600 139.600 296.400 ;
        RECT 142.000 295.800 144.400 296.600 ;
        RECT 130.800 293.600 131.600 295.200 ;
        RECT 132.400 294.800 133.200 295.000 ;
        RECT 132.400 294.200 136.800 294.800 ;
        RECT 136.000 294.000 136.800 294.200 ;
        RECT 118.000 287.400 118.800 293.000 ;
        RECT 127.400 292.600 129.400 293.400 ;
        RECT 133.200 292.600 136.400 293.400 ;
        RECT 138.800 292.800 139.600 295.600 ;
        RECT 143.600 295.200 144.400 295.800 ;
        RECT 143.600 294.600 145.400 295.200 ;
        RECT 144.600 293.400 145.400 294.600 ;
        RECT 148.400 294.600 149.200 299.800 ;
        RECT 150.000 296.000 150.800 299.800 ;
        RECT 153.800 296.400 154.600 299.800 ;
        RECT 150.000 295.200 151.000 296.000 ;
        RECT 153.800 295.800 155.600 296.400 ;
        RECT 158.000 295.800 158.800 299.800 ;
        RECT 159.600 296.000 160.400 299.800 ;
        RECT 162.800 296.000 163.600 299.800 ;
        RECT 159.600 295.800 163.600 296.000 ;
        RECT 148.400 294.000 149.600 294.600 ;
        RECT 144.600 292.600 148.400 293.400 ;
        RECT 119.400 292.000 120.200 292.200 ;
        RECT 124.400 292.000 125.200 292.400 ;
        RECT 142.000 292.000 142.800 292.600 ;
        RECT 149.000 292.000 149.600 294.000 ;
        RECT 119.400 291.400 142.800 292.000 ;
        RECT 148.800 291.400 149.600 292.000 ;
        RECT 148.800 289.600 149.400 291.400 ;
        RECT 150.200 290.800 151.000 295.200 ;
        RECT 153.200 294.300 154.000 294.400 ;
        RECT 154.800 294.300 155.600 295.800 ;
        RECT 153.200 293.700 155.600 294.300 ;
        RECT 153.200 293.600 154.000 293.700 ;
        RECT 127.600 289.400 128.400 289.600 ;
        RECT 123.000 289.000 128.400 289.400 ;
        RECT 122.200 288.800 128.400 289.000 ;
        RECT 129.400 289.000 138.000 289.600 ;
        RECT 119.600 288.000 121.200 288.800 ;
        RECT 122.200 288.200 123.600 288.800 ;
        RECT 129.400 288.200 130.000 289.000 ;
        RECT 137.200 288.800 138.000 289.000 ;
        RECT 140.400 289.000 149.400 289.600 ;
        RECT 140.400 288.800 141.200 289.000 ;
        RECT 120.600 287.600 121.200 288.000 ;
        RECT 124.200 287.600 130.000 288.200 ;
        RECT 130.600 287.600 133.200 288.400 ;
        RECT 118.000 286.800 120.000 287.400 ;
        RECT 120.600 286.800 124.800 287.600 ;
        RECT 119.400 286.200 120.000 286.800 ;
        RECT 119.400 285.600 120.400 286.200 ;
        RECT 119.600 282.200 120.400 285.600 ;
        RECT 122.800 282.200 123.600 286.800 ;
        RECT 126.000 282.200 126.800 285.000 ;
        RECT 127.600 282.200 128.400 285.000 ;
        RECT 129.200 282.200 130.000 287.000 ;
        RECT 132.400 282.200 133.200 287.000 ;
        RECT 135.600 282.200 136.400 288.400 ;
        RECT 143.600 287.600 146.200 288.400 ;
        RECT 138.800 286.800 143.000 287.600 ;
        RECT 137.200 282.200 138.000 285.000 ;
        RECT 138.800 282.200 139.600 285.000 ;
        RECT 140.400 282.200 141.200 285.000 ;
        RECT 143.600 282.200 144.400 287.600 ;
        RECT 148.800 287.400 149.400 289.000 ;
        RECT 146.800 286.800 149.400 287.400 ;
        RECT 150.000 290.000 151.000 290.800 ;
        RECT 146.800 282.200 147.600 286.800 ;
        RECT 150.000 282.200 150.800 290.000 ;
        RECT 153.200 288.800 154.000 290.400 ;
        RECT 154.800 282.200 155.600 293.700 ;
        RECT 156.400 294.300 157.200 295.200 ;
        RECT 158.200 294.400 158.800 295.800 ;
        RECT 159.800 295.400 163.400 295.800 ;
        RECT 162.000 294.400 162.800 294.800 ;
        RECT 158.000 294.300 160.600 294.400 ;
        RECT 156.400 293.700 160.600 294.300 ;
        RECT 162.000 293.800 163.600 294.400 ;
        RECT 156.400 293.600 157.200 293.700 ;
        RECT 158.000 293.600 160.600 293.700 ;
        RECT 162.800 293.600 163.600 293.800 ;
        RECT 164.400 293.800 165.200 299.800 ;
        RECT 170.800 296.600 171.600 299.800 ;
        RECT 172.400 297.000 173.200 299.800 ;
        RECT 174.000 297.000 174.800 299.800 ;
        RECT 175.600 297.000 176.400 299.800 ;
        RECT 178.800 297.000 179.600 299.800 ;
        RECT 182.000 297.000 182.800 299.800 ;
        RECT 183.600 297.000 184.400 299.800 ;
        RECT 185.200 297.000 186.000 299.800 ;
        RECT 186.800 297.000 187.600 299.800 ;
        RECT 169.000 295.800 171.600 296.600 ;
        RECT 188.400 296.600 189.200 299.800 ;
        RECT 175.000 295.800 179.600 296.400 ;
        RECT 169.000 295.200 169.800 295.800 ;
        RECT 166.800 294.400 169.800 295.200 ;
        RECT 158.000 290.200 158.800 290.400 ;
        RECT 160.000 290.200 160.600 293.600 ;
        RECT 161.200 291.600 162.000 293.200 ;
        RECT 164.400 293.000 173.200 293.800 ;
        RECT 175.000 293.400 175.800 295.800 ;
        RECT 178.800 295.600 179.600 295.800 ;
        RECT 180.400 295.600 182.000 296.400 ;
        RECT 185.000 295.600 186.000 296.400 ;
        RECT 188.400 295.800 190.800 296.600 ;
        RECT 177.200 293.600 178.000 295.200 ;
        RECT 178.800 294.800 179.600 295.000 ;
        RECT 178.800 294.200 183.200 294.800 ;
        RECT 182.400 294.000 183.200 294.200 ;
        RECT 158.000 289.600 159.400 290.200 ;
        RECT 160.000 289.600 161.000 290.200 ;
        RECT 158.800 288.400 159.400 289.600 ;
        RECT 156.400 288.300 157.200 288.400 ;
        RECT 158.800 288.300 159.600 288.400 ;
        RECT 156.400 287.700 159.600 288.300 ;
        RECT 156.400 287.600 157.200 287.700 ;
        RECT 158.800 287.600 159.600 287.700 ;
        RECT 160.200 282.200 161.000 289.600 ;
        RECT 164.400 287.400 165.200 293.000 ;
        RECT 173.800 292.600 175.800 293.400 ;
        RECT 179.600 292.600 182.800 293.400 ;
        RECT 185.200 292.800 186.000 295.600 ;
        RECT 190.000 295.200 190.800 295.800 ;
        RECT 190.000 294.600 191.800 295.200 ;
        RECT 191.000 293.400 191.800 294.600 ;
        RECT 194.800 294.600 195.600 299.800 ;
        RECT 196.400 296.000 197.200 299.800 ;
        RECT 199.600 296.000 200.400 299.800 ;
        RECT 202.800 296.000 203.600 299.800 ;
        RECT 196.400 295.200 197.400 296.000 ;
        RECT 199.600 295.800 203.600 296.000 ;
        RECT 204.400 295.800 205.200 299.800 ;
        RECT 199.800 295.400 203.400 295.800 ;
        RECT 194.800 294.000 196.000 294.600 ;
        RECT 191.000 292.600 194.800 293.400 ;
        RECT 165.800 292.000 166.600 292.200 ;
        RECT 170.800 292.000 171.600 292.400 ;
        RECT 188.400 292.000 189.200 292.600 ;
        RECT 195.400 292.000 196.000 294.000 ;
        RECT 165.800 291.400 189.200 292.000 ;
        RECT 195.200 291.400 196.000 292.000 ;
        RECT 195.200 289.600 195.800 291.400 ;
        RECT 196.600 290.800 197.400 295.200 ;
        RECT 200.400 294.400 201.200 294.800 ;
        RECT 204.400 294.400 205.000 295.800 ;
        RECT 199.600 293.800 201.200 294.400 ;
        RECT 199.600 293.600 200.400 293.800 ;
        RECT 202.600 293.600 205.200 294.400 ;
        RECT 206.000 293.800 206.800 299.800 ;
        RECT 212.400 296.600 213.200 299.800 ;
        RECT 214.000 297.000 214.800 299.800 ;
        RECT 215.600 297.000 216.400 299.800 ;
        RECT 217.200 297.000 218.000 299.800 ;
        RECT 220.400 297.000 221.200 299.800 ;
        RECT 223.600 297.000 224.400 299.800 ;
        RECT 225.200 297.000 226.000 299.800 ;
        RECT 226.800 297.000 227.600 299.800 ;
        RECT 228.400 297.000 229.200 299.800 ;
        RECT 210.600 295.800 213.200 296.600 ;
        RECT 230.000 296.600 230.800 299.800 ;
        RECT 216.600 295.800 221.200 296.400 ;
        RECT 210.600 295.200 211.400 295.800 ;
        RECT 208.400 294.400 211.400 295.200 ;
        RECT 201.200 291.600 202.000 293.200 ;
        RECT 174.000 289.400 174.800 289.600 ;
        RECT 169.400 289.000 174.800 289.400 ;
        RECT 168.600 288.800 174.800 289.000 ;
        RECT 175.800 289.000 184.400 289.600 ;
        RECT 166.000 288.000 167.600 288.800 ;
        RECT 168.600 288.200 170.000 288.800 ;
        RECT 175.800 288.200 176.400 289.000 ;
        RECT 183.600 288.800 184.400 289.000 ;
        RECT 186.800 289.000 195.800 289.600 ;
        RECT 186.800 288.800 187.600 289.000 ;
        RECT 167.000 287.600 167.600 288.000 ;
        RECT 170.600 287.600 176.400 288.200 ;
        RECT 177.000 287.600 179.600 288.400 ;
        RECT 164.400 286.800 166.400 287.400 ;
        RECT 167.000 286.800 171.200 287.600 ;
        RECT 165.800 286.200 166.400 286.800 ;
        RECT 165.800 285.600 166.800 286.200 ;
        RECT 166.000 282.200 166.800 285.600 ;
        RECT 169.200 282.200 170.000 286.800 ;
        RECT 172.400 282.200 173.200 285.000 ;
        RECT 174.000 282.200 174.800 285.000 ;
        RECT 175.600 282.200 176.400 287.000 ;
        RECT 178.800 282.200 179.600 287.000 ;
        RECT 182.000 282.200 182.800 288.400 ;
        RECT 190.000 287.600 192.600 288.400 ;
        RECT 185.200 286.800 189.400 287.600 ;
        RECT 183.600 282.200 184.400 285.000 ;
        RECT 185.200 282.200 186.000 285.000 ;
        RECT 186.800 282.200 187.600 285.000 ;
        RECT 190.000 282.200 190.800 287.600 ;
        RECT 195.200 287.400 195.800 289.000 ;
        RECT 193.200 286.800 195.800 287.400 ;
        RECT 196.400 290.000 197.400 290.800 ;
        RECT 202.600 290.200 203.200 293.600 ;
        RECT 206.000 293.000 214.800 293.800 ;
        RECT 216.600 293.400 217.400 295.800 ;
        RECT 220.400 295.600 221.200 295.800 ;
        RECT 222.000 295.600 223.600 296.400 ;
        RECT 226.600 295.600 227.600 296.400 ;
        RECT 230.000 295.800 232.400 296.600 ;
        RECT 218.800 293.600 219.600 295.200 ;
        RECT 220.400 294.800 221.200 295.000 ;
        RECT 220.400 294.200 224.800 294.800 ;
        RECT 224.000 294.000 224.800 294.200 ;
        RECT 204.400 290.200 205.200 290.400 ;
        RECT 193.200 282.200 194.000 286.800 ;
        RECT 196.400 282.200 197.200 290.000 ;
        RECT 202.200 289.600 203.200 290.200 ;
        RECT 203.800 289.600 205.200 290.200 ;
        RECT 202.200 282.200 203.000 289.600 ;
        RECT 203.800 288.400 204.400 289.600 ;
        RECT 203.600 287.600 204.400 288.400 ;
        RECT 206.000 287.400 206.800 293.000 ;
        RECT 215.400 292.600 217.400 293.400 ;
        RECT 221.200 292.600 224.400 293.400 ;
        RECT 226.800 292.800 227.600 295.600 ;
        RECT 231.600 295.200 232.400 295.800 ;
        RECT 231.600 294.600 233.400 295.200 ;
        RECT 232.600 293.400 233.400 294.600 ;
        RECT 236.400 294.600 237.200 299.800 ;
        RECT 238.000 296.000 238.800 299.800 ;
        RECT 238.000 295.200 239.000 296.000 ;
        RECT 236.400 294.000 237.600 294.600 ;
        RECT 232.600 292.600 236.400 293.400 ;
        RECT 207.400 292.000 208.200 292.200 ;
        RECT 212.400 292.000 213.200 292.400 ;
        RECT 218.800 292.000 219.600 292.400 ;
        RECT 230.000 292.000 230.800 292.600 ;
        RECT 237.000 292.000 237.600 294.000 ;
        RECT 207.400 291.400 230.800 292.000 ;
        RECT 236.800 291.400 237.600 292.000 ;
        RECT 238.200 294.300 239.000 295.200 ;
        RECT 241.200 294.300 242.000 295.200 ;
        RECT 238.200 293.700 242.000 294.300 ;
        RECT 236.800 289.600 237.400 291.400 ;
        RECT 238.200 290.800 239.000 293.700 ;
        RECT 241.200 293.600 242.000 293.700 ;
        RECT 215.600 289.400 216.400 289.600 ;
        RECT 211.000 289.000 216.400 289.400 ;
        RECT 210.200 288.800 216.400 289.000 ;
        RECT 217.400 289.000 226.000 289.600 ;
        RECT 207.600 288.000 209.200 288.800 ;
        RECT 210.200 288.200 211.600 288.800 ;
        RECT 217.400 288.200 218.000 289.000 ;
        RECT 225.200 288.800 226.000 289.000 ;
        RECT 228.400 289.000 237.400 289.600 ;
        RECT 228.400 288.800 229.200 289.000 ;
        RECT 208.600 287.600 209.200 288.000 ;
        RECT 212.200 287.600 218.000 288.200 ;
        RECT 218.600 287.600 221.200 288.400 ;
        RECT 206.000 286.800 208.000 287.400 ;
        RECT 208.600 286.800 212.800 287.600 ;
        RECT 207.400 286.200 208.000 286.800 ;
        RECT 207.400 285.600 208.400 286.200 ;
        RECT 207.600 282.200 208.400 285.600 ;
        RECT 210.800 282.200 211.600 286.800 ;
        RECT 214.000 282.200 214.800 285.000 ;
        RECT 215.600 282.200 216.400 285.000 ;
        RECT 217.200 282.200 218.000 287.000 ;
        RECT 220.400 282.200 221.200 287.000 ;
        RECT 223.600 282.200 224.400 288.400 ;
        RECT 231.600 287.600 234.200 288.400 ;
        RECT 226.800 286.800 231.000 287.600 ;
        RECT 225.200 282.200 226.000 285.000 ;
        RECT 226.800 282.200 227.600 285.000 ;
        RECT 228.400 282.200 229.200 285.000 ;
        RECT 231.600 282.200 232.400 287.600 ;
        RECT 236.800 287.400 237.400 289.000 ;
        RECT 234.800 286.800 237.400 287.400 ;
        RECT 238.000 290.000 239.000 290.800 ;
        RECT 234.800 282.200 235.600 286.800 ;
        RECT 238.000 282.200 238.800 290.000 ;
        RECT 242.800 282.200 243.600 299.800 ;
        RECT 247.000 296.400 247.800 299.800 ;
        RECT 251.800 296.400 252.600 299.800 ;
        RECT 246.000 295.800 247.800 296.400 ;
        RECT 250.800 295.800 252.600 296.400 ;
        RECT 244.400 293.600 245.200 295.200 ;
        RECT 246.000 294.300 246.800 295.800 ;
        RECT 249.200 294.300 250.000 295.200 ;
        RECT 246.000 293.700 250.000 294.300 ;
        RECT 246.000 282.200 246.800 293.700 ;
        RECT 249.200 293.600 250.000 293.700 ;
        RECT 247.600 288.800 248.400 290.400 ;
        RECT 250.800 282.200 251.600 295.800 ;
        RECT 258.800 293.800 259.600 299.800 ;
        RECT 265.200 296.600 266.000 299.800 ;
        RECT 266.800 297.000 267.600 299.800 ;
        RECT 268.400 297.000 269.200 299.800 ;
        RECT 270.000 297.000 270.800 299.800 ;
        RECT 273.200 297.000 274.000 299.800 ;
        RECT 276.400 297.000 277.200 299.800 ;
        RECT 278.000 297.000 278.800 299.800 ;
        RECT 279.600 297.000 280.400 299.800 ;
        RECT 281.200 297.000 282.000 299.800 ;
        RECT 263.400 295.800 266.000 296.600 ;
        RECT 282.800 296.600 283.600 299.800 ;
        RECT 269.400 295.800 274.000 296.400 ;
        RECT 263.400 295.200 264.200 295.800 ;
        RECT 261.200 294.400 264.200 295.200 ;
        RECT 258.800 293.000 267.600 293.800 ;
        RECT 269.400 293.400 270.200 295.800 ;
        RECT 273.200 295.600 274.000 295.800 ;
        RECT 274.800 295.600 276.400 296.400 ;
        RECT 279.400 295.600 280.400 296.400 ;
        RECT 282.800 295.800 285.200 296.600 ;
        RECT 271.600 293.600 272.400 295.200 ;
        RECT 273.200 294.800 274.000 295.000 ;
        RECT 273.200 294.200 277.600 294.800 ;
        RECT 276.800 294.000 277.600 294.200 ;
        RECT 252.400 288.800 253.200 290.400 ;
        RECT 258.800 287.400 259.600 293.000 ;
        RECT 268.200 292.600 270.200 293.400 ;
        RECT 274.000 292.600 277.200 293.400 ;
        RECT 279.600 292.800 280.400 295.600 ;
        RECT 284.400 295.200 285.200 295.800 ;
        RECT 284.400 294.600 286.200 295.200 ;
        RECT 285.400 293.400 286.200 294.600 ;
        RECT 289.200 294.600 290.000 299.800 ;
        RECT 290.800 296.000 291.600 299.800 ;
        RECT 290.800 295.200 291.800 296.000 ;
        RECT 289.200 294.000 290.400 294.600 ;
        RECT 285.400 292.600 289.200 293.400 ;
        RECT 260.200 292.000 261.000 292.200 ;
        RECT 265.200 292.000 266.000 292.400 ;
        RECT 282.800 292.000 283.600 292.600 ;
        RECT 289.800 292.000 290.400 294.000 ;
        RECT 260.200 291.400 283.600 292.000 ;
        RECT 289.600 291.400 290.400 292.000 ;
        RECT 289.600 289.600 290.200 291.400 ;
        RECT 291.000 290.800 291.800 295.200 ;
        RECT 297.600 294.200 298.400 299.800 ;
        RECT 300.400 295.200 301.200 299.800 ;
        RECT 300.400 294.600 302.600 295.200 ;
        RECT 297.600 293.800 299.400 294.200 ;
        RECT 297.800 293.600 299.400 293.800 ;
        RECT 295.600 291.600 297.200 292.400 ;
        RECT 268.400 289.400 269.200 289.600 ;
        RECT 263.800 289.000 269.200 289.400 ;
        RECT 263.000 288.800 269.200 289.000 ;
        RECT 270.200 289.000 278.800 289.600 ;
        RECT 260.400 288.000 262.000 288.800 ;
        RECT 263.000 288.200 264.400 288.800 ;
        RECT 270.200 288.200 270.800 289.000 ;
        RECT 278.000 288.800 278.800 289.000 ;
        RECT 281.200 289.000 290.200 289.600 ;
        RECT 281.200 288.800 282.000 289.000 ;
        RECT 261.400 287.600 262.000 288.000 ;
        RECT 265.000 287.600 270.800 288.200 ;
        RECT 271.400 287.600 274.000 288.400 ;
        RECT 258.800 286.800 260.800 287.400 ;
        RECT 261.400 286.800 265.600 287.600 ;
        RECT 260.200 286.200 260.800 286.800 ;
        RECT 260.200 285.600 261.200 286.200 ;
        RECT 260.400 282.200 261.200 285.600 ;
        RECT 263.600 282.200 264.400 286.800 ;
        RECT 266.800 282.200 267.600 285.000 ;
        RECT 268.400 282.200 269.200 285.000 ;
        RECT 270.000 282.200 270.800 287.000 ;
        RECT 273.200 282.200 274.000 287.000 ;
        RECT 276.400 282.200 277.200 288.400 ;
        RECT 284.400 287.600 287.000 288.400 ;
        RECT 279.600 286.800 283.800 287.600 ;
        RECT 278.000 282.200 278.800 285.000 ;
        RECT 279.600 282.200 280.400 285.000 ;
        RECT 281.200 282.200 282.000 285.000 ;
        RECT 284.400 282.200 285.200 287.600 ;
        RECT 289.600 287.400 290.200 289.000 ;
        RECT 287.600 286.800 290.200 287.400 ;
        RECT 290.800 290.000 291.800 290.800 ;
        RECT 298.800 290.400 299.400 293.600 ;
        RECT 300.400 291.600 301.200 293.200 ;
        RECT 302.000 291.600 302.600 294.600 ;
        RECT 303.600 292.400 304.400 299.800 ;
        RECT 306.400 294.200 307.200 299.800 ;
        RECT 312.800 294.200 313.600 299.800 ;
        RECT 319.200 294.200 320.000 299.800 ;
        RECT 325.000 296.400 325.800 299.800 ;
        RECT 330.400 298.400 331.200 299.800 ;
        RECT 330.400 297.600 331.600 298.400 ;
        RECT 325.000 295.800 326.800 296.400 ;
        RECT 302.000 290.800 303.200 291.600 ;
        RECT 287.600 282.200 288.400 286.800 ;
        RECT 290.800 282.200 291.600 290.000 ;
        RECT 298.800 289.600 299.600 290.400 ;
        RECT 302.000 290.200 302.600 290.800 ;
        RECT 303.800 290.200 304.400 292.400 ;
        RECT 305.400 293.800 307.200 294.200 ;
        RECT 311.800 293.800 313.600 294.200 ;
        RECT 318.200 293.800 320.000 294.200 ;
        RECT 305.400 293.600 307.000 293.800 ;
        RECT 311.800 293.600 313.400 293.800 ;
        RECT 318.200 293.600 319.800 293.800 ;
        RECT 305.400 290.400 306.000 293.600 ;
        RECT 307.600 291.600 309.200 292.400 ;
        RECT 311.800 290.400 312.400 293.600 ;
        RECT 314.000 291.600 315.600 292.400 ;
        RECT 318.200 290.400 318.800 293.600 ;
        RECT 320.400 291.600 322.000 292.400 ;
        RECT 300.400 289.600 302.600 290.200 ;
        RECT 297.200 287.600 298.000 289.200 ;
        RECT 298.800 287.000 299.400 289.600 ;
        RECT 295.800 286.400 299.400 287.000 ;
        RECT 295.800 286.200 296.400 286.400 ;
        RECT 295.600 282.200 296.400 286.200 ;
        RECT 298.800 286.200 299.400 286.400 ;
        RECT 298.800 282.200 299.600 286.200 ;
        RECT 300.400 282.200 301.200 289.600 ;
        RECT 303.600 282.200 304.400 290.200 ;
        RECT 305.200 289.600 306.000 290.400 ;
        RECT 311.600 289.600 312.400 290.400 ;
        RECT 318.000 289.600 318.800 290.400 ;
        RECT 322.800 289.600 323.600 291.200 ;
        RECT 305.400 287.000 306.000 289.600 ;
        RECT 306.800 287.600 307.600 289.200 ;
        RECT 311.800 287.000 312.400 289.600 ;
        RECT 313.200 287.600 314.000 289.200 ;
        RECT 318.200 287.000 318.800 289.600 ;
        RECT 319.600 288.300 320.400 289.200 ;
        RECT 324.400 288.800 325.200 290.400 ;
        RECT 322.800 288.300 323.600 288.400 ;
        RECT 319.600 287.700 323.600 288.300 ;
        RECT 319.600 287.600 320.400 287.700 ;
        RECT 322.800 287.600 323.600 287.700 ;
        RECT 305.400 286.400 309.000 287.000 ;
        RECT 305.400 286.200 306.000 286.400 ;
        RECT 305.200 282.200 306.000 286.200 ;
        RECT 308.400 286.200 309.000 286.400 ;
        RECT 311.800 286.400 315.400 287.000 ;
        RECT 311.800 286.200 312.400 286.400 ;
        RECT 308.400 282.200 309.200 286.200 ;
        RECT 311.600 282.200 312.400 286.200 ;
        RECT 314.800 286.200 315.400 286.400 ;
        RECT 318.200 286.400 321.800 287.000 ;
        RECT 318.200 286.200 318.800 286.400 ;
        RECT 314.800 282.200 315.600 286.200 ;
        RECT 318.000 282.200 318.800 286.200 ;
        RECT 321.200 282.200 322.000 286.400 ;
        RECT 326.000 282.200 326.800 295.800 ;
        RECT 327.600 293.600 328.400 295.200 ;
        RECT 330.400 294.200 331.200 297.600 ;
        RECT 329.400 293.800 331.200 294.200 ;
        RECT 339.200 294.200 340.000 299.800 ;
        RECT 343.200 294.200 344.000 299.800 ;
        RECT 339.200 293.800 341.000 294.200 ;
        RECT 329.400 293.600 331.000 293.800 ;
        RECT 339.400 293.600 341.000 293.800 ;
        RECT 329.400 290.400 330.000 293.600 ;
        RECT 329.200 289.600 330.000 290.400 ;
        RECT 334.000 290.300 334.800 291.200 ;
        RECT 335.600 290.300 336.400 291.200 ;
        RECT 340.400 290.400 341.000 293.600 ;
        RECT 342.200 293.800 344.000 294.200 ;
        RECT 352.000 294.200 352.800 299.800 ;
        RECT 358.600 296.400 359.400 299.000 ;
        RECT 362.800 297.000 363.600 299.000 ;
        RECT 358.600 296.000 360.400 296.400 ;
        RECT 357.800 295.600 360.400 296.000 ;
        RECT 357.800 295.400 359.400 295.600 ;
        RECT 357.800 295.000 358.600 295.400 ;
        RECT 357.800 294.400 358.400 295.000 ;
        RECT 363.000 294.800 363.600 297.000 ;
        RECT 352.000 293.800 353.800 294.200 ;
        RECT 342.200 293.600 343.800 293.800 ;
        RECT 352.200 293.600 353.800 293.800 ;
        RECT 356.400 293.600 358.400 294.400 ;
        RECT 359.400 294.200 363.600 294.800 ;
        RECT 359.400 293.800 360.400 294.200 ;
        RECT 342.200 290.400 342.800 293.600 ;
        RECT 344.400 291.600 346.000 292.400 ;
        RECT 337.200 290.300 338.000 290.400 ;
        RECT 334.000 289.700 338.000 290.300 ;
        RECT 334.000 289.600 334.800 289.700 ;
        RECT 335.600 289.600 336.400 289.700 ;
        RECT 337.200 289.600 338.000 289.700 ;
        RECT 340.400 289.600 341.200 290.400 ;
        RECT 342.000 289.600 342.800 290.400 ;
        RECT 346.800 290.300 347.600 291.200 ;
        RECT 348.400 290.300 349.200 291.200 ;
        RECT 346.800 289.700 349.200 290.300 ;
        RECT 346.800 289.600 347.600 289.700 ;
        RECT 348.400 289.600 349.200 289.700 ;
        RECT 353.200 290.400 353.800 293.600 ;
        RECT 356.400 290.800 357.200 292.400 ;
        RECT 353.200 289.600 354.000 290.400 ;
        RECT 357.800 289.800 358.400 293.600 ;
        RECT 359.000 293.000 360.400 293.800 ;
        RECT 359.800 291.000 360.400 293.000 ;
        RECT 361.200 291.600 362.000 293.200 ;
        RECT 362.800 291.600 363.600 293.200 ;
        RECT 359.800 290.400 363.600 291.000 ;
        RECT 329.400 287.000 330.000 289.600 ;
        RECT 330.800 288.300 331.600 289.200 ;
        RECT 332.400 288.300 333.200 288.400 ;
        RECT 330.800 287.700 333.200 288.300 ;
        RECT 330.800 287.600 331.600 287.700 ;
        RECT 332.400 287.600 333.200 287.700 ;
        RECT 338.800 287.600 339.600 289.200 ;
        RECT 340.400 287.000 341.000 289.600 ;
        RECT 329.400 286.400 333.000 287.000 ;
        RECT 329.400 286.200 330.000 286.400 ;
        RECT 329.200 282.200 330.000 286.200 ;
        RECT 332.400 286.200 333.000 286.400 ;
        RECT 337.400 286.400 341.000 287.000 ;
        RECT 337.400 286.200 338.000 286.400 ;
        RECT 332.400 282.200 333.200 286.200 ;
        RECT 337.200 282.200 338.000 286.200 ;
        RECT 340.400 286.200 341.000 286.400 ;
        RECT 342.200 287.000 342.800 289.600 ;
        RECT 343.600 287.600 344.400 289.200 ;
        RECT 348.400 288.300 349.200 288.400 ;
        RECT 345.300 287.700 349.200 288.300 ;
        RECT 345.300 287.000 345.900 287.700 ;
        RECT 348.400 287.600 349.200 287.700 ;
        RECT 351.600 287.600 352.400 289.200 ;
        RECT 353.200 287.000 353.800 289.600 ;
        RECT 357.800 289.200 359.400 289.800 ;
        RECT 342.200 286.400 345.900 287.000 ;
        RECT 342.200 286.200 342.800 286.400 ;
        RECT 340.400 282.200 341.200 286.200 ;
        RECT 342.000 282.200 342.800 286.200 ;
        RECT 345.200 286.200 345.900 286.400 ;
        RECT 350.200 286.400 353.800 287.000 ;
        RECT 350.200 286.200 350.800 286.400 ;
        RECT 345.200 282.200 346.000 286.200 ;
        RECT 350.000 282.200 350.800 286.200 ;
        RECT 353.200 286.200 353.800 286.400 ;
        RECT 353.200 282.200 354.000 286.200 ;
        RECT 358.600 282.200 359.400 289.200 ;
        RECT 363.000 287.000 363.600 290.400 ;
        RECT 362.800 283.000 363.600 287.000 ;
        RECT 364.400 282.200 365.200 299.800 ;
        RECT 366.000 296.300 366.800 297.200 ;
        RECT 369.200 296.300 370.000 299.800 ;
        RECT 366.000 295.700 370.000 296.300 ;
        RECT 366.000 295.600 366.800 295.700 ;
        RECT 369.000 295.200 370.000 295.700 ;
        RECT 369.000 290.800 369.800 295.200 ;
        RECT 370.800 294.600 371.600 299.800 ;
        RECT 377.200 296.600 378.000 299.800 ;
        RECT 378.800 297.000 379.600 299.800 ;
        RECT 380.400 297.000 381.200 299.800 ;
        RECT 382.000 297.000 382.800 299.800 ;
        RECT 383.600 297.000 384.400 299.800 ;
        RECT 386.800 297.000 387.600 299.800 ;
        RECT 390.000 297.000 390.800 299.800 ;
        RECT 391.600 297.000 392.400 299.800 ;
        RECT 393.200 297.000 394.000 299.800 ;
        RECT 375.600 295.800 378.000 296.600 ;
        RECT 394.800 296.600 395.600 299.800 ;
        RECT 375.600 295.200 376.400 295.800 ;
        RECT 370.400 294.000 371.600 294.600 ;
        RECT 374.600 294.600 376.400 295.200 ;
        RECT 380.400 295.600 381.400 296.400 ;
        RECT 384.400 295.600 386.000 296.400 ;
        RECT 386.800 295.800 391.400 296.400 ;
        RECT 394.800 295.800 397.400 296.600 ;
        RECT 386.800 295.600 387.600 295.800 ;
        RECT 370.400 292.000 371.000 294.000 ;
        RECT 374.600 293.400 375.400 294.600 ;
        RECT 371.600 292.600 375.400 293.400 ;
        RECT 380.400 292.800 381.200 295.600 ;
        RECT 386.800 294.800 387.600 295.000 ;
        RECT 383.200 294.200 387.600 294.800 ;
        RECT 383.200 294.000 384.000 294.200 ;
        RECT 388.400 293.600 389.200 295.200 ;
        RECT 390.600 293.400 391.400 295.800 ;
        RECT 396.600 295.200 397.400 295.800 ;
        RECT 396.600 294.400 399.600 295.200 ;
        RECT 401.200 293.800 402.000 299.800 ;
        RECT 402.800 297.000 403.600 299.000 ;
        RECT 407.000 298.400 407.800 299.000 ;
        RECT 407.000 297.600 408.400 298.400 ;
        RECT 402.800 294.800 403.400 297.000 ;
        RECT 407.000 296.000 407.800 297.600 ;
        RECT 407.000 295.400 408.600 296.000 ;
        RECT 407.800 295.000 408.600 295.400 ;
        RECT 402.800 294.200 407.000 294.800 ;
        RECT 383.600 292.600 386.800 293.400 ;
        RECT 390.600 292.600 392.600 293.400 ;
        RECT 393.200 293.000 402.000 293.800 ;
        RECT 406.000 293.800 407.000 294.200 ;
        RECT 408.000 294.400 408.600 295.000 ;
        RECT 377.200 292.000 378.000 292.600 ;
        RECT 394.800 292.000 395.600 292.400 ;
        RECT 399.800 292.000 400.600 292.200 ;
        RECT 370.400 291.400 371.200 292.000 ;
        RECT 377.200 291.400 400.600 292.000 ;
        RECT 369.000 290.000 370.000 290.800 ;
        RECT 369.200 282.200 370.000 290.000 ;
        RECT 370.600 289.600 371.200 291.400 ;
        RECT 370.600 289.000 379.600 289.600 ;
        RECT 370.600 287.400 371.200 289.000 ;
        RECT 378.800 288.800 379.600 289.000 ;
        RECT 382.000 289.000 390.600 289.600 ;
        RECT 382.000 288.800 382.800 289.000 ;
        RECT 373.800 287.600 376.400 288.400 ;
        RECT 370.600 286.800 373.200 287.400 ;
        RECT 372.400 282.200 373.200 286.800 ;
        RECT 375.600 282.200 376.400 287.600 ;
        RECT 377.000 286.800 381.200 287.600 ;
        RECT 378.800 282.200 379.600 285.000 ;
        RECT 380.400 282.200 381.200 285.000 ;
        RECT 382.000 282.200 382.800 285.000 ;
        RECT 383.600 282.200 384.400 288.400 ;
        RECT 386.800 287.600 389.400 288.400 ;
        RECT 390.000 288.200 390.600 289.000 ;
        RECT 391.600 289.400 392.400 289.600 ;
        RECT 391.600 289.000 397.000 289.400 ;
        RECT 391.600 288.800 397.800 289.000 ;
        RECT 396.400 288.200 397.800 288.800 ;
        RECT 390.000 287.600 395.800 288.200 ;
        RECT 398.800 288.000 400.400 288.800 ;
        RECT 398.800 287.600 399.400 288.000 ;
        RECT 386.800 282.200 387.600 287.000 ;
        RECT 390.000 282.200 390.800 287.000 ;
        RECT 395.200 286.800 399.400 287.600 ;
        RECT 401.200 287.400 402.000 293.000 ;
        RECT 402.800 291.600 403.600 293.200 ;
        RECT 404.400 291.600 405.200 293.200 ;
        RECT 406.000 293.000 407.400 293.800 ;
        RECT 408.000 293.600 410.000 294.400 ;
        RECT 406.000 291.000 406.600 293.000 ;
        RECT 400.000 286.800 402.000 287.400 ;
        RECT 402.800 290.400 406.600 291.000 ;
        RECT 402.800 287.000 403.400 290.400 ;
        RECT 408.000 289.800 408.600 293.600 ;
        RECT 409.200 292.300 410.000 292.400 ;
        RECT 412.400 292.300 413.200 299.800 ;
        RECT 414.000 295.600 414.800 297.200 ;
        RECT 409.200 291.700 413.200 292.300 ;
        RECT 409.200 290.800 410.000 291.700 ;
        RECT 407.000 289.200 408.600 289.800 ;
        RECT 391.600 282.200 392.400 285.000 ;
        RECT 393.200 282.200 394.000 285.000 ;
        RECT 396.400 282.200 397.200 286.800 ;
        RECT 400.000 286.200 400.600 286.800 ;
        RECT 399.600 285.600 400.600 286.200 ;
        RECT 399.600 282.200 400.400 285.600 ;
        RECT 402.800 283.000 403.600 287.000 ;
        RECT 407.000 282.200 407.800 289.200 ;
        RECT 412.400 282.200 413.200 291.700 ;
        RECT 420.400 293.800 421.200 299.800 ;
        RECT 426.800 296.600 427.600 299.800 ;
        RECT 428.400 297.000 429.200 299.800 ;
        RECT 430.000 297.000 430.800 299.800 ;
        RECT 431.600 297.000 432.400 299.800 ;
        RECT 434.800 297.000 435.600 299.800 ;
        RECT 438.000 297.000 438.800 299.800 ;
        RECT 439.600 297.000 440.400 299.800 ;
        RECT 441.200 297.000 442.000 299.800 ;
        RECT 442.800 297.000 443.600 299.800 ;
        RECT 425.000 295.800 427.600 296.600 ;
        RECT 444.400 296.600 445.200 299.800 ;
        RECT 431.000 295.800 435.600 296.400 ;
        RECT 425.000 295.200 425.800 295.800 ;
        RECT 422.800 294.400 425.800 295.200 ;
        RECT 420.400 293.000 429.200 293.800 ;
        RECT 431.000 293.400 431.800 295.800 ;
        RECT 434.800 295.600 435.600 295.800 ;
        RECT 436.400 295.600 438.000 296.400 ;
        RECT 441.000 295.600 442.000 296.400 ;
        RECT 444.400 295.800 446.800 296.600 ;
        RECT 433.200 293.600 434.000 295.200 ;
        RECT 434.800 294.800 435.600 295.000 ;
        RECT 434.800 294.200 439.200 294.800 ;
        RECT 438.400 294.000 439.200 294.200 ;
        RECT 420.400 287.400 421.200 293.000 ;
        RECT 429.800 292.600 431.800 293.400 ;
        RECT 435.600 292.600 438.800 293.400 ;
        RECT 441.200 292.800 442.000 295.600 ;
        RECT 446.000 295.200 446.800 295.800 ;
        RECT 446.000 294.600 447.800 295.200 ;
        RECT 447.000 293.400 447.800 294.600 ;
        RECT 450.800 294.600 451.600 299.800 ;
        RECT 452.400 296.000 453.200 299.800 ;
        RECT 452.400 295.200 453.400 296.000 ;
        RECT 455.600 295.800 456.400 299.800 ;
        RECT 457.200 296.000 458.000 299.800 ;
        RECT 460.400 296.000 461.200 299.800 ;
        RECT 457.200 295.800 461.200 296.000 ;
        RECT 450.800 294.000 452.000 294.600 ;
        RECT 447.000 292.600 450.800 293.400 ;
        RECT 421.800 292.000 422.600 292.200 ;
        RECT 426.800 292.000 427.600 292.400 ;
        RECT 433.200 292.000 434.000 292.400 ;
        RECT 444.400 292.000 445.200 292.600 ;
        RECT 451.400 292.000 452.000 294.000 ;
        RECT 421.800 291.400 445.200 292.000 ;
        RECT 451.200 291.400 452.000 292.000 ;
        RECT 451.200 289.600 451.800 291.400 ;
        RECT 452.600 290.800 453.400 295.200 ;
        RECT 455.800 294.400 456.400 295.800 ;
        RECT 457.400 295.400 461.000 295.800 ;
        RECT 459.600 294.400 460.400 294.800 ;
        RECT 454.000 294.300 454.800 294.400 ;
        RECT 455.600 294.300 458.200 294.400 ;
        RECT 454.000 293.700 458.200 294.300 ;
        RECT 459.600 294.300 461.200 294.400 ;
        RECT 462.000 294.300 462.800 299.800 ;
        RECT 463.600 295.600 464.400 297.200 ;
        RECT 465.200 296.000 466.000 299.800 ;
        RECT 468.400 296.000 469.200 299.800 ;
        RECT 465.200 295.800 469.200 296.000 ;
        RECT 470.000 295.800 470.800 299.800 ;
        RECT 475.400 296.400 476.200 299.000 ;
        RECT 479.600 297.000 480.400 299.000 ;
        RECT 475.400 296.000 477.200 296.400 ;
        RECT 465.400 295.400 469.000 295.800 ;
        RECT 466.000 294.400 466.800 294.800 ;
        RECT 470.000 294.400 470.600 295.800 ;
        RECT 474.600 295.600 477.200 296.000 ;
        RECT 474.600 295.400 476.200 295.600 ;
        RECT 474.600 295.000 475.400 295.400 ;
        RECT 474.600 294.400 475.200 295.000 ;
        RECT 479.800 294.800 480.400 297.000 ;
        RECT 481.200 296.000 482.000 299.800 ;
        RECT 484.400 296.000 485.200 299.800 ;
        RECT 481.200 295.800 485.200 296.000 ;
        RECT 486.000 295.800 486.800 299.800 ;
        RECT 481.400 295.400 485.000 295.800 ;
        RECT 459.600 293.800 462.800 294.300 ;
        RECT 454.000 293.600 454.800 293.700 ;
        RECT 455.600 293.600 458.200 293.700 ;
        RECT 460.400 293.700 462.800 293.800 ;
        RECT 460.400 293.600 461.200 293.700 ;
        RECT 430.000 289.400 430.800 289.600 ;
        RECT 425.400 289.000 430.800 289.400 ;
        RECT 424.600 288.800 430.800 289.000 ;
        RECT 431.800 289.000 440.400 289.600 ;
        RECT 422.000 288.000 423.600 288.800 ;
        RECT 424.600 288.200 426.000 288.800 ;
        RECT 431.800 288.200 432.400 289.000 ;
        RECT 439.600 288.800 440.400 289.000 ;
        RECT 442.800 289.000 451.800 289.600 ;
        RECT 442.800 288.800 443.600 289.000 ;
        RECT 423.000 287.600 423.600 288.000 ;
        RECT 426.600 287.600 432.400 288.200 ;
        RECT 433.000 287.600 435.600 288.400 ;
        RECT 420.400 286.800 422.400 287.400 ;
        RECT 423.000 286.800 427.200 287.600 ;
        RECT 421.800 286.200 422.400 286.800 ;
        RECT 421.800 285.600 422.800 286.200 ;
        RECT 422.000 282.200 422.800 285.600 ;
        RECT 425.200 282.200 426.000 286.800 ;
        RECT 428.400 282.200 429.200 285.000 ;
        RECT 430.000 282.200 430.800 285.000 ;
        RECT 431.600 282.200 432.400 287.000 ;
        RECT 434.800 282.200 435.600 287.000 ;
        RECT 438.000 282.200 438.800 288.400 ;
        RECT 446.000 287.600 448.600 288.400 ;
        RECT 441.200 286.800 445.400 287.600 ;
        RECT 439.600 282.200 440.400 285.000 ;
        RECT 441.200 282.200 442.000 285.000 ;
        RECT 442.800 282.200 443.600 285.000 ;
        RECT 446.000 282.200 446.800 287.600 ;
        RECT 451.200 287.400 451.800 289.000 ;
        RECT 449.200 286.800 451.800 287.400 ;
        RECT 452.400 290.000 453.400 290.800 ;
        RECT 455.600 290.200 456.400 290.400 ;
        RECT 457.600 290.200 458.200 293.600 ;
        RECT 458.800 291.600 459.600 293.200 ;
        RECT 449.200 282.200 450.000 286.800 ;
        RECT 452.400 282.200 453.200 290.000 ;
        RECT 455.600 289.600 457.000 290.200 ;
        RECT 457.600 289.600 458.600 290.200 ;
        RECT 456.400 288.400 457.000 289.600 ;
        RECT 456.400 287.600 457.200 288.400 ;
        RECT 457.800 282.200 458.600 289.600 ;
        RECT 462.000 282.200 462.800 293.700 ;
        RECT 465.200 293.800 466.800 294.400 ;
        RECT 468.200 294.300 470.800 294.400 ;
        RECT 471.600 294.300 472.400 294.400 ;
        RECT 465.200 293.600 466.000 293.800 ;
        RECT 468.200 293.700 472.400 294.300 ;
        RECT 468.200 293.600 470.800 293.700 ;
        RECT 471.600 293.600 472.400 293.700 ;
        RECT 473.200 293.600 475.200 294.400 ;
        RECT 476.200 294.200 480.400 294.800 ;
        RECT 482.000 294.400 482.800 294.800 ;
        RECT 486.000 294.400 486.600 295.800 ;
        RECT 487.600 295.400 488.400 299.800 ;
        RECT 491.800 298.400 493.000 299.800 ;
        RECT 491.800 297.800 493.200 298.400 ;
        RECT 496.400 297.800 497.200 299.800 ;
        RECT 500.800 298.400 501.600 299.800 ;
        RECT 500.800 297.800 502.800 298.400 ;
        RECT 492.400 297.000 493.200 297.800 ;
        RECT 496.600 297.200 497.200 297.800 ;
        RECT 496.600 296.600 499.400 297.200 ;
        RECT 498.600 296.400 499.400 296.600 ;
        RECT 500.400 296.400 501.200 297.200 ;
        RECT 502.000 297.000 502.800 297.800 ;
        RECT 490.600 295.400 491.400 295.600 ;
        RECT 487.600 294.800 491.400 295.400 ;
        RECT 476.200 293.800 477.200 294.200 ;
        RECT 463.600 292.300 464.400 292.400 ;
        RECT 466.800 292.300 467.600 293.200 ;
        RECT 463.600 291.700 467.600 292.300 ;
        RECT 463.600 291.600 464.400 291.700 ;
        RECT 466.800 291.600 467.600 291.700 ;
        RECT 468.200 290.200 468.800 293.600 ;
        RECT 473.200 290.800 474.000 292.400 ;
        RECT 470.000 290.200 470.800 290.400 ;
        RECT 467.800 289.600 468.800 290.200 ;
        RECT 469.400 289.600 470.800 290.200 ;
        RECT 474.600 289.800 475.200 293.600 ;
        RECT 475.800 293.000 477.200 293.800 ;
        RECT 481.200 293.800 482.800 294.400 ;
        RECT 481.200 293.600 482.000 293.800 ;
        RECT 484.200 293.600 486.800 294.400 ;
        RECT 476.600 291.000 477.200 293.000 ;
        RECT 478.000 291.600 478.800 293.200 ;
        RECT 479.600 291.600 480.400 293.200 ;
        RECT 482.800 291.600 483.600 293.200 ;
        RECT 476.600 290.400 480.400 291.000 ;
        RECT 467.800 282.200 468.600 289.600 ;
        RECT 469.400 288.400 470.000 289.600 ;
        RECT 474.600 289.200 476.200 289.800 ;
        RECT 469.200 287.600 470.000 288.400 ;
        RECT 475.400 282.200 476.200 289.200 ;
        RECT 479.800 287.000 480.400 290.400 ;
        RECT 484.200 290.200 484.800 293.600 ;
        RECT 487.600 291.400 488.400 294.800 ;
        RECT 500.400 294.400 501.000 296.400 ;
        RECT 505.200 295.000 506.000 299.800 ;
        RECT 506.800 295.600 507.600 297.200 ;
        RECT 494.600 294.200 495.400 294.400 ;
        RECT 500.400 294.200 501.200 294.400 ;
        RECT 503.600 294.200 505.200 294.400 ;
        RECT 494.200 293.600 505.200 294.200 ;
        RECT 492.400 292.800 493.200 293.000 ;
        RECT 489.400 292.200 493.200 292.800 ;
        RECT 489.400 292.000 490.200 292.200 ;
        RECT 491.000 291.400 491.800 291.600 ;
        RECT 487.600 290.800 491.800 291.400 ;
        RECT 486.000 290.200 486.800 290.400 ;
        RECT 479.600 283.000 480.400 287.000 ;
        RECT 483.800 289.600 484.800 290.200 ;
        RECT 485.400 289.600 486.800 290.200 ;
        RECT 483.800 282.200 484.600 289.600 ;
        RECT 485.400 288.400 486.000 289.600 ;
        RECT 485.200 287.600 486.000 288.400 ;
        RECT 487.600 282.200 488.400 290.800 ;
        RECT 494.200 290.400 494.800 293.600 ;
        RECT 501.400 293.400 502.200 293.600 ;
        RECT 503.000 292.400 503.800 292.600 ;
        RECT 497.200 292.300 498.000 292.400 ;
        RECT 498.800 292.300 503.800 292.400 ;
        RECT 497.200 291.800 503.800 292.300 ;
        RECT 497.200 291.700 499.600 291.800 ;
        RECT 497.200 291.600 498.000 291.700 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 500.400 291.000 506.000 291.200 ;
        RECT 500.200 290.800 506.000 291.000 ;
        RECT 492.400 289.800 494.800 290.400 ;
        RECT 496.200 290.600 506.000 290.800 ;
        RECT 496.200 290.200 501.000 290.600 ;
        RECT 492.400 288.800 493.000 289.800 ;
        RECT 491.600 288.000 493.000 288.800 ;
        RECT 494.600 289.000 495.400 289.200 ;
        RECT 496.200 289.000 496.800 290.200 ;
        RECT 494.600 288.400 496.800 289.000 ;
        RECT 497.400 289.000 502.800 289.600 ;
        RECT 497.400 288.800 498.200 289.000 ;
        RECT 502.000 288.800 502.800 289.000 ;
        RECT 495.800 287.400 496.600 287.600 ;
        RECT 498.600 287.400 499.400 287.600 ;
        RECT 492.400 286.200 493.200 287.000 ;
        RECT 495.800 286.800 499.400 287.400 ;
        RECT 496.600 286.200 497.200 286.800 ;
        RECT 502.000 286.200 502.800 287.000 ;
        RECT 491.800 282.200 493.000 286.200 ;
        RECT 496.400 282.200 497.200 286.200 ;
        RECT 500.800 285.600 502.800 286.200 ;
        RECT 500.800 282.200 501.600 285.600 ;
        RECT 505.200 282.200 506.000 290.600 ;
        RECT 508.400 282.200 509.200 299.800 ;
        RECT 513.800 296.000 514.600 299.000 ;
        RECT 518.000 297.000 518.800 299.000 ;
        RECT 513.000 295.400 514.600 296.000 ;
        RECT 513.000 295.000 513.800 295.400 ;
        RECT 513.000 294.400 513.600 295.000 ;
        RECT 518.200 294.800 518.800 297.000 ;
        RECT 519.600 295.800 520.400 299.800 ;
        RECT 521.200 296.000 522.000 299.800 ;
        RECT 524.400 296.000 525.200 299.800 ;
        RECT 521.200 295.800 525.200 296.000 ;
        RECT 526.000 296.000 526.800 299.800 ;
        RECT 529.200 296.000 530.000 299.800 ;
        RECT 526.000 295.800 530.000 296.000 ;
        RECT 530.800 295.800 531.600 299.800 ;
        RECT 532.400 297.000 533.200 299.000 ;
        RECT 511.600 293.600 513.600 294.400 ;
        RECT 514.600 294.200 518.800 294.800 ;
        RECT 519.800 294.400 520.400 295.800 ;
        RECT 521.400 295.400 525.000 295.800 ;
        RECT 526.200 295.400 529.800 295.800 ;
        RECT 523.600 294.400 524.400 294.800 ;
        RECT 526.800 294.400 527.600 294.800 ;
        RECT 530.800 294.400 531.400 295.800 ;
        RECT 532.400 294.800 533.000 297.000 ;
        RECT 536.600 296.000 537.400 299.000 ;
        RECT 536.600 295.400 538.200 296.000 ;
        RECT 542.000 295.800 542.800 299.800 ;
        RECT 543.600 296.000 544.400 299.800 ;
        RECT 546.800 296.000 547.600 299.800 ;
        RECT 543.600 295.800 547.600 296.000 ;
        RECT 537.400 295.000 538.200 295.400 ;
        RECT 514.600 293.800 515.600 294.200 ;
        RECT 511.600 290.800 512.400 292.400 ;
        RECT 513.000 289.800 513.600 293.600 ;
        RECT 514.200 293.000 515.600 293.800 ;
        RECT 519.600 293.600 522.200 294.400 ;
        RECT 523.600 294.300 525.200 294.400 ;
        RECT 526.000 294.300 527.600 294.400 ;
        RECT 523.600 293.800 527.600 294.300 ;
        RECT 524.400 293.700 526.800 293.800 ;
        RECT 524.400 293.600 525.200 293.700 ;
        RECT 526.000 293.600 526.800 293.700 ;
        RECT 529.000 293.600 531.600 294.400 ;
        RECT 532.400 294.200 536.600 294.800 ;
        RECT 535.600 293.800 536.600 294.200 ;
        RECT 537.600 294.400 538.200 295.000 ;
        RECT 542.200 294.400 542.800 295.800 ;
        RECT 543.800 295.400 547.400 295.800 ;
        RECT 546.000 294.400 546.800 294.800 ;
        RECT 515.000 291.000 515.600 293.000 ;
        RECT 516.400 291.600 517.200 293.200 ;
        RECT 518.000 291.600 518.800 293.200 ;
        RECT 521.600 292.400 522.200 293.600 ;
        RECT 521.200 291.600 522.200 292.400 ;
        RECT 522.800 292.300 523.600 293.200 ;
        RECT 527.600 292.300 528.400 293.200 ;
        RECT 522.800 291.700 528.400 292.300 ;
        RECT 522.800 291.600 523.600 291.700 ;
        RECT 527.600 291.600 528.400 291.700 ;
        RECT 515.000 290.400 518.800 291.000 ;
        RECT 513.000 289.200 514.600 289.800 ;
        RECT 513.800 284.400 514.600 289.200 ;
        RECT 518.200 287.000 518.800 290.400 ;
        RECT 519.600 290.200 520.400 290.400 ;
        RECT 521.600 290.200 522.200 291.600 ;
        RECT 529.000 290.200 529.600 293.600 ;
        RECT 532.400 291.600 533.200 293.200 ;
        RECT 534.000 291.600 534.800 293.200 ;
        RECT 535.600 293.000 537.000 293.800 ;
        RECT 537.600 293.600 539.600 294.400 ;
        RECT 542.000 293.600 544.600 294.400 ;
        RECT 546.000 294.300 547.600 294.400 ;
        RECT 548.400 294.300 549.200 299.800 ;
        RECT 550.000 295.600 550.800 297.200 ;
        RECT 551.600 295.200 552.400 299.800 ;
        RECT 554.800 296.400 555.600 299.800 ;
        RECT 554.800 295.800 555.800 296.400 ;
        RECT 551.600 294.600 554.200 295.200 ;
        RECT 546.000 293.800 549.200 294.300 ;
        RECT 546.800 293.700 549.200 293.800 ;
        RECT 546.800 293.600 547.600 293.700 ;
        RECT 535.600 291.000 536.200 293.000 ;
        RECT 532.400 290.400 536.200 291.000 ;
        RECT 530.800 290.200 531.600 290.400 ;
        RECT 519.600 289.600 521.000 290.200 ;
        RECT 521.600 289.600 522.600 290.200 ;
        RECT 520.400 288.400 521.000 289.600 ;
        RECT 520.400 287.600 521.200 288.400 ;
        RECT 513.800 283.600 515.600 284.400 ;
        RECT 513.800 282.200 514.600 283.600 ;
        RECT 518.000 283.000 518.800 287.000 ;
        RECT 521.800 282.200 522.600 289.600 ;
        RECT 528.600 289.600 529.600 290.200 ;
        RECT 530.200 289.600 531.600 290.200 ;
        RECT 528.600 284.400 529.400 289.600 ;
        RECT 530.200 288.400 530.800 289.600 ;
        RECT 530.000 287.600 530.800 288.400 ;
        RECT 527.600 283.600 529.400 284.400 ;
        RECT 528.600 282.200 529.400 283.600 ;
        RECT 532.400 287.000 533.000 290.400 ;
        RECT 537.600 289.800 538.200 293.600 ;
        RECT 538.800 290.800 539.600 292.400 ;
        RECT 536.600 289.200 538.200 289.800 ;
        RECT 542.000 290.200 542.800 290.400 ;
        RECT 544.000 290.200 544.600 293.600 ;
        RECT 545.200 291.600 546.000 293.200 ;
        RECT 542.000 289.600 543.400 290.200 ;
        RECT 544.000 289.600 545.000 290.200 ;
        RECT 532.400 283.000 533.200 287.000 ;
        RECT 536.600 284.400 537.400 289.200 ;
        RECT 542.800 288.400 543.400 289.600 ;
        RECT 542.800 287.600 543.600 288.400 ;
        RECT 535.600 283.600 537.400 284.400 ;
        RECT 536.600 282.200 537.400 283.600 ;
        RECT 544.200 282.200 545.000 289.600 ;
        RECT 548.400 282.200 549.200 293.700 ;
        RECT 551.800 292.400 552.600 293.200 ;
        RECT 551.600 291.600 552.600 292.400 ;
        RECT 553.600 293.000 554.200 294.600 ;
        RECT 555.200 294.400 555.800 295.800 ;
        RECT 558.000 295.000 558.800 299.800 ;
        RECT 562.400 298.400 563.200 299.800 ;
        RECT 561.200 297.800 563.200 298.400 ;
        RECT 566.800 297.800 567.600 299.800 ;
        RECT 571.000 298.400 572.200 299.800 ;
        RECT 570.800 297.800 572.200 298.400 ;
        RECT 575.600 298.300 576.400 299.800 ;
        RECT 580.400 298.300 581.200 298.400 ;
        RECT 561.200 297.000 562.000 297.800 ;
        RECT 566.800 297.200 567.400 297.800 ;
        RECT 562.800 296.400 563.600 297.200 ;
        RECT 564.600 296.600 567.400 297.200 ;
        RECT 570.800 297.000 571.600 297.800 ;
        RECT 575.600 297.700 581.200 298.300 ;
        RECT 564.600 296.400 565.400 296.600 ;
        RECT 554.800 293.600 555.800 294.400 ;
        RECT 558.800 294.200 560.400 294.400 ;
        RECT 563.000 294.200 563.600 296.400 ;
        RECT 572.600 295.400 573.400 295.600 ;
        RECT 575.600 295.400 576.400 297.700 ;
        RECT 580.400 297.600 581.200 297.700 ;
        RECT 572.600 294.800 576.400 295.400 ;
        RECT 568.600 294.200 569.400 294.400 ;
        RECT 558.800 293.600 569.800 294.200 ;
        RECT 553.600 292.200 554.600 293.000 ;
        RECT 553.600 290.200 554.200 292.200 ;
        RECT 555.200 290.200 555.800 293.600 ;
        RECT 561.800 293.400 562.600 293.600 ;
        RECT 560.200 292.400 561.000 292.600 ;
        RECT 569.200 292.400 569.800 293.600 ;
        RECT 570.800 292.800 571.600 293.000 ;
        RECT 560.200 291.800 565.200 292.400 ;
        RECT 564.400 291.600 565.200 291.800 ;
        RECT 569.200 291.600 570.000 292.400 ;
        RECT 570.800 292.200 574.600 292.800 ;
        RECT 573.800 292.000 574.600 292.200 ;
        RECT 551.600 289.600 554.200 290.200 ;
        RECT 551.600 282.200 552.400 289.600 ;
        RECT 554.800 289.200 555.800 290.200 ;
        RECT 558.000 291.000 563.600 291.200 ;
        RECT 558.000 290.800 563.800 291.000 ;
        RECT 558.000 290.600 567.800 290.800 ;
        RECT 554.800 282.200 555.600 289.200 ;
        RECT 558.000 282.200 558.800 290.600 ;
        RECT 563.000 290.200 567.800 290.600 ;
        RECT 561.200 289.000 566.600 289.600 ;
        RECT 561.200 288.800 562.000 289.000 ;
        RECT 565.800 288.800 566.600 289.000 ;
        RECT 567.200 289.000 567.800 290.200 ;
        RECT 569.200 290.400 569.800 291.600 ;
        RECT 572.200 291.400 573.000 291.600 ;
        RECT 575.600 291.400 576.400 294.800 ;
        RECT 582.000 297.000 582.800 299.000 ;
        RECT 582.000 294.800 582.600 297.000 ;
        RECT 586.200 296.000 587.000 299.000 ;
        RECT 591.600 297.000 592.400 299.000 ;
        RECT 586.200 295.400 587.800 296.000 ;
        RECT 587.000 295.000 587.800 295.400 ;
        RECT 582.000 294.200 586.200 294.800 ;
        RECT 585.200 293.800 586.200 294.200 ;
        RECT 587.200 294.400 587.800 295.000 ;
        RECT 591.600 294.800 592.200 297.000 ;
        RECT 595.800 296.000 596.600 299.000 ;
        RECT 601.200 296.000 602.000 299.800 ;
        RECT 604.400 296.000 605.200 299.800 ;
        RECT 595.800 295.400 597.400 296.000 ;
        RECT 601.200 295.800 605.200 296.000 ;
        RECT 606.000 295.800 606.800 299.800 ;
        RECT 607.600 295.800 608.400 299.800 ;
        RECT 609.200 296.000 610.000 299.800 ;
        RECT 612.400 296.000 613.200 299.800 ;
        RECT 609.200 295.800 613.200 296.000 ;
        RECT 614.000 295.800 614.800 299.800 ;
        RECT 615.600 296.000 616.400 299.800 ;
        RECT 618.800 296.000 619.600 299.800 ;
        RECT 615.600 295.800 619.600 296.000 ;
        RECT 601.400 295.400 605.000 295.800 ;
        RECT 596.600 295.000 597.400 295.400 ;
        RECT 582.000 291.600 582.800 293.200 ;
        RECT 583.600 291.600 584.400 293.200 ;
        RECT 585.200 293.000 586.600 293.800 ;
        RECT 587.200 293.600 589.200 294.400 ;
        RECT 591.600 294.200 595.800 294.800 ;
        RECT 594.800 293.800 595.800 294.200 ;
        RECT 596.800 294.400 597.400 295.000 ;
        RECT 602.000 294.400 602.800 294.800 ;
        RECT 606.000 294.400 606.600 295.800 ;
        RECT 607.800 294.400 608.400 295.800 ;
        RECT 609.400 295.400 613.000 295.800 ;
        RECT 611.600 294.400 612.400 294.800 ;
        RECT 614.200 294.400 614.800 295.800 ;
        RECT 615.800 295.400 619.400 295.800 ;
        RECT 620.400 295.600 621.200 299.800 ;
        RECT 622.000 296.000 622.800 299.800 ;
        RECT 625.200 296.000 626.000 299.800 ;
        RECT 622.000 295.800 626.000 296.000 ;
        RECT 627.400 296.400 628.200 299.800 ;
        RECT 627.400 295.800 629.200 296.400 ;
        RECT 618.000 294.400 618.800 294.800 ;
        RECT 620.600 294.400 621.200 295.600 ;
        RECT 622.200 295.400 625.800 295.800 ;
        RECT 624.400 294.400 625.200 294.800 ;
        RECT 596.800 294.300 598.800 294.400 ;
        RECT 572.200 290.800 576.400 291.400 ;
        RECT 585.200 291.000 585.800 293.000 ;
        RECT 569.200 289.800 571.600 290.400 ;
        RECT 568.600 289.000 569.400 289.200 ;
        RECT 567.200 288.400 569.400 289.000 ;
        RECT 571.000 288.800 571.600 289.800 ;
        RECT 571.000 288.000 572.400 288.800 ;
        RECT 564.600 287.400 565.400 287.600 ;
        RECT 567.400 287.400 568.200 287.600 ;
        RECT 561.200 286.200 562.000 287.000 ;
        RECT 564.600 286.800 568.200 287.400 ;
        RECT 566.800 286.200 567.400 286.800 ;
        RECT 570.800 286.200 571.600 287.000 ;
        RECT 561.200 285.600 563.200 286.200 ;
        RECT 562.400 282.200 563.200 285.600 ;
        RECT 566.800 282.200 567.600 286.200 ;
        RECT 571.000 282.200 572.200 286.200 ;
        RECT 575.600 282.200 576.400 290.800 ;
        RECT 582.000 290.400 585.800 291.000 ;
        RECT 582.000 287.000 582.600 290.400 ;
        RECT 587.200 289.800 587.800 293.600 ;
        RECT 588.400 290.800 589.200 292.400 ;
        RECT 591.600 291.600 592.400 293.200 ;
        RECT 593.200 291.600 594.000 293.200 ;
        RECT 594.800 293.000 596.200 293.800 ;
        RECT 596.800 293.700 600.300 294.300 ;
        RECT 596.800 293.600 598.800 293.700 ;
        RECT 594.800 291.000 595.400 293.000 ;
        RECT 586.200 289.200 587.800 289.800 ;
        RECT 591.600 290.400 595.400 291.000 ;
        RECT 586.200 288.400 587.000 289.200 ;
        RECT 586.200 287.600 587.600 288.400 ;
        RECT 582.000 283.000 582.800 287.000 ;
        RECT 586.200 282.200 587.000 287.600 ;
        RECT 591.600 287.000 592.200 290.400 ;
        RECT 596.800 289.800 597.400 293.600 ;
        RECT 598.000 290.800 598.800 292.400 ;
        RECT 599.700 292.300 600.300 293.700 ;
        RECT 601.200 293.800 602.800 294.400 ;
        RECT 601.200 293.600 602.000 293.800 ;
        RECT 604.200 293.600 606.800 294.400 ;
        RECT 607.600 293.600 610.200 294.400 ;
        RECT 611.600 293.800 613.200 294.400 ;
        RECT 612.400 293.600 613.200 293.800 ;
        RECT 614.000 293.600 616.600 294.400 ;
        RECT 618.000 293.800 619.600 294.400 ;
        RECT 618.800 293.600 619.600 293.800 ;
        RECT 620.400 293.600 623.000 294.400 ;
        RECT 624.400 293.800 626.000 294.400 ;
        RECT 625.200 293.600 626.000 293.800 ;
        RECT 602.800 292.300 603.600 293.200 ;
        RECT 599.700 291.700 603.600 292.300 ;
        RECT 602.800 291.600 603.600 291.700 ;
        RECT 604.200 290.200 604.800 293.600 ;
        RECT 609.600 292.300 610.200 293.600 ;
        RECT 606.100 291.700 610.200 292.300 ;
        RECT 606.100 290.400 606.700 291.700 ;
        RECT 606.000 290.200 606.800 290.400 ;
        RECT 595.800 289.200 597.400 289.800 ;
        RECT 603.800 289.600 604.800 290.200 ;
        RECT 605.400 289.600 606.800 290.200 ;
        RECT 607.600 290.200 608.400 290.400 ;
        RECT 609.600 290.200 610.200 291.700 ;
        RECT 610.800 291.600 611.600 293.200 ;
        RECT 614.000 290.200 614.800 290.400 ;
        RECT 616.000 290.200 616.600 293.600 ;
        RECT 617.200 291.600 618.000 293.200 ;
        RECT 620.400 290.200 621.200 290.400 ;
        RECT 622.400 290.200 623.000 293.600 ;
        RECT 623.600 291.600 624.400 293.200 ;
        RECT 625.200 292.300 626.000 292.400 ;
        RECT 628.400 292.300 629.200 295.800 ;
        RECT 630.000 293.600 630.800 295.200 ;
        RECT 625.200 291.700 629.200 292.300 ;
        RECT 625.200 291.600 626.000 291.700 ;
        RECT 607.600 289.600 609.000 290.200 ;
        RECT 609.600 289.600 610.600 290.200 ;
        RECT 614.000 289.600 615.400 290.200 ;
        RECT 616.000 289.600 617.000 290.200 ;
        RECT 620.400 289.600 621.800 290.200 ;
        RECT 622.400 289.600 623.400 290.200 ;
        RECT 591.600 283.000 592.400 287.000 ;
        RECT 595.800 282.200 596.600 289.200 ;
        RECT 603.800 286.400 604.600 289.600 ;
        RECT 605.400 288.400 606.000 289.600 ;
        RECT 605.200 287.600 606.000 288.400 ;
        RECT 608.400 288.400 609.000 289.600 ;
        RECT 608.400 287.600 609.200 288.400 ;
        RECT 602.800 285.600 604.600 286.400 ;
        RECT 603.800 282.200 604.600 285.600 ;
        RECT 609.800 282.200 610.600 289.600 ;
        RECT 614.800 288.400 615.400 289.600 ;
        RECT 614.800 287.600 615.600 288.400 ;
        RECT 616.200 282.200 617.000 289.600 ;
        RECT 621.200 288.400 621.800 289.600 ;
        RECT 621.200 287.600 622.000 288.400 ;
        RECT 622.600 282.200 623.400 289.600 ;
        RECT 626.800 288.800 627.600 290.400 ;
        RECT 628.400 282.200 629.200 291.700 ;
        RECT 631.600 282.200 632.400 299.800 ;
        RECT 633.200 295.600 634.000 297.200 ;
        RECT 634.800 297.000 635.600 299.000 ;
        RECT 639.000 298.400 639.800 299.000 ;
        RECT 639.000 297.600 640.400 298.400 ;
        RECT 634.800 294.800 635.400 297.000 ;
        RECT 639.000 296.000 639.800 297.600 ;
        RECT 644.400 296.000 645.200 299.800 ;
        RECT 647.600 296.000 648.400 299.800 ;
        RECT 639.000 295.400 640.600 296.000 ;
        RECT 644.400 295.800 648.400 296.000 ;
        RECT 649.200 295.800 650.000 299.800 ;
        RECT 644.600 295.400 648.200 295.800 ;
        RECT 639.800 295.000 640.600 295.400 ;
        RECT 634.800 294.200 639.000 294.800 ;
        RECT 638.000 293.800 639.000 294.200 ;
        RECT 640.000 294.400 640.600 295.000 ;
        RECT 645.200 294.400 646.000 294.800 ;
        RECT 649.200 294.400 649.800 295.800 ;
        RECT 650.800 295.400 651.600 299.800 ;
        RECT 655.000 298.400 656.200 299.800 ;
        RECT 655.000 297.800 656.400 298.400 ;
        RECT 659.600 297.800 660.400 299.800 ;
        RECT 664.000 298.400 664.800 299.800 ;
        RECT 664.000 297.800 666.000 298.400 ;
        RECT 655.600 297.000 656.400 297.800 ;
        RECT 659.800 297.200 660.400 297.800 ;
        RECT 659.800 296.600 662.600 297.200 ;
        RECT 661.800 296.400 662.600 296.600 ;
        RECT 663.600 296.400 664.400 297.200 ;
        RECT 665.200 297.000 666.000 297.800 ;
        RECT 653.800 295.400 654.600 295.600 ;
        RECT 650.800 294.800 654.600 295.400 ;
        RECT 634.800 291.600 635.600 293.200 ;
        RECT 636.400 291.600 637.200 293.200 ;
        RECT 638.000 293.000 639.400 293.800 ;
        RECT 640.000 293.600 642.000 294.400 ;
        RECT 644.400 293.800 646.000 294.400 ;
        RECT 644.400 293.600 645.200 293.800 ;
        RECT 647.400 293.600 650.000 294.400 ;
        RECT 638.000 291.000 638.600 293.000 ;
        RECT 634.800 290.400 638.600 291.000 ;
        RECT 634.800 287.000 635.400 290.400 ;
        RECT 640.000 289.800 640.600 293.600 ;
        RECT 641.200 290.800 642.000 292.400 ;
        RECT 646.000 291.600 646.800 293.200 ;
        RECT 647.400 290.200 648.000 293.600 ;
        RECT 650.800 291.400 651.600 294.800 ;
        RECT 657.800 294.200 658.600 294.400 ;
        RECT 663.600 294.200 664.200 296.400 ;
        RECT 668.400 295.000 669.200 299.800 ;
        RECT 671.600 295.200 672.400 299.800 ;
        RECT 674.800 295.200 675.600 299.800 ;
        RECT 678.000 295.200 678.800 299.800 ;
        RECT 681.200 295.200 682.000 299.800 ;
        RECT 671.600 294.400 673.400 295.200 ;
        RECT 674.800 294.400 677.000 295.200 ;
        RECT 678.000 294.400 680.200 295.200 ;
        RECT 681.200 294.400 683.600 295.200 ;
        RECT 666.800 294.200 668.400 294.400 ;
        RECT 657.400 293.600 668.400 294.200 ;
        RECT 670.000 293.800 670.800 294.400 ;
        RECT 672.600 293.800 673.400 294.400 ;
        RECT 676.200 293.800 677.000 294.400 ;
        RECT 679.400 293.800 680.200 294.400 ;
        RECT 655.600 292.800 656.400 293.000 ;
        RECT 652.600 292.200 656.400 292.800 ;
        RECT 652.600 292.000 653.400 292.200 ;
        RECT 654.200 291.400 655.000 291.600 ;
        RECT 650.800 290.800 655.000 291.400 ;
        RECT 649.200 290.300 650.000 290.400 ;
        RECT 650.800 290.300 651.600 290.800 ;
        RECT 657.400 290.400 658.000 293.600 ;
        RECT 664.600 293.400 665.400 293.600 ;
        RECT 670.000 293.000 671.800 293.800 ;
        RECT 672.600 293.000 675.200 293.800 ;
        RECT 676.200 293.000 678.600 293.800 ;
        RECT 679.400 293.000 682.000 293.800 ;
        RECT 666.200 292.400 667.000 292.600 ;
        RECT 662.000 291.800 667.000 292.400 ;
        RECT 662.000 291.600 662.800 291.800 ;
        RECT 672.600 291.600 673.400 293.000 ;
        RECT 676.200 291.600 677.000 293.000 ;
        RECT 679.400 291.600 680.200 293.000 ;
        RECT 682.800 291.600 683.600 294.400 ;
        RECT 663.600 291.000 669.200 291.200 ;
        RECT 663.400 290.800 669.200 291.000 ;
        RECT 649.200 290.200 651.600 290.300 ;
        RECT 639.000 289.200 640.600 289.800 ;
        RECT 647.000 289.600 648.000 290.200 ;
        RECT 648.600 289.700 651.600 290.200 ;
        RECT 648.600 289.600 650.000 289.700 ;
        RECT 634.800 283.000 635.600 287.000 ;
        RECT 639.000 282.200 639.800 289.200 ;
        RECT 647.000 282.200 647.800 289.600 ;
        RECT 648.600 288.400 649.200 289.600 ;
        RECT 648.400 287.600 649.200 288.400 ;
        RECT 650.800 282.200 651.600 289.700 ;
        RECT 655.600 289.800 658.000 290.400 ;
        RECT 659.400 290.600 669.200 290.800 ;
        RECT 659.400 290.200 664.200 290.600 ;
        RECT 655.600 288.800 656.200 289.800 ;
        RECT 654.800 288.000 656.200 288.800 ;
        RECT 657.800 289.000 658.600 289.200 ;
        RECT 659.400 289.000 660.000 290.200 ;
        RECT 657.800 288.400 660.000 289.000 ;
        RECT 660.600 289.000 666.000 289.600 ;
        RECT 660.600 288.800 661.400 289.000 ;
        RECT 665.200 288.800 666.000 289.000 ;
        RECT 659.000 287.400 659.800 287.600 ;
        RECT 661.800 287.400 662.600 287.600 ;
        RECT 655.600 286.200 656.400 287.000 ;
        RECT 659.000 286.800 662.600 287.400 ;
        RECT 659.800 286.200 660.400 286.800 ;
        RECT 665.200 286.200 666.000 287.000 ;
        RECT 655.000 282.200 656.200 286.200 ;
        RECT 659.600 282.200 660.400 286.200 ;
        RECT 664.000 285.600 666.000 286.200 ;
        RECT 664.000 282.200 664.800 285.600 ;
        RECT 668.400 282.200 669.200 290.600 ;
        RECT 671.600 290.800 673.400 291.600 ;
        RECT 674.800 290.800 677.000 291.600 ;
        RECT 678.000 290.800 680.200 291.600 ;
        RECT 681.200 290.800 683.600 291.600 ;
        RECT 671.600 282.200 672.400 290.800 ;
        RECT 674.800 282.200 675.600 290.800 ;
        RECT 678.000 282.200 678.800 290.800 ;
        RECT 681.200 282.200 682.000 290.800 ;
        RECT 2.800 276.400 3.600 279.800 ;
        RECT 2.600 275.800 3.600 276.400 ;
        RECT 2.600 275.200 3.200 275.800 ;
        RECT 6.000 275.200 6.800 279.800 ;
        RECT 9.200 277.000 10.000 279.800 ;
        RECT 10.800 277.000 11.600 279.800 ;
        RECT 1.200 274.600 3.200 275.200 ;
        RECT 1.200 269.000 2.000 274.600 ;
        RECT 3.800 274.400 8.000 275.200 ;
        RECT 12.400 275.000 13.200 279.800 ;
        RECT 15.600 275.000 16.400 279.800 ;
        RECT 3.800 274.000 4.400 274.400 ;
        RECT 2.800 273.200 4.400 274.000 ;
        RECT 7.400 273.800 13.200 274.400 ;
        RECT 5.400 273.200 6.800 273.800 ;
        RECT 5.400 273.000 11.600 273.200 ;
        RECT 6.200 272.600 11.600 273.000 ;
        RECT 10.800 272.400 11.600 272.600 ;
        RECT 12.600 273.000 13.200 273.800 ;
        RECT 13.800 273.600 16.400 274.400 ;
        RECT 18.800 273.600 19.600 279.800 ;
        RECT 20.400 277.000 21.200 279.800 ;
        RECT 22.000 277.000 22.800 279.800 ;
        RECT 23.600 277.000 24.400 279.800 ;
        RECT 22.000 274.400 26.200 275.200 ;
        RECT 26.800 274.400 27.600 279.800 ;
        RECT 30.000 275.200 30.800 279.800 ;
        RECT 30.000 274.600 32.600 275.200 ;
        RECT 26.800 273.600 29.400 274.400 ;
        RECT 20.400 273.000 21.200 273.200 ;
        RECT 12.600 272.400 21.200 273.000 ;
        RECT 23.600 273.000 24.400 273.200 ;
        RECT 32.000 273.000 32.600 274.600 ;
        RECT 23.600 272.400 32.600 273.000 ;
        RECT 32.000 270.600 32.600 272.400 ;
        RECT 33.200 272.000 34.000 279.800 ;
        RECT 33.200 271.200 34.200 272.000 ;
        RECT 38.000 271.200 38.800 279.800 ;
        RECT 41.200 271.200 42.000 279.800 ;
        RECT 44.400 271.200 45.200 279.800 ;
        RECT 47.600 271.200 48.400 279.800 ;
        RECT 51.600 273.600 52.400 274.400 ;
        RECT 51.600 272.400 52.200 273.600 ;
        RECT 53.000 272.400 53.800 279.800 ;
        RECT 50.800 271.800 52.200 272.400 ;
        RECT 52.800 271.800 53.800 272.400 ;
        RECT 50.800 271.600 51.600 271.800 ;
        RECT 2.600 270.000 26.000 270.600 ;
        RECT 32.000 270.000 32.800 270.600 ;
        RECT 2.600 269.800 3.400 270.000 ;
        RECT 7.600 269.600 8.400 270.000 ;
        RECT 25.200 269.400 26.000 270.000 ;
        RECT 1.200 268.200 10.000 269.000 ;
        RECT 10.600 268.600 12.600 269.400 ;
        RECT 16.400 268.600 19.600 269.400 ;
        RECT 1.200 262.200 2.000 268.200 ;
        RECT 3.600 266.800 6.600 267.600 ;
        RECT 5.800 266.200 6.600 266.800 ;
        RECT 11.800 266.200 12.600 268.600 ;
        RECT 14.000 266.800 14.800 268.400 ;
        RECT 19.200 267.800 20.000 268.000 ;
        RECT 15.600 267.200 20.000 267.800 ;
        RECT 15.600 267.000 16.400 267.200 ;
        RECT 22.000 266.400 22.800 269.200 ;
        RECT 27.800 268.600 31.600 269.400 ;
        RECT 27.800 267.400 28.600 268.600 ;
        RECT 32.200 268.000 32.800 270.000 ;
        RECT 15.600 266.200 16.400 266.400 ;
        RECT 5.800 265.400 8.400 266.200 ;
        RECT 11.800 265.600 16.400 266.200 ;
        RECT 17.200 265.600 18.800 266.400 ;
        RECT 21.800 265.600 22.800 266.400 ;
        RECT 26.800 266.800 28.600 267.400 ;
        RECT 31.600 267.400 32.800 268.000 ;
        RECT 26.800 266.200 27.600 266.800 ;
        RECT 7.600 262.200 8.400 265.400 ;
        RECT 25.200 265.400 27.600 266.200 ;
        RECT 9.200 262.200 10.000 265.000 ;
        RECT 10.800 262.200 11.600 265.000 ;
        RECT 12.400 262.200 13.200 265.000 ;
        RECT 15.600 262.200 16.400 265.000 ;
        RECT 18.800 262.200 19.600 265.000 ;
        RECT 20.400 262.200 21.200 265.000 ;
        RECT 22.000 262.200 22.800 265.000 ;
        RECT 23.600 262.200 24.400 265.000 ;
        RECT 25.200 262.200 26.000 265.400 ;
        RECT 31.600 262.200 32.400 267.400 ;
        RECT 33.400 266.800 34.200 271.200 ;
        RECT 36.400 270.400 38.800 271.200 ;
        RECT 39.800 270.400 42.000 271.200 ;
        RECT 43.000 270.400 45.200 271.200 ;
        RECT 46.600 270.400 48.400 271.200 ;
        RECT 36.400 267.600 37.200 270.400 ;
        RECT 39.800 269.000 40.600 270.400 ;
        RECT 43.000 269.000 43.800 270.400 ;
        RECT 46.600 269.000 47.400 270.400 ;
        RECT 38.000 268.200 40.600 269.000 ;
        RECT 41.400 268.200 43.800 269.000 ;
        RECT 44.800 268.200 47.400 269.000 ;
        RECT 48.200 268.200 50.000 269.000 ;
        RECT 52.800 268.400 53.400 271.800 ;
        RECT 54.000 268.800 54.800 270.400 ;
        RECT 58.800 270.300 59.600 279.800 ;
        RECT 63.000 272.400 63.800 279.800 ;
        RECT 64.400 273.600 65.200 274.400 ;
        RECT 64.600 272.400 65.200 273.600 ;
        RECT 63.000 271.800 64.000 272.400 ;
        RECT 64.600 271.800 66.000 272.400 ;
        RECT 68.400 272.000 69.200 279.800 ;
        RECT 71.600 275.200 72.400 279.800 ;
        RECT 62.000 270.300 62.800 270.400 ;
        RECT 58.800 269.700 62.800 270.300 ;
        RECT 39.800 267.600 40.600 268.200 ;
        RECT 43.000 267.600 43.800 268.200 ;
        RECT 46.600 267.600 47.400 268.200 ;
        RECT 49.200 267.600 50.000 268.200 ;
        RECT 50.800 267.600 53.400 268.400 ;
        RECT 55.600 268.200 56.400 268.400 ;
        RECT 54.800 267.600 56.400 268.200 ;
        RECT 36.400 266.800 38.800 267.600 ;
        RECT 39.800 266.800 42.000 267.600 ;
        RECT 43.000 266.800 45.200 267.600 ;
        RECT 46.600 266.800 48.400 267.600 ;
        RECT 33.200 266.000 34.200 266.800 ;
        RECT 33.200 262.200 34.000 266.000 ;
        RECT 38.000 262.200 38.800 266.800 ;
        RECT 41.200 262.200 42.000 266.800 ;
        RECT 44.400 262.200 45.200 266.800 ;
        RECT 47.600 262.200 48.400 266.800 ;
        RECT 51.000 266.200 51.600 267.600 ;
        RECT 54.800 267.200 55.600 267.600 ;
        RECT 52.600 266.200 56.200 266.600 ;
        RECT 50.800 262.200 51.600 266.200 ;
        RECT 52.400 266.000 56.400 266.200 ;
        RECT 52.400 262.200 53.200 266.000 ;
        RECT 55.600 262.200 56.400 266.000 ;
        RECT 57.200 264.800 58.000 266.400 ;
        RECT 58.800 262.200 59.600 269.700 ;
        RECT 62.000 268.800 62.800 269.700 ;
        RECT 63.400 268.400 64.000 271.800 ;
        RECT 65.200 271.600 66.000 271.800 ;
        RECT 68.200 271.200 69.200 272.000 ;
        RECT 69.800 274.600 72.400 275.200 ;
        RECT 69.800 273.000 70.400 274.600 ;
        RECT 74.800 274.400 75.600 279.800 ;
        RECT 78.000 277.000 78.800 279.800 ;
        RECT 79.600 277.000 80.400 279.800 ;
        RECT 81.200 277.000 82.000 279.800 ;
        RECT 76.200 274.400 80.400 275.200 ;
        RECT 73.000 273.600 75.600 274.400 ;
        RECT 82.800 273.600 83.600 279.800 ;
        RECT 86.000 275.000 86.800 279.800 ;
        RECT 89.200 275.000 90.000 279.800 ;
        RECT 90.800 277.000 91.600 279.800 ;
        RECT 92.400 277.000 93.200 279.800 ;
        RECT 95.600 275.200 96.400 279.800 ;
        RECT 98.800 276.400 99.600 279.800 ;
        RECT 98.800 275.800 99.800 276.400 ;
        RECT 99.200 275.200 99.800 275.800 ;
        RECT 94.400 274.400 98.600 275.200 ;
        RECT 99.200 274.600 101.200 275.200 ;
        RECT 86.000 273.600 88.600 274.400 ;
        RECT 89.200 273.800 95.000 274.400 ;
        RECT 98.000 274.000 98.600 274.400 ;
        RECT 78.000 273.000 78.800 273.200 ;
        RECT 69.800 272.400 78.800 273.000 ;
        RECT 81.200 273.000 82.000 273.200 ;
        RECT 89.200 273.000 89.800 273.800 ;
        RECT 95.600 273.200 97.000 273.800 ;
        RECT 98.000 273.200 99.600 274.000 ;
        RECT 81.200 272.400 89.800 273.000 ;
        RECT 90.800 273.000 97.000 273.200 ;
        RECT 90.800 272.600 96.200 273.000 ;
        RECT 90.800 272.400 91.600 272.600 ;
        RECT 60.400 268.200 61.200 268.400 ;
        RECT 60.400 267.600 62.000 268.200 ;
        RECT 63.400 267.600 66.000 268.400 ;
        RECT 61.200 267.200 62.000 267.600 ;
        RECT 60.600 266.200 64.200 266.600 ;
        RECT 65.200 266.200 65.800 267.600 ;
        RECT 68.200 266.800 69.000 271.200 ;
        RECT 69.800 270.600 70.400 272.400 ;
        RECT 69.600 270.000 70.400 270.600 ;
        RECT 76.400 270.000 99.800 270.600 ;
        RECT 69.600 268.000 70.200 270.000 ;
        RECT 76.400 269.400 77.200 270.000 ;
        RECT 94.000 269.600 94.800 270.000 ;
        RECT 97.200 269.600 98.000 270.000 ;
        RECT 99.000 269.800 99.800 270.000 ;
        RECT 70.800 268.600 74.600 269.400 ;
        RECT 69.600 267.400 70.800 268.000 ;
        RECT 60.400 266.000 64.400 266.200 ;
        RECT 60.400 262.200 61.200 266.000 ;
        RECT 63.600 262.200 64.400 266.000 ;
        RECT 65.200 262.200 66.000 266.200 ;
        RECT 68.200 266.000 69.200 266.800 ;
        RECT 68.400 262.200 69.200 266.000 ;
        RECT 70.000 262.200 70.800 267.400 ;
        RECT 73.800 267.400 74.600 268.600 ;
        RECT 73.800 266.800 75.600 267.400 ;
        RECT 74.800 266.200 75.600 266.800 ;
        RECT 79.600 266.400 80.400 269.200 ;
        RECT 82.800 268.600 86.000 269.400 ;
        RECT 89.800 268.600 91.800 269.400 ;
        RECT 100.400 269.000 101.200 274.600 ;
        RECT 82.400 267.800 83.200 268.000 ;
        RECT 82.400 267.200 86.800 267.800 ;
        RECT 86.000 267.000 86.800 267.200 ;
        RECT 87.600 266.800 88.400 268.400 ;
        RECT 74.800 265.400 77.200 266.200 ;
        RECT 79.600 265.600 80.600 266.400 ;
        RECT 83.600 265.600 85.200 266.400 ;
        RECT 86.000 266.200 86.800 266.400 ;
        RECT 89.800 266.200 90.600 268.600 ;
        RECT 92.400 268.200 101.200 269.000 ;
        RECT 95.800 266.800 98.800 267.600 ;
        RECT 95.800 266.200 96.600 266.800 ;
        RECT 86.000 265.600 90.600 266.200 ;
        RECT 76.400 262.200 77.200 265.400 ;
        RECT 94.000 265.400 96.600 266.200 ;
        RECT 78.000 262.200 78.800 265.000 ;
        RECT 79.600 262.200 80.400 265.000 ;
        RECT 81.200 262.200 82.000 265.000 ;
        RECT 82.800 262.200 83.600 265.000 ;
        RECT 86.000 262.200 86.800 265.000 ;
        RECT 89.200 262.200 90.000 265.000 ;
        RECT 90.800 262.200 91.600 265.000 ;
        RECT 92.400 262.200 93.200 265.000 ;
        RECT 94.000 262.200 94.800 265.400 ;
        RECT 100.400 262.200 101.200 268.200 ;
        RECT 102.000 262.200 102.800 279.800 ;
        RECT 103.600 264.800 104.400 266.400 ;
        RECT 105.200 262.200 106.000 279.800 ;
        RECT 108.400 271.600 109.200 273.200 ;
        RECT 110.000 266.400 110.800 279.800 ;
        RECT 119.600 271.200 120.400 279.800 ;
        RECT 122.800 271.200 123.600 279.800 ;
        RECT 126.000 271.200 126.800 279.800 ;
        RECT 129.200 271.200 130.000 279.800 ;
        RECT 118.000 270.400 120.400 271.200 ;
        RECT 121.400 270.400 123.600 271.200 ;
        RECT 124.600 270.400 126.800 271.200 ;
        RECT 128.200 270.400 130.000 271.200 ;
        RECT 111.600 266.800 112.400 268.400 ;
        RECT 118.000 267.600 118.800 270.400 ;
        RECT 121.400 269.000 122.200 270.400 ;
        RECT 124.600 269.000 125.400 270.400 ;
        RECT 128.200 269.000 129.000 270.400 ;
        RECT 119.600 268.200 122.200 269.000 ;
        RECT 123.000 268.200 125.400 269.000 ;
        RECT 126.400 268.200 129.000 269.000 ;
        RECT 129.800 268.200 131.600 269.000 ;
        RECT 121.400 267.600 122.200 268.200 ;
        RECT 124.600 267.600 125.400 268.200 ;
        RECT 128.200 267.600 129.000 268.200 ;
        RECT 130.800 267.600 131.600 268.200 ;
        RECT 118.000 266.800 120.400 267.600 ;
        RECT 121.400 266.800 123.600 267.600 ;
        RECT 124.600 266.800 126.800 267.600 ;
        RECT 128.200 266.800 130.000 267.600 ;
        RECT 106.800 264.800 107.600 266.400 ;
        RECT 108.400 265.600 110.800 266.400 ;
        RECT 109.000 262.200 109.800 265.600 ;
        RECT 119.600 262.200 120.400 266.800 ;
        RECT 122.800 262.200 123.600 266.800 ;
        RECT 126.000 262.200 126.800 266.800 ;
        RECT 129.200 262.200 130.000 266.800 ;
        RECT 132.400 262.200 133.200 279.800 ;
        RECT 137.200 272.000 138.000 279.800 ;
        RECT 140.400 275.200 141.200 279.800 ;
        RECT 137.000 271.200 138.000 272.000 ;
        RECT 138.600 274.600 141.200 275.200 ;
        RECT 138.600 273.000 139.200 274.600 ;
        RECT 143.600 274.400 144.400 279.800 ;
        RECT 146.800 277.000 147.600 279.800 ;
        RECT 148.400 277.000 149.200 279.800 ;
        RECT 150.000 277.000 150.800 279.800 ;
        RECT 145.000 274.400 149.200 275.200 ;
        RECT 141.800 273.600 144.400 274.400 ;
        RECT 151.600 273.600 152.400 279.800 ;
        RECT 154.800 275.000 155.600 279.800 ;
        RECT 158.000 275.000 158.800 279.800 ;
        RECT 159.600 277.000 160.400 279.800 ;
        RECT 161.200 277.000 162.000 279.800 ;
        RECT 164.400 275.200 165.200 279.800 ;
        RECT 167.600 276.400 168.400 279.800 ;
        RECT 167.600 275.800 168.600 276.400 ;
        RECT 168.000 275.200 168.600 275.800 ;
        RECT 163.200 274.400 167.400 275.200 ;
        RECT 168.000 274.600 170.000 275.200 ;
        RECT 154.800 273.600 157.400 274.400 ;
        RECT 158.000 273.800 163.800 274.400 ;
        RECT 166.800 274.000 167.400 274.400 ;
        RECT 146.800 273.000 147.600 273.200 ;
        RECT 138.600 272.400 147.600 273.000 ;
        RECT 150.000 273.000 150.800 273.200 ;
        RECT 158.000 273.000 158.600 273.800 ;
        RECT 164.400 273.200 165.800 273.800 ;
        RECT 166.800 273.200 168.400 274.000 ;
        RECT 150.000 272.400 158.600 273.000 ;
        RECT 159.600 273.000 165.800 273.200 ;
        RECT 159.600 272.600 165.000 273.000 ;
        RECT 159.600 272.400 160.400 272.600 ;
        RECT 137.000 266.800 137.800 271.200 ;
        RECT 138.600 270.600 139.200 272.400 ;
        RECT 138.400 270.000 139.200 270.600 ;
        RECT 145.200 270.000 168.600 270.600 ;
        RECT 138.400 268.000 139.000 270.000 ;
        RECT 145.200 269.400 146.000 270.000 ;
        RECT 162.800 269.600 163.600 270.000 ;
        RECT 164.400 269.600 165.200 270.000 ;
        RECT 167.800 269.800 168.600 270.000 ;
        RECT 139.600 268.600 143.400 269.400 ;
        RECT 138.400 267.400 139.600 268.000 ;
        RECT 134.000 264.800 134.800 266.400 ;
        RECT 137.000 266.000 138.000 266.800 ;
        RECT 137.200 262.200 138.000 266.000 ;
        RECT 138.800 262.200 139.600 267.400 ;
        RECT 142.600 267.400 143.400 268.600 ;
        RECT 142.600 266.800 144.400 267.400 ;
        RECT 143.600 266.200 144.400 266.800 ;
        RECT 148.400 266.400 149.200 269.200 ;
        RECT 151.600 268.600 154.800 269.400 ;
        RECT 158.600 268.600 160.600 269.400 ;
        RECT 169.200 269.000 170.000 274.600 ;
        RECT 170.800 271.600 171.600 273.200 ;
        RECT 151.200 267.800 152.000 268.000 ;
        RECT 151.200 267.200 155.600 267.800 ;
        RECT 154.800 267.000 155.600 267.200 ;
        RECT 156.400 266.800 157.200 268.400 ;
        RECT 143.600 265.400 146.000 266.200 ;
        RECT 148.400 265.600 149.400 266.400 ;
        RECT 152.400 265.600 154.000 266.400 ;
        RECT 154.800 266.200 155.600 266.400 ;
        RECT 158.600 266.200 159.400 268.600 ;
        RECT 161.200 268.200 170.000 269.000 ;
        RECT 164.600 266.800 167.600 267.600 ;
        RECT 164.600 266.200 165.400 266.800 ;
        RECT 154.800 265.600 159.400 266.200 ;
        RECT 145.200 262.200 146.000 265.400 ;
        RECT 162.800 265.400 165.400 266.200 ;
        RECT 146.800 262.200 147.600 265.000 ;
        RECT 148.400 262.200 149.200 265.000 ;
        RECT 150.000 262.200 150.800 265.000 ;
        RECT 151.600 262.200 152.400 265.000 ;
        RECT 154.800 262.200 155.600 265.000 ;
        RECT 158.000 262.200 158.800 265.000 ;
        RECT 159.600 262.200 160.400 265.000 ;
        RECT 161.200 262.200 162.000 265.000 ;
        RECT 162.800 262.200 163.600 265.400 ;
        RECT 169.200 262.200 170.000 268.200 ;
        RECT 170.800 268.300 171.600 268.400 ;
        RECT 172.400 268.300 173.200 279.800 ;
        RECT 176.400 273.600 177.200 274.400 ;
        RECT 176.400 272.400 177.000 273.600 ;
        RECT 177.800 272.400 178.600 279.800 ;
        RECT 183.600 272.800 184.400 279.800 ;
        RECT 174.000 272.300 174.800 272.400 ;
        RECT 175.600 272.300 177.000 272.400 ;
        RECT 174.000 271.800 177.000 272.300 ;
        RECT 177.600 271.800 178.600 272.400 ;
        RECT 183.400 271.800 184.400 272.800 ;
        RECT 186.800 272.400 187.600 279.800 ;
        RECT 185.000 271.800 187.600 272.400 ;
        RECT 190.000 272.000 190.800 279.800 ;
        RECT 193.200 275.200 194.000 279.800 ;
        RECT 174.000 271.700 176.400 271.800 ;
        RECT 174.000 271.600 174.800 271.700 ;
        RECT 175.600 271.600 176.400 271.700 ;
        RECT 177.600 268.400 178.200 271.800 ;
        RECT 178.800 268.800 179.600 270.400 ;
        RECT 183.400 268.400 184.000 271.800 ;
        RECT 185.000 269.800 185.600 271.800 ;
        RECT 184.600 269.000 185.600 269.800 ;
        RECT 170.800 267.700 173.200 268.300 ;
        RECT 170.800 267.600 171.600 267.700 ;
        RECT 172.400 266.200 173.200 267.700 ;
        RECT 174.000 268.300 174.800 268.400 ;
        RECT 175.600 268.300 178.200 268.400 ;
        RECT 174.000 267.700 178.200 268.300 ;
        RECT 180.400 268.200 181.200 268.400 ;
        RECT 174.000 266.800 174.800 267.700 ;
        RECT 175.600 267.600 178.200 267.700 ;
        RECT 179.600 267.600 181.200 268.200 ;
        RECT 183.400 267.600 184.400 268.400 ;
        RECT 175.800 266.200 176.400 267.600 ;
        RECT 179.600 267.200 180.400 267.600 ;
        RECT 177.400 266.200 181.000 266.600 ;
        RECT 183.400 266.200 184.000 267.600 ;
        RECT 185.000 267.400 185.600 269.000 ;
        RECT 189.800 271.200 190.800 272.000 ;
        RECT 191.400 274.600 194.000 275.200 ;
        RECT 191.400 273.000 192.000 274.600 ;
        RECT 196.400 274.400 197.200 279.800 ;
        RECT 199.600 277.000 200.400 279.800 ;
        RECT 201.200 277.000 202.000 279.800 ;
        RECT 202.800 277.000 203.600 279.800 ;
        RECT 197.800 274.400 202.000 275.200 ;
        RECT 194.600 273.600 197.200 274.400 ;
        RECT 204.400 273.600 205.200 279.800 ;
        RECT 207.600 275.000 208.400 279.800 ;
        RECT 210.800 275.000 211.600 279.800 ;
        RECT 212.400 277.000 213.200 279.800 ;
        RECT 214.000 277.000 214.800 279.800 ;
        RECT 217.200 275.200 218.000 279.800 ;
        RECT 220.400 276.400 221.200 279.800 ;
        RECT 224.200 278.400 225.000 279.800 ;
        RECT 223.600 277.600 225.000 278.400 ;
        RECT 220.400 275.800 221.400 276.400 ;
        RECT 220.800 275.200 221.400 275.800 ;
        RECT 216.000 274.400 220.200 275.200 ;
        RECT 220.800 274.600 222.800 275.200 ;
        RECT 207.600 273.600 210.200 274.400 ;
        RECT 210.800 273.800 216.600 274.400 ;
        RECT 219.600 274.000 220.200 274.400 ;
        RECT 199.600 273.000 200.400 273.200 ;
        RECT 191.400 272.400 200.400 273.000 ;
        RECT 202.800 273.000 203.600 273.200 ;
        RECT 210.800 273.000 211.400 273.800 ;
        RECT 217.200 273.200 218.600 273.800 ;
        RECT 219.600 273.200 221.200 274.000 ;
        RECT 202.800 272.400 211.400 273.000 ;
        RECT 212.400 273.000 218.600 273.200 ;
        RECT 212.400 272.600 217.800 273.000 ;
        RECT 212.400 272.400 213.200 272.600 ;
        RECT 185.000 266.800 187.600 267.400 ;
        RECT 171.400 265.600 173.200 266.200 ;
        RECT 171.400 262.200 172.200 265.600 ;
        RECT 175.600 262.200 176.400 266.200 ;
        RECT 177.200 266.000 181.200 266.200 ;
        RECT 177.200 262.200 178.000 266.000 ;
        RECT 180.400 262.200 181.200 266.000 ;
        RECT 183.400 265.600 184.400 266.200 ;
        RECT 183.600 262.200 184.400 265.600 ;
        RECT 186.800 262.200 187.600 266.800 ;
        RECT 189.800 266.800 190.600 271.200 ;
        RECT 191.400 270.600 192.000 272.400 ;
        RECT 191.200 270.000 192.000 270.600 ;
        RECT 198.000 270.000 221.400 270.600 ;
        RECT 191.200 268.000 191.800 270.000 ;
        RECT 198.000 269.400 198.800 270.000 ;
        RECT 215.600 269.600 216.400 270.000 ;
        RECT 218.800 269.600 219.600 270.000 ;
        RECT 220.600 269.800 221.400 270.000 ;
        RECT 192.400 268.600 196.200 269.400 ;
        RECT 191.200 267.400 192.400 268.000 ;
        RECT 189.800 266.000 190.800 266.800 ;
        RECT 190.000 262.200 190.800 266.000 ;
        RECT 191.600 262.200 192.400 267.400 ;
        RECT 195.400 267.400 196.200 268.600 ;
        RECT 195.400 266.800 197.200 267.400 ;
        RECT 196.400 266.200 197.200 266.800 ;
        RECT 201.200 266.400 202.000 269.200 ;
        RECT 204.400 268.600 207.600 269.400 ;
        RECT 211.400 268.600 213.400 269.400 ;
        RECT 222.000 269.000 222.800 274.600 ;
        RECT 224.200 272.600 225.000 277.600 ;
        RECT 224.200 271.800 226.000 272.600 ;
        RECT 230.000 272.000 230.800 279.800 ;
        RECT 233.200 275.200 234.000 279.800 ;
        RECT 223.600 269.600 224.400 271.200 ;
        RECT 204.000 267.800 204.800 268.000 ;
        RECT 204.000 267.200 208.400 267.800 ;
        RECT 207.600 267.000 208.400 267.200 ;
        RECT 209.200 266.800 210.000 268.400 ;
        RECT 196.400 265.400 198.800 266.200 ;
        RECT 201.200 265.600 202.200 266.400 ;
        RECT 205.200 265.600 206.800 266.400 ;
        RECT 207.600 266.200 208.400 266.400 ;
        RECT 211.400 266.200 212.200 268.600 ;
        RECT 214.000 268.200 222.800 269.000 ;
        RECT 217.400 266.800 220.400 267.600 ;
        RECT 217.400 266.200 218.200 266.800 ;
        RECT 207.600 265.600 212.200 266.200 ;
        RECT 198.000 262.200 198.800 265.400 ;
        RECT 215.600 265.400 218.200 266.200 ;
        RECT 199.600 262.200 200.400 265.000 ;
        RECT 201.200 262.200 202.000 265.000 ;
        RECT 202.800 262.200 203.600 265.000 ;
        RECT 204.400 262.200 205.200 265.000 ;
        RECT 207.600 262.200 208.400 265.000 ;
        RECT 210.800 262.200 211.600 265.000 ;
        RECT 212.400 262.200 213.200 265.000 ;
        RECT 214.000 262.200 214.800 265.000 ;
        RECT 215.600 262.200 216.400 265.400 ;
        RECT 222.000 262.200 222.800 268.200 ;
        RECT 225.200 268.400 225.800 271.800 ;
        RECT 229.800 271.200 230.800 272.000 ;
        RECT 231.400 274.600 234.000 275.200 ;
        RECT 231.400 273.000 232.000 274.600 ;
        RECT 236.400 274.400 237.200 279.800 ;
        RECT 239.600 277.000 240.400 279.800 ;
        RECT 241.200 277.000 242.000 279.800 ;
        RECT 242.800 277.000 243.600 279.800 ;
        RECT 237.800 274.400 242.000 275.200 ;
        RECT 234.600 273.600 237.200 274.400 ;
        RECT 244.400 273.600 245.200 279.800 ;
        RECT 247.600 275.000 248.400 279.800 ;
        RECT 250.800 275.000 251.600 279.800 ;
        RECT 252.400 277.000 253.200 279.800 ;
        RECT 254.000 277.000 254.800 279.800 ;
        RECT 257.200 275.200 258.000 279.800 ;
        RECT 260.400 276.400 261.200 279.800 ;
        RECT 260.400 275.800 261.400 276.400 ;
        RECT 260.800 275.200 261.400 275.800 ;
        RECT 256.000 274.400 260.200 275.200 ;
        RECT 260.800 274.600 262.800 275.200 ;
        RECT 247.600 273.600 250.200 274.400 ;
        RECT 250.800 273.800 256.600 274.400 ;
        RECT 259.600 274.000 260.200 274.400 ;
        RECT 239.600 273.000 240.400 273.200 ;
        RECT 231.400 272.400 240.400 273.000 ;
        RECT 242.800 273.000 243.600 273.200 ;
        RECT 250.800 273.000 251.400 273.800 ;
        RECT 257.200 273.200 258.600 273.800 ;
        RECT 259.600 273.200 261.200 274.000 ;
        RECT 242.800 272.400 251.400 273.000 ;
        RECT 252.400 273.000 258.600 273.200 ;
        RECT 252.400 272.600 257.800 273.000 ;
        RECT 252.400 272.400 253.200 272.600 ;
        RECT 225.200 267.600 226.000 268.400 ;
        RECT 225.200 264.200 225.800 267.600 ;
        RECT 229.800 266.800 230.600 271.200 ;
        RECT 231.400 270.600 232.000 272.400 ;
        RECT 231.200 270.000 232.000 270.600 ;
        RECT 238.000 270.000 261.400 270.600 ;
        RECT 231.200 268.000 231.800 270.000 ;
        RECT 238.000 269.400 238.800 270.000 ;
        RECT 255.600 269.600 256.400 270.000 ;
        RECT 258.800 269.600 259.600 270.000 ;
        RECT 260.600 269.800 261.400 270.000 ;
        RECT 232.400 268.600 236.200 269.400 ;
        RECT 231.200 267.400 232.400 268.000 ;
        RECT 226.800 266.300 227.600 266.400 ;
        RECT 228.400 266.300 229.200 266.400 ;
        RECT 226.800 265.700 229.200 266.300 ;
        RECT 229.800 266.000 230.800 266.800 ;
        RECT 226.800 264.800 227.600 265.700 ;
        RECT 228.400 265.600 229.200 265.700 ;
        RECT 225.200 262.200 226.000 264.200 ;
        RECT 230.000 262.200 230.800 266.000 ;
        RECT 231.600 262.200 232.400 267.400 ;
        RECT 235.400 267.400 236.200 268.600 ;
        RECT 235.400 266.800 237.200 267.400 ;
        RECT 236.400 266.200 237.200 266.800 ;
        RECT 241.200 266.400 242.000 269.200 ;
        RECT 244.400 268.600 247.600 269.400 ;
        RECT 251.400 268.600 253.400 269.400 ;
        RECT 262.000 269.000 262.800 274.600 ;
        RECT 268.400 272.400 269.200 279.800 ;
        RECT 271.600 272.800 272.400 279.800 ;
        RECT 274.800 275.800 275.600 279.800 ;
        RECT 275.000 275.600 275.600 275.800 ;
        RECT 278.000 275.800 278.800 279.800 ;
        RECT 278.000 275.600 278.600 275.800 ;
        RECT 275.000 275.000 278.600 275.600 ;
        RECT 268.400 271.800 271.000 272.400 ;
        RECT 271.600 271.800 272.600 272.800 ;
        RECT 275.000 272.400 275.600 275.000 ;
        RECT 276.400 272.800 277.200 274.400 ;
        RECT 282.000 273.600 282.800 274.400 ;
        RECT 282.000 272.400 282.600 273.600 ;
        RECT 283.400 272.400 284.200 279.800 ;
        RECT 290.200 278.400 291.000 279.800 ;
        RECT 289.200 277.600 291.000 278.400 ;
        RECT 290.200 272.400 291.000 277.600 ;
        RECT 295.600 276.400 296.400 279.800 ;
        RECT 295.400 275.800 296.400 276.400 ;
        RECT 295.400 275.200 296.000 275.800 ;
        RECT 298.800 275.200 299.600 279.800 ;
        RECT 302.000 277.000 302.800 279.800 ;
        RECT 303.600 277.000 304.400 279.800 ;
        RECT 294.000 274.600 296.000 275.200 ;
        RECT 291.600 273.600 292.400 274.400 ;
        RECT 291.800 272.400 292.400 273.600 ;
        RECT 268.400 269.600 269.400 270.400 ;
        RECT 244.000 267.800 244.800 268.000 ;
        RECT 244.000 267.200 248.400 267.800 ;
        RECT 247.600 267.000 248.400 267.200 ;
        RECT 249.200 266.800 250.000 268.400 ;
        RECT 236.400 265.400 238.800 266.200 ;
        RECT 241.200 265.600 242.200 266.400 ;
        RECT 245.200 265.600 246.800 266.400 ;
        RECT 247.600 266.200 248.400 266.400 ;
        RECT 251.400 266.200 252.200 268.600 ;
        RECT 254.000 268.200 262.800 269.000 ;
        RECT 268.600 268.800 269.400 269.600 ;
        RECT 270.400 269.800 271.000 271.800 ;
        RECT 270.400 269.000 271.400 269.800 ;
        RECT 257.400 266.800 260.400 267.600 ;
        RECT 257.400 266.200 258.200 266.800 ;
        RECT 247.600 265.600 252.200 266.200 ;
        RECT 238.000 262.200 238.800 265.400 ;
        RECT 255.600 265.400 258.200 266.200 ;
        RECT 239.600 262.200 240.400 265.000 ;
        RECT 241.200 262.200 242.000 265.000 ;
        RECT 242.800 262.200 243.600 265.000 ;
        RECT 244.400 262.200 245.200 265.000 ;
        RECT 247.600 262.200 248.400 265.000 ;
        RECT 250.800 262.200 251.600 265.000 ;
        RECT 252.400 262.200 253.200 265.000 ;
        RECT 254.000 262.200 254.800 265.000 ;
        RECT 255.600 262.200 256.400 265.400 ;
        RECT 262.000 262.200 262.800 268.200 ;
        RECT 270.400 267.400 271.000 269.000 ;
        RECT 272.000 268.400 272.600 271.800 ;
        RECT 274.800 271.600 275.600 272.400 ;
        RECT 281.200 271.800 282.600 272.400 ;
        RECT 281.200 271.600 282.000 271.800 ;
        RECT 283.200 271.600 285.200 272.400 ;
        RECT 290.200 271.800 291.200 272.400 ;
        RECT 291.800 271.800 293.200 272.400 ;
        RECT 271.600 267.600 272.600 268.400 ;
        RECT 275.000 268.400 275.600 271.600 ;
        RECT 277.200 269.600 278.800 270.400 ;
        RECT 283.200 268.400 283.800 271.600 ;
        RECT 284.400 268.800 285.200 270.400 ;
        RECT 286.000 270.300 286.800 270.400 ;
        RECT 289.200 270.300 290.000 270.400 ;
        RECT 286.000 269.700 290.000 270.300 ;
        RECT 286.000 269.600 286.800 269.700 ;
        RECT 289.200 268.800 290.000 269.700 ;
        RECT 290.600 268.400 291.200 271.800 ;
        RECT 292.400 271.600 293.200 271.800 ;
        RECT 294.000 269.000 294.800 274.600 ;
        RECT 296.600 274.400 300.800 275.200 ;
        RECT 305.200 275.000 306.000 279.800 ;
        RECT 308.400 275.000 309.200 279.800 ;
        RECT 296.600 274.000 297.200 274.400 ;
        RECT 295.600 273.200 297.200 274.000 ;
        RECT 300.200 273.800 306.000 274.400 ;
        RECT 298.200 273.200 299.600 273.800 ;
        RECT 298.200 273.000 304.400 273.200 ;
        RECT 299.000 272.600 304.400 273.000 ;
        RECT 303.600 272.400 304.400 272.600 ;
        RECT 305.400 273.000 306.000 273.800 ;
        RECT 306.600 273.600 309.200 274.400 ;
        RECT 311.600 273.600 312.400 279.800 ;
        RECT 313.200 277.000 314.000 279.800 ;
        RECT 314.800 277.000 315.600 279.800 ;
        RECT 316.400 277.000 317.200 279.800 ;
        RECT 314.800 274.400 319.000 275.200 ;
        RECT 319.600 274.400 320.400 279.800 ;
        RECT 322.800 275.200 323.600 279.800 ;
        RECT 322.800 274.600 325.400 275.200 ;
        RECT 319.600 273.600 322.200 274.400 ;
        RECT 313.200 273.000 314.000 273.200 ;
        RECT 305.400 272.400 314.000 273.000 ;
        RECT 316.400 273.000 317.200 273.200 ;
        RECT 324.800 273.000 325.400 274.600 ;
        RECT 316.400 272.400 325.400 273.000 ;
        RECT 324.800 270.600 325.400 272.400 ;
        RECT 326.000 272.000 326.800 279.800 ;
        RECT 326.000 271.200 327.000 272.000 ;
        RECT 295.400 270.000 318.800 270.600 ;
        RECT 324.800 270.000 325.600 270.600 ;
        RECT 295.400 269.800 296.200 270.000 ;
        RECT 297.200 269.600 298.000 270.000 ;
        RECT 300.400 269.600 301.200 270.000 ;
        RECT 318.000 269.400 318.800 270.000 ;
        RECT 275.000 268.200 276.600 268.400 ;
        RECT 275.000 267.800 276.800 268.200 ;
        RECT 268.400 266.800 271.000 267.400 ;
        RECT 268.400 262.200 269.200 266.800 ;
        RECT 272.000 266.200 272.600 267.600 ;
        RECT 271.600 265.600 272.600 266.200 ;
        RECT 271.600 262.200 272.400 265.600 ;
        RECT 276.000 262.200 276.800 267.800 ;
        RECT 281.200 267.600 283.800 268.400 ;
        RECT 286.000 268.200 286.800 268.400 ;
        RECT 285.200 267.600 286.800 268.200 ;
        RECT 287.600 268.200 288.400 268.400 ;
        RECT 287.600 267.600 289.200 268.200 ;
        RECT 290.600 267.600 293.200 268.400 ;
        RECT 294.000 268.200 302.800 269.000 ;
        RECT 303.400 268.600 305.400 269.400 ;
        RECT 309.200 268.600 312.400 269.400 ;
        RECT 281.400 266.200 282.000 267.600 ;
        RECT 285.200 267.200 286.000 267.600 ;
        RECT 288.400 267.200 289.200 267.600 ;
        RECT 283.000 266.200 286.600 266.600 ;
        RECT 287.800 266.200 291.400 266.600 ;
        RECT 292.400 266.200 293.000 267.600 ;
        RECT 281.200 262.200 282.000 266.200 ;
        RECT 282.800 266.000 286.800 266.200 ;
        RECT 282.800 262.200 283.600 266.000 ;
        RECT 286.000 262.200 286.800 266.000 ;
        RECT 287.600 266.000 291.600 266.200 ;
        RECT 287.600 262.200 288.400 266.000 ;
        RECT 290.800 262.200 291.600 266.000 ;
        RECT 292.400 262.200 293.200 266.200 ;
        RECT 294.000 262.200 294.800 268.200 ;
        RECT 296.400 266.800 299.400 267.600 ;
        RECT 298.600 266.200 299.400 266.800 ;
        RECT 304.600 266.200 305.400 268.600 ;
        RECT 306.800 266.800 307.600 268.400 ;
        RECT 312.000 267.800 312.800 268.000 ;
        RECT 308.400 267.200 312.800 267.800 ;
        RECT 308.400 267.000 309.200 267.200 ;
        RECT 314.800 266.400 315.600 269.200 ;
        RECT 320.600 268.600 324.400 269.400 ;
        RECT 320.600 267.400 321.400 268.600 ;
        RECT 325.000 268.000 325.600 270.000 ;
        RECT 308.400 266.200 309.200 266.400 ;
        RECT 298.600 265.400 301.200 266.200 ;
        RECT 304.600 265.600 309.200 266.200 ;
        RECT 310.000 265.600 311.600 266.400 ;
        RECT 314.600 265.600 315.600 266.400 ;
        RECT 319.600 266.800 321.400 267.400 ;
        RECT 324.400 267.400 325.600 268.000 ;
        RECT 319.600 266.200 320.400 266.800 ;
        RECT 300.400 262.200 301.200 265.400 ;
        RECT 318.000 265.400 320.400 266.200 ;
        RECT 302.000 262.200 302.800 265.000 ;
        RECT 303.600 262.200 304.400 265.000 ;
        RECT 305.200 262.200 306.000 265.000 ;
        RECT 308.400 262.200 309.200 265.000 ;
        RECT 311.600 262.200 312.400 265.000 ;
        RECT 313.200 262.200 314.000 265.000 ;
        RECT 314.800 262.200 315.600 265.000 ;
        RECT 316.400 262.200 317.200 265.000 ;
        RECT 318.000 262.200 318.800 265.400 ;
        RECT 324.400 262.200 325.200 267.400 ;
        RECT 326.200 266.800 327.000 271.200 ;
        RECT 326.000 266.000 327.000 266.800 ;
        RECT 330.800 266.200 331.600 279.800 ;
        RECT 332.400 271.600 333.200 273.200 ;
        RECT 326.000 262.200 326.800 266.000 ;
        RECT 330.800 265.600 332.600 266.200 ;
        RECT 331.800 264.400 332.600 265.600 ;
        RECT 331.800 263.600 333.200 264.400 ;
        RECT 331.800 262.200 332.600 263.600 ;
        RECT 334.000 262.200 334.800 279.800 ;
        RECT 335.600 268.300 336.400 268.400 ;
        RECT 337.200 268.300 338.000 268.400 ;
        RECT 335.600 267.700 338.000 268.300 ;
        RECT 335.600 266.800 336.400 267.700 ;
        RECT 337.200 266.800 338.000 267.700 ;
        RECT 338.800 268.300 339.600 279.800 ;
        RECT 340.400 271.600 341.200 273.200 ;
        RECT 342.000 268.300 342.800 268.400 ;
        RECT 338.800 267.700 342.800 268.300 ;
        RECT 338.800 266.200 339.600 267.700 ;
        RECT 342.000 266.800 342.800 267.700 ;
        RECT 343.600 266.200 344.400 279.800 ;
        RECT 347.600 273.600 348.400 274.400 ;
        RECT 345.200 271.600 346.000 273.200 ;
        RECT 347.600 272.400 348.200 273.600 ;
        RECT 349.000 272.400 349.800 279.800 ;
        RECT 346.800 271.800 348.200 272.400 ;
        RECT 348.800 271.800 349.800 272.400 ;
        RECT 346.800 271.600 347.600 271.800 ;
        RECT 348.800 268.400 349.400 271.800 ;
        RECT 350.000 268.800 350.800 270.400 ;
        RECT 346.800 267.600 349.400 268.400 ;
        RECT 351.600 268.300 352.400 268.400 ;
        RECT 353.200 268.300 354.000 279.800 ;
        RECT 359.000 278.400 359.800 279.800 ;
        RECT 358.000 277.600 359.800 278.400 ;
        RECT 359.000 272.400 359.800 277.600 ;
        RECT 360.400 273.600 361.200 274.400 ;
        RECT 360.600 272.400 361.200 273.600 ;
        RECT 363.600 273.600 364.400 274.400 ;
        RECT 363.600 272.400 364.200 273.600 ;
        RECT 365.000 272.400 365.800 279.800 ;
        RECT 359.000 271.800 360.000 272.400 ;
        RECT 360.600 271.800 362.000 272.400 ;
        RECT 358.000 268.800 358.800 270.400 ;
        RECT 359.400 268.400 360.000 271.800 ;
        RECT 361.200 271.600 362.000 271.800 ;
        RECT 362.800 271.800 364.200 272.400 ;
        RECT 364.800 271.800 365.800 272.400 ;
        RECT 362.800 271.600 363.600 271.800 ;
        RECT 361.200 270.300 362.000 270.400 ;
        RECT 364.800 270.300 365.400 271.800 ;
        RECT 361.200 269.700 365.400 270.300 ;
        RECT 361.200 269.600 362.000 269.700 ;
        RECT 364.800 268.400 365.400 269.700 ;
        RECT 366.000 270.300 366.800 270.400 ;
        RECT 367.600 270.300 368.400 270.400 ;
        RECT 366.000 269.700 368.400 270.300 ;
        RECT 366.000 268.800 366.800 269.700 ;
        RECT 367.600 269.600 368.400 269.700 ;
        RECT 351.600 268.200 354.000 268.300 ;
        RECT 350.800 267.700 354.000 268.200 ;
        RECT 350.800 267.600 352.400 267.700 ;
        RECT 347.000 266.200 347.600 267.600 ;
        RECT 350.800 267.200 351.600 267.600 ;
        RECT 348.600 266.200 352.200 266.600 ;
        RECT 338.800 265.600 340.600 266.200 ;
        RECT 343.600 265.600 345.400 266.200 ;
        RECT 339.800 262.200 340.600 265.600 ;
        RECT 344.600 262.200 345.400 265.600 ;
        RECT 346.800 262.200 347.600 266.200 ;
        RECT 348.400 266.000 352.400 266.200 ;
        RECT 348.400 262.200 349.200 266.000 ;
        RECT 351.600 262.200 352.400 266.000 ;
        RECT 353.200 262.200 354.000 267.700 ;
        RECT 354.800 268.300 355.600 268.400 ;
        RECT 356.400 268.300 357.200 268.400 ;
        RECT 354.800 268.200 357.200 268.300 ;
        RECT 354.800 267.700 358.000 268.200 ;
        RECT 354.800 267.600 355.600 267.700 ;
        RECT 356.400 267.600 358.000 267.700 ;
        RECT 359.400 267.600 362.000 268.400 ;
        RECT 362.800 267.600 365.400 268.400 ;
        RECT 367.600 268.300 368.400 268.400 ;
        RECT 369.200 268.300 370.000 279.800 ;
        RECT 367.600 268.200 370.000 268.300 ;
        RECT 366.800 267.700 370.000 268.200 ;
        RECT 366.800 267.600 368.400 267.700 ;
        RECT 357.200 267.200 358.000 267.600 ;
        RECT 354.800 264.800 355.600 266.400 ;
        RECT 356.600 266.200 360.200 266.600 ;
        RECT 361.200 266.200 361.800 267.600 ;
        RECT 363.000 266.200 363.600 267.600 ;
        RECT 366.800 267.200 367.600 267.600 ;
        RECT 364.600 266.200 368.200 266.600 ;
        RECT 356.400 266.000 360.400 266.200 ;
        RECT 356.400 262.200 357.200 266.000 ;
        RECT 359.600 262.200 360.400 266.000 ;
        RECT 361.200 262.200 362.000 266.200 ;
        RECT 362.800 262.200 363.600 266.200 ;
        RECT 364.400 266.000 368.400 266.200 ;
        RECT 364.400 262.200 365.200 266.000 ;
        RECT 367.600 262.200 368.400 266.000 ;
        RECT 369.200 262.200 370.000 267.700 ;
        RECT 370.800 268.300 371.600 268.400 ;
        RECT 372.400 268.300 373.200 268.400 ;
        RECT 370.800 267.700 373.200 268.300 ;
        RECT 370.800 267.600 371.600 267.700 ;
        RECT 372.400 266.800 373.200 267.700 ;
        RECT 370.800 264.800 371.600 266.400 ;
        RECT 374.000 266.200 374.800 279.800 ;
        RECT 378.800 275.800 379.600 279.800 ;
        RECT 379.000 275.600 379.600 275.800 ;
        RECT 382.000 275.800 382.800 279.800 ;
        RECT 382.000 275.600 382.600 275.800 ;
        RECT 379.000 275.000 382.600 275.600 ;
        RECT 375.600 271.600 376.400 273.200 ;
        RECT 382.000 272.400 382.600 275.000 ;
        RECT 377.200 270.800 378.000 272.400 ;
        RECT 382.000 271.600 382.800 272.400 ;
        RECT 378.800 269.600 380.400 270.400 ;
        RECT 382.000 268.400 382.600 271.600 ;
        RECT 385.200 271.200 386.000 279.800 ;
        RECT 388.400 271.200 389.200 279.800 ;
        RECT 391.600 272.400 392.400 279.800 ;
        RECT 394.800 272.800 395.600 279.800 ;
        RECT 391.600 271.800 394.200 272.400 ;
        RECT 394.800 271.800 395.800 272.800 ;
        RECT 398.000 272.400 398.800 279.800 ;
        RECT 401.200 274.300 402.000 279.800 ;
        RECT 404.400 275.800 405.200 279.800 ;
        RECT 404.600 275.600 405.200 275.800 ;
        RECT 407.600 275.800 408.400 279.800 ;
        RECT 407.600 275.600 408.200 275.800 ;
        RECT 404.600 275.000 408.200 275.600 ;
        RECT 401.200 273.700 403.500 274.300 ;
        RECT 398.000 271.800 400.200 272.400 ;
        RECT 401.200 271.800 402.000 273.700 ;
        RECT 402.900 272.400 403.500 273.700 ;
        RECT 406.000 272.800 406.800 274.400 ;
        RECT 407.600 272.400 408.200 275.000 ;
        RECT 409.200 275.000 410.000 279.000 ;
        RECT 385.200 270.400 389.200 271.200 ;
        RECT 381.000 268.200 382.600 268.400 ;
        RECT 380.800 267.800 382.600 268.200 ;
        RECT 374.000 265.600 375.800 266.200 ;
        RECT 375.000 264.400 375.800 265.600 ;
        RECT 374.000 263.600 375.800 264.400 ;
        RECT 375.000 262.200 375.800 263.600 ;
        RECT 380.800 262.200 381.600 267.800 ;
        RECT 388.400 267.600 389.200 270.400 ;
        RECT 390.000 270.300 390.800 270.400 ;
        RECT 391.600 270.300 392.600 270.400 ;
        RECT 390.000 269.700 392.600 270.300 ;
        RECT 390.000 269.600 390.800 269.700 ;
        RECT 391.600 269.600 392.600 269.700 ;
        RECT 391.800 268.800 392.600 269.600 ;
        RECT 393.600 269.800 394.200 271.800 ;
        RECT 393.600 269.000 394.600 269.800 ;
        RECT 385.200 266.800 389.200 267.600 ;
        RECT 393.600 267.400 394.200 269.000 ;
        RECT 395.200 268.400 395.800 271.800 ;
        RECT 399.600 271.200 400.200 271.800 ;
        RECT 399.600 270.400 400.800 271.200 ;
        RECT 398.000 268.800 398.800 270.400 ;
        RECT 394.800 267.600 395.800 268.400 ;
        RECT 385.200 262.200 386.000 266.800 ;
        RECT 388.400 262.200 389.200 266.800 ;
        RECT 391.600 266.800 394.200 267.400 ;
        RECT 391.600 262.200 392.400 266.800 ;
        RECT 395.200 266.200 395.800 267.600 ;
        RECT 399.600 267.400 400.200 270.400 ;
        RECT 401.400 269.600 402.000 271.800 ;
        RECT 402.800 270.800 403.600 272.400 ;
        RECT 407.600 271.600 408.400 272.400 ;
        RECT 409.200 271.600 409.800 275.000 ;
        RECT 413.400 272.800 414.200 279.800 ;
        RECT 413.400 272.200 415.000 272.800 ;
        RECT 394.800 265.600 395.800 266.200 ;
        RECT 398.000 266.800 400.200 267.400 ;
        RECT 394.800 262.200 395.600 265.600 ;
        RECT 398.000 262.200 398.800 266.800 ;
        RECT 401.200 262.200 402.000 269.600 ;
        RECT 407.600 268.400 408.200 271.600 ;
        RECT 409.200 271.000 413.000 271.600 ;
        RECT 409.200 268.800 410.000 270.400 ;
        RECT 410.800 268.800 411.600 270.400 ;
        RECT 412.400 269.000 413.000 271.000 ;
        RECT 406.600 268.200 408.200 268.400 ;
        RECT 406.400 267.800 408.200 268.200 ;
        RECT 412.400 268.200 413.800 269.000 ;
        RECT 414.400 268.400 415.000 272.200 ;
        RECT 415.600 270.300 416.400 271.200 ;
        RECT 423.600 270.300 424.400 279.800 ;
        RECT 428.400 276.400 429.200 279.800 ;
        RECT 428.200 275.800 429.200 276.400 ;
        RECT 428.200 275.200 428.800 275.800 ;
        RECT 431.600 275.200 432.400 279.800 ;
        RECT 434.800 277.000 435.600 279.800 ;
        RECT 436.400 277.000 437.200 279.800 ;
        RECT 415.600 269.700 424.400 270.300 ;
        RECT 415.600 269.600 416.400 269.700 ;
        RECT 412.400 267.800 413.400 268.200 ;
        RECT 404.400 264.300 405.200 264.400 ;
        RECT 406.400 264.300 407.200 267.800 ;
        RECT 404.400 263.700 407.200 264.300 ;
        RECT 404.400 263.600 405.200 263.700 ;
        RECT 406.400 262.200 407.200 263.700 ;
        RECT 409.200 267.200 413.400 267.800 ;
        RECT 414.400 267.600 416.400 268.400 ;
        RECT 409.200 265.000 409.800 267.200 ;
        RECT 414.400 267.000 415.000 267.600 ;
        RECT 414.200 266.600 415.000 267.000 ;
        RECT 413.400 266.000 415.000 266.600 ;
        RECT 409.200 263.000 410.000 265.000 ;
        RECT 413.400 264.400 414.200 266.000 ;
        RECT 413.400 263.600 414.800 264.400 ;
        RECT 413.400 263.000 414.200 263.600 ;
        RECT 423.600 262.200 424.400 269.700 ;
        RECT 426.800 274.600 428.800 275.200 ;
        RECT 426.800 269.000 427.600 274.600 ;
        RECT 429.400 274.400 433.600 275.200 ;
        RECT 438.000 275.000 438.800 279.800 ;
        RECT 441.200 275.000 442.000 279.800 ;
        RECT 429.400 274.000 430.000 274.400 ;
        RECT 428.400 273.200 430.000 274.000 ;
        RECT 433.000 273.800 438.800 274.400 ;
        RECT 431.000 273.200 432.400 273.800 ;
        RECT 431.000 273.000 437.200 273.200 ;
        RECT 431.800 272.600 437.200 273.000 ;
        RECT 436.400 272.400 437.200 272.600 ;
        RECT 438.200 273.000 438.800 273.800 ;
        RECT 439.400 273.600 442.000 274.400 ;
        RECT 444.400 273.600 445.200 279.800 ;
        RECT 446.000 277.000 446.800 279.800 ;
        RECT 447.600 277.000 448.400 279.800 ;
        RECT 449.200 277.000 450.000 279.800 ;
        RECT 447.600 274.400 451.800 275.200 ;
        RECT 452.400 274.400 453.200 279.800 ;
        RECT 455.600 275.200 456.400 279.800 ;
        RECT 455.600 274.600 458.200 275.200 ;
        RECT 452.400 273.600 455.000 274.400 ;
        RECT 446.000 273.000 446.800 273.200 ;
        RECT 438.200 272.400 446.800 273.000 ;
        RECT 449.200 273.000 450.000 273.200 ;
        RECT 457.600 273.000 458.200 274.600 ;
        RECT 449.200 272.400 458.200 273.000 ;
        RECT 457.600 270.600 458.200 272.400 ;
        RECT 458.800 272.000 459.600 279.800 ;
        RECT 458.800 271.200 459.800 272.000 ;
        RECT 428.200 270.000 451.600 270.600 ;
        RECT 457.600 270.000 458.400 270.600 ;
        RECT 428.200 269.800 429.000 270.000 ;
        RECT 433.200 269.600 434.000 270.000 ;
        RECT 450.800 269.400 451.600 270.000 ;
        RECT 426.800 268.200 435.600 269.000 ;
        RECT 436.200 268.600 438.200 269.400 ;
        RECT 442.000 268.600 445.200 269.400 ;
        RECT 425.200 264.800 426.000 266.400 ;
        RECT 426.800 262.200 427.600 268.200 ;
        RECT 429.200 266.800 432.200 267.600 ;
        RECT 431.400 266.200 432.200 266.800 ;
        RECT 437.400 266.200 438.200 268.600 ;
        RECT 439.600 266.800 440.400 268.400 ;
        RECT 444.800 267.800 445.600 268.000 ;
        RECT 441.200 267.200 445.600 267.800 ;
        RECT 441.200 267.000 442.000 267.200 ;
        RECT 447.600 266.400 448.400 269.200 ;
        RECT 453.400 268.600 457.200 269.400 ;
        RECT 453.400 267.400 454.200 268.600 ;
        RECT 457.800 268.000 458.400 270.000 ;
        RECT 441.200 266.200 442.000 266.400 ;
        RECT 431.400 265.400 434.000 266.200 ;
        RECT 437.400 265.600 442.000 266.200 ;
        RECT 442.800 265.600 444.400 266.400 ;
        RECT 447.400 265.600 448.400 266.400 ;
        RECT 452.400 266.800 454.200 267.400 ;
        RECT 457.200 267.400 458.400 268.000 ;
        RECT 452.400 266.200 453.200 266.800 ;
        RECT 433.200 262.200 434.000 265.400 ;
        RECT 450.800 265.400 453.200 266.200 ;
        RECT 434.800 262.200 435.600 265.000 ;
        RECT 436.400 262.200 437.200 265.000 ;
        RECT 438.000 262.200 438.800 265.000 ;
        RECT 441.200 262.200 442.000 265.000 ;
        RECT 444.400 262.200 445.200 265.000 ;
        RECT 446.000 262.200 446.800 265.000 ;
        RECT 447.600 262.200 448.400 265.000 ;
        RECT 449.200 262.200 450.000 265.000 ;
        RECT 450.800 262.200 451.600 265.400 ;
        RECT 457.200 262.200 458.000 267.400 ;
        RECT 459.000 266.800 459.800 271.200 ;
        RECT 458.800 266.300 459.800 266.800 ;
        RECT 462.000 266.300 462.800 266.400 ;
        RECT 458.800 265.700 462.800 266.300 ;
        RECT 458.800 262.200 459.600 265.700 ;
        RECT 462.000 264.800 462.800 265.700 ;
        RECT 463.600 262.200 464.400 279.800 ;
        RECT 466.800 276.400 467.600 279.800 ;
        RECT 466.600 275.800 467.600 276.400 ;
        RECT 466.600 275.200 467.200 275.800 ;
        RECT 470.000 275.200 470.800 279.800 ;
        RECT 473.200 277.000 474.000 279.800 ;
        RECT 474.800 277.000 475.600 279.800 ;
        RECT 465.200 274.600 467.200 275.200 ;
        RECT 465.200 269.000 466.000 274.600 ;
        RECT 467.800 274.400 472.000 275.200 ;
        RECT 476.400 275.000 477.200 279.800 ;
        RECT 479.600 275.000 480.400 279.800 ;
        RECT 467.800 274.000 468.400 274.400 ;
        RECT 466.800 273.200 468.400 274.000 ;
        RECT 471.400 273.800 477.200 274.400 ;
        RECT 469.400 273.200 470.800 273.800 ;
        RECT 469.400 273.000 475.600 273.200 ;
        RECT 470.200 272.600 475.600 273.000 ;
        RECT 474.800 272.400 475.600 272.600 ;
        RECT 476.600 273.000 477.200 273.800 ;
        RECT 477.800 273.600 480.400 274.400 ;
        RECT 482.800 273.600 483.600 279.800 ;
        RECT 484.400 277.000 485.200 279.800 ;
        RECT 486.000 277.000 486.800 279.800 ;
        RECT 487.600 277.000 488.400 279.800 ;
        RECT 486.000 274.400 490.200 275.200 ;
        RECT 490.800 274.400 491.600 279.800 ;
        RECT 494.000 275.200 494.800 279.800 ;
        RECT 494.000 274.600 496.600 275.200 ;
        RECT 490.800 273.600 493.400 274.400 ;
        RECT 484.400 273.000 485.200 273.200 ;
        RECT 476.600 272.400 485.200 273.000 ;
        RECT 487.600 273.000 488.400 273.200 ;
        RECT 496.000 273.000 496.600 274.600 ;
        RECT 487.600 272.400 496.600 273.000 ;
        RECT 496.000 270.600 496.600 272.400 ;
        RECT 497.200 272.000 498.000 279.800 ;
        RECT 497.200 271.200 498.200 272.000 ;
        RECT 466.600 270.000 490.000 270.600 ;
        RECT 496.000 270.000 496.800 270.600 ;
        RECT 466.600 269.800 467.400 270.000 ;
        RECT 468.400 269.600 469.200 270.000 ;
        RECT 471.600 269.600 472.400 270.000 ;
        RECT 489.200 269.400 490.000 270.000 ;
        RECT 465.200 268.200 474.000 269.000 ;
        RECT 474.600 268.600 476.600 269.400 ;
        RECT 480.400 268.600 483.600 269.400 ;
        RECT 465.200 262.200 466.000 268.200 ;
        RECT 467.600 266.800 470.600 267.600 ;
        RECT 469.800 266.200 470.600 266.800 ;
        RECT 475.800 266.200 476.600 268.600 ;
        RECT 478.000 266.800 478.800 268.400 ;
        RECT 483.200 267.800 484.000 268.000 ;
        RECT 479.600 267.200 484.000 267.800 ;
        RECT 479.600 267.000 480.400 267.200 ;
        RECT 486.000 266.400 486.800 269.200 ;
        RECT 491.800 268.600 495.600 269.400 ;
        RECT 491.800 267.400 492.600 268.600 ;
        RECT 496.200 268.000 496.800 270.000 ;
        RECT 479.600 266.200 480.400 266.400 ;
        RECT 469.800 265.400 472.400 266.200 ;
        RECT 475.800 265.600 480.400 266.200 ;
        RECT 481.200 265.600 482.800 266.400 ;
        RECT 485.800 265.600 486.800 266.400 ;
        RECT 490.800 266.800 492.600 267.400 ;
        RECT 495.600 267.400 496.800 268.000 ;
        RECT 490.800 266.200 491.600 266.800 ;
        RECT 471.600 262.200 472.400 265.400 ;
        RECT 489.200 265.400 491.600 266.200 ;
        RECT 473.200 262.200 474.000 265.000 ;
        RECT 474.800 262.200 475.600 265.000 ;
        RECT 476.400 262.200 477.200 265.000 ;
        RECT 479.600 262.200 480.400 265.000 ;
        RECT 482.800 262.200 483.600 265.000 ;
        RECT 484.400 262.200 485.200 265.000 ;
        RECT 486.000 262.200 486.800 265.000 ;
        RECT 487.600 262.200 488.400 265.000 ;
        RECT 489.200 262.200 490.000 265.400 ;
        RECT 495.600 262.200 496.400 267.400 ;
        RECT 497.400 266.800 498.200 271.200 ;
        RECT 497.200 266.300 498.200 266.800 ;
        RECT 500.400 266.300 501.200 266.400 ;
        RECT 497.200 265.700 501.200 266.300 ;
        RECT 497.200 262.200 498.000 265.700 ;
        RECT 500.400 264.800 501.200 265.700 ;
        RECT 502.000 262.200 502.800 279.800 ;
        RECT 503.600 262.200 504.400 279.800 ;
        RECT 508.400 271.200 509.200 279.800 ;
        RECT 511.600 271.200 512.400 279.800 ;
        RECT 514.800 271.200 515.600 279.800 ;
        RECT 518.000 271.200 518.800 279.800 ;
        RECT 522.000 273.600 522.800 274.400 ;
        RECT 522.000 272.400 522.600 273.600 ;
        RECT 523.400 272.400 524.200 279.800 ;
        RECT 529.200 272.800 530.000 279.800 ;
        RECT 521.200 271.800 522.600 272.400 ;
        RECT 523.200 271.800 524.200 272.400 ;
        RECT 529.000 271.800 530.000 272.800 ;
        RECT 532.400 272.400 533.200 279.800 ;
        RECT 530.600 271.800 533.200 272.400 ;
        RECT 536.600 272.400 537.400 279.800 ;
        RECT 538.000 273.600 538.800 274.400 ;
        RECT 538.200 272.400 538.800 273.600 ;
        RECT 536.600 271.800 537.600 272.400 ;
        RECT 538.200 271.800 539.600 272.400 ;
        RECT 521.200 271.600 522.000 271.800 ;
        RECT 508.400 270.400 510.200 271.200 ;
        RECT 511.600 270.400 513.800 271.200 ;
        RECT 514.800 270.400 517.000 271.200 ;
        RECT 518.000 270.400 520.400 271.200 ;
        RECT 509.400 269.000 510.200 270.400 ;
        RECT 513.000 269.000 513.800 270.400 ;
        RECT 516.200 269.000 517.000 270.400 ;
        RECT 506.800 268.200 508.600 269.000 ;
        RECT 509.400 268.200 512.000 269.000 ;
        RECT 513.000 268.200 515.400 269.000 ;
        RECT 516.200 268.200 518.800 269.000 ;
        RECT 506.800 267.600 507.600 268.200 ;
        RECT 509.400 267.600 510.200 268.200 ;
        RECT 513.000 267.600 513.800 268.200 ;
        RECT 516.200 267.600 517.000 268.200 ;
        RECT 519.600 267.600 520.400 270.400 ;
        RECT 523.200 268.400 523.800 271.800 ;
        RECT 524.400 268.800 525.200 270.400 ;
        RECT 529.000 268.400 529.600 271.800 ;
        RECT 530.600 269.800 531.200 271.800 ;
        RECT 530.200 269.000 531.200 269.800 ;
        RECT 521.200 267.600 523.800 268.400 ;
        RECT 526.000 268.300 526.800 268.400 ;
        RECT 529.000 268.300 530.000 268.400 ;
        RECT 526.000 268.200 530.000 268.300 ;
        RECT 525.200 267.700 530.000 268.200 ;
        RECT 525.200 267.600 526.800 267.700 ;
        RECT 529.000 267.600 530.000 267.700 ;
        RECT 508.400 266.800 510.200 267.600 ;
        RECT 511.600 266.800 513.800 267.600 ;
        RECT 514.800 266.800 517.000 267.600 ;
        RECT 518.000 266.800 520.400 267.600 ;
        RECT 505.200 264.800 506.000 266.400 ;
        RECT 508.400 262.200 509.200 266.800 ;
        RECT 511.600 262.200 512.400 266.800 ;
        RECT 514.800 262.200 515.600 266.800 ;
        RECT 518.000 262.200 518.800 266.800 ;
        RECT 521.400 266.200 522.000 267.600 ;
        RECT 525.200 267.200 526.000 267.600 ;
        RECT 523.000 266.200 526.600 266.600 ;
        RECT 529.000 266.200 529.600 267.600 ;
        RECT 530.600 267.400 531.200 269.000 ;
        RECT 532.200 269.600 533.200 270.400 ;
        RECT 532.200 268.800 533.000 269.600 ;
        RECT 535.600 268.800 536.400 270.400 ;
        RECT 537.000 270.300 537.600 271.800 ;
        RECT 538.800 271.600 539.600 271.800 ;
        RECT 540.400 271.400 541.200 279.800 ;
        RECT 544.800 276.400 545.600 279.800 ;
        RECT 543.600 275.800 545.600 276.400 ;
        RECT 549.200 275.800 550.000 279.800 ;
        RECT 553.400 275.800 554.600 279.800 ;
        RECT 543.600 275.000 544.400 275.800 ;
        RECT 549.200 275.200 549.800 275.800 ;
        RECT 547.000 274.600 550.600 275.200 ;
        RECT 553.200 275.000 554.000 275.800 ;
        RECT 547.000 274.400 547.800 274.600 ;
        RECT 549.800 274.400 550.600 274.600 ;
        RECT 543.600 273.000 544.400 273.200 ;
        RECT 548.200 273.000 549.000 273.200 ;
        RECT 543.600 272.400 549.000 273.000 ;
        RECT 549.600 273.000 551.800 273.600 ;
        RECT 549.600 271.800 550.200 273.000 ;
        RECT 551.000 272.800 551.800 273.000 ;
        RECT 553.400 273.200 554.800 274.000 ;
        RECT 553.400 272.200 554.000 273.200 ;
        RECT 545.400 271.400 550.200 271.800 ;
        RECT 540.400 271.200 550.200 271.400 ;
        RECT 551.600 271.600 554.000 272.200 ;
        RECT 540.400 271.000 546.200 271.200 ;
        RECT 540.400 270.800 546.000 271.000 ;
        RECT 538.800 270.300 539.600 270.400 ;
        RECT 537.000 269.700 539.600 270.300 ;
        RECT 546.800 270.200 547.600 270.400 ;
        RECT 537.000 268.400 537.600 269.700 ;
        RECT 538.800 269.600 539.600 269.700 ;
        RECT 542.600 269.600 547.600 270.200 ;
        RECT 542.600 269.400 543.400 269.600 ;
        RECT 545.200 269.400 546.000 269.600 ;
        RECT 544.200 268.400 545.000 268.600 ;
        RECT 551.600 268.400 552.200 271.600 ;
        RECT 558.000 271.200 558.800 279.800 ;
        RECT 559.600 271.600 560.400 273.200 ;
        RECT 554.600 270.600 558.800 271.200 ;
        RECT 554.600 270.400 555.400 270.600 ;
        RECT 556.200 269.800 557.000 270.000 ;
        RECT 553.200 269.200 557.000 269.800 ;
        RECT 553.200 269.000 554.000 269.200 ;
        RECT 534.000 268.200 534.800 268.400 ;
        RECT 534.000 267.600 535.600 268.200 ;
        RECT 537.000 267.600 539.600 268.400 ;
        RECT 541.200 267.800 552.200 268.400 ;
        RECT 541.200 267.600 542.800 267.800 ;
        RECT 530.600 266.800 533.200 267.400 ;
        RECT 534.800 267.200 535.600 267.600 ;
        RECT 521.200 262.200 522.000 266.200 ;
        RECT 522.800 266.000 526.800 266.200 ;
        RECT 522.800 262.200 523.600 266.000 ;
        RECT 526.000 262.200 526.800 266.000 ;
        RECT 529.000 265.600 530.000 266.200 ;
        RECT 529.200 262.200 530.000 265.600 ;
        RECT 532.400 262.200 533.200 266.800 ;
        RECT 534.200 266.200 537.800 266.600 ;
        RECT 538.800 266.200 539.400 267.600 ;
        RECT 534.000 266.000 538.000 266.200 ;
        RECT 534.000 262.200 534.800 266.000 ;
        RECT 537.200 262.200 538.000 266.000 ;
        RECT 538.800 262.200 539.600 266.200 ;
        RECT 540.400 262.200 541.200 267.000 ;
        RECT 545.400 265.600 546.000 267.800 ;
        RECT 551.000 267.600 551.800 267.800 ;
        RECT 558.000 267.200 558.800 270.600 ;
        RECT 555.000 266.600 558.800 267.200 ;
        RECT 555.000 266.400 555.800 266.600 ;
        RECT 543.600 264.200 544.400 265.000 ;
        RECT 545.200 264.800 546.000 265.600 ;
        RECT 547.000 265.400 547.800 265.600 ;
        RECT 547.000 264.800 549.800 265.400 ;
        RECT 549.200 264.200 549.800 264.800 ;
        RECT 553.200 264.200 554.000 265.000 ;
        RECT 543.600 263.600 545.600 264.200 ;
        RECT 544.800 262.200 545.600 263.600 ;
        RECT 549.200 262.200 550.000 264.200 ;
        RECT 553.200 263.600 554.600 264.200 ;
        RECT 553.400 262.200 554.600 263.600 ;
        RECT 558.000 262.200 558.800 266.600 ;
        RECT 561.200 266.200 562.000 279.800 ;
        RECT 568.200 272.800 569.000 279.800 ;
        RECT 572.400 275.000 573.200 279.000 ;
        RECT 567.400 272.200 569.000 272.800 ;
        RECT 562.800 270.300 563.600 270.400 ;
        RECT 566.000 270.300 566.800 271.200 ;
        RECT 562.800 269.700 566.800 270.300 ;
        RECT 562.800 269.600 563.600 269.700 ;
        RECT 566.000 269.600 566.800 269.700 ;
        RECT 567.400 268.400 568.000 272.200 ;
        RECT 572.600 271.600 573.200 275.000 ;
        RECT 582.600 276.400 583.400 279.800 ;
        RECT 582.600 275.600 584.400 276.400 ;
        RECT 582.600 272.800 583.400 275.600 ;
        RECT 586.800 275.000 587.600 279.000 ;
        RECT 569.400 271.000 573.200 271.600 ;
        RECT 581.800 272.200 583.400 272.800 ;
        RECT 569.400 269.000 570.000 271.000 ;
        RECT 562.800 266.800 563.600 268.400 ;
        RECT 566.000 267.600 568.000 268.400 ;
        RECT 568.600 268.200 570.000 269.000 ;
        RECT 570.800 268.800 571.600 270.400 ;
        RECT 572.400 268.800 573.200 270.400 ;
        RECT 580.400 269.600 581.200 271.200 ;
        RECT 581.800 268.400 582.400 272.200 ;
        RECT 587.000 271.600 587.600 275.000 ;
        RECT 589.200 273.600 590.000 274.400 ;
        RECT 589.200 272.400 589.800 273.600 ;
        RECT 590.600 272.400 591.400 279.800 ;
        RECT 595.600 273.600 596.400 274.400 ;
        RECT 595.600 272.400 596.200 273.600 ;
        RECT 597.000 272.400 597.800 279.800 ;
        RECT 588.400 271.800 589.800 272.400 ;
        RECT 588.400 271.600 589.200 271.800 ;
        RECT 590.400 271.600 592.400 272.400 ;
        RECT 594.800 271.800 596.200 272.400 ;
        RECT 596.800 271.800 597.800 272.400 ;
        RECT 601.200 272.400 602.000 279.800 ;
        RECT 604.400 272.800 605.200 279.800 ;
        RECT 601.200 271.800 603.800 272.400 ;
        RECT 604.400 271.800 605.400 272.800 ;
        RECT 610.200 272.400 611.000 279.800 ;
        RECT 611.600 273.600 612.400 274.400 ;
        RECT 611.800 272.400 612.400 273.600 ;
        RECT 614.800 273.600 615.600 274.400 ;
        RECT 614.800 272.400 615.400 273.600 ;
        RECT 616.200 272.400 617.000 279.800 ;
        RECT 610.200 271.800 611.200 272.400 ;
        RECT 611.800 271.800 613.200 272.400 ;
        RECT 594.800 271.600 595.600 271.800 ;
        RECT 583.800 271.000 587.600 271.600 ;
        RECT 583.800 269.000 584.400 271.000 ;
        RECT 567.400 267.000 568.000 267.600 ;
        RECT 569.000 267.800 570.000 268.200 ;
        RECT 569.000 267.200 573.200 267.800 ;
        RECT 580.400 267.600 582.400 268.400 ;
        RECT 583.000 268.200 584.400 269.000 ;
        RECT 585.200 268.800 586.000 270.400 ;
        RECT 586.800 268.800 587.600 270.400 ;
        RECT 590.400 268.400 591.000 271.600 ;
        RECT 591.600 270.300 592.400 270.400 ;
        RECT 594.800 270.300 595.600 270.400 ;
        RECT 591.600 269.700 595.600 270.300 ;
        RECT 591.600 268.800 592.400 269.700 ;
        RECT 594.800 269.600 595.600 269.700 ;
        RECT 596.800 268.400 597.400 271.800 ;
        RECT 598.000 268.800 598.800 270.400 ;
        RECT 599.600 270.300 600.400 270.400 ;
        RECT 601.200 270.300 602.200 270.400 ;
        RECT 599.600 269.700 602.200 270.300 ;
        RECT 599.600 269.600 600.400 269.700 ;
        RECT 601.200 269.600 602.200 269.700 ;
        RECT 601.400 268.800 602.200 269.600 ;
        RECT 603.200 269.800 603.800 271.800 ;
        RECT 603.200 269.000 604.200 269.800 ;
        RECT 560.200 265.600 562.000 266.200 ;
        RECT 567.400 266.600 568.200 267.000 ;
        RECT 567.400 266.000 569.000 266.600 ;
        RECT 560.200 262.200 561.000 265.600 ;
        RECT 568.200 264.400 569.000 266.000 ;
        RECT 572.600 265.000 573.200 267.200 ;
        RECT 581.800 267.000 582.400 267.600 ;
        RECT 583.400 267.800 584.400 268.200 ;
        RECT 583.400 267.200 587.600 267.800 ;
        RECT 588.400 267.600 591.000 268.400 ;
        RECT 593.200 268.200 594.000 268.400 ;
        RECT 592.400 267.600 594.000 268.200 ;
        RECT 594.800 267.600 597.400 268.400 ;
        RECT 599.600 268.200 600.400 268.400 ;
        RECT 598.800 267.600 600.400 268.200 ;
        RECT 581.800 266.600 582.600 267.000 ;
        RECT 581.800 266.000 583.400 266.600 ;
        RECT 567.600 263.600 569.000 264.400 ;
        RECT 568.200 263.000 569.000 263.600 ;
        RECT 572.400 263.000 573.200 265.000 ;
        RECT 582.600 263.000 583.400 266.000 ;
        RECT 587.000 265.000 587.600 267.200 ;
        RECT 588.600 266.200 589.200 267.600 ;
        RECT 592.400 267.200 593.200 267.600 ;
        RECT 590.200 266.200 593.800 266.600 ;
        RECT 595.000 266.200 595.600 267.600 ;
        RECT 598.800 267.200 599.600 267.600 ;
        RECT 603.200 267.400 603.800 269.000 ;
        RECT 604.800 268.400 605.400 271.800 ;
        RECT 609.200 268.800 610.000 270.400 ;
        RECT 610.600 270.300 611.200 271.800 ;
        RECT 612.400 271.600 613.200 271.800 ;
        RECT 614.000 271.800 615.400 272.400 ;
        RECT 616.000 271.800 617.000 272.400 ;
        RECT 614.000 271.600 614.800 271.800 ;
        RECT 614.100 270.300 614.700 271.600 ;
        RECT 610.600 269.700 614.700 270.300 ;
        RECT 610.600 268.400 611.200 269.700 ;
        RECT 616.000 268.400 616.600 271.800 ;
        RECT 617.200 268.800 618.000 270.400 ;
        RECT 604.400 267.600 605.400 268.400 ;
        RECT 607.600 268.200 608.400 268.400 ;
        RECT 607.600 267.600 609.200 268.200 ;
        RECT 610.600 267.600 613.200 268.400 ;
        RECT 614.000 267.600 616.600 268.400 ;
        RECT 618.800 268.200 619.600 268.400 ;
        RECT 618.000 267.600 619.600 268.200 ;
        RECT 601.200 266.800 603.800 267.400 ;
        RECT 596.600 266.200 600.200 266.600 ;
        RECT 586.800 263.000 587.600 265.000 ;
        RECT 588.400 262.200 589.200 266.200 ;
        RECT 590.000 266.000 594.000 266.200 ;
        RECT 590.000 262.200 590.800 266.000 ;
        RECT 593.200 262.200 594.000 266.000 ;
        RECT 594.800 262.200 595.600 266.200 ;
        RECT 596.400 266.000 600.400 266.200 ;
        RECT 596.400 262.200 597.200 266.000 ;
        RECT 599.600 262.200 600.400 266.000 ;
        RECT 601.200 262.200 602.000 266.800 ;
        RECT 604.800 266.200 605.400 267.600 ;
        RECT 608.400 267.200 609.200 267.600 ;
        RECT 607.800 266.200 611.400 266.600 ;
        RECT 612.400 266.200 613.000 267.600 ;
        RECT 614.200 266.200 614.800 267.600 ;
        RECT 618.000 267.200 618.800 267.600 ;
        RECT 615.800 266.200 619.400 266.600 ;
        RECT 604.400 265.600 605.400 266.200 ;
        RECT 607.600 266.000 611.600 266.200 ;
        RECT 604.400 262.200 605.200 265.600 ;
        RECT 607.600 262.200 608.400 266.000 ;
        RECT 610.800 262.200 611.600 266.000 ;
        RECT 612.400 262.200 613.200 266.200 ;
        RECT 614.000 262.200 614.800 266.200 ;
        RECT 615.600 266.000 619.600 266.200 ;
        RECT 615.600 262.200 616.400 266.000 ;
        RECT 618.800 262.200 619.600 266.000 ;
        RECT 620.400 262.200 621.200 279.800 ;
        RECT 623.600 271.600 624.400 273.200 ;
        RECT 622.000 264.800 622.800 266.400 ;
        RECT 625.200 266.200 626.000 279.800 ;
        RECT 628.400 275.000 629.200 279.000 ;
        RECT 628.400 271.600 629.000 275.000 ;
        RECT 632.600 272.800 633.400 279.800 ;
        RECT 632.600 272.200 634.200 272.800 ;
        RECT 628.400 271.000 632.200 271.600 ;
        RECT 628.400 268.800 629.200 270.400 ;
        RECT 630.000 268.800 630.800 270.400 ;
        RECT 631.600 269.000 632.200 271.000 ;
        RECT 626.800 266.800 627.600 268.400 ;
        RECT 631.600 268.200 633.000 269.000 ;
        RECT 633.600 268.400 634.200 272.200 ;
        RECT 640.600 272.400 641.400 279.800 ;
        RECT 647.000 274.400 647.800 279.800 ;
        RECT 642.000 273.600 642.800 274.400 ;
        RECT 646.000 273.600 647.800 274.400 ;
        RECT 648.400 273.600 649.200 274.400 ;
        RECT 642.200 272.400 642.800 273.600 ;
        RECT 647.000 272.400 647.800 273.600 ;
        RECT 648.600 272.400 649.200 273.600 ;
        RECT 654.600 272.800 655.400 279.800 ;
        RECT 658.800 275.000 659.600 279.000 ;
        RECT 640.600 271.800 641.600 272.400 ;
        RECT 642.200 271.800 643.600 272.400 ;
        RECT 647.000 271.800 648.000 272.400 ;
        RECT 648.600 271.800 650.000 272.400 ;
        RECT 634.800 269.600 635.600 271.200 ;
        RECT 639.600 268.800 640.400 270.400 ;
        RECT 641.000 268.400 641.600 271.800 ;
        RECT 642.800 271.600 643.600 271.800 ;
        RECT 646.000 268.800 646.800 270.400 ;
        RECT 647.400 268.400 648.000 271.800 ;
        RECT 649.200 271.600 650.000 271.800 ;
        RECT 653.800 272.200 655.400 272.800 ;
        RECT 653.800 271.600 654.800 272.200 ;
        RECT 659.000 271.600 659.600 275.000 ;
        RECT 662.600 274.400 663.400 279.800 ;
        RECT 661.200 273.600 662.000 274.400 ;
        RECT 662.600 273.600 664.400 274.400 ;
        RECT 661.200 272.400 661.800 273.600 ;
        RECT 662.600 272.400 663.400 273.600 ;
        RECT 660.400 271.800 661.800 272.400 ;
        RECT 662.400 271.800 663.400 272.400 ;
        RECT 660.400 271.600 661.200 271.800 ;
        RECT 652.400 269.600 653.200 271.200 ;
        RECT 653.800 268.400 654.400 271.600 ;
        RECT 655.800 271.000 659.600 271.600 ;
        RECT 655.800 269.000 656.400 271.000 ;
        RECT 631.600 267.800 632.600 268.200 ;
        RECT 628.400 267.200 632.600 267.800 ;
        RECT 633.600 267.600 635.600 268.400 ;
        RECT 636.400 268.300 637.200 268.400 ;
        RECT 638.000 268.300 638.800 268.400 ;
        RECT 636.400 268.200 638.800 268.300 ;
        RECT 636.400 267.700 639.600 268.200 ;
        RECT 636.400 267.600 637.200 267.700 ;
        RECT 638.000 267.600 639.600 267.700 ;
        RECT 641.000 267.600 643.600 268.400 ;
        RECT 644.400 268.200 645.200 268.400 ;
        RECT 644.400 267.600 646.000 268.200 ;
        RECT 647.400 267.600 650.000 268.400 ;
        RECT 652.400 267.600 654.400 268.400 ;
        RECT 655.000 268.200 656.400 269.000 ;
        RECT 657.200 268.800 658.000 270.400 ;
        RECT 658.800 268.800 659.600 270.400 ;
        RECT 662.400 268.400 663.000 271.800 ;
        RECT 666.800 271.200 667.600 279.800 ;
        RECT 671.000 275.800 672.200 279.800 ;
        RECT 675.600 275.800 676.400 279.800 ;
        RECT 680.000 276.400 680.800 279.800 ;
        RECT 680.000 275.800 682.000 276.400 ;
        RECT 671.600 275.000 672.400 275.800 ;
        RECT 675.800 275.200 676.400 275.800 ;
        RECT 675.000 274.600 678.600 275.200 ;
        RECT 681.200 275.000 682.000 275.800 ;
        RECT 675.000 274.400 675.800 274.600 ;
        RECT 677.800 274.400 678.600 274.600 ;
        RECT 670.800 273.200 672.200 274.000 ;
        RECT 671.600 272.200 672.200 273.200 ;
        RECT 673.800 273.000 676.000 273.600 ;
        RECT 673.800 272.800 674.600 273.000 ;
        RECT 671.600 271.600 674.000 272.200 ;
        RECT 666.800 270.600 671.000 271.200 ;
        RECT 663.600 268.800 664.400 270.400 ;
        RECT 624.200 265.600 626.000 266.200 ;
        RECT 624.200 262.200 625.000 265.600 ;
        RECT 628.400 265.000 629.000 267.200 ;
        RECT 633.600 267.000 634.200 267.600 ;
        RECT 638.800 267.200 639.600 267.600 ;
        RECT 633.400 266.600 634.200 267.000 ;
        RECT 632.600 266.000 634.200 266.600 ;
        RECT 638.200 266.200 641.800 266.600 ;
        RECT 642.800 266.200 643.400 267.600 ;
        RECT 645.200 267.200 646.000 267.600 ;
        RECT 644.600 266.200 648.200 266.600 ;
        RECT 649.200 266.200 649.800 267.600 ;
        RECT 653.800 267.000 654.400 267.600 ;
        RECT 655.400 267.800 656.400 268.200 ;
        RECT 655.400 267.200 659.600 267.800 ;
        RECT 660.400 267.600 663.000 268.400 ;
        RECT 665.200 268.200 666.000 268.400 ;
        RECT 664.400 267.600 666.000 268.200 ;
        RECT 653.800 266.600 654.600 267.000 ;
        RECT 638.000 266.000 642.000 266.200 ;
        RECT 628.400 263.000 629.200 265.000 ;
        RECT 632.600 264.400 633.400 266.000 ;
        RECT 631.600 263.600 633.400 264.400 ;
        RECT 632.600 263.000 633.400 263.600 ;
        RECT 638.000 262.200 638.800 266.000 ;
        RECT 641.200 262.200 642.000 266.000 ;
        RECT 642.800 262.200 643.600 266.200 ;
        RECT 644.400 266.000 648.400 266.200 ;
        RECT 644.400 262.200 645.200 266.000 ;
        RECT 647.600 262.200 648.400 266.000 ;
        RECT 649.200 262.200 650.000 266.200 ;
        RECT 653.800 266.000 655.400 266.600 ;
        RECT 654.600 263.000 655.400 266.000 ;
        RECT 659.000 265.000 659.600 267.200 ;
        RECT 660.600 266.200 661.200 267.600 ;
        RECT 664.400 267.200 665.200 267.600 ;
        RECT 666.800 267.200 667.600 270.600 ;
        RECT 670.200 270.400 671.000 270.600 ;
        RECT 673.400 270.400 674.000 271.600 ;
        RECT 675.400 271.800 676.000 273.000 ;
        RECT 676.600 273.000 677.400 273.200 ;
        RECT 681.200 273.000 682.000 273.200 ;
        RECT 676.600 272.400 682.000 273.000 ;
        RECT 675.400 271.400 680.200 271.800 ;
        RECT 684.400 271.400 685.200 279.800 ;
        RECT 675.400 271.200 685.200 271.400 ;
        RECT 679.400 271.000 685.200 271.200 ;
        RECT 679.600 270.800 685.200 271.000 ;
        RECT 668.600 269.800 669.400 270.000 ;
        RECT 668.600 269.200 672.400 269.800 ;
        RECT 673.200 269.600 674.000 270.400 ;
        RECT 676.400 270.300 677.200 270.400 ;
        RECT 678.000 270.300 678.800 270.400 ;
        RECT 676.400 270.200 678.800 270.300 ;
        RECT 676.400 269.700 683.000 270.200 ;
        RECT 676.400 269.600 677.200 269.700 ;
        RECT 678.000 269.600 683.000 269.700 ;
        RECT 671.600 269.000 672.400 269.200 ;
        RECT 673.400 268.400 674.000 269.600 ;
        RECT 682.200 269.400 683.000 269.600 ;
        RECT 680.600 268.400 681.400 268.600 ;
        RECT 673.400 267.800 684.400 268.400 ;
        RECT 673.800 267.600 674.600 267.800 ;
        RECT 666.800 266.600 670.600 267.200 ;
        RECT 662.200 266.200 665.800 266.600 ;
        RECT 658.800 263.000 659.600 265.000 ;
        RECT 660.400 262.200 661.200 266.200 ;
        RECT 662.000 266.000 666.000 266.200 ;
        RECT 662.000 262.200 662.800 266.000 ;
        RECT 665.200 262.200 666.000 266.000 ;
        RECT 666.800 262.200 667.600 266.600 ;
        RECT 669.800 266.400 670.600 266.600 ;
        RECT 679.600 265.600 680.200 267.800 ;
        RECT 682.800 267.600 684.400 267.800 ;
        RECT 677.800 265.400 678.600 265.600 ;
        RECT 671.600 264.200 672.400 265.000 ;
        RECT 675.800 264.800 678.600 265.400 ;
        RECT 679.600 264.800 680.400 265.600 ;
        RECT 675.800 264.200 676.400 264.800 ;
        RECT 681.200 264.200 682.000 265.000 ;
        RECT 671.000 263.600 672.400 264.200 ;
        RECT 671.000 262.200 672.200 263.600 ;
        RECT 675.600 262.200 676.400 264.200 ;
        RECT 680.000 263.600 682.000 264.200 ;
        RECT 680.000 262.200 680.800 263.600 ;
        RECT 684.400 262.200 685.200 267.000 ;
        RECT 4.400 255.200 5.200 259.800 ;
        RECT 9.200 255.200 10.000 259.800 ;
        RECT 10.800 255.600 11.600 257.200 ;
        RECT 3.000 254.600 5.200 255.200 ;
        RECT 7.800 254.600 10.000 255.200 ;
        RECT 3.000 251.600 3.600 254.600 ;
        RECT 4.400 251.600 5.200 253.200 ;
        RECT 7.800 251.600 8.400 254.600 ;
        RECT 9.200 252.300 10.000 253.200 ;
        RECT 10.800 252.300 11.600 252.400 ;
        RECT 9.200 251.700 11.600 252.300 ;
        RECT 9.200 251.600 10.000 251.700 ;
        RECT 10.800 251.600 11.600 251.700 ;
        RECT 2.400 250.800 3.600 251.600 ;
        RECT 7.200 250.800 8.400 251.600 ;
        RECT 3.000 250.200 3.600 250.800 ;
        RECT 7.800 250.200 8.400 250.800 ;
        RECT 3.000 249.600 5.200 250.200 ;
        RECT 7.800 249.600 10.000 250.200 ;
        RECT 4.400 242.200 5.200 249.600 ;
        RECT 9.200 242.200 10.000 249.600 ;
        RECT 12.400 242.200 13.200 259.800 ;
        RECT 14.000 256.300 14.800 256.400 ;
        RECT 15.600 256.300 16.400 259.800 ;
        RECT 14.000 255.700 16.400 256.300 ;
        RECT 14.000 255.600 14.800 255.700 ;
        RECT 15.400 255.200 16.400 255.700 ;
        RECT 15.400 250.800 16.200 255.200 ;
        RECT 17.200 254.600 18.000 259.800 ;
        RECT 23.600 256.600 24.400 259.800 ;
        RECT 25.200 257.000 26.000 259.800 ;
        RECT 26.800 257.000 27.600 259.800 ;
        RECT 28.400 257.000 29.200 259.800 ;
        RECT 30.000 257.000 30.800 259.800 ;
        RECT 33.200 257.000 34.000 259.800 ;
        RECT 36.400 257.000 37.200 259.800 ;
        RECT 38.000 257.000 38.800 259.800 ;
        RECT 39.600 257.000 40.400 259.800 ;
        RECT 22.000 255.800 24.400 256.600 ;
        RECT 41.200 256.600 42.000 259.800 ;
        RECT 22.000 255.200 22.800 255.800 ;
        RECT 16.800 254.000 18.000 254.600 ;
        RECT 21.000 254.600 22.800 255.200 ;
        RECT 26.800 255.600 27.800 256.400 ;
        RECT 30.800 255.600 32.400 256.400 ;
        RECT 33.200 255.800 37.800 256.400 ;
        RECT 41.200 255.800 43.800 256.600 ;
        RECT 33.200 255.600 34.000 255.800 ;
        RECT 16.800 252.000 17.400 254.000 ;
        RECT 21.000 253.400 21.800 254.600 ;
        RECT 18.000 252.600 21.800 253.400 ;
        RECT 26.800 252.800 27.600 255.600 ;
        RECT 33.200 254.800 34.000 255.000 ;
        RECT 29.600 254.200 34.000 254.800 ;
        RECT 29.600 254.000 30.400 254.200 ;
        RECT 34.800 253.600 35.600 255.200 ;
        RECT 37.000 253.400 37.800 255.800 ;
        RECT 43.000 255.200 43.800 255.800 ;
        RECT 43.000 254.400 46.000 255.200 ;
        RECT 47.600 253.800 48.400 259.800 ;
        RECT 50.800 256.000 51.600 259.800 ;
        RECT 30.000 252.600 33.200 253.400 ;
        RECT 37.000 252.600 39.000 253.400 ;
        RECT 39.600 253.000 48.400 253.800 ;
        RECT 23.600 252.000 24.400 252.600 ;
        RECT 41.200 252.000 42.000 252.400 ;
        RECT 44.400 252.000 45.200 252.400 ;
        RECT 46.200 252.000 47.000 252.200 ;
        RECT 16.800 251.400 17.600 252.000 ;
        RECT 23.600 251.400 47.000 252.000 ;
        RECT 15.400 250.000 16.400 250.800 ;
        RECT 15.600 242.200 16.400 250.000 ;
        RECT 17.000 249.600 17.600 251.400 ;
        RECT 17.000 249.000 26.000 249.600 ;
        RECT 17.000 247.400 17.600 249.000 ;
        RECT 25.200 248.800 26.000 249.000 ;
        RECT 28.400 249.000 37.000 249.600 ;
        RECT 28.400 248.800 29.200 249.000 ;
        RECT 20.200 247.600 22.800 248.400 ;
        RECT 17.000 246.800 19.600 247.400 ;
        RECT 18.800 242.200 19.600 246.800 ;
        RECT 22.000 242.200 22.800 247.600 ;
        RECT 23.400 246.800 27.600 247.600 ;
        RECT 25.200 242.200 26.000 245.000 ;
        RECT 26.800 242.200 27.600 245.000 ;
        RECT 28.400 242.200 29.200 245.000 ;
        RECT 30.000 242.200 30.800 248.400 ;
        RECT 33.200 247.600 35.800 248.400 ;
        RECT 36.400 248.200 37.000 249.000 ;
        RECT 38.000 249.400 38.800 249.600 ;
        RECT 38.000 249.000 43.400 249.400 ;
        RECT 38.000 248.800 44.200 249.000 ;
        RECT 42.800 248.200 44.200 248.800 ;
        RECT 36.400 247.600 42.200 248.200 ;
        RECT 45.200 248.000 46.800 248.800 ;
        RECT 45.200 247.600 45.800 248.000 ;
        RECT 33.200 242.200 34.000 247.000 ;
        RECT 36.400 242.200 37.200 247.000 ;
        RECT 41.600 246.800 45.800 247.600 ;
        RECT 47.600 247.400 48.400 253.000 ;
        RECT 50.600 255.200 51.600 256.000 ;
        RECT 50.600 250.800 51.400 255.200 ;
        RECT 52.400 254.600 53.200 259.800 ;
        RECT 58.800 256.600 59.600 259.800 ;
        RECT 60.400 257.000 61.200 259.800 ;
        RECT 62.000 257.000 62.800 259.800 ;
        RECT 63.600 257.000 64.400 259.800 ;
        RECT 65.200 257.000 66.000 259.800 ;
        RECT 68.400 257.000 69.200 259.800 ;
        RECT 71.600 257.000 72.400 259.800 ;
        RECT 73.200 257.000 74.000 259.800 ;
        RECT 74.800 257.000 75.600 259.800 ;
        RECT 57.200 255.800 59.600 256.600 ;
        RECT 76.400 256.600 77.200 259.800 ;
        RECT 57.200 255.200 58.000 255.800 ;
        RECT 52.000 254.000 53.200 254.600 ;
        RECT 56.200 254.600 58.000 255.200 ;
        RECT 62.000 255.600 63.000 256.400 ;
        RECT 66.000 255.600 67.600 256.400 ;
        RECT 68.400 255.800 73.000 256.400 ;
        RECT 76.400 255.800 79.000 256.600 ;
        RECT 68.400 255.600 69.200 255.800 ;
        RECT 52.000 252.000 52.600 254.000 ;
        RECT 56.200 253.400 57.000 254.600 ;
        RECT 53.200 252.600 57.000 253.400 ;
        RECT 62.000 252.800 62.800 255.600 ;
        RECT 68.400 254.800 69.200 255.000 ;
        RECT 64.800 254.200 69.200 254.800 ;
        RECT 64.800 254.000 65.600 254.200 ;
        RECT 70.000 253.600 70.800 255.200 ;
        RECT 72.200 253.400 73.000 255.800 ;
        RECT 78.200 255.200 79.000 255.800 ;
        RECT 78.200 254.400 81.200 255.200 ;
        RECT 82.800 253.800 83.600 259.800 ;
        RECT 65.200 252.600 68.400 253.400 ;
        RECT 72.200 252.600 74.200 253.400 ;
        RECT 74.800 253.000 83.600 253.800 ;
        RECT 58.800 252.000 59.600 252.600 ;
        RECT 76.400 252.000 77.200 252.400 ;
        RECT 81.400 252.000 82.200 252.200 ;
        RECT 52.000 251.400 52.800 252.000 ;
        RECT 58.800 251.400 82.200 252.000 ;
        RECT 50.600 250.000 51.600 250.800 ;
        RECT 46.400 246.800 48.400 247.400 ;
        RECT 38.000 242.200 38.800 245.000 ;
        RECT 39.600 242.200 40.400 245.000 ;
        RECT 42.800 242.200 43.600 246.800 ;
        RECT 46.400 246.200 47.000 246.800 ;
        RECT 46.000 245.600 47.000 246.200 ;
        RECT 46.000 242.200 46.800 245.600 ;
        RECT 50.800 242.200 51.600 250.000 ;
        RECT 52.200 249.600 52.800 251.400 ;
        RECT 52.200 249.000 61.200 249.600 ;
        RECT 52.200 247.400 52.800 249.000 ;
        RECT 60.400 248.800 61.200 249.000 ;
        RECT 63.600 249.000 72.200 249.600 ;
        RECT 63.600 248.800 64.400 249.000 ;
        RECT 55.400 247.600 58.000 248.400 ;
        RECT 52.200 246.800 54.800 247.400 ;
        RECT 54.000 242.200 54.800 246.800 ;
        RECT 57.200 242.200 58.000 247.600 ;
        RECT 58.600 246.800 62.800 247.600 ;
        RECT 60.400 242.200 61.200 245.000 ;
        RECT 62.000 242.200 62.800 245.000 ;
        RECT 63.600 242.200 64.400 245.000 ;
        RECT 65.200 242.200 66.000 248.400 ;
        RECT 68.400 247.600 71.000 248.400 ;
        RECT 71.600 248.200 72.200 249.000 ;
        RECT 73.200 249.400 74.000 249.600 ;
        RECT 73.200 249.000 78.600 249.400 ;
        RECT 73.200 248.800 79.400 249.000 ;
        RECT 78.000 248.200 79.400 248.800 ;
        RECT 71.600 247.600 77.400 248.200 ;
        RECT 80.400 248.000 82.000 248.800 ;
        RECT 80.400 247.600 81.000 248.000 ;
        RECT 68.400 242.200 69.200 247.000 ;
        RECT 71.600 242.200 72.400 247.000 ;
        RECT 76.800 246.800 81.000 247.600 ;
        RECT 82.800 247.400 83.600 253.000 ;
        RECT 81.600 246.800 83.600 247.400 ;
        RECT 73.200 242.200 74.000 245.000 ;
        RECT 74.800 242.200 75.600 245.000 ;
        RECT 78.000 242.200 78.800 246.800 ;
        RECT 81.600 246.200 82.200 246.800 ;
        RECT 81.200 245.600 82.200 246.200 ;
        RECT 81.200 242.200 82.000 245.600 ;
        RECT 84.400 242.200 85.200 259.800 ;
        RECT 86.000 256.300 86.800 257.200 ;
        RECT 89.200 256.300 90.000 259.800 ;
        RECT 86.000 255.700 90.000 256.300 ;
        RECT 86.000 255.600 86.800 255.700 ;
        RECT 89.000 255.200 90.000 255.700 ;
        RECT 89.000 250.800 89.800 255.200 ;
        RECT 90.800 254.600 91.600 259.800 ;
        RECT 97.200 256.600 98.000 259.800 ;
        RECT 98.800 257.000 99.600 259.800 ;
        RECT 100.400 257.000 101.200 259.800 ;
        RECT 102.000 257.000 102.800 259.800 ;
        RECT 103.600 257.000 104.400 259.800 ;
        RECT 106.800 257.000 107.600 259.800 ;
        RECT 110.000 257.000 110.800 259.800 ;
        RECT 111.600 257.000 112.400 259.800 ;
        RECT 113.200 257.000 114.000 259.800 ;
        RECT 95.600 255.800 98.000 256.600 ;
        RECT 114.800 256.600 115.600 259.800 ;
        RECT 95.600 255.200 96.400 255.800 ;
        RECT 90.400 254.000 91.600 254.600 ;
        RECT 94.600 254.600 96.400 255.200 ;
        RECT 100.400 255.600 101.400 256.400 ;
        RECT 104.400 255.600 106.000 256.400 ;
        RECT 106.800 255.800 111.400 256.400 ;
        RECT 114.800 255.800 117.400 256.600 ;
        RECT 106.800 255.600 107.600 255.800 ;
        RECT 90.400 252.000 91.000 254.000 ;
        RECT 94.600 253.400 95.400 254.600 ;
        RECT 91.600 252.600 95.400 253.400 ;
        RECT 100.400 252.800 101.200 255.600 ;
        RECT 106.800 254.800 107.600 255.000 ;
        RECT 103.200 254.200 107.600 254.800 ;
        RECT 103.200 254.000 104.000 254.200 ;
        RECT 108.400 253.600 109.200 255.200 ;
        RECT 110.600 253.400 111.400 255.800 ;
        RECT 116.600 255.200 117.400 255.800 ;
        RECT 116.600 254.400 119.600 255.200 ;
        RECT 121.200 253.800 122.000 259.800 ;
        RECT 129.200 255.200 130.000 259.800 ;
        RECT 132.400 255.200 133.200 259.800 ;
        RECT 135.600 255.200 136.400 259.800 ;
        RECT 138.800 255.200 139.600 259.800 ;
        RECT 103.600 252.600 106.800 253.400 ;
        RECT 110.600 252.600 112.600 253.400 ;
        RECT 113.200 253.000 122.000 253.800 ;
        RECT 97.200 252.000 98.000 252.600 ;
        RECT 114.800 252.000 115.600 252.400 ;
        RECT 118.000 252.000 118.800 252.400 ;
        RECT 119.800 252.000 120.600 252.200 ;
        RECT 90.400 251.400 91.200 252.000 ;
        RECT 97.200 251.400 120.600 252.000 ;
        RECT 89.000 250.000 90.000 250.800 ;
        RECT 89.200 242.200 90.000 250.000 ;
        RECT 90.600 249.600 91.200 251.400 ;
        RECT 90.600 249.000 99.600 249.600 ;
        RECT 90.600 247.400 91.200 249.000 ;
        RECT 98.800 248.800 99.600 249.000 ;
        RECT 102.000 249.000 110.600 249.600 ;
        RECT 102.000 248.800 102.800 249.000 ;
        RECT 93.800 247.600 96.400 248.400 ;
        RECT 90.600 246.800 93.200 247.400 ;
        RECT 92.400 242.200 93.200 246.800 ;
        RECT 95.600 242.200 96.400 247.600 ;
        RECT 97.000 246.800 101.200 247.600 ;
        RECT 98.800 242.200 99.600 245.000 ;
        RECT 100.400 242.200 101.200 245.000 ;
        RECT 102.000 242.200 102.800 245.000 ;
        RECT 103.600 242.200 104.400 248.400 ;
        RECT 106.800 247.600 109.400 248.400 ;
        RECT 110.000 248.200 110.600 249.000 ;
        RECT 111.600 249.400 112.400 249.600 ;
        RECT 111.600 249.000 117.000 249.400 ;
        RECT 111.600 248.800 117.800 249.000 ;
        RECT 116.400 248.200 117.800 248.800 ;
        RECT 110.000 247.600 115.800 248.200 ;
        RECT 118.800 248.000 120.400 248.800 ;
        RECT 118.800 247.600 119.400 248.000 ;
        RECT 106.800 242.200 107.600 247.000 ;
        RECT 110.000 242.200 110.800 247.000 ;
        RECT 115.200 246.800 119.400 247.600 ;
        RECT 121.200 247.400 122.000 253.000 ;
        RECT 127.600 254.400 130.000 255.200 ;
        RECT 131.000 254.400 133.200 255.200 ;
        RECT 134.200 254.400 136.400 255.200 ;
        RECT 137.800 254.400 139.600 255.200 ;
        RECT 143.600 255.200 144.400 259.800 ;
        RECT 146.800 255.200 147.600 259.800 ;
        RECT 150.000 255.200 150.800 259.800 ;
        RECT 153.200 255.200 154.000 259.800 ;
        RECT 156.400 255.600 157.200 257.200 ;
        RECT 143.600 254.400 145.400 255.200 ;
        RECT 146.800 254.400 149.000 255.200 ;
        RECT 150.000 254.400 152.200 255.200 ;
        RECT 153.200 254.400 155.600 255.200 ;
        RECT 127.600 251.600 128.400 254.400 ;
        RECT 131.000 253.800 131.800 254.400 ;
        RECT 134.200 253.800 135.000 254.400 ;
        RECT 137.800 253.800 138.600 254.400 ;
        RECT 140.400 254.300 141.200 254.400 ;
        RECT 142.000 254.300 142.800 254.400 ;
        RECT 140.400 253.800 142.800 254.300 ;
        RECT 144.600 253.800 145.400 254.400 ;
        RECT 148.200 253.800 149.000 254.400 ;
        RECT 151.400 253.800 152.200 254.400 ;
        RECT 129.200 253.000 131.800 253.800 ;
        RECT 132.600 253.000 135.000 253.800 ;
        RECT 136.000 253.000 138.600 253.800 ;
        RECT 139.400 253.700 143.800 253.800 ;
        RECT 139.400 253.000 141.200 253.700 ;
        RECT 142.000 253.000 143.800 253.700 ;
        RECT 144.600 253.000 147.200 253.800 ;
        RECT 148.200 253.000 150.600 253.800 ;
        RECT 151.400 253.000 154.000 253.800 ;
        RECT 131.000 251.600 131.800 253.000 ;
        RECT 134.200 251.600 135.000 253.000 ;
        RECT 137.800 251.600 138.600 253.000 ;
        RECT 144.600 251.600 145.400 253.000 ;
        RECT 148.200 251.600 149.000 253.000 ;
        RECT 151.400 251.600 152.200 253.000 ;
        RECT 154.800 251.600 155.600 254.400 ;
        RECT 127.600 250.800 130.000 251.600 ;
        RECT 131.000 250.800 133.200 251.600 ;
        RECT 134.200 250.800 136.400 251.600 ;
        RECT 137.800 250.800 139.600 251.600 ;
        RECT 120.000 246.800 122.000 247.400 ;
        RECT 111.600 242.200 112.400 245.000 ;
        RECT 113.200 242.200 114.000 245.000 ;
        RECT 116.400 242.200 117.200 246.800 ;
        RECT 120.000 246.200 120.600 246.800 ;
        RECT 119.600 245.600 120.600 246.200 ;
        RECT 119.600 242.200 120.400 245.600 ;
        RECT 129.200 242.200 130.000 250.800 ;
        RECT 132.400 242.200 133.200 250.800 ;
        RECT 135.600 242.200 136.400 250.800 ;
        RECT 138.800 242.200 139.600 250.800 ;
        RECT 143.600 250.800 145.400 251.600 ;
        RECT 146.800 250.800 149.000 251.600 ;
        RECT 150.000 250.800 152.200 251.600 ;
        RECT 153.200 250.800 155.600 251.600 ;
        RECT 158.000 252.300 158.800 259.800 ;
        RECT 163.400 256.000 164.200 259.000 ;
        RECT 167.600 257.000 168.400 259.000 ;
        RECT 162.600 255.400 164.200 256.000 ;
        RECT 162.600 255.000 163.400 255.400 ;
        RECT 162.600 254.400 163.200 255.000 ;
        RECT 167.800 254.800 168.400 257.000 ;
        RECT 169.200 255.600 170.000 257.200 ;
        RECT 159.600 254.300 160.400 254.400 ;
        RECT 161.200 254.300 163.200 254.400 ;
        RECT 159.600 253.700 163.200 254.300 ;
        RECT 164.200 254.200 168.400 254.800 ;
        RECT 164.200 253.800 165.200 254.200 ;
        RECT 159.600 253.600 160.400 253.700 ;
        RECT 161.200 253.600 163.200 253.700 ;
        RECT 161.200 252.300 162.000 252.400 ;
        RECT 158.000 251.700 162.000 252.300 ;
        RECT 143.600 242.200 144.400 250.800 ;
        RECT 146.800 242.200 147.600 250.800 ;
        RECT 150.000 242.200 150.800 250.800 ;
        RECT 153.200 242.200 154.000 250.800 ;
        RECT 158.000 242.200 158.800 251.700 ;
        RECT 161.200 250.800 162.000 251.700 ;
        RECT 162.600 249.800 163.200 253.600 ;
        RECT 163.800 253.000 165.200 253.800 ;
        RECT 164.600 251.000 165.200 253.000 ;
        RECT 166.000 251.600 166.800 253.200 ;
        RECT 167.600 251.600 168.400 253.200 ;
        RECT 170.800 252.300 171.600 259.800 ;
        RECT 176.200 256.000 177.000 259.000 ;
        RECT 180.400 257.000 181.200 259.000 ;
        RECT 175.400 255.400 177.000 256.000 ;
        RECT 175.400 255.000 176.200 255.400 ;
        RECT 175.400 254.400 176.000 255.000 ;
        RECT 180.600 254.800 181.200 257.000 ;
        RECT 182.000 255.600 182.800 257.200 ;
        RECT 174.000 253.600 176.000 254.400 ;
        RECT 177.000 254.200 181.200 254.800 ;
        RECT 177.000 253.800 178.000 254.200 ;
        RECT 174.000 252.300 174.800 252.400 ;
        RECT 170.800 251.700 174.800 252.300 ;
        RECT 164.600 250.400 168.400 251.000 ;
        RECT 162.600 249.200 164.200 249.800 ;
        RECT 163.400 242.200 164.200 249.200 ;
        RECT 167.800 247.000 168.400 250.400 ;
        RECT 167.600 243.000 168.400 247.000 ;
        RECT 170.800 242.200 171.600 251.700 ;
        RECT 174.000 250.800 174.800 251.700 ;
        RECT 175.400 249.800 176.000 253.600 ;
        RECT 176.600 253.000 178.000 253.800 ;
        RECT 177.400 251.000 178.000 253.000 ;
        RECT 178.800 251.600 179.600 253.200 ;
        RECT 180.400 251.600 181.200 253.200 ;
        RECT 177.400 250.400 181.200 251.000 ;
        RECT 175.400 249.200 177.000 249.800 ;
        RECT 176.200 244.400 177.000 249.200 ;
        RECT 180.600 247.000 181.200 250.400 ;
        RECT 175.600 243.600 177.000 244.400 ;
        RECT 176.200 242.200 177.000 243.600 ;
        RECT 180.400 243.000 181.200 247.000 ;
        RECT 183.600 242.200 184.400 259.800 ;
        RECT 185.200 253.800 186.000 259.800 ;
        RECT 191.600 256.600 192.400 259.800 ;
        RECT 193.200 257.000 194.000 259.800 ;
        RECT 194.800 257.000 195.600 259.800 ;
        RECT 196.400 257.000 197.200 259.800 ;
        RECT 199.600 257.000 200.400 259.800 ;
        RECT 202.800 257.000 203.600 259.800 ;
        RECT 204.400 257.000 205.200 259.800 ;
        RECT 206.000 257.000 206.800 259.800 ;
        RECT 207.600 257.000 208.400 259.800 ;
        RECT 189.800 255.800 192.400 256.600 ;
        RECT 209.200 256.600 210.000 259.800 ;
        RECT 195.800 255.800 200.400 256.400 ;
        RECT 189.800 255.200 190.600 255.800 ;
        RECT 187.600 254.400 190.600 255.200 ;
        RECT 185.200 253.000 194.000 253.800 ;
        RECT 195.800 253.400 196.600 255.800 ;
        RECT 199.600 255.600 200.400 255.800 ;
        RECT 201.200 255.600 202.800 256.400 ;
        RECT 205.800 255.600 206.800 256.400 ;
        RECT 209.200 255.800 211.600 256.600 ;
        RECT 198.000 253.600 198.800 255.200 ;
        RECT 199.600 254.800 200.400 255.000 ;
        RECT 199.600 254.200 204.000 254.800 ;
        RECT 203.200 254.000 204.000 254.200 ;
        RECT 185.200 247.400 186.000 253.000 ;
        RECT 194.600 252.600 196.600 253.400 ;
        RECT 200.400 252.600 203.600 253.400 ;
        RECT 206.000 252.800 206.800 255.600 ;
        RECT 210.800 255.200 211.600 255.800 ;
        RECT 210.800 254.600 212.600 255.200 ;
        RECT 211.800 253.400 212.600 254.600 ;
        RECT 215.600 254.600 216.400 259.800 ;
        RECT 217.200 256.000 218.000 259.800 ;
        RECT 217.200 255.200 218.200 256.000 ;
        RECT 220.400 255.600 221.200 257.200 ;
        RECT 215.600 254.000 216.800 254.600 ;
        RECT 211.800 252.600 215.600 253.400 ;
        RECT 186.800 252.200 187.600 252.400 ;
        RECT 186.600 252.000 187.600 252.200 ;
        RECT 191.600 252.000 192.400 252.400 ;
        RECT 209.200 252.000 210.000 252.600 ;
        RECT 216.200 252.000 216.800 254.000 ;
        RECT 186.600 251.400 210.000 252.000 ;
        RECT 216.000 251.400 216.800 252.000 ;
        RECT 216.000 249.600 216.600 251.400 ;
        RECT 217.400 250.800 218.200 255.200 ;
        RECT 194.800 249.400 195.600 249.600 ;
        RECT 190.200 249.000 195.600 249.400 ;
        RECT 189.400 248.800 195.600 249.000 ;
        RECT 196.600 249.000 205.200 249.600 ;
        RECT 186.800 248.000 188.400 248.800 ;
        RECT 189.400 248.200 190.800 248.800 ;
        RECT 196.600 248.200 197.200 249.000 ;
        RECT 204.400 248.800 205.200 249.000 ;
        RECT 207.600 249.000 216.600 249.600 ;
        RECT 207.600 248.800 208.400 249.000 ;
        RECT 187.800 247.600 188.400 248.000 ;
        RECT 191.400 247.600 197.200 248.200 ;
        RECT 197.800 247.600 200.400 248.400 ;
        RECT 185.200 246.800 187.200 247.400 ;
        RECT 187.800 246.800 192.000 247.600 ;
        RECT 186.600 246.200 187.200 246.800 ;
        RECT 186.600 245.600 187.600 246.200 ;
        RECT 186.800 242.200 187.600 245.600 ;
        RECT 190.000 242.200 190.800 246.800 ;
        RECT 193.200 242.200 194.000 245.000 ;
        RECT 194.800 242.200 195.600 245.000 ;
        RECT 196.400 242.200 197.200 247.000 ;
        RECT 199.600 242.200 200.400 247.000 ;
        RECT 202.800 242.200 203.600 248.400 ;
        RECT 210.800 247.600 213.400 248.400 ;
        RECT 206.000 246.800 210.200 247.600 ;
        RECT 204.400 242.200 205.200 245.000 ;
        RECT 206.000 242.200 206.800 245.000 ;
        RECT 207.600 242.200 208.400 245.000 ;
        RECT 210.800 242.200 211.600 247.600 ;
        RECT 216.000 247.400 216.600 249.000 ;
        RECT 214.000 246.800 216.600 247.400 ;
        RECT 217.200 250.000 218.200 250.800 ;
        RECT 214.000 242.200 214.800 246.800 ;
        RECT 217.200 242.200 218.000 250.000 ;
        RECT 222.000 242.200 222.800 259.800 ;
        RECT 225.200 256.000 226.000 259.800 ;
        RECT 225.000 255.200 226.000 256.000 ;
        RECT 225.000 250.800 225.800 255.200 ;
        RECT 226.800 254.600 227.600 259.800 ;
        RECT 233.200 256.600 234.000 259.800 ;
        RECT 234.800 257.000 235.600 259.800 ;
        RECT 236.400 257.000 237.200 259.800 ;
        RECT 238.000 257.000 238.800 259.800 ;
        RECT 239.600 257.000 240.400 259.800 ;
        RECT 242.800 257.000 243.600 259.800 ;
        RECT 246.000 257.000 246.800 259.800 ;
        RECT 247.600 257.000 248.400 259.800 ;
        RECT 249.200 257.000 250.000 259.800 ;
        RECT 231.600 255.800 234.000 256.600 ;
        RECT 250.800 256.600 251.600 259.800 ;
        RECT 231.600 255.200 232.400 255.800 ;
        RECT 226.400 254.000 227.600 254.600 ;
        RECT 230.600 254.600 232.400 255.200 ;
        RECT 236.400 255.600 237.400 256.400 ;
        RECT 240.400 255.600 242.000 256.400 ;
        RECT 242.800 255.800 247.400 256.400 ;
        RECT 250.800 255.800 253.400 256.600 ;
        RECT 242.800 255.600 243.600 255.800 ;
        RECT 226.400 252.000 227.000 254.000 ;
        RECT 230.600 253.400 231.400 254.600 ;
        RECT 227.600 252.600 231.400 253.400 ;
        RECT 236.400 252.800 237.200 255.600 ;
        RECT 242.800 254.800 243.600 255.000 ;
        RECT 239.200 254.200 243.600 254.800 ;
        RECT 239.200 254.000 240.000 254.200 ;
        RECT 244.400 253.600 245.200 255.200 ;
        RECT 246.600 253.400 247.400 255.800 ;
        RECT 252.600 255.200 253.400 255.800 ;
        RECT 252.600 254.400 255.600 255.200 ;
        RECT 257.200 253.800 258.000 259.800 ;
        RECT 258.800 255.600 259.600 257.200 ;
        RECT 239.600 252.600 242.800 253.400 ;
        RECT 246.600 252.600 248.600 253.400 ;
        RECT 249.200 253.000 258.000 253.800 ;
        RECT 233.200 252.000 234.000 252.600 ;
        RECT 244.400 252.000 245.200 252.400 ;
        RECT 250.800 252.000 251.600 252.400 ;
        RECT 255.800 252.000 256.600 252.200 ;
        RECT 226.400 251.400 227.200 252.000 ;
        RECT 233.200 251.400 256.600 252.000 ;
        RECT 225.000 250.000 226.000 250.800 ;
        RECT 225.200 242.200 226.000 250.000 ;
        RECT 226.600 249.600 227.200 251.400 ;
        RECT 226.600 249.000 235.600 249.600 ;
        RECT 226.600 247.400 227.200 249.000 ;
        RECT 234.800 248.800 235.600 249.000 ;
        RECT 238.000 249.000 246.600 249.600 ;
        RECT 238.000 248.800 238.800 249.000 ;
        RECT 229.800 247.600 232.400 248.400 ;
        RECT 226.600 246.800 229.200 247.400 ;
        RECT 228.400 242.200 229.200 246.800 ;
        RECT 231.600 242.200 232.400 247.600 ;
        RECT 233.000 246.800 237.200 247.600 ;
        RECT 234.800 242.200 235.600 245.000 ;
        RECT 236.400 242.200 237.200 245.000 ;
        RECT 238.000 242.200 238.800 245.000 ;
        RECT 239.600 242.200 240.400 248.400 ;
        RECT 242.800 247.600 245.400 248.400 ;
        RECT 246.000 248.200 246.600 249.000 ;
        RECT 247.600 249.400 248.400 249.600 ;
        RECT 247.600 249.000 253.000 249.400 ;
        RECT 247.600 248.800 253.800 249.000 ;
        RECT 252.400 248.200 253.800 248.800 ;
        RECT 246.000 247.600 251.800 248.200 ;
        RECT 254.800 248.000 256.400 248.800 ;
        RECT 254.800 247.600 255.400 248.000 ;
        RECT 242.800 242.200 243.600 247.000 ;
        RECT 246.000 242.200 246.800 247.000 ;
        RECT 251.200 246.800 255.400 247.600 ;
        RECT 257.200 247.400 258.000 253.000 ;
        RECT 256.000 246.800 258.000 247.400 ;
        RECT 260.400 254.300 261.200 259.800 ;
        RECT 266.800 256.000 267.600 259.800 ;
        RECT 270.000 256.000 270.800 259.800 ;
        RECT 266.800 255.800 270.800 256.000 ;
        RECT 271.600 255.800 272.400 259.800 ;
        RECT 274.800 256.000 275.600 259.800 ;
        RECT 267.000 255.400 270.600 255.800 ;
        RECT 267.600 254.400 268.400 254.800 ;
        RECT 271.600 254.400 272.200 255.800 ;
        RECT 274.600 255.200 275.600 256.000 ;
        RECT 266.800 254.300 268.400 254.400 ;
        RECT 260.400 253.800 268.400 254.300 ;
        RECT 260.400 253.700 267.600 253.800 ;
        RECT 247.600 242.200 248.400 245.000 ;
        RECT 249.200 242.200 250.000 245.000 ;
        RECT 252.400 242.200 253.200 246.800 ;
        RECT 256.000 246.200 256.600 246.800 ;
        RECT 255.600 245.600 256.600 246.200 ;
        RECT 255.600 242.200 256.400 245.600 ;
        RECT 260.400 242.200 261.200 253.700 ;
        RECT 266.800 253.600 267.600 253.700 ;
        RECT 269.800 253.600 272.400 254.400 ;
        RECT 268.400 251.600 269.200 253.200 ;
        RECT 269.800 250.200 270.400 253.600 ;
        RECT 274.600 250.800 275.400 255.200 ;
        RECT 276.400 254.600 277.200 259.800 ;
        RECT 282.800 256.600 283.600 259.800 ;
        RECT 284.400 257.000 285.200 259.800 ;
        RECT 286.000 257.000 286.800 259.800 ;
        RECT 287.600 257.000 288.400 259.800 ;
        RECT 289.200 257.000 290.000 259.800 ;
        RECT 292.400 257.000 293.200 259.800 ;
        RECT 295.600 257.000 296.400 259.800 ;
        RECT 297.200 257.000 298.000 259.800 ;
        RECT 298.800 257.000 299.600 259.800 ;
        RECT 281.200 255.800 283.600 256.600 ;
        RECT 300.400 256.600 301.200 259.800 ;
        RECT 281.200 255.200 282.000 255.800 ;
        RECT 276.000 254.000 277.200 254.600 ;
        RECT 280.200 254.600 282.000 255.200 ;
        RECT 286.000 255.600 287.000 256.400 ;
        RECT 290.000 255.600 291.600 256.400 ;
        RECT 292.400 255.800 297.000 256.400 ;
        RECT 300.400 255.800 303.000 256.600 ;
        RECT 292.400 255.600 293.200 255.800 ;
        RECT 276.000 252.000 276.600 254.000 ;
        RECT 280.200 253.400 281.000 254.600 ;
        RECT 277.200 252.600 281.000 253.400 ;
        RECT 286.000 252.800 286.800 255.600 ;
        RECT 292.400 254.800 293.200 255.000 ;
        RECT 288.800 254.200 293.200 254.800 ;
        RECT 288.800 254.000 289.600 254.200 ;
        RECT 294.000 253.600 294.800 255.200 ;
        RECT 296.200 253.400 297.000 255.800 ;
        RECT 302.200 255.200 303.000 255.800 ;
        RECT 302.200 254.400 305.200 255.200 ;
        RECT 306.800 253.800 307.600 259.800 ;
        RECT 312.000 254.200 312.800 259.800 ;
        RECT 318.400 254.200 319.200 259.800 ;
        RECT 321.200 255.800 322.000 259.800 ;
        RECT 322.800 256.000 323.600 259.800 ;
        RECT 326.000 256.000 326.800 259.800 ;
        RECT 322.800 255.800 326.800 256.000 ;
        RECT 327.600 259.200 331.600 259.800 ;
        RECT 327.600 255.800 328.400 259.200 ;
        RECT 321.400 254.400 322.000 255.800 ;
        RECT 323.000 255.400 326.600 255.800 ;
        RECT 329.200 255.600 330.000 258.600 ;
        RECT 330.800 256.000 331.600 259.200 ;
        RECT 334.000 256.000 334.800 259.800 ;
        RECT 338.200 256.400 339.000 259.800 ;
        RECT 330.800 255.800 334.800 256.000 ;
        RECT 337.200 255.800 339.000 256.400 ;
        RECT 325.200 254.400 326.000 254.800 ;
        RECT 329.200 254.400 329.800 255.600 ;
        RECT 331.000 255.400 334.600 255.800 ;
        RECT 333.200 254.400 334.000 254.800 ;
        RECT 312.000 253.800 313.800 254.200 ;
        RECT 318.400 253.800 320.200 254.200 ;
        RECT 289.200 252.600 292.400 253.400 ;
        RECT 296.200 252.600 298.200 253.400 ;
        RECT 298.800 253.000 307.600 253.800 ;
        RECT 312.200 253.600 313.800 253.800 ;
        RECT 318.600 253.600 320.200 253.800 ;
        RECT 321.200 253.600 323.800 254.400 ;
        RECT 325.200 253.800 326.800 254.400 ;
        RECT 326.000 253.600 326.800 253.800 ;
        RECT 282.800 252.000 283.600 252.600 ;
        RECT 300.400 252.000 301.200 252.400 ;
        RECT 302.000 252.000 302.800 252.400 ;
        RECT 305.400 252.000 306.200 252.200 ;
        RECT 276.000 251.400 276.800 252.000 ;
        RECT 282.800 251.400 306.200 252.000 ;
        RECT 271.600 250.200 272.400 250.400 ;
        RECT 269.400 249.600 270.400 250.200 ;
        RECT 271.000 249.600 272.400 250.200 ;
        RECT 274.600 250.000 275.600 250.800 ;
        RECT 269.400 242.200 270.200 249.600 ;
        RECT 271.000 248.400 271.600 249.600 ;
        RECT 270.800 247.600 271.600 248.400 ;
        RECT 274.800 242.200 275.600 250.000 ;
        RECT 276.200 249.600 276.800 251.400 ;
        RECT 276.200 249.000 285.200 249.600 ;
        RECT 276.200 247.400 276.800 249.000 ;
        RECT 284.400 248.800 285.200 249.000 ;
        RECT 287.600 249.000 296.200 249.600 ;
        RECT 287.600 248.800 288.400 249.000 ;
        RECT 279.400 247.600 282.000 248.400 ;
        RECT 276.200 246.800 278.800 247.400 ;
        RECT 278.000 242.200 278.800 246.800 ;
        RECT 281.200 242.200 282.000 247.600 ;
        RECT 282.600 246.800 286.800 247.600 ;
        RECT 284.400 242.200 285.200 245.000 ;
        RECT 286.000 242.200 286.800 245.000 ;
        RECT 287.600 242.200 288.400 245.000 ;
        RECT 289.200 242.200 290.000 248.400 ;
        RECT 292.400 247.600 295.000 248.400 ;
        RECT 295.600 248.200 296.200 249.000 ;
        RECT 297.200 249.400 298.000 249.600 ;
        RECT 297.200 249.000 302.600 249.400 ;
        RECT 297.200 248.800 303.400 249.000 ;
        RECT 302.000 248.200 303.400 248.800 ;
        RECT 295.600 247.600 301.400 248.200 ;
        RECT 304.400 248.000 306.000 248.800 ;
        RECT 304.400 247.600 305.000 248.000 ;
        RECT 292.400 242.200 293.200 247.000 ;
        RECT 295.600 242.200 296.400 247.000 ;
        RECT 300.800 246.800 305.000 247.600 ;
        RECT 306.800 247.400 307.600 253.000 ;
        RECT 310.000 251.600 311.600 252.400 ;
        RECT 313.200 250.400 313.800 253.600 ;
        RECT 316.400 251.600 318.000 252.400 ;
        RECT 319.600 250.400 320.200 253.600 ;
        RECT 323.200 250.400 323.800 253.600 ;
        RECT 324.400 251.600 325.200 253.200 ;
        RECT 327.600 252.800 328.400 254.400 ;
        RECT 329.200 253.800 331.600 254.400 ;
        RECT 333.200 253.800 334.800 254.400 ;
        RECT 330.800 253.600 331.600 253.800 ;
        RECT 334.000 253.600 334.800 253.800 ;
        RECT 335.600 253.600 336.400 255.200 ;
        RECT 329.200 251.600 330.000 253.200 ;
        RECT 313.200 249.600 314.000 250.400 ;
        RECT 319.600 249.600 320.400 250.400 ;
        RECT 321.200 250.200 322.000 250.400 ;
        RECT 321.200 249.600 322.600 250.200 ;
        RECT 323.200 249.600 325.200 250.400 ;
        RECT 331.000 250.200 331.600 253.600 ;
        RECT 332.400 251.600 333.200 253.200 ;
        RECT 311.600 247.600 312.400 249.200 ;
        RECT 305.600 246.800 307.600 247.400 ;
        RECT 313.200 247.000 313.800 249.600 ;
        RECT 318.000 247.600 318.800 249.200 ;
        RECT 319.600 247.000 320.200 249.600 ;
        RECT 322.000 248.400 322.600 249.600 ;
        RECT 322.000 247.600 322.800 248.400 ;
        RECT 297.200 242.200 298.000 245.000 ;
        RECT 298.800 242.200 299.600 245.000 ;
        RECT 302.000 242.200 302.800 246.800 ;
        RECT 305.600 246.200 306.200 246.800 ;
        RECT 310.200 246.400 313.800 247.000 ;
        RECT 310.200 246.200 310.800 246.400 ;
        RECT 305.200 245.600 306.200 246.200 ;
        RECT 305.200 242.200 306.000 245.600 ;
        RECT 310.000 242.200 310.800 246.200 ;
        RECT 313.200 246.200 313.800 246.400 ;
        RECT 316.600 246.400 320.200 247.000 ;
        RECT 316.600 246.200 317.200 246.400 ;
        RECT 313.200 242.200 314.000 246.200 ;
        RECT 316.400 242.200 317.200 246.200 ;
        RECT 319.600 246.200 320.200 246.400 ;
        RECT 319.600 242.200 320.400 246.200 ;
        RECT 323.400 242.200 324.200 249.600 ;
        RECT 330.200 242.200 332.200 250.200 ;
        RECT 337.200 242.200 338.000 255.800 ;
        RECT 342.000 255.200 342.800 259.800 ;
        RECT 345.200 255.200 346.000 259.800 ;
        RECT 348.400 255.200 349.200 259.800 ;
        RECT 351.600 255.200 352.400 259.800 ;
        RECT 354.800 255.800 355.600 259.800 ;
        RECT 356.400 256.000 357.200 259.800 ;
        RECT 359.600 256.000 360.400 259.800 ;
        RECT 356.400 255.800 360.400 256.000 ;
        RECT 361.200 256.000 362.000 259.800 ;
        RECT 364.400 259.200 368.400 259.800 ;
        RECT 364.400 256.000 365.200 259.200 ;
        RECT 361.200 255.800 365.200 256.000 ;
        RECT 366.000 255.800 366.800 258.600 ;
        RECT 367.600 255.800 368.400 259.200 ;
        RECT 371.800 256.400 372.600 259.800 ;
        RECT 370.800 255.800 372.600 256.400 ;
        RECT 374.000 256.000 374.800 259.800 ;
        RECT 377.200 256.000 378.000 259.800 ;
        RECT 374.000 255.800 378.000 256.000 ;
        RECT 378.800 255.800 379.600 259.800 ;
        RECT 382.000 257.800 382.800 259.800 ;
        RECT 340.400 254.400 342.800 255.200 ;
        RECT 343.800 254.400 346.000 255.200 ;
        RECT 347.000 254.400 349.200 255.200 ;
        RECT 350.600 254.400 352.400 255.200 ;
        RECT 355.000 254.400 355.600 255.800 ;
        RECT 356.600 255.400 360.200 255.800 ;
        RECT 361.400 255.400 365.000 255.800 ;
        RECT 358.800 254.400 359.600 254.800 ;
        RECT 362.000 254.400 362.800 254.800 ;
        RECT 366.200 254.400 366.800 255.800 ;
        RECT 340.400 251.600 341.200 254.400 ;
        RECT 343.800 253.800 344.600 254.400 ;
        RECT 347.000 253.800 347.800 254.400 ;
        RECT 350.600 253.800 351.400 254.400 ;
        RECT 353.200 253.800 354.000 254.400 ;
        RECT 342.000 253.000 344.600 253.800 ;
        RECT 345.400 253.000 347.800 253.800 ;
        RECT 348.800 253.000 351.400 253.800 ;
        RECT 352.200 253.000 354.000 253.800 ;
        RECT 354.800 253.600 357.400 254.400 ;
        RECT 358.800 253.800 360.400 254.400 ;
        RECT 359.600 253.600 360.400 253.800 ;
        RECT 361.200 253.800 362.800 254.400 ;
        RECT 364.400 253.800 366.800 254.400 ;
        RECT 361.200 253.600 362.000 253.800 ;
        RECT 364.400 253.600 365.200 253.800 ;
        RECT 343.800 251.600 344.600 253.000 ;
        RECT 347.000 251.600 347.800 253.000 ;
        RECT 350.600 251.600 351.400 253.000 ;
        RECT 340.400 250.800 342.800 251.600 ;
        RECT 343.800 250.800 346.000 251.600 ;
        RECT 347.000 250.800 349.200 251.600 ;
        RECT 350.600 250.800 352.400 251.600 ;
        RECT 338.800 248.800 339.600 250.400 ;
        RECT 342.000 242.200 342.800 250.800 ;
        RECT 345.200 242.200 346.000 250.800 ;
        RECT 348.400 242.200 349.200 250.800 ;
        RECT 351.600 242.200 352.400 250.800 ;
        RECT 356.800 250.400 357.400 253.600 ;
        RECT 359.600 252.300 360.400 252.400 ;
        RECT 362.800 252.300 363.600 253.200 ;
        RECT 359.600 251.700 363.600 252.300 ;
        RECT 359.600 251.600 360.400 251.700 ;
        RECT 362.800 251.600 363.600 251.700 ;
        RECT 354.800 250.200 355.600 250.400 ;
        RECT 354.800 249.600 356.200 250.200 ;
        RECT 356.800 249.600 358.800 250.400 ;
        RECT 364.400 250.200 365.000 253.600 ;
        RECT 366.000 251.600 366.800 253.200 ;
        RECT 367.600 252.800 368.400 254.400 ;
        RECT 369.200 253.600 370.000 255.200 ;
        RECT 355.600 248.400 356.200 249.600 ;
        RECT 355.600 247.600 356.400 248.400 ;
        RECT 357.000 242.200 357.800 249.600 ;
        RECT 363.800 244.400 365.800 250.200 ;
        RECT 362.800 243.600 365.800 244.400 ;
        RECT 363.800 242.200 365.800 243.600 ;
        RECT 370.800 242.200 371.600 255.800 ;
        RECT 374.200 255.400 377.800 255.800 ;
        RECT 374.800 254.400 375.600 254.800 ;
        RECT 378.800 254.400 379.400 255.800 ;
        RECT 380.400 255.600 381.200 257.200 ;
        RECT 382.200 254.400 382.800 257.800 ;
        RECT 374.000 253.800 375.600 254.400 ;
        RECT 374.000 253.600 374.800 253.800 ;
        RECT 377.000 253.600 379.600 254.400 ;
        RECT 380.400 254.300 381.200 254.400 ;
        RECT 382.000 254.300 382.800 254.400 ;
        RECT 380.400 253.700 382.800 254.300 ;
        RECT 388.800 254.200 389.600 259.800 ;
        RECT 388.800 253.800 390.600 254.200 ;
        RECT 380.400 253.600 381.200 253.700 ;
        RECT 382.000 253.600 382.800 253.700 ;
        RECT 389.000 253.600 390.600 253.800 ;
        RECT 372.400 252.300 373.200 252.400 ;
        RECT 375.600 252.300 376.400 253.200 ;
        RECT 372.400 251.700 376.400 252.300 ;
        RECT 372.400 251.600 373.200 251.700 ;
        RECT 375.600 251.600 376.400 251.700 ;
        RECT 372.400 248.800 373.200 250.400 ;
        RECT 377.000 250.200 377.600 253.600 ;
        RECT 378.800 250.200 379.600 250.400 ;
        RECT 382.200 250.200 382.800 253.600 ;
        RECT 383.600 250.800 384.400 252.400 ;
        RECT 386.800 251.600 388.400 252.400 ;
        RECT 376.600 249.600 377.600 250.200 ;
        RECT 378.200 249.600 379.600 250.200 ;
        RECT 376.600 244.400 377.400 249.600 ;
        RECT 378.200 248.400 378.800 249.600 ;
        RECT 382.000 249.400 383.800 250.200 ;
        RECT 385.200 249.600 386.000 251.200 ;
        RECT 390.000 250.400 390.600 253.600 ;
        RECT 390.000 249.600 390.800 250.400 ;
        RECT 378.000 247.600 378.800 248.400 ;
        RECT 375.600 243.600 377.400 244.400 ;
        RECT 376.600 242.200 377.400 243.600 ;
        RECT 383.000 242.200 383.800 249.400 ;
        RECT 388.400 247.600 389.200 249.200 ;
        RECT 390.000 247.000 390.600 249.600 ;
        RECT 387.000 246.400 390.600 247.000 ;
        RECT 387.000 246.200 387.600 246.400 ;
        RECT 386.800 242.200 387.600 246.200 ;
        RECT 390.000 242.200 390.800 246.400 ;
        RECT 391.600 242.200 392.400 259.800 ;
        RECT 395.400 258.400 396.200 259.800 ;
        RECT 394.800 257.600 396.200 258.400 ;
        RECT 395.400 256.400 396.200 257.600 ;
        RECT 395.400 255.800 397.200 256.400 ;
        RECT 393.200 250.300 394.000 250.400 ;
        RECT 394.800 250.300 395.600 250.400 ;
        RECT 393.200 249.700 395.600 250.300 ;
        RECT 393.200 249.600 394.000 249.700 ;
        RECT 394.800 248.800 395.600 249.700 ;
        RECT 396.400 242.200 397.200 255.800 ;
        RECT 399.600 255.200 400.400 259.800 ;
        RECT 402.800 256.400 403.600 259.800 ;
        RECT 402.800 255.800 403.800 256.400 ;
        RECT 398.000 253.600 398.800 255.200 ;
        RECT 399.600 254.600 402.200 255.200 ;
        RECT 399.800 252.400 400.600 253.200 ;
        RECT 399.600 251.600 400.600 252.400 ;
        RECT 401.600 253.000 402.200 254.600 ;
        RECT 403.200 254.400 403.800 255.800 ;
        RECT 402.800 253.600 403.800 254.400 ;
        RECT 401.600 252.200 402.600 253.000 ;
        RECT 401.600 250.200 402.200 252.200 ;
        RECT 403.200 250.200 403.800 253.600 ;
        RECT 399.600 249.600 402.200 250.200 ;
        RECT 399.600 242.200 400.400 249.600 ;
        RECT 402.800 249.200 403.800 250.200 ;
        RECT 406.000 255.800 406.800 259.800 ;
        RECT 409.200 257.800 410.000 259.800 ;
        RECT 406.000 252.400 406.600 255.800 ;
        RECT 409.200 255.600 409.800 257.800 ;
        RECT 410.800 255.600 411.600 257.200 ;
        RECT 407.400 255.000 409.800 255.600 ;
        RECT 406.000 251.600 406.800 252.400 ;
        RECT 407.400 252.000 408.000 255.000 ;
        RECT 416.000 254.200 416.800 259.800 ;
        RECT 416.000 253.800 417.800 254.200 ;
        RECT 416.200 253.600 417.800 253.800 ;
        RECT 406.000 250.200 406.600 251.600 ;
        RECT 407.400 251.400 408.200 252.000 ;
        RECT 407.400 251.200 411.600 251.400 ;
        RECT 407.600 250.800 411.600 251.200 ;
        RECT 406.000 249.600 407.400 250.200 ;
        RECT 402.800 242.200 403.600 249.200 ;
        RECT 406.600 242.200 407.400 249.600 ;
        RECT 410.800 242.200 411.600 250.800 ;
        RECT 412.400 249.600 413.200 251.200 ;
        RECT 417.200 250.400 417.800 253.600 ;
        RECT 423.600 253.800 424.400 259.800 ;
        RECT 430.000 256.600 430.800 259.800 ;
        RECT 431.600 257.000 432.400 259.800 ;
        RECT 433.200 257.000 434.000 259.800 ;
        RECT 434.800 257.000 435.600 259.800 ;
        RECT 438.000 257.000 438.800 259.800 ;
        RECT 441.200 257.000 442.000 259.800 ;
        RECT 442.800 257.000 443.600 259.800 ;
        RECT 444.400 257.000 445.200 259.800 ;
        RECT 446.000 257.000 446.800 259.800 ;
        RECT 428.200 255.800 430.800 256.600 ;
        RECT 447.600 256.600 448.400 259.800 ;
        RECT 434.200 255.800 438.800 256.400 ;
        RECT 428.200 255.200 429.000 255.800 ;
        RECT 426.000 254.400 429.000 255.200 ;
        RECT 423.600 253.000 432.400 253.800 ;
        RECT 434.200 253.400 435.000 255.800 ;
        RECT 438.000 255.600 438.800 255.800 ;
        RECT 439.600 255.600 441.200 256.400 ;
        RECT 444.200 255.600 445.200 256.400 ;
        RECT 447.600 255.800 450.000 256.600 ;
        RECT 436.400 253.600 437.200 255.200 ;
        RECT 438.000 254.800 438.800 255.000 ;
        RECT 438.000 254.200 442.400 254.800 ;
        RECT 441.600 254.000 442.400 254.200 ;
        RECT 417.200 249.600 418.000 250.400 ;
        RECT 415.600 247.600 416.400 249.200 ;
        RECT 417.200 247.000 417.800 249.600 ;
        RECT 414.200 246.400 417.800 247.000 ;
        RECT 423.600 247.400 424.400 253.000 ;
        RECT 433.000 252.600 435.000 253.400 ;
        RECT 438.800 252.600 442.000 253.400 ;
        RECT 444.400 252.800 445.200 255.600 ;
        RECT 449.200 255.200 450.000 255.800 ;
        RECT 449.200 254.600 451.000 255.200 ;
        RECT 450.200 253.400 451.000 254.600 ;
        RECT 454.000 254.600 454.800 259.800 ;
        RECT 455.600 256.000 456.400 259.800 ;
        RECT 458.800 257.000 459.600 259.000 ;
        RECT 463.000 258.400 463.800 259.000 ;
        RECT 463.000 257.600 464.400 258.400 ;
        RECT 455.600 255.200 456.600 256.000 ;
        RECT 454.000 254.000 455.200 254.600 ;
        RECT 450.200 252.600 454.000 253.400 ;
        RECT 425.000 252.000 425.800 252.200 ;
        RECT 426.800 252.000 427.600 252.400 ;
        RECT 430.000 252.000 430.800 252.400 ;
        RECT 447.600 252.000 448.400 252.600 ;
        RECT 454.600 252.000 455.200 254.000 ;
        RECT 425.000 251.400 448.400 252.000 ;
        RECT 454.400 251.400 455.200 252.000 ;
        RECT 454.400 249.600 455.000 251.400 ;
        RECT 455.800 250.800 456.600 255.200 ;
        RECT 458.800 254.800 459.400 257.000 ;
        RECT 463.000 256.000 463.800 257.600 ;
        RECT 463.000 255.400 464.600 256.000 ;
        RECT 463.800 255.000 464.600 255.400 ;
        RECT 458.800 254.200 463.000 254.800 ;
        RECT 462.000 253.800 463.000 254.200 ;
        RECT 464.000 254.400 464.600 255.000 ;
        RECT 457.200 252.300 458.000 252.400 ;
        RECT 458.800 252.300 459.600 253.200 ;
        RECT 457.200 251.700 459.600 252.300 ;
        RECT 457.200 251.600 458.000 251.700 ;
        RECT 458.800 251.600 459.600 251.700 ;
        RECT 460.400 251.600 461.200 253.200 ;
        RECT 462.000 253.000 463.400 253.800 ;
        RECT 464.000 253.600 466.000 254.400 ;
        RECT 462.000 251.000 462.600 253.000 ;
        RECT 433.200 249.400 434.000 249.600 ;
        RECT 428.600 249.000 434.000 249.400 ;
        RECT 427.800 248.800 434.000 249.000 ;
        RECT 435.000 249.000 443.600 249.600 ;
        RECT 425.200 248.000 426.800 248.800 ;
        RECT 427.800 248.200 429.200 248.800 ;
        RECT 435.000 248.200 435.600 249.000 ;
        RECT 442.800 248.800 443.600 249.000 ;
        RECT 446.000 249.000 455.000 249.600 ;
        RECT 446.000 248.800 446.800 249.000 ;
        RECT 426.200 247.600 426.800 248.000 ;
        RECT 429.800 247.600 435.600 248.200 ;
        RECT 436.200 247.600 438.800 248.400 ;
        RECT 423.600 246.800 425.600 247.400 ;
        RECT 426.200 246.800 430.400 247.600 ;
        RECT 414.000 242.200 414.800 246.400 ;
        RECT 417.200 246.200 417.800 246.400 ;
        RECT 425.000 246.200 425.600 246.800 ;
        RECT 417.200 242.200 418.000 246.200 ;
        RECT 425.000 245.600 426.000 246.200 ;
        RECT 425.200 242.200 426.000 245.600 ;
        RECT 428.400 242.200 429.200 246.800 ;
        RECT 431.600 242.200 432.400 245.000 ;
        RECT 433.200 242.200 434.000 245.000 ;
        RECT 434.800 242.200 435.600 247.000 ;
        RECT 438.000 242.200 438.800 247.000 ;
        RECT 441.200 242.200 442.000 248.400 ;
        RECT 449.200 247.600 451.800 248.400 ;
        RECT 444.400 246.800 448.600 247.600 ;
        RECT 442.800 242.200 443.600 245.000 ;
        RECT 444.400 242.200 445.200 245.000 ;
        RECT 446.000 242.200 446.800 245.000 ;
        RECT 449.200 242.200 450.000 247.600 ;
        RECT 454.400 247.400 455.000 249.000 ;
        RECT 452.400 246.800 455.000 247.400 ;
        RECT 455.600 250.000 456.600 250.800 ;
        RECT 458.800 250.400 462.600 251.000 ;
        RECT 452.400 242.200 453.200 246.800 ;
        RECT 455.600 242.200 456.400 250.000 ;
        RECT 458.800 247.000 459.400 250.400 ;
        RECT 464.000 249.800 464.600 253.600 ;
        RECT 465.200 252.300 466.000 252.400 ;
        RECT 468.400 252.300 469.200 259.800 ;
        RECT 470.000 255.600 470.800 257.200 ;
        RECT 473.200 255.200 474.000 259.800 ;
        RECT 476.400 255.200 477.200 259.800 ;
        RECT 479.600 255.200 480.400 259.800 ;
        RECT 482.800 255.200 483.600 259.800 ;
        RECT 465.200 251.700 469.200 252.300 ;
        RECT 465.200 250.800 466.000 251.700 ;
        RECT 463.000 249.200 464.600 249.800 ;
        RECT 458.800 243.000 459.600 247.000 ;
        RECT 463.000 242.200 463.800 249.200 ;
        RECT 468.400 242.200 469.200 251.700 ;
        RECT 471.600 254.400 474.000 255.200 ;
        RECT 475.000 254.400 477.200 255.200 ;
        RECT 478.200 254.400 480.400 255.200 ;
        RECT 481.800 254.400 483.600 255.200 ;
        RECT 486.000 257.000 486.800 259.000 ;
        RECT 490.200 258.400 491.000 259.000 ;
        RECT 489.200 257.600 491.000 258.400 ;
        RECT 486.000 254.800 486.600 257.000 ;
        RECT 490.200 256.000 491.000 257.600 ;
        RECT 490.200 255.400 491.800 256.000 ;
        RECT 491.000 255.000 491.800 255.400 ;
        RECT 471.600 251.600 472.400 254.400 ;
        RECT 475.000 253.800 475.800 254.400 ;
        RECT 478.200 253.800 479.000 254.400 ;
        RECT 481.800 253.800 482.600 254.400 ;
        RECT 484.400 253.800 485.200 254.400 ;
        RECT 486.000 254.200 490.200 254.800 ;
        RECT 473.200 253.000 475.800 253.800 ;
        RECT 476.600 253.000 479.000 253.800 ;
        RECT 480.000 253.000 482.600 253.800 ;
        RECT 483.400 253.000 485.200 253.800 ;
        RECT 489.200 253.800 490.200 254.200 ;
        RECT 491.200 254.400 491.800 255.000 ;
        RECT 475.000 251.600 475.800 253.000 ;
        RECT 478.200 251.600 479.000 253.000 ;
        RECT 481.800 251.600 482.600 253.000 ;
        RECT 486.000 251.600 486.800 253.200 ;
        RECT 487.600 251.600 488.400 253.200 ;
        RECT 489.200 253.000 490.600 253.800 ;
        RECT 491.200 253.600 493.200 254.400 ;
        RECT 471.600 250.800 474.000 251.600 ;
        RECT 475.000 250.800 477.200 251.600 ;
        RECT 478.200 250.800 480.400 251.600 ;
        RECT 481.800 250.800 483.600 251.600 ;
        RECT 489.200 251.000 489.800 253.000 ;
        RECT 473.200 242.200 474.000 250.800 ;
        RECT 476.400 242.200 477.200 250.800 ;
        RECT 479.600 242.200 480.400 250.800 ;
        RECT 482.800 242.200 483.600 250.800 ;
        RECT 486.000 250.400 489.800 251.000 ;
        RECT 486.000 247.000 486.600 250.400 ;
        RECT 491.200 249.800 491.800 253.600 ;
        RECT 492.400 252.300 493.200 252.400 ;
        RECT 495.600 252.300 496.400 259.800 ;
        RECT 497.200 255.600 498.000 257.200 ;
        RECT 498.800 257.000 499.600 259.000 ;
        RECT 498.800 254.800 499.400 257.000 ;
        RECT 503.000 256.000 503.800 259.000 ;
        RECT 503.000 255.400 504.600 256.000 ;
        RECT 503.800 255.000 504.600 255.400 ;
        RECT 498.800 254.200 503.000 254.800 ;
        RECT 502.000 253.800 503.000 254.200 ;
        RECT 504.000 254.400 504.600 255.000 ;
        RECT 504.000 254.300 506.000 254.400 ;
        RECT 506.800 254.300 507.600 254.400 ;
        RECT 492.400 251.700 496.400 252.300 ;
        RECT 492.400 250.800 493.200 251.700 ;
        RECT 490.200 249.200 491.800 249.800 ;
        RECT 486.000 243.000 486.800 247.000 ;
        RECT 490.200 242.200 491.000 249.200 ;
        RECT 495.600 242.200 496.400 251.700 ;
        RECT 498.800 251.600 499.600 253.200 ;
        RECT 500.400 251.600 501.200 253.200 ;
        RECT 502.000 253.000 503.400 253.800 ;
        RECT 504.000 253.700 507.600 254.300 ;
        RECT 504.000 253.600 506.000 253.700 ;
        RECT 506.800 253.600 507.600 253.700 ;
        RECT 502.000 251.000 502.600 253.000 ;
        RECT 498.800 250.400 502.600 251.000 ;
        RECT 498.800 247.000 499.400 250.400 ;
        RECT 504.000 249.800 504.600 253.600 ;
        RECT 505.200 252.300 506.000 252.400 ;
        RECT 508.400 252.300 509.200 259.800 ;
        RECT 510.000 255.600 510.800 257.200 ;
        RECT 505.200 251.700 509.200 252.300 ;
        RECT 505.200 250.800 506.000 251.700 ;
        RECT 503.000 249.200 504.600 249.800 ;
        RECT 498.800 243.000 499.600 247.000 ;
        RECT 503.000 242.200 503.800 249.200 ;
        RECT 508.400 242.200 509.200 251.700 ;
        RECT 511.600 253.800 512.400 259.800 ;
        RECT 518.000 256.600 518.800 259.800 ;
        RECT 519.600 257.000 520.400 259.800 ;
        RECT 521.200 257.000 522.000 259.800 ;
        RECT 522.800 257.000 523.600 259.800 ;
        RECT 526.000 257.000 526.800 259.800 ;
        RECT 529.200 257.000 530.000 259.800 ;
        RECT 530.800 257.000 531.600 259.800 ;
        RECT 532.400 257.000 533.200 259.800 ;
        RECT 534.000 257.000 534.800 259.800 ;
        RECT 516.200 255.800 518.800 256.600 ;
        RECT 535.600 256.600 536.400 259.800 ;
        RECT 522.200 255.800 526.800 256.400 ;
        RECT 516.200 255.200 517.000 255.800 ;
        RECT 514.000 254.400 517.000 255.200 ;
        RECT 511.600 253.000 520.400 253.800 ;
        RECT 522.200 253.400 523.000 255.800 ;
        RECT 526.000 255.600 526.800 255.800 ;
        RECT 527.600 255.600 529.200 256.400 ;
        RECT 532.200 255.600 533.200 256.400 ;
        RECT 535.600 255.800 538.000 256.600 ;
        RECT 524.400 253.600 525.200 255.200 ;
        RECT 526.000 254.800 526.800 255.000 ;
        RECT 526.000 254.200 530.400 254.800 ;
        RECT 529.600 254.000 530.400 254.200 ;
        RECT 511.600 247.400 512.400 253.000 ;
        RECT 521.000 252.600 523.000 253.400 ;
        RECT 526.800 252.600 530.000 253.400 ;
        RECT 532.400 252.800 533.200 255.600 ;
        RECT 537.200 255.200 538.000 255.800 ;
        RECT 537.200 254.600 539.000 255.200 ;
        RECT 538.200 253.400 539.000 254.600 ;
        RECT 542.000 254.600 542.800 259.800 ;
        RECT 543.600 256.000 544.400 259.800 ;
        RECT 543.600 255.200 544.600 256.000 ;
        RECT 542.000 254.000 543.200 254.600 ;
        RECT 538.200 252.600 542.000 253.400 ;
        RECT 513.000 252.000 513.800 252.200 ;
        RECT 514.800 252.000 515.600 252.400 ;
        RECT 518.000 252.000 518.800 252.400 ;
        RECT 535.600 252.000 536.400 252.600 ;
        RECT 542.600 252.000 543.200 254.000 ;
        RECT 513.000 251.400 536.400 252.000 ;
        RECT 542.400 251.400 543.200 252.000 ;
        RECT 542.400 249.600 543.000 251.400 ;
        RECT 543.800 250.800 544.600 255.200 ;
        RECT 521.200 249.400 522.000 249.600 ;
        RECT 516.600 249.000 522.000 249.400 ;
        RECT 515.800 248.800 522.000 249.000 ;
        RECT 523.000 249.000 531.600 249.600 ;
        RECT 513.200 248.000 514.800 248.800 ;
        RECT 515.800 248.200 517.200 248.800 ;
        RECT 523.000 248.200 523.600 249.000 ;
        RECT 530.800 248.800 531.600 249.000 ;
        RECT 534.000 249.000 543.000 249.600 ;
        RECT 534.000 248.800 534.800 249.000 ;
        RECT 514.200 247.600 514.800 248.000 ;
        RECT 517.800 247.600 523.600 248.200 ;
        RECT 524.200 247.600 526.800 248.400 ;
        RECT 511.600 246.800 513.600 247.400 ;
        RECT 514.200 246.800 518.400 247.600 ;
        RECT 513.000 246.200 513.600 246.800 ;
        RECT 513.000 245.600 514.000 246.200 ;
        RECT 513.200 242.200 514.000 245.600 ;
        RECT 516.400 242.200 517.200 246.800 ;
        RECT 519.600 242.200 520.400 245.000 ;
        RECT 521.200 242.200 522.000 245.000 ;
        RECT 522.800 242.200 523.600 247.000 ;
        RECT 526.000 242.200 526.800 247.000 ;
        RECT 529.200 242.200 530.000 248.400 ;
        RECT 537.200 247.600 539.800 248.400 ;
        RECT 532.400 246.800 536.600 247.600 ;
        RECT 530.800 242.200 531.600 245.000 ;
        RECT 532.400 242.200 533.200 245.000 ;
        RECT 534.000 242.200 534.800 245.000 ;
        RECT 537.200 242.200 538.000 247.600 ;
        RECT 542.400 247.400 543.000 249.000 ;
        RECT 540.400 246.800 543.000 247.400 ;
        RECT 543.600 250.000 544.600 250.800 ;
        RECT 546.800 255.400 547.600 259.800 ;
        RECT 551.000 258.400 552.200 259.800 ;
        RECT 551.000 257.800 552.400 258.400 ;
        RECT 555.600 257.800 556.400 259.800 ;
        RECT 560.000 258.400 560.800 259.800 ;
        RECT 560.000 257.800 562.000 258.400 ;
        RECT 551.600 257.000 552.400 257.800 ;
        RECT 555.800 257.200 556.400 257.800 ;
        RECT 555.800 256.600 558.600 257.200 ;
        RECT 557.800 256.400 558.600 256.600 ;
        RECT 559.600 255.600 560.400 257.200 ;
        RECT 561.200 257.000 562.000 257.800 ;
        RECT 549.800 255.400 550.600 255.600 ;
        RECT 546.800 254.800 550.600 255.400 ;
        RECT 546.800 251.400 547.600 254.800 ;
        RECT 553.800 254.200 554.600 254.400 ;
        RECT 559.600 254.200 560.200 255.600 ;
        RECT 564.400 255.000 565.200 259.800 ;
        RECT 566.000 256.000 566.800 259.800 ;
        RECT 569.200 256.000 570.000 259.800 ;
        RECT 566.000 255.800 570.000 256.000 ;
        RECT 570.800 255.800 571.600 259.800 ;
        RECT 577.200 255.800 578.000 259.800 ;
        RECT 578.800 256.000 579.600 259.800 ;
        RECT 582.000 256.000 582.800 259.800 ;
        RECT 578.800 255.800 582.800 256.000 ;
        RECT 566.200 255.400 569.800 255.800 ;
        RECT 566.800 254.400 567.600 254.800 ;
        RECT 570.800 254.400 571.400 255.800 ;
        RECT 577.400 254.400 578.000 255.800 ;
        RECT 579.000 255.400 582.600 255.800 ;
        RECT 583.600 255.000 584.400 259.800 ;
        RECT 588.000 258.400 588.800 259.800 ;
        RECT 586.800 257.800 588.800 258.400 ;
        RECT 592.400 257.800 593.200 259.800 ;
        RECT 596.600 258.400 597.800 259.800 ;
        RECT 596.400 257.800 597.800 258.400 ;
        RECT 586.800 257.000 587.600 257.800 ;
        RECT 592.400 257.200 593.000 257.800 ;
        RECT 588.400 255.600 589.200 257.200 ;
        RECT 590.200 256.600 593.000 257.200 ;
        RECT 596.400 257.000 597.200 257.800 ;
        RECT 590.200 256.400 591.000 256.600 ;
        RECT 581.200 254.400 582.000 254.800 ;
        RECT 562.800 254.200 564.400 254.400 ;
        RECT 553.400 253.600 564.400 254.200 ;
        RECT 566.000 253.800 567.600 254.400 ;
        RECT 569.000 254.300 571.600 254.400 ;
        RECT 575.600 254.300 576.400 254.400 ;
        RECT 566.000 253.600 566.800 253.800 ;
        RECT 569.000 253.700 576.400 254.300 ;
        RECT 569.000 253.600 571.600 253.700 ;
        RECT 575.600 253.600 576.400 253.700 ;
        RECT 577.200 253.600 579.800 254.400 ;
        RECT 581.200 253.800 582.800 254.400 ;
        RECT 582.000 253.600 582.800 253.800 ;
        RECT 584.400 254.200 586.000 254.400 ;
        RECT 588.600 254.200 589.200 255.600 ;
        RECT 598.200 255.400 599.000 255.600 ;
        RECT 601.200 255.400 602.000 259.800 ;
        RECT 598.200 254.800 602.000 255.400 ;
        RECT 594.200 254.200 595.000 254.400 ;
        RECT 584.400 253.600 595.400 254.200 ;
        RECT 551.600 252.800 552.400 253.000 ;
        RECT 548.600 252.200 552.400 252.800 ;
        RECT 548.600 252.000 549.400 252.200 ;
        RECT 550.200 251.400 551.000 251.600 ;
        RECT 546.800 250.800 551.000 251.400 ;
        RECT 540.400 242.200 541.200 246.800 ;
        RECT 543.600 242.200 544.400 250.000 ;
        RECT 546.800 242.200 547.600 250.800 ;
        RECT 553.400 250.400 554.000 253.600 ;
        RECT 560.600 253.400 561.400 253.600 ;
        RECT 562.200 252.400 563.000 252.600 ;
        RECT 558.000 251.800 563.000 252.400 ;
        RECT 558.000 251.600 558.800 251.800 ;
        RECT 567.600 251.600 568.400 253.200 ;
        RECT 559.600 251.000 565.200 251.200 ;
        RECT 559.400 250.800 565.200 251.000 ;
        RECT 551.600 249.800 554.000 250.400 ;
        RECT 555.400 250.600 565.200 250.800 ;
        RECT 555.400 250.200 560.200 250.600 ;
        RECT 551.600 248.800 552.200 249.800 ;
        RECT 550.800 248.000 552.200 248.800 ;
        RECT 553.800 249.000 554.600 249.200 ;
        RECT 555.400 249.000 556.000 250.200 ;
        RECT 553.800 248.400 556.000 249.000 ;
        RECT 556.600 249.000 562.000 249.600 ;
        RECT 556.600 248.800 557.400 249.000 ;
        RECT 561.200 248.800 562.000 249.000 ;
        RECT 555.000 247.400 555.800 247.600 ;
        RECT 557.800 247.400 558.600 247.600 ;
        RECT 551.600 246.200 552.400 247.000 ;
        RECT 555.000 246.800 558.600 247.400 ;
        RECT 555.800 246.200 556.400 246.800 ;
        RECT 561.200 246.200 562.000 247.000 ;
        RECT 551.000 242.200 552.200 246.200 ;
        RECT 555.600 242.200 556.400 246.200 ;
        RECT 560.000 245.600 562.000 246.200 ;
        RECT 560.000 242.200 560.800 245.600 ;
        RECT 564.400 242.200 565.200 250.600 ;
        RECT 569.000 250.200 569.600 253.600 ;
        RECT 579.200 252.300 579.800 253.600 ;
        RECT 587.400 253.400 588.200 253.600 ;
        RECT 570.900 251.700 579.800 252.300 ;
        RECT 570.900 250.400 571.500 251.700 ;
        RECT 570.800 250.200 571.600 250.400 ;
        RECT 568.600 249.600 569.600 250.200 ;
        RECT 570.200 249.600 571.600 250.200 ;
        RECT 577.200 250.200 578.000 250.400 ;
        RECT 579.200 250.200 579.800 251.700 ;
        RECT 580.400 251.600 581.200 253.200 ;
        RECT 585.800 252.400 586.600 252.600 ;
        RECT 588.400 252.400 589.200 252.600 ;
        RECT 585.800 251.800 590.800 252.400 ;
        RECT 590.000 251.600 590.800 251.800 ;
        RECT 583.600 251.000 589.200 251.200 ;
        RECT 583.600 250.800 589.400 251.000 ;
        RECT 583.600 250.600 593.400 250.800 ;
        RECT 577.200 249.600 578.600 250.200 ;
        RECT 579.200 249.600 580.200 250.200 ;
        RECT 568.600 242.200 569.400 249.600 ;
        RECT 570.200 248.400 570.800 249.600 ;
        RECT 570.000 247.600 570.800 248.400 ;
        RECT 578.000 248.400 578.600 249.600 ;
        RECT 578.000 247.600 578.800 248.400 ;
        RECT 579.400 242.200 580.200 249.600 ;
        RECT 583.600 242.200 584.400 250.600 ;
        RECT 588.600 250.200 593.400 250.600 ;
        RECT 586.800 249.000 592.200 249.600 ;
        RECT 586.800 248.800 587.600 249.000 ;
        RECT 591.400 248.800 592.200 249.000 ;
        RECT 592.800 249.000 593.400 250.200 ;
        RECT 594.800 250.400 595.400 253.600 ;
        RECT 596.400 252.800 597.200 253.000 ;
        RECT 596.400 252.200 600.200 252.800 ;
        RECT 599.400 252.000 600.200 252.200 ;
        RECT 597.800 251.400 598.600 251.600 ;
        RECT 601.200 251.400 602.000 254.800 ;
        RECT 597.800 250.800 602.000 251.400 ;
        RECT 594.800 249.800 597.200 250.400 ;
        RECT 594.200 249.000 595.000 249.200 ;
        RECT 592.800 248.400 595.000 249.000 ;
        RECT 596.600 248.800 597.200 249.800 ;
        RECT 596.600 248.000 598.000 248.800 ;
        RECT 590.200 247.400 591.000 247.600 ;
        RECT 593.000 247.400 593.800 247.600 ;
        RECT 586.800 246.200 587.600 247.000 ;
        RECT 590.200 246.800 593.800 247.400 ;
        RECT 592.400 246.200 593.000 246.800 ;
        RECT 596.400 246.200 597.200 247.000 ;
        RECT 586.800 245.600 588.800 246.200 ;
        RECT 588.000 242.200 588.800 245.600 ;
        RECT 592.400 242.200 593.200 246.200 ;
        RECT 596.600 242.200 597.800 246.200 ;
        RECT 601.200 242.200 602.000 250.800 ;
        RECT 602.800 255.400 603.600 259.800 ;
        RECT 607.000 258.400 608.200 259.800 ;
        RECT 607.000 257.800 608.400 258.400 ;
        RECT 611.600 257.800 612.400 259.800 ;
        RECT 616.000 258.400 616.800 259.800 ;
        RECT 616.000 257.800 618.000 258.400 ;
        RECT 607.600 257.000 608.400 257.800 ;
        RECT 611.800 257.200 612.400 257.800 ;
        RECT 611.800 256.600 614.600 257.200 ;
        RECT 613.800 256.400 614.600 256.600 ;
        RECT 615.600 256.400 616.400 257.200 ;
        RECT 617.200 257.000 618.000 257.800 ;
        RECT 605.800 255.400 606.600 255.600 ;
        RECT 602.800 254.800 606.600 255.400 ;
        RECT 602.800 251.400 603.600 254.800 ;
        RECT 609.800 254.200 610.600 254.400 ;
        RECT 615.600 254.200 616.200 256.400 ;
        RECT 620.400 255.000 621.200 259.800 ;
        RECT 622.000 255.400 622.800 259.800 ;
        RECT 626.200 258.400 627.400 259.800 ;
        RECT 626.200 257.800 627.600 258.400 ;
        RECT 630.800 257.800 631.600 259.800 ;
        RECT 635.200 258.400 636.000 259.800 ;
        RECT 635.200 257.800 637.200 258.400 ;
        RECT 626.800 257.000 627.600 257.800 ;
        RECT 631.000 257.200 631.600 257.800 ;
        RECT 631.000 256.600 633.800 257.200 ;
        RECT 633.000 256.400 633.800 256.600 ;
        RECT 634.800 256.400 635.600 257.200 ;
        RECT 636.400 257.000 637.200 257.800 ;
        RECT 625.000 255.400 625.800 255.600 ;
        RECT 622.000 254.800 625.800 255.400 ;
        RECT 618.800 254.200 620.400 254.400 ;
        RECT 609.400 253.600 620.400 254.200 ;
        RECT 607.600 252.800 608.400 253.000 ;
        RECT 604.600 252.200 608.400 252.800 ;
        RECT 604.600 252.000 605.400 252.200 ;
        RECT 606.200 251.400 607.000 251.600 ;
        RECT 602.800 250.800 607.000 251.400 ;
        RECT 602.800 242.200 603.600 250.800 ;
        RECT 609.400 250.400 610.000 253.600 ;
        RECT 616.600 253.400 617.400 253.600 ;
        RECT 618.200 252.400 619.000 252.600 ;
        RECT 612.400 252.300 613.200 252.400 ;
        RECT 614.000 252.300 619.000 252.400 ;
        RECT 612.400 251.800 619.000 252.300 ;
        RECT 612.400 251.700 614.800 251.800 ;
        RECT 612.400 251.600 613.200 251.700 ;
        RECT 614.000 251.600 614.800 251.700 ;
        RECT 622.000 251.400 622.800 254.800 ;
        RECT 629.000 254.200 629.800 254.400 ;
        RECT 634.800 254.200 635.400 256.400 ;
        RECT 639.600 255.000 640.400 259.800 ;
        RECT 641.200 255.800 642.000 259.800 ;
        RECT 642.800 256.000 643.600 259.800 ;
        RECT 646.000 256.000 646.800 259.800 ;
        RECT 642.800 255.800 646.800 256.000 ;
        RECT 647.600 255.800 648.400 259.800 ;
        RECT 649.200 256.000 650.000 259.800 ;
        RECT 652.400 256.000 653.200 259.800 ;
        RECT 657.800 256.000 658.600 259.000 ;
        RECT 662.000 257.000 662.800 259.000 ;
        RECT 649.200 255.800 653.200 256.000 ;
        RECT 641.400 254.400 642.000 255.800 ;
        RECT 643.000 255.400 646.600 255.800 ;
        RECT 645.200 254.400 646.000 254.800 ;
        RECT 647.800 254.400 648.400 255.800 ;
        RECT 649.400 255.400 653.000 255.800 ;
        RECT 657.000 255.400 658.600 256.000 ;
        RECT 657.000 255.000 657.800 255.400 ;
        RECT 651.600 254.400 652.400 254.800 ;
        RECT 657.000 254.400 657.600 255.000 ;
        RECT 662.200 254.800 662.800 257.000 ;
        RECT 663.600 256.000 664.400 259.800 ;
        RECT 666.800 256.000 667.600 259.800 ;
        RECT 663.600 255.800 667.600 256.000 ;
        RECT 668.400 255.800 669.200 259.800 ;
        RECT 663.800 255.400 667.400 255.800 ;
        RECT 638.000 254.200 639.600 254.400 ;
        RECT 628.600 253.600 639.600 254.200 ;
        RECT 641.200 253.600 643.800 254.400 ;
        RECT 645.200 253.800 646.800 254.400 ;
        RECT 646.000 253.600 646.800 253.800 ;
        RECT 647.600 253.600 650.200 254.400 ;
        RECT 651.600 253.800 653.200 254.400 ;
        RECT 652.400 253.600 653.200 253.800 ;
        RECT 655.600 253.600 657.600 254.400 ;
        RECT 658.600 254.200 662.800 254.800 ;
        RECT 664.400 254.400 665.200 254.800 ;
        RECT 668.400 254.400 669.000 255.800 ;
        RECT 670.000 255.000 670.800 259.800 ;
        RECT 674.400 258.400 675.200 259.800 ;
        RECT 673.200 257.800 675.200 258.400 ;
        RECT 678.800 257.800 679.600 259.800 ;
        RECT 683.000 258.400 684.200 259.800 ;
        RECT 682.800 257.800 684.200 258.400 ;
        RECT 673.200 257.000 674.000 257.800 ;
        RECT 678.800 257.200 679.400 257.800 ;
        RECT 674.800 256.400 675.600 257.200 ;
        RECT 676.600 256.600 679.400 257.200 ;
        RECT 682.800 257.000 683.600 257.800 ;
        RECT 676.600 256.400 677.400 256.600 ;
        RECT 658.600 253.800 659.600 254.200 ;
        RECT 626.800 252.800 627.600 253.000 ;
        RECT 623.800 252.200 627.600 252.800 ;
        RECT 628.600 252.400 629.200 253.600 ;
        RECT 635.800 253.400 636.600 253.600 ;
        RECT 637.400 252.400 638.200 252.600 ;
        RECT 623.800 252.000 624.600 252.200 ;
        RECT 628.400 251.600 629.200 252.400 ;
        RECT 633.200 251.800 638.200 252.400 ;
        RECT 633.200 251.600 634.000 251.800 ;
        RECT 625.400 251.400 626.200 251.600 ;
        RECT 615.600 251.000 621.200 251.200 ;
        RECT 615.400 250.800 621.200 251.000 ;
        RECT 607.600 249.800 610.000 250.400 ;
        RECT 611.400 250.600 621.200 250.800 ;
        RECT 611.400 250.200 616.200 250.600 ;
        RECT 607.600 248.800 608.200 249.800 ;
        RECT 606.800 248.000 608.200 248.800 ;
        RECT 609.800 249.000 610.600 249.200 ;
        RECT 611.400 249.000 612.000 250.200 ;
        RECT 609.800 248.400 612.000 249.000 ;
        RECT 612.600 249.000 618.000 249.600 ;
        RECT 612.600 248.800 613.400 249.000 ;
        RECT 617.200 248.800 618.000 249.000 ;
        RECT 611.000 247.400 611.800 247.600 ;
        RECT 613.800 247.400 614.600 247.600 ;
        RECT 607.600 246.200 608.400 247.000 ;
        RECT 611.000 246.800 614.600 247.400 ;
        RECT 611.800 246.200 612.400 246.800 ;
        RECT 617.200 246.200 618.000 247.000 ;
        RECT 607.000 242.200 608.200 246.200 ;
        RECT 611.600 242.200 612.400 246.200 ;
        RECT 616.000 245.600 618.000 246.200 ;
        RECT 616.000 242.200 616.800 245.600 ;
        RECT 620.400 242.200 621.200 250.600 ;
        RECT 622.000 250.800 626.200 251.400 ;
        RECT 622.000 242.200 622.800 250.800 ;
        RECT 628.600 250.400 629.200 251.600 ;
        RECT 634.800 251.000 640.400 251.200 ;
        RECT 634.600 250.800 640.400 251.000 ;
        RECT 626.800 249.800 629.200 250.400 ;
        RECT 630.600 250.600 640.400 250.800 ;
        RECT 630.600 250.200 635.400 250.600 ;
        RECT 626.800 248.800 627.400 249.800 ;
        RECT 626.000 248.000 627.400 248.800 ;
        RECT 629.000 249.000 629.800 249.200 ;
        RECT 630.600 249.000 631.200 250.200 ;
        RECT 629.000 248.400 631.200 249.000 ;
        RECT 631.800 249.000 637.200 249.600 ;
        RECT 631.800 248.800 632.600 249.000 ;
        RECT 636.400 248.800 637.200 249.000 ;
        RECT 630.200 247.400 631.000 247.600 ;
        RECT 633.000 247.400 633.800 247.600 ;
        RECT 626.800 246.200 627.600 247.000 ;
        RECT 630.200 246.800 633.800 247.400 ;
        RECT 631.000 246.200 631.600 246.800 ;
        RECT 636.400 246.200 637.200 247.000 ;
        RECT 626.200 242.200 627.400 246.200 ;
        RECT 630.800 242.200 631.600 246.200 ;
        RECT 635.200 245.600 637.200 246.200 ;
        RECT 635.200 242.200 636.000 245.600 ;
        RECT 639.600 242.200 640.400 250.600 ;
        RECT 641.200 250.200 642.000 250.400 ;
        RECT 643.200 250.200 643.800 253.600 ;
        RECT 644.400 251.600 645.200 253.200 ;
        RECT 646.000 252.300 646.800 252.400 ;
        RECT 649.600 252.300 650.200 253.600 ;
        RECT 646.000 251.700 650.200 252.300 ;
        RECT 646.000 251.600 646.800 251.700 ;
        RECT 647.600 250.200 648.400 250.400 ;
        RECT 649.600 250.200 650.200 251.700 ;
        RECT 650.800 252.300 651.600 253.200 ;
        RECT 657.000 252.400 657.600 253.600 ;
        RECT 658.200 253.000 659.600 253.800 ;
        RECT 663.600 253.800 665.200 254.400 ;
        RECT 663.600 253.600 664.400 253.800 ;
        RECT 666.600 253.600 669.200 254.400 ;
        RECT 670.800 254.200 672.400 254.400 ;
        RECT 675.000 254.200 675.600 256.400 ;
        RECT 684.600 255.400 685.400 255.600 ;
        RECT 687.600 255.400 688.400 259.800 ;
        RECT 684.600 254.800 688.400 255.400 ;
        RECT 680.600 254.200 681.400 254.400 ;
        RECT 670.800 253.600 681.800 254.200 ;
        RECT 652.400 252.300 653.200 252.400 ;
        RECT 650.800 251.700 653.200 252.300 ;
        RECT 650.800 251.600 651.600 251.700 ;
        RECT 652.400 251.600 653.200 251.700 ;
        RECT 655.600 250.800 656.400 252.400 ;
        RECT 657.000 251.600 658.000 252.400 ;
        RECT 641.200 249.600 642.600 250.200 ;
        RECT 643.200 249.600 644.200 250.200 ;
        RECT 647.600 249.600 649.000 250.200 ;
        RECT 649.600 249.600 650.600 250.200 ;
        RECT 642.000 248.400 642.600 249.600 ;
        RECT 643.400 248.400 644.200 249.600 ;
        RECT 648.400 248.400 649.000 249.600 ;
        RECT 642.000 247.600 642.800 248.400 ;
        RECT 643.400 247.600 645.200 248.400 ;
        RECT 648.400 247.600 649.200 248.400 ;
        RECT 643.400 242.200 644.200 247.600 ;
        RECT 649.800 242.200 650.600 249.600 ;
        RECT 657.000 249.800 657.600 251.600 ;
        RECT 659.000 251.000 659.600 253.000 ;
        RECT 660.400 251.600 661.200 253.200 ;
        RECT 662.000 251.600 662.800 253.200 ;
        RECT 665.200 251.600 666.000 253.200 ;
        RECT 666.600 252.300 667.200 253.600 ;
        RECT 673.800 253.400 674.600 253.600 ;
        RECT 672.200 252.400 673.000 252.600 ;
        RECT 674.800 252.400 675.600 252.600 ;
        RECT 668.400 252.300 669.200 252.400 ;
        RECT 666.600 251.700 669.200 252.300 ;
        RECT 672.200 251.800 677.200 252.400 ;
        RECT 659.000 250.400 662.800 251.000 ;
        RECT 657.000 249.200 658.600 249.800 ;
        RECT 657.800 242.200 658.600 249.200 ;
        RECT 662.200 247.000 662.800 250.400 ;
        RECT 666.600 250.200 667.200 251.700 ;
        RECT 668.400 251.600 669.200 251.700 ;
        RECT 676.400 251.600 677.200 251.800 ;
        RECT 670.000 251.000 675.600 251.200 ;
        RECT 670.000 250.800 675.800 251.000 ;
        RECT 670.000 250.600 679.800 250.800 ;
        RECT 668.400 250.200 669.200 250.400 ;
        RECT 662.000 243.000 662.800 247.000 ;
        RECT 666.200 249.600 667.200 250.200 ;
        RECT 667.800 249.600 669.200 250.200 ;
        RECT 666.200 242.200 667.000 249.600 ;
        RECT 667.800 248.400 668.400 249.600 ;
        RECT 667.600 247.600 668.400 248.400 ;
        RECT 670.000 242.200 670.800 250.600 ;
        RECT 675.000 250.200 679.800 250.600 ;
        RECT 673.200 249.000 678.600 249.600 ;
        RECT 673.200 248.800 674.000 249.000 ;
        RECT 677.800 248.800 678.600 249.000 ;
        RECT 679.200 249.000 679.800 250.200 ;
        RECT 681.200 250.400 681.800 253.600 ;
        RECT 682.800 252.800 683.600 253.000 ;
        RECT 682.800 252.200 686.600 252.800 ;
        RECT 685.800 252.000 686.600 252.200 ;
        RECT 684.200 251.400 685.000 251.600 ;
        RECT 687.600 251.400 688.400 254.800 ;
        RECT 684.200 250.800 688.400 251.400 ;
        RECT 681.200 249.800 683.600 250.400 ;
        RECT 680.600 249.000 681.400 249.200 ;
        RECT 679.200 248.400 681.400 249.000 ;
        RECT 683.000 248.800 683.600 249.800 ;
        RECT 683.000 248.000 684.400 248.800 ;
        RECT 676.600 247.400 677.400 247.600 ;
        RECT 679.400 247.400 680.200 247.600 ;
        RECT 673.200 246.200 674.000 247.000 ;
        RECT 676.600 246.800 680.200 247.400 ;
        RECT 678.800 246.200 679.400 246.800 ;
        RECT 682.800 246.200 683.600 247.000 ;
        RECT 673.200 245.600 675.200 246.200 ;
        RECT 674.400 242.200 675.200 245.600 ;
        RECT 678.800 242.200 679.600 246.200 ;
        RECT 683.000 242.200 684.200 246.200 ;
        RECT 687.600 242.200 688.400 250.800 ;
        RECT 2.800 231.200 3.600 239.800 ;
        RECT 6.000 231.200 6.800 239.800 ;
        RECT 9.200 231.200 10.000 239.800 ;
        RECT 12.400 231.200 13.200 239.800 ;
        RECT 1.200 230.400 3.600 231.200 ;
        RECT 4.600 230.400 6.800 231.200 ;
        RECT 7.800 230.400 10.000 231.200 ;
        RECT 11.400 230.400 13.200 231.200 ;
        RECT 1.200 227.600 2.000 230.400 ;
        RECT 4.600 229.000 5.400 230.400 ;
        RECT 7.800 229.000 8.600 230.400 ;
        RECT 11.400 229.000 12.200 230.400 ;
        RECT 15.600 230.300 16.400 239.800 ;
        RECT 18.800 230.300 19.600 230.400 ;
        RECT 15.600 229.700 19.600 230.300 ;
        RECT 2.800 228.200 5.400 229.000 ;
        RECT 6.200 228.200 8.600 229.000 ;
        RECT 9.600 228.200 12.200 229.000 ;
        RECT 13.000 228.200 14.800 229.000 ;
        RECT 4.600 227.600 5.400 228.200 ;
        RECT 7.800 227.600 8.600 228.200 ;
        RECT 11.400 227.600 12.200 228.200 ;
        RECT 14.000 227.600 14.800 228.200 ;
        RECT 1.200 226.800 3.600 227.600 ;
        RECT 4.600 226.800 6.800 227.600 ;
        RECT 7.800 226.800 10.000 227.600 ;
        RECT 11.400 226.800 13.200 227.600 ;
        RECT 2.800 222.200 3.600 226.800 ;
        RECT 6.000 222.200 6.800 226.800 ;
        RECT 9.200 222.200 10.000 226.800 ;
        RECT 12.400 222.200 13.200 226.800 ;
        RECT 15.600 222.200 16.400 229.700 ;
        RECT 18.800 229.600 19.600 229.700 ;
        RECT 17.200 226.300 18.000 226.400 ;
        RECT 18.800 226.300 19.600 226.400 ;
        RECT 17.200 225.700 19.600 226.300 ;
        RECT 17.200 224.800 18.000 225.700 ;
        RECT 18.800 224.800 19.600 225.700 ;
        RECT 20.400 222.200 21.200 239.800 ;
        RECT 23.600 232.000 24.400 239.800 ;
        RECT 26.800 235.200 27.600 239.800 ;
        RECT 23.400 231.200 24.400 232.000 ;
        RECT 25.000 234.600 27.600 235.200 ;
        RECT 25.000 233.000 25.600 234.600 ;
        RECT 30.000 234.400 30.800 239.800 ;
        RECT 33.200 237.000 34.000 239.800 ;
        RECT 34.800 237.000 35.600 239.800 ;
        RECT 36.400 237.000 37.200 239.800 ;
        RECT 31.400 234.400 35.600 235.200 ;
        RECT 28.200 233.600 30.800 234.400 ;
        RECT 38.000 233.600 38.800 239.800 ;
        RECT 41.200 235.000 42.000 239.800 ;
        RECT 44.400 235.000 45.200 239.800 ;
        RECT 46.000 237.000 46.800 239.800 ;
        RECT 47.600 237.000 48.400 239.800 ;
        RECT 50.800 235.200 51.600 239.800 ;
        RECT 54.000 236.400 54.800 239.800 ;
        RECT 54.000 235.800 55.000 236.400 ;
        RECT 54.400 235.200 55.000 235.800 ;
        RECT 49.600 234.400 53.800 235.200 ;
        RECT 54.400 234.600 56.400 235.200 ;
        RECT 41.200 233.600 43.800 234.400 ;
        RECT 44.400 233.800 50.200 234.400 ;
        RECT 53.200 234.000 53.800 234.400 ;
        RECT 33.200 233.000 34.000 233.200 ;
        RECT 25.000 232.400 34.000 233.000 ;
        RECT 36.400 233.000 37.200 233.200 ;
        RECT 44.400 233.000 45.000 233.800 ;
        RECT 50.800 233.200 52.200 233.800 ;
        RECT 53.200 233.200 54.800 234.000 ;
        RECT 36.400 232.400 45.000 233.000 ;
        RECT 46.000 233.000 52.200 233.200 ;
        RECT 46.000 232.600 51.400 233.000 ;
        RECT 46.000 232.400 46.800 232.600 ;
        RECT 23.400 226.800 24.200 231.200 ;
        RECT 25.000 230.600 25.600 232.400 ;
        RECT 24.800 230.000 25.600 230.600 ;
        RECT 31.600 230.000 55.000 230.600 ;
        RECT 24.800 228.000 25.400 230.000 ;
        RECT 31.600 229.400 32.400 230.000 ;
        RECT 49.200 229.600 50.000 230.000 ;
        RECT 52.400 229.600 53.200 230.000 ;
        RECT 54.200 229.800 55.000 230.000 ;
        RECT 26.000 228.600 29.800 229.400 ;
        RECT 24.800 227.400 26.000 228.000 ;
        RECT 23.400 226.000 24.400 226.800 ;
        RECT 23.600 222.200 24.400 226.000 ;
        RECT 25.200 222.200 26.000 227.400 ;
        RECT 29.000 227.400 29.800 228.600 ;
        RECT 29.000 226.800 30.800 227.400 ;
        RECT 30.000 226.200 30.800 226.800 ;
        RECT 34.800 226.400 35.600 229.200 ;
        RECT 38.000 228.600 41.200 229.400 ;
        RECT 45.000 228.600 47.000 229.400 ;
        RECT 55.600 229.000 56.400 234.600 ;
        RECT 61.000 232.800 61.800 239.800 ;
        RECT 65.200 235.000 66.000 239.000 ;
        RECT 60.200 232.200 61.800 232.800 ;
        RECT 58.800 229.600 59.600 231.200 ;
        RECT 37.600 227.800 38.400 228.000 ;
        RECT 37.600 227.200 42.000 227.800 ;
        RECT 41.200 227.000 42.000 227.200 ;
        RECT 42.800 226.800 43.600 228.400 ;
        RECT 30.000 225.400 32.400 226.200 ;
        RECT 34.800 225.600 35.800 226.400 ;
        RECT 38.800 225.600 40.400 226.400 ;
        RECT 41.200 226.200 42.000 226.400 ;
        RECT 45.000 226.200 45.800 228.600 ;
        RECT 47.600 228.200 56.400 229.000 ;
        RECT 60.200 228.400 60.800 232.200 ;
        RECT 65.400 231.600 66.000 235.000 ;
        RECT 69.400 232.600 70.200 239.800 ;
        RECT 68.400 231.800 70.200 232.600 ;
        RECT 71.600 231.800 72.400 239.800 ;
        RECT 73.200 232.400 74.000 239.800 ;
        RECT 76.400 232.400 77.200 239.800 ;
        RECT 73.200 231.800 77.200 232.400 ;
        RECT 78.000 235.000 78.800 239.000 ;
        RECT 82.200 238.400 83.000 239.800 ;
        RECT 82.200 237.600 83.600 238.400 ;
        RECT 62.200 231.000 66.000 231.600 ;
        RECT 62.200 229.000 62.800 231.000 ;
        RECT 51.000 226.800 54.000 227.600 ;
        RECT 51.000 226.200 51.800 226.800 ;
        RECT 41.200 225.600 45.800 226.200 ;
        RECT 31.600 222.200 32.400 225.400 ;
        RECT 49.200 225.400 51.800 226.200 ;
        RECT 33.200 222.200 34.000 225.000 ;
        RECT 34.800 222.200 35.600 225.000 ;
        RECT 36.400 222.200 37.200 225.000 ;
        RECT 38.000 222.200 38.800 225.000 ;
        RECT 41.200 222.200 42.000 225.000 ;
        RECT 44.400 222.200 45.200 225.000 ;
        RECT 46.000 222.200 46.800 225.000 ;
        RECT 47.600 222.200 48.400 225.000 ;
        RECT 49.200 222.200 50.000 225.400 ;
        RECT 55.600 222.200 56.400 228.200 ;
        RECT 57.200 228.300 58.000 228.400 ;
        RECT 58.800 228.300 60.800 228.400 ;
        RECT 57.200 227.700 60.800 228.300 ;
        RECT 61.400 228.200 62.800 229.000 ;
        RECT 63.600 228.800 64.400 230.400 ;
        RECT 65.200 228.800 66.000 230.400 ;
        RECT 68.600 228.400 69.200 231.800 ;
        RECT 70.000 229.600 70.800 231.200 ;
        RECT 71.800 230.400 72.400 231.800 ;
        RECT 78.000 231.600 78.600 235.000 ;
        RECT 82.200 232.800 83.000 237.600 ;
        RECT 89.200 236.400 90.000 239.800 ;
        RECT 89.000 235.800 90.000 236.400 ;
        RECT 89.000 235.200 89.600 235.800 ;
        RECT 92.400 235.200 93.200 239.800 ;
        RECT 95.600 237.000 96.400 239.800 ;
        RECT 97.200 237.000 98.000 239.800 ;
        RECT 87.600 234.600 89.600 235.200 ;
        RECT 82.200 232.200 83.800 232.800 ;
        RECT 78.000 231.000 81.800 231.600 ;
        RECT 75.600 230.400 76.400 230.800 ;
        RECT 71.600 229.800 74.000 230.400 ;
        RECT 75.600 229.800 77.200 230.400 ;
        RECT 71.600 229.600 72.400 229.800 ;
        RECT 57.200 227.600 58.000 227.700 ;
        RECT 58.800 227.600 60.800 227.700 ;
        RECT 60.200 227.000 60.800 227.600 ;
        RECT 61.800 227.800 62.800 228.200 ;
        RECT 61.800 227.200 66.000 227.800 ;
        RECT 68.400 227.600 69.200 228.400 ;
        RECT 60.200 226.600 61.000 227.000 ;
        RECT 60.200 226.000 61.800 226.600 ;
        RECT 61.000 223.000 61.800 226.000 ;
        RECT 65.400 225.000 66.000 227.200 ;
        RECT 65.200 223.000 66.000 225.000 ;
        RECT 66.800 224.800 67.600 226.400 ;
        RECT 68.600 226.300 69.200 227.600 ;
        RECT 71.600 226.300 72.400 226.400 ;
        RECT 68.500 225.700 72.400 226.300 ;
        RECT 73.400 226.200 74.000 229.800 ;
        RECT 76.400 229.600 77.200 229.800 ;
        RECT 74.800 227.600 75.600 229.200 ;
        RECT 78.000 228.800 78.800 230.400 ;
        RECT 79.600 228.800 80.400 230.400 ;
        RECT 81.200 229.000 81.800 231.000 ;
        RECT 81.200 228.200 82.600 229.000 ;
        RECT 83.200 228.400 83.800 232.200 ;
        RECT 84.400 229.600 85.200 231.200 ;
        RECT 87.600 229.000 88.400 234.600 ;
        RECT 90.200 234.400 94.400 235.200 ;
        RECT 98.800 235.000 99.600 239.800 ;
        RECT 102.000 235.000 102.800 239.800 ;
        RECT 90.200 234.000 90.800 234.400 ;
        RECT 89.200 233.200 90.800 234.000 ;
        RECT 93.800 233.800 99.600 234.400 ;
        RECT 91.800 233.200 93.200 233.800 ;
        RECT 91.800 233.000 98.000 233.200 ;
        RECT 92.600 232.600 98.000 233.000 ;
        RECT 97.200 232.400 98.000 232.600 ;
        RECT 99.000 233.000 99.600 233.800 ;
        RECT 100.200 233.600 102.800 234.400 ;
        RECT 105.200 233.600 106.000 239.800 ;
        RECT 106.800 237.000 107.600 239.800 ;
        RECT 108.400 237.000 109.200 239.800 ;
        RECT 110.000 237.000 110.800 239.800 ;
        RECT 108.400 234.400 112.600 235.200 ;
        RECT 113.200 234.400 114.000 239.800 ;
        RECT 116.400 235.200 117.200 239.800 ;
        RECT 116.400 234.600 119.000 235.200 ;
        RECT 113.200 233.600 115.800 234.400 ;
        RECT 106.800 233.000 107.600 233.200 ;
        RECT 99.000 232.400 107.600 233.000 ;
        RECT 110.000 233.000 110.800 233.200 ;
        RECT 118.400 233.000 119.000 234.600 ;
        RECT 110.000 232.400 119.000 233.000 ;
        RECT 118.400 230.600 119.000 232.400 ;
        RECT 119.600 232.000 120.400 239.800 ;
        RECT 128.200 232.600 129.000 239.800 ;
        RECT 119.600 231.200 120.600 232.000 ;
        RECT 128.200 231.800 130.000 232.600 ;
        RECT 132.400 231.800 133.200 239.800 ;
        RECT 134.000 232.400 134.800 239.800 ;
        RECT 137.200 232.400 138.000 239.800 ;
        RECT 134.000 231.800 138.000 232.400 ;
        RECT 140.400 232.000 141.200 239.800 ;
        RECT 143.600 235.200 144.400 239.800 ;
        RECT 89.000 230.000 112.400 230.600 ;
        RECT 118.400 230.000 119.200 230.600 ;
        RECT 89.000 229.800 89.800 230.000 ;
        RECT 90.800 229.600 91.600 230.000 ;
        RECT 94.000 229.600 94.800 230.000 ;
        RECT 111.600 229.400 112.400 230.000 ;
        RECT 81.200 227.800 82.200 228.200 ;
        RECT 68.600 224.200 69.200 225.700 ;
        RECT 71.600 225.600 72.400 225.700 ;
        RECT 71.800 224.800 72.600 225.600 ;
        RECT 68.400 222.200 69.200 224.200 ;
        RECT 73.200 222.200 74.000 226.200 ;
        RECT 78.000 227.200 82.200 227.800 ;
        RECT 83.200 227.600 85.200 228.400 ;
        RECT 87.600 228.200 96.400 229.000 ;
        RECT 97.000 228.600 99.000 229.400 ;
        RECT 102.800 228.600 106.000 229.400 ;
        RECT 78.000 225.000 78.600 227.200 ;
        RECT 83.200 227.000 83.800 227.600 ;
        RECT 83.000 226.600 83.800 227.000 ;
        RECT 82.200 226.000 83.800 226.600 ;
        RECT 78.000 223.000 78.800 225.000 ;
        RECT 82.200 223.000 83.000 226.000 ;
        RECT 87.600 222.200 88.400 228.200 ;
        RECT 90.000 226.800 93.000 227.600 ;
        RECT 92.200 226.200 93.000 226.800 ;
        RECT 98.200 226.200 99.000 228.600 ;
        RECT 100.400 226.800 101.200 228.400 ;
        RECT 105.600 227.800 106.400 228.000 ;
        RECT 102.000 227.200 106.400 227.800 ;
        RECT 102.000 227.000 102.800 227.200 ;
        RECT 108.400 226.400 109.200 229.200 ;
        RECT 114.200 228.600 118.000 229.400 ;
        RECT 114.200 227.400 115.000 228.600 ;
        RECT 118.600 228.000 119.200 230.000 ;
        RECT 102.000 226.200 102.800 226.400 ;
        RECT 92.200 225.400 94.800 226.200 ;
        RECT 98.200 225.600 102.800 226.200 ;
        RECT 103.600 225.600 105.200 226.400 ;
        RECT 108.200 225.600 109.200 226.400 ;
        RECT 113.200 226.800 115.000 227.400 ;
        RECT 118.000 227.400 119.200 228.000 ;
        RECT 113.200 226.200 114.000 226.800 ;
        RECT 94.000 222.200 94.800 225.400 ;
        RECT 111.600 225.400 114.000 226.200 ;
        RECT 95.600 222.200 96.400 225.000 ;
        RECT 97.200 222.200 98.000 225.000 ;
        RECT 98.800 222.200 99.600 225.000 ;
        RECT 102.000 222.200 102.800 225.000 ;
        RECT 105.200 222.200 106.000 225.000 ;
        RECT 106.800 222.200 107.600 225.000 ;
        RECT 108.400 222.200 109.200 225.000 ;
        RECT 110.000 222.200 110.800 225.000 ;
        RECT 111.600 222.200 112.400 225.400 ;
        RECT 118.000 222.200 118.800 227.400 ;
        RECT 119.800 226.800 120.600 231.200 ;
        RECT 127.600 229.600 128.400 231.200 ;
        RECT 119.600 226.000 120.600 226.800 ;
        RECT 129.200 228.400 129.800 231.800 ;
        RECT 132.600 230.400 133.200 231.800 ;
        RECT 140.200 231.200 141.200 232.000 ;
        RECT 141.800 234.600 144.400 235.200 ;
        RECT 141.800 233.000 142.400 234.600 ;
        RECT 146.800 234.400 147.600 239.800 ;
        RECT 150.000 237.000 150.800 239.800 ;
        RECT 151.600 237.000 152.400 239.800 ;
        RECT 153.200 237.000 154.000 239.800 ;
        RECT 148.200 234.400 152.400 235.200 ;
        RECT 145.000 233.600 147.600 234.400 ;
        RECT 154.800 233.600 155.600 239.800 ;
        RECT 158.000 235.000 158.800 239.800 ;
        RECT 161.200 235.000 162.000 239.800 ;
        RECT 162.800 237.000 163.600 239.800 ;
        RECT 164.400 237.000 165.200 239.800 ;
        RECT 167.600 235.200 168.400 239.800 ;
        RECT 170.800 236.400 171.600 239.800 ;
        RECT 170.800 235.800 171.800 236.400 ;
        RECT 171.200 235.200 171.800 235.800 ;
        RECT 166.400 234.400 170.600 235.200 ;
        RECT 171.200 234.600 173.200 235.200 ;
        RECT 158.000 233.600 160.600 234.400 ;
        RECT 161.200 233.800 167.000 234.400 ;
        RECT 170.000 234.000 170.600 234.400 ;
        RECT 150.000 233.000 150.800 233.200 ;
        RECT 141.800 232.400 150.800 233.000 ;
        RECT 153.200 233.000 154.000 233.200 ;
        RECT 161.200 233.000 161.800 233.800 ;
        RECT 167.600 233.200 169.000 233.800 ;
        RECT 170.000 233.200 171.600 234.000 ;
        RECT 153.200 232.400 161.800 233.000 ;
        RECT 162.800 233.000 169.000 233.200 ;
        RECT 162.800 232.600 168.200 233.000 ;
        RECT 162.800 232.400 163.600 232.600 ;
        RECT 136.400 230.400 137.200 230.800 ;
        RECT 132.400 229.800 134.800 230.400 ;
        RECT 136.400 229.800 138.000 230.400 ;
        RECT 132.400 229.600 133.200 229.800 ;
        RECT 129.200 228.300 130.000 228.400 ;
        RECT 129.200 227.700 133.100 228.300 ;
        RECT 129.200 227.600 130.000 227.700 ;
        RECT 119.600 222.200 120.400 226.000 ;
        RECT 129.200 224.200 129.800 227.600 ;
        RECT 132.500 226.400 133.100 227.700 ;
        RECT 130.800 224.800 131.600 226.400 ;
        RECT 132.400 225.600 133.200 226.400 ;
        RECT 134.200 226.200 134.800 229.800 ;
        RECT 137.200 229.600 138.000 229.800 ;
        RECT 135.600 227.600 136.400 229.200 ;
        RECT 132.600 224.800 133.400 225.600 ;
        RECT 129.200 222.200 130.000 224.200 ;
        RECT 134.000 222.200 134.800 226.200 ;
        RECT 140.200 226.800 141.000 231.200 ;
        RECT 141.800 230.600 142.400 232.400 ;
        RECT 141.600 230.000 142.400 230.600 ;
        RECT 148.400 230.000 171.800 230.600 ;
        RECT 141.600 228.000 142.200 230.000 ;
        RECT 148.400 229.400 149.200 230.000 ;
        RECT 166.000 229.600 166.800 230.000 ;
        RECT 167.600 229.600 168.400 230.000 ;
        RECT 171.000 229.800 171.800 230.000 ;
        RECT 142.800 228.600 146.600 229.400 ;
        RECT 141.600 227.400 142.800 228.000 ;
        RECT 140.200 226.000 141.200 226.800 ;
        RECT 140.400 222.200 141.200 226.000 ;
        RECT 142.000 222.200 142.800 227.400 ;
        RECT 145.800 227.400 146.600 228.600 ;
        RECT 145.800 226.800 147.600 227.400 ;
        RECT 146.800 226.200 147.600 226.800 ;
        RECT 151.600 226.400 152.400 229.200 ;
        RECT 154.800 228.600 158.000 229.400 ;
        RECT 161.800 228.600 163.800 229.400 ;
        RECT 172.400 229.000 173.200 234.600 ;
        RECT 154.400 227.800 155.200 228.000 ;
        RECT 154.400 227.200 158.800 227.800 ;
        RECT 158.000 227.000 158.800 227.200 ;
        RECT 159.600 226.800 160.400 228.400 ;
        RECT 146.800 225.400 149.200 226.200 ;
        RECT 151.600 225.600 152.600 226.400 ;
        RECT 155.600 225.600 157.200 226.400 ;
        RECT 158.000 226.200 158.800 226.400 ;
        RECT 161.800 226.200 162.600 228.600 ;
        RECT 164.400 228.200 173.200 229.000 ;
        RECT 167.800 226.800 170.800 227.600 ;
        RECT 167.800 226.200 168.600 226.800 ;
        RECT 158.000 225.600 162.600 226.200 ;
        RECT 148.400 222.200 149.200 225.400 ;
        RECT 166.000 225.400 168.600 226.200 ;
        RECT 150.000 222.200 150.800 225.000 ;
        RECT 151.600 222.200 152.400 225.000 ;
        RECT 153.200 222.200 154.000 225.000 ;
        RECT 154.800 222.200 155.600 225.000 ;
        RECT 158.000 222.200 158.800 225.000 ;
        RECT 161.200 222.200 162.000 225.000 ;
        RECT 162.800 222.200 163.600 225.000 ;
        RECT 164.400 222.200 165.200 225.000 ;
        RECT 166.000 222.200 166.800 225.400 ;
        RECT 172.400 222.200 173.200 228.200 ;
        RECT 175.600 230.300 176.400 239.800 ;
        RECT 181.000 232.800 181.800 239.800 ;
        RECT 185.200 235.000 186.000 239.000 ;
        RECT 180.200 232.200 181.800 232.800 ;
        RECT 178.800 230.300 179.600 231.200 ;
        RECT 175.600 229.700 179.600 230.300 ;
        RECT 174.000 224.800 174.800 226.400 ;
        RECT 175.600 222.200 176.400 229.700 ;
        RECT 178.800 229.600 179.600 229.700 ;
        RECT 180.200 228.400 180.800 232.200 ;
        RECT 185.400 231.600 186.000 235.000 ;
        RECT 188.400 232.000 189.200 239.800 ;
        RECT 191.600 235.200 192.400 239.800 ;
        RECT 182.200 231.000 186.000 231.600 ;
        RECT 188.200 231.200 189.200 232.000 ;
        RECT 189.800 234.600 192.400 235.200 ;
        RECT 189.800 233.000 190.400 234.600 ;
        RECT 194.800 234.400 195.600 239.800 ;
        RECT 198.000 237.000 198.800 239.800 ;
        RECT 199.600 237.000 200.400 239.800 ;
        RECT 201.200 237.000 202.000 239.800 ;
        RECT 196.200 234.400 200.400 235.200 ;
        RECT 193.000 233.600 195.600 234.400 ;
        RECT 202.800 233.600 203.600 239.800 ;
        RECT 206.000 235.000 206.800 239.800 ;
        RECT 209.200 235.000 210.000 239.800 ;
        RECT 210.800 237.000 211.600 239.800 ;
        RECT 212.400 237.000 213.200 239.800 ;
        RECT 215.600 235.200 216.400 239.800 ;
        RECT 218.800 236.400 219.600 239.800 ;
        RECT 225.800 238.400 226.600 239.800 ;
        RECT 225.800 237.600 227.600 238.400 ;
        RECT 218.800 235.800 219.800 236.400 ;
        RECT 219.200 235.200 219.800 235.800 ;
        RECT 214.400 234.400 218.600 235.200 ;
        RECT 219.200 234.600 221.200 235.200 ;
        RECT 206.000 233.600 208.600 234.400 ;
        RECT 209.200 233.800 215.000 234.400 ;
        RECT 218.000 234.000 218.600 234.400 ;
        RECT 198.000 233.000 198.800 233.200 ;
        RECT 189.800 232.400 198.800 233.000 ;
        RECT 201.200 233.000 202.000 233.200 ;
        RECT 209.200 233.000 209.800 233.800 ;
        RECT 215.600 233.200 217.000 233.800 ;
        RECT 218.000 233.200 219.600 234.000 ;
        RECT 201.200 232.400 209.800 233.000 ;
        RECT 210.800 233.000 217.000 233.200 ;
        RECT 210.800 232.600 216.200 233.000 ;
        RECT 210.800 232.400 211.600 232.600 ;
        RECT 182.200 229.000 182.800 231.000 ;
        RECT 178.800 227.600 180.800 228.400 ;
        RECT 181.400 228.200 182.800 229.000 ;
        RECT 183.600 228.800 184.400 230.400 ;
        RECT 185.200 228.800 186.000 230.400 ;
        RECT 180.200 227.000 180.800 227.600 ;
        RECT 181.800 227.800 182.800 228.200 ;
        RECT 181.800 227.200 186.000 227.800 ;
        RECT 180.200 226.600 181.000 227.000 ;
        RECT 180.200 226.000 181.800 226.600 ;
        RECT 181.000 224.400 181.800 226.000 ;
        RECT 185.400 225.000 186.000 227.200 ;
        RECT 188.200 226.800 189.000 231.200 ;
        RECT 189.800 230.600 190.400 232.400 ;
        RECT 189.600 230.000 190.400 230.600 ;
        RECT 196.400 230.000 219.800 230.600 ;
        RECT 189.600 228.000 190.200 230.000 ;
        RECT 196.400 229.400 197.200 230.000 ;
        RECT 214.000 229.600 214.800 230.000 ;
        RECT 217.200 229.600 218.000 230.000 ;
        RECT 219.000 229.800 219.800 230.000 ;
        RECT 190.800 228.600 194.600 229.400 ;
        RECT 189.600 227.400 190.800 228.000 ;
        RECT 188.200 226.000 189.200 226.800 ;
        RECT 180.400 223.600 181.800 224.400 ;
        RECT 181.000 223.000 181.800 223.600 ;
        RECT 185.200 223.000 186.000 225.000 ;
        RECT 188.400 222.200 189.200 226.000 ;
        RECT 190.000 222.200 190.800 227.400 ;
        RECT 193.800 227.400 194.600 228.600 ;
        RECT 193.800 226.800 195.600 227.400 ;
        RECT 194.800 226.200 195.600 226.800 ;
        RECT 199.600 226.400 200.400 229.200 ;
        RECT 202.800 228.600 206.000 229.400 ;
        RECT 209.800 228.600 211.800 229.400 ;
        RECT 220.400 229.000 221.200 234.600 ;
        RECT 225.800 232.800 226.600 237.600 ;
        RECT 230.000 235.000 230.800 239.000 ;
        RECT 225.000 232.200 226.600 232.800 ;
        RECT 222.000 230.300 222.800 230.400 ;
        RECT 223.600 230.300 224.400 231.200 ;
        RECT 222.000 229.700 224.400 230.300 ;
        RECT 222.000 229.600 222.800 229.700 ;
        RECT 223.600 229.600 224.400 229.700 ;
        RECT 202.400 227.800 203.200 228.000 ;
        RECT 202.400 227.200 206.800 227.800 ;
        RECT 206.000 227.000 206.800 227.200 ;
        RECT 207.600 226.800 208.400 228.400 ;
        RECT 194.800 225.400 197.200 226.200 ;
        RECT 199.600 225.600 200.600 226.400 ;
        RECT 203.600 225.600 205.200 226.400 ;
        RECT 206.000 226.200 206.800 226.400 ;
        RECT 209.800 226.200 210.600 228.600 ;
        RECT 212.400 228.200 221.200 229.000 ;
        RECT 225.000 228.400 225.600 232.200 ;
        RECT 230.200 231.600 230.800 235.000 ;
        RECT 232.400 233.600 233.200 234.400 ;
        RECT 232.400 232.400 233.000 233.600 ;
        RECT 233.800 232.400 234.600 239.800 ;
        RECT 239.600 236.400 240.400 239.800 ;
        RECT 239.400 235.800 240.400 236.400 ;
        RECT 239.400 235.200 240.000 235.800 ;
        RECT 242.800 235.200 243.600 239.800 ;
        RECT 246.000 237.000 246.800 239.800 ;
        RECT 247.600 237.000 248.400 239.800 ;
        RECT 231.600 231.800 233.000 232.400 ;
        RECT 233.600 231.800 234.600 232.400 ;
        RECT 238.000 234.600 240.000 235.200 ;
        RECT 231.600 231.600 232.400 231.800 ;
        RECT 227.000 231.000 230.800 231.600 ;
        RECT 227.000 229.000 227.600 231.000 ;
        RECT 233.600 230.400 234.200 231.800 ;
        RECT 215.800 226.800 218.800 227.600 ;
        RECT 215.800 226.200 216.600 226.800 ;
        RECT 206.000 225.600 210.600 226.200 ;
        RECT 196.400 222.200 197.200 225.400 ;
        RECT 214.000 225.400 216.600 226.200 ;
        RECT 198.000 222.200 198.800 225.000 ;
        RECT 199.600 222.200 200.400 225.000 ;
        RECT 201.200 222.200 202.000 225.000 ;
        RECT 202.800 222.200 203.600 225.000 ;
        RECT 206.000 222.200 206.800 225.000 ;
        RECT 209.200 222.200 210.000 225.000 ;
        RECT 210.800 222.200 211.600 225.000 ;
        RECT 212.400 222.200 213.200 225.000 ;
        RECT 214.000 222.200 214.800 225.400 ;
        RECT 220.400 222.200 221.200 228.200 ;
        RECT 223.600 227.600 225.600 228.400 ;
        RECT 226.200 228.200 227.600 229.000 ;
        RECT 228.400 228.800 229.200 230.400 ;
        RECT 230.000 228.800 230.800 230.400 ;
        RECT 233.200 229.600 234.200 230.400 ;
        RECT 233.600 228.400 234.200 229.600 ;
        RECT 234.800 228.800 235.600 230.400 ;
        RECT 238.000 229.000 238.800 234.600 ;
        RECT 240.600 234.400 244.800 235.200 ;
        RECT 249.200 235.000 250.000 239.800 ;
        RECT 252.400 235.000 253.200 239.800 ;
        RECT 240.600 234.000 241.200 234.400 ;
        RECT 239.600 233.200 241.200 234.000 ;
        RECT 244.200 233.800 250.000 234.400 ;
        RECT 242.200 233.200 243.600 233.800 ;
        RECT 242.200 233.000 248.400 233.200 ;
        RECT 243.000 232.600 248.400 233.000 ;
        RECT 247.600 232.400 248.400 232.600 ;
        RECT 249.400 233.000 250.000 233.800 ;
        RECT 250.600 233.600 253.200 234.400 ;
        RECT 255.600 233.600 256.400 239.800 ;
        RECT 257.200 237.000 258.000 239.800 ;
        RECT 258.800 237.000 259.600 239.800 ;
        RECT 260.400 237.000 261.200 239.800 ;
        RECT 258.800 234.400 263.000 235.200 ;
        RECT 263.600 234.400 264.400 239.800 ;
        RECT 266.800 235.200 267.600 239.800 ;
        RECT 266.800 234.600 269.400 235.200 ;
        RECT 263.600 233.600 266.200 234.400 ;
        RECT 257.200 233.000 258.000 233.200 ;
        RECT 249.400 232.400 258.000 233.000 ;
        RECT 260.400 233.000 261.200 233.200 ;
        RECT 268.800 233.000 269.400 234.600 ;
        RECT 260.400 232.400 269.400 233.000 ;
        RECT 268.800 230.600 269.400 232.400 ;
        RECT 270.000 232.000 270.800 239.800 ;
        RECT 278.600 232.400 279.400 239.800 ;
        RECT 270.000 231.200 271.000 232.000 ;
        RECT 239.400 230.000 262.800 230.600 ;
        RECT 268.800 230.000 269.600 230.600 ;
        RECT 239.400 229.800 240.400 230.000 ;
        RECT 239.600 229.600 240.400 229.800 ;
        RECT 244.400 229.600 245.200 230.000 ;
        RECT 262.000 229.400 262.800 230.000 ;
        RECT 225.000 227.000 225.600 227.600 ;
        RECT 226.600 227.800 227.600 228.200 ;
        RECT 226.600 227.200 230.800 227.800 ;
        RECT 231.600 227.600 234.200 228.400 ;
        RECT 236.400 228.200 237.200 228.400 ;
        RECT 235.600 227.600 237.200 228.200 ;
        RECT 238.000 228.200 246.800 229.000 ;
        RECT 247.400 228.600 249.400 229.400 ;
        RECT 253.200 228.600 256.400 229.400 ;
        RECT 225.000 226.600 225.800 227.000 ;
        RECT 225.000 226.000 226.600 226.600 ;
        RECT 225.800 223.000 226.600 226.000 ;
        RECT 230.200 225.000 230.800 227.200 ;
        RECT 231.800 226.200 232.400 227.600 ;
        RECT 235.600 227.200 236.400 227.600 ;
        RECT 233.400 226.200 237.000 226.600 ;
        RECT 230.000 223.000 230.800 225.000 ;
        RECT 231.600 222.200 232.400 226.200 ;
        RECT 233.200 226.000 237.200 226.200 ;
        RECT 233.200 222.200 234.000 226.000 ;
        RECT 236.400 222.200 237.200 226.000 ;
        RECT 238.000 222.200 238.800 228.200 ;
        RECT 240.400 226.800 243.400 227.600 ;
        RECT 242.600 226.200 243.400 226.800 ;
        RECT 248.600 226.200 249.400 228.600 ;
        RECT 250.800 226.800 251.600 228.400 ;
        RECT 256.000 227.800 256.800 228.000 ;
        RECT 252.400 227.200 256.800 227.800 ;
        RECT 252.400 227.000 253.200 227.200 ;
        RECT 258.800 226.400 259.600 229.200 ;
        RECT 264.600 228.600 268.400 229.400 ;
        RECT 264.600 227.400 265.400 228.600 ;
        RECT 269.000 228.000 269.600 230.000 ;
        RECT 252.400 226.200 253.200 226.400 ;
        RECT 242.600 225.400 245.200 226.200 ;
        RECT 248.600 225.600 253.200 226.200 ;
        RECT 254.000 225.600 255.600 226.400 ;
        RECT 258.600 225.600 259.600 226.400 ;
        RECT 263.600 226.800 265.400 227.400 ;
        RECT 268.400 227.400 269.600 228.000 ;
        RECT 263.600 226.200 264.400 226.800 ;
        RECT 244.400 222.200 245.200 225.400 ;
        RECT 262.000 225.400 264.400 226.200 ;
        RECT 246.000 222.200 246.800 225.000 ;
        RECT 247.600 222.200 248.400 225.000 ;
        RECT 249.200 222.200 250.000 225.000 ;
        RECT 252.400 222.200 253.200 225.000 ;
        RECT 255.600 222.200 256.400 225.000 ;
        RECT 257.200 222.200 258.000 225.000 ;
        RECT 258.800 222.200 259.600 225.000 ;
        RECT 260.400 222.200 261.200 225.000 ;
        RECT 262.000 222.200 262.800 225.400 ;
        RECT 268.400 222.200 269.200 227.400 ;
        RECT 270.200 226.800 271.000 231.200 ;
        RECT 270.000 226.000 271.000 226.800 ;
        RECT 278.000 231.800 279.400 232.400 ;
        RECT 278.000 230.400 278.600 231.800 ;
        RECT 282.800 231.200 283.600 239.800 ;
        RECT 279.600 230.800 283.600 231.200 ;
        RECT 279.400 230.600 283.600 230.800 ;
        RECT 278.000 229.600 278.800 230.400 ;
        RECT 279.400 230.000 280.200 230.600 ;
        RECT 278.000 226.200 278.600 229.600 ;
        RECT 279.400 227.000 280.000 230.000 ;
        RECT 279.400 226.400 281.800 227.000 ;
        RECT 270.000 222.200 270.800 226.000 ;
        RECT 273.200 224.300 274.000 224.400 ;
        RECT 278.000 224.300 278.800 226.200 ;
        RECT 273.200 223.700 278.800 224.300 ;
        RECT 273.200 223.600 274.000 223.700 ;
        RECT 278.000 222.200 278.800 223.700 ;
        RECT 281.200 224.200 281.800 226.400 ;
        RECT 282.800 224.800 283.600 226.400 ;
        RECT 281.200 222.200 282.000 224.200 ;
        RECT 284.400 222.200 285.200 239.800 ;
        RECT 289.200 234.300 290.000 239.800 ;
        RECT 290.800 234.300 291.600 234.400 ;
        RECT 289.200 233.700 291.600 234.300 ;
        RECT 287.600 226.800 288.400 228.400 ;
        RECT 286.000 224.800 286.800 226.400 ;
        RECT 289.200 222.200 290.000 233.700 ;
        RECT 290.800 233.600 291.600 233.700 ;
        RECT 290.800 226.800 291.600 228.400 ;
        RECT 292.400 226.200 293.200 239.800 ;
        RECT 296.400 233.600 297.200 234.400 ;
        RECT 294.000 231.600 294.800 233.200 ;
        RECT 296.400 232.400 297.000 233.600 ;
        RECT 297.800 232.400 298.600 239.800 ;
        RECT 295.600 231.800 297.000 232.400 ;
        RECT 297.600 231.800 298.600 232.400 ;
        RECT 295.600 231.600 296.400 231.800 ;
        RECT 297.600 228.400 298.200 231.800 ;
        RECT 298.800 230.300 299.600 230.400 ;
        RECT 300.400 230.300 301.200 230.400 ;
        RECT 298.800 229.700 301.200 230.300 ;
        RECT 298.800 228.800 299.600 229.700 ;
        RECT 300.400 229.600 301.200 229.700 ;
        RECT 295.600 227.600 298.200 228.400 ;
        RECT 300.400 228.200 301.200 228.400 ;
        RECT 299.600 227.600 301.200 228.200 ;
        RECT 303.600 228.300 304.400 239.800 ;
        RECT 307.800 232.400 308.600 239.800 ;
        RECT 309.200 233.600 310.000 234.400 ;
        RECT 309.400 232.400 310.000 233.600 ;
        RECT 314.200 232.400 315.000 239.800 ;
        RECT 319.600 236.400 320.400 239.800 ;
        RECT 319.400 235.800 320.400 236.400 ;
        RECT 319.400 235.200 320.000 235.800 ;
        RECT 322.800 235.200 323.600 239.800 ;
        RECT 326.000 237.000 326.800 239.800 ;
        RECT 327.600 237.000 328.400 239.800 ;
        RECT 318.000 234.600 320.000 235.200 ;
        RECT 315.600 233.600 316.400 234.400 ;
        RECT 315.800 232.400 316.400 233.600 ;
        RECT 307.800 231.800 308.800 232.400 ;
        RECT 309.400 231.800 310.800 232.400 ;
        RECT 314.200 231.800 315.200 232.400 ;
        RECT 315.800 231.800 317.200 232.400 ;
        RECT 306.800 228.800 307.600 230.400 ;
        RECT 308.200 228.400 308.800 231.800 ;
        RECT 310.000 231.600 310.800 231.800 ;
        RECT 313.200 228.800 314.000 230.400 ;
        RECT 314.600 230.300 315.200 231.800 ;
        RECT 316.400 231.600 317.200 231.800 ;
        RECT 316.400 230.300 317.200 230.400 ;
        RECT 314.600 229.700 317.200 230.300 ;
        RECT 314.600 228.400 315.200 229.700 ;
        RECT 316.400 229.600 317.200 229.700 ;
        RECT 318.000 229.000 318.800 234.600 ;
        RECT 320.600 234.400 324.800 235.200 ;
        RECT 329.200 235.000 330.000 239.800 ;
        RECT 332.400 235.000 333.200 239.800 ;
        RECT 320.600 234.000 321.200 234.400 ;
        RECT 319.600 233.200 321.200 234.000 ;
        RECT 324.200 233.800 330.000 234.400 ;
        RECT 322.200 233.200 323.600 233.800 ;
        RECT 322.200 233.000 328.400 233.200 ;
        RECT 323.000 232.600 328.400 233.000 ;
        RECT 327.600 232.400 328.400 232.600 ;
        RECT 329.400 233.000 330.000 233.800 ;
        RECT 330.600 233.600 333.200 234.400 ;
        RECT 335.600 233.600 336.400 239.800 ;
        RECT 337.200 237.000 338.000 239.800 ;
        RECT 338.800 237.000 339.600 239.800 ;
        RECT 340.400 237.000 341.200 239.800 ;
        RECT 338.800 234.400 343.000 235.200 ;
        RECT 343.600 234.400 344.400 239.800 ;
        RECT 346.800 235.200 347.600 239.800 ;
        RECT 346.800 234.600 349.400 235.200 ;
        RECT 343.600 233.600 346.200 234.400 ;
        RECT 337.200 233.000 338.000 233.200 ;
        RECT 329.400 232.400 338.000 233.000 ;
        RECT 340.400 233.000 341.200 233.200 ;
        RECT 348.800 233.000 349.400 234.600 ;
        RECT 340.400 232.400 349.400 233.000 ;
        RECT 348.800 230.600 349.400 232.400 ;
        RECT 350.000 232.000 350.800 239.800 ;
        RECT 350.000 231.200 351.000 232.000 ;
        RECT 319.400 230.000 342.800 230.600 ;
        RECT 348.800 230.000 349.600 230.600 ;
        RECT 319.400 229.800 320.200 230.000 ;
        RECT 322.800 229.600 323.600 230.000 ;
        RECT 324.400 229.600 325.200 230.000 ;
        RECT 342.000 229.400 342.800 230.000 ;
        RECT 305.200 228.300 306.000 228.400 ;
        RECT 303.600 228.200 306.000 228.300 ;
        RECT 303.600 227.700 306.800 228.200 ;
        RECT 295.800 226.200 296.400 227.600 ;
        RECT 299.600 227.200 300.400 227.600 ;
        RECT 297.400 226.200 301.000 226.600 ;
        RECT 292.400 225.600 294.200 226.200 ;
        RECT 293.400 224.400 294.200 225.600 ;
        RECT 293.400 223.600 294.800 224.400 ;
        RECT 293.400 222.200 294.200 223.600 ;
        RECT 295.600 222.200 296.400 226.200 ;
        RECT 297.200 226.000 301.200 226.200 ;
        RECT 297.200 222.200 298.000 226.000 ;
        RECT 300.400 222.200 301.200 226.000 ;
        RECT 302.000 224.800 302.800 226.400 ;
        RECT 303.600 222.200 304.400 227.700 ;
        RECT 305.200 227.600 306.800 227.700 ;
        RECT 308.200 227.600 310.800 228.400 ;
        RECT 311.600 228.200 312.400 228.400 ;
        RECT 311.600 227.600 313.200 228.200 ;
        RECT 314.600 227.600 317.200 228.400 ;
        RECT 318.000 228.200 326.800 229.000 ;
        RECT 327.400 228.600 329.400 229.400 ;
        RECT 333.200 228.600 336.400 229.400 ;
        RECT 306.000 227.200 306.800 227.600 ;
        RECT 305.400 226.200 309.000 226.600 ;
        RECT 310.000 226.200 310.600 227.600 ;
        RECT 312.400 227.200 313.200 227.600 ;
        RECT 311.800 226.200 315.400 226.600 ;
        RECT 316.400 226.200 317.000 227.600 ;
        RECT 305.200 226.000 309.200 226.200 ;
        RECT 305.200 222.200 306.000 226.000 ;
        RECT 308.400 222.200 309.200 226.000 ;
        RECT 310.000 222.200 310.800 226.200 ;
        RECT 311.600 226.000 315.600 226.200 ;
        RECT 311.600 222.200 312.400 226.000 ;
        RECT 314.800 222.200 315.600 226.000 ;
        RECT 316.400 222.200 317.200 226.200 ;
        RECT 318.000 222.200 318.800 228.200 ;
        RECT 320.400 226.800 323.400 227.600 ;
        RECT 322.600 226.200 323.400 226.800 ;
        RECT 328.600 226.200 329.400 228.600 ;
        RECT 330.800 226.800 331.600 228.400 ;
        RECT 336.000 227.800 336.800 228.000 ;
        RECT 332.400 227.200 336.800 227.800 ;
        RECT 332.400 227.000 333.200 227.200 ;
        RECT 338.800 226.400 339.600 229.200 ;
        RECT 344.600 228.600 348.400 229.400 ;
        RECT 344.600 227.400 345.400 228.600 ;
        RECT 349.000 228.000 349.600 230.000 ;
        RECT 332.400 226.200 333.200 226.400 ;
        RECT 322.600 225.400 325.200 226.200 ;
        RECT 328.600 225.600 333.200 226.200 ;
        RECT 334.000 225.600 335.600 226.400 ;
        RECT 338.600 225.600 339.600 226.400 ;
        RECT 343.600 226.800 345.400 227.400 ;
        RECT 348.400 227.400 349.600 228.000 ;
        RECT 343.600 226.200 344.400 226.800 ;
        RECT 324.400 222.200 325.200 225.400 ;
        RECT 342.000 225.400 344.400 226.200 ;
        RECT 326.000 222.200 326.800 225.000 ;
        RECT 327.600 222.200 328.400 225.000 ;
        RECT 329.200 222.200 330.000 225.000 ;
        RECT 332.400 222.200 333.200 225.000 ;
        RECT 335.600 222.200 336.400 225.000 ;
        RECT 337.200 222.200 338.000 225.000 ;
        RECT 338.800 222.200 339.600 225.000 ;
        RECT 340.400 222.200 341.200 225.000 ;
        RECT 342.000 222.200 342.800 225.400 ;
        RECT 348.400 222.200 349.200 227.400 ;
        RECT 350.200 226.800 351.000 231.200 ;
        RECT 353.200 226.800 354.000 228.400 ;
        RECT 350.000 226.300 351.000 226.800 ;
        RECT 351.600 226.300 352.400 226.400 ;
        RECT 350.000 225.700 352.400 226.300 ;
        RECT 350.000 222.200 350.800 225.700 ;
        RECT 351.600 225.600 352.400 225.700 ;
        RECT 354.800 222.200 355.600 239.800 ;
        RECT 356.400 226.800 357.200 228.400 ;
        RECT 358.000 226.200 358.800 239.800 ;
        RECT 362.000 233.600 362.800 234.400 ;
        RECT 359.600 231.600 360.400 233.200 ;
        RECT 362.000 232.400 362.600 233.600 ;
        RECT 363.400 232.400 364.200 239.800 ;
        RECT 361.200 231.800 362.600 232.400 ;
        RECT 363.200 231.800 364.200 232.400 ;
        RECT 367.600 232.400 368.400 239.800 ;
        RECT 370.800 232.800 371.600 239.800 ;
        RECT 374.000 235.800 374.800 239.800 ;
        RECT 374.200 235.600 374.800 235.800 ;
        RECT 377.200 235.800 378.000 239.800 ;
        RECT 380.400 235.800 381.200 239.800 ;
        RECT 377.200 235.600 377.800 235.800 ;
        RECT 374.200 235.000 377.800 235.600 ;
        RECT 380.600 235.600 381.200 235.800 ;
        RECT 383.600 235.800 384.400 239.800 ;
        RECT 388.400 236.400 389.200 239.800 ;
        RECT 388.200 235.800 389.200 236.400 ;
        RECT 383.600 235.600 384.200 235.800 ;
        RECT 380.600 235.000 384.200 235.600 ;
        RECT 388.200 235.200 388.800 235.800 ;
        RECT 391.600 235.200 392.400 239.800 ;
        RECT 394.800 237.000 395.600 239.800 ;
        RECT 396.400 237.000 397.200 239.800 ;
        RECT 367.600 231.800 370.200 232.400 ;
        RECT 370.800 231.800 371.800 232.800 ;
        RECT 374.200 232.400 374.800 235.000 ;
        RECT 375.600 232.800 376.400 234.400 ;
        RECT 380.600 232.400 381.200 235.000 ;
        RECT 386.800 234.600 388.800 235.200 ;
        RECT 382.000 232.800 382.800 234.400 ;
        RECT 361.200 231.600 362.000 231.800 ;
        RECT 359.700 230.300 360.300 231.600 ;
        RECT 363.200 230.300 363.800 231.800 ;
        RECT 359.700 229.700 363.800 230.300 ;
        RECT 363.200 228.400 363.800 229.700 ;
        RECT 364.400 228.800 365.200 230.400 ;
        RECT 367.600 229.600 368.600 230.400 ;
        RECT 367.800 228.800 368.600 229.600 ;
        RECT 369.600 229.800 370.200 231.800 ;
        RECT 369.600 229.000 370.600 229.800 ;
        RECT 361.200 227.600 363.800 228.400 ;
        RECT 366.000 228.200 366.800 228.400 ;
        RECT 365.200 227.600 366.800 228.200 ;
        RECT 361.400 226.200 362.000 227.600 ;
        RECT 365.200 227.200 366.000 227.600 ;
        RECT 369.600 227.400 370.200 229.000 ;
        RECT 371.200 228.400 371.800 231.800 ;
        RECT 374.000 231.600 374.800 232.400 ;
        RECT 374.200 228.400 374.800 231.600 ;
        RECT 378.800 230.800 379.600 232.400 ;
        RECT 380.400 231.600 381.200 232.400 ;
        RECT 376.400 229.600 378.000 230.400 ;
        RECT 380.600 228.400 381.200 231.600 ;
        RECT 385.200 230.800 386.000 232.400 ;
        RECT 382.800 229.600 384.400 230.400 ;
        RECT 386.800 229.000 387.600 234.600 ;
        RECT 389.400 234.400 393.600 235.200 ;
        RECT 398.000 235.000 398.800 239.800 ;
        RECT 401.200 235.000 402.000 239.800 ;
        RECT 389.400 234.000 390.000 234.400 ;
        RECT 388.400 233.200 390.000 234.000 ;
        RECT 393.000 233.800 398.800 234.400 ;
        RECT 391.000 233.200 392.400 233.800 ;
        RECT 391.000 233.000 397.200 233.200 ;
        RECT 391.800 232.600 397.200 233.000 ;
        RECT 396.400 232.400 397.200 232.600 ;
        RECT 398.200 233.000 398.800 233.800 ;
        RECT 399.400 233.600 402.000 234.400 ;
        RECT 404.400 233.600 405.200 239.800 ;
        RECT 406.000 237.000 406.800 239.800 ;
        RECT 407.600 237.000 408.400 239.800 ;
        RECT 409.200 237.000 410.000 239.800 ;
        RECT 407.600 234.400 411.800 235.200 ;
        RECT 412.400 234.400 413.200 239.800 ;
        RECT 415.600 235.200 416.400 239.800 ;
        RECT 415.600 234.600 418.200 235.200 ;
        RECT 412.400 233.600 415.000 234.400 ;
        RECT 406.000 233.000 406.800 233.200 ;
        RECT 398.200 232.400 406.800 233.000 ;
        RECT 409.200 233.000 410.000 233.200 ;
        RECT 417.600 233.000 418.200 234.600 ;
        RECT 409.200 232.400 418.200 233.000 ;
        RECT 417.600 230.600 418.200 232.400 ;
        RECT 418.800 232.000 419.600 239.800 ;
        RECT 426.800 235.000 427.600 239.000 ;
        RECT 418.800 231.200 419.800 232.000 ;
        RECT 388.200 230.000 411.600 230.600 ;
        RECT 417.600 230.000 418.400 230.600 ;
        RECT 388.200 229.800 389.000 230.000 ;
        RECT 390.000 229.600 390.800 230.000 ;
        RECT 393.200 229.600 394.000 230.000 ;
        RECT 410.800 229.400 411.600 230.000 ;
        RECT 370.800 228.300 371.800 228.400 ;
        RECT 372.400 228.300 373.200 228.400 ;
        RECT 370.800 227.700 373.200 228.300 ;
        RECT 374.200 228.200 375.800 228.400 ;
        RECT 380.600 228.200 382.200 228.400 ;
        RECT 386.800 228.200 395.600 229.000 ;
        RECT 396.200 228.600 398.200 229.400 ;
        RECT 402.000 228.600 405.200 229.400 ;
        RECT 374.200 227.800 376.000 228.200 ;
        RECT 380.600 227.800 382.400 228.200 ;
        RECT 370.800 227.600 371.800 227.700 ;
        RECT 372.400 227.600 373.200 227.700 ;
        RECT 367.600 226.800 370.200 227.400 ;
        RECT 363.000 226.200 366.600 226.600 ;
        RECT 358.000 225.600 359.800 226.200 ;
        RECT 359.000 224.400 359.800 225.600 ;
        RECT 359.000 223.600 360.400 224.400 ;
        RECT 359.000 222.200 359.800 223.600 ;
        RECT 361.200 222.200 362.000 226.200 ;
        RECT 362.800 226.000 366.800 226.200 ;
        RECT 362.800 222.200 363.600 226.000 ;
        RECT 366.000 222.200 366.800 226.000 ;
        RECT 367.600 222.200 368.400 226.800 ;
        RECT 371.200 226.200 371.800 227.600 ;
        RECT 370.800 225.600 371.800 226.200 ;
        RECT 370.800 222.200 371.600 225.600 ;
        RECT 375.200 222.200 376.000 227.800 ;
        RECT 381.600 222.200 382.400 227.800 ;
        RECT 386.800 222.200 387.600 228.200 ;
        RECT 389.200 226.800 392.200 227.600 ;
        RECT 391.400 226.200 392.200 226.800 ;
        RECT 397.400 226.200 398.200 228.600 ;
        RECT 399.600 226.800 400.400 228.400 ;
        RECT 404.800 227.800 405.600 228.000 ;
        RECT 401.200 227.200 405.600 227.800 ;
        RECT 401.200 227.000 402.000 227.200 ;
        RECT 407.600 226.400 408.400 229.200 ;
        RECT 413.400 228.600 417.200 229.400 ;
        RECT 413.400 227.400 414.200 228.600 ;
        RECT 417.800 228.000 418.400 230.000 ;
        RECT 401.200 226.200 402.000 226.400 ;
        RECT 391.400 225.400 394.000 226.200 ;
        RECT 397.400 225.600 402.000 226.200 ;
        RECT 402.800 225.600 404.400 226.400 ;
        RECT 407.400 225.600 408.400 226.400 ;
        RECT 412.400 226.800 414.200 227.400 ;
        RECT 417.200 227.400 418.400 228.000 ;
        RECT 412.400 226.200 413.200 226.800 ;
        RECT 393.200 222.200 394.000 225.400 ;
        RECT 410.800 225.400 413.200 226.200 ;
        RECT 394.800 222.200 395.600 225.000 ;
        RECT 396.400 222.200 397.200 225.000 ;
        RECT 398.000 222.200 398.800 225.000 ;
        RECT 401.200 222.200 402.000 225.000 ;
        RECT 404.400 222.200 405.200 225.000 ;
        RECT 406.000 222.200 406.800 225.000 ;
        RECT 407.600 222.200 408.400 225.000 ;
        RECT 409.200 222.200 410.000 225.000 ;
        RECT 410.800 222.200 411.600 225.400 ;
        RECT 417.200 222.200 418.000 227.400 ;
        RECT 419.000 226.800 419.800 231.200 ;
        RECT 426.800 231.600 427.400 235.000 ;
        RECT 431.000 232.800 431.800 239.800 ;
        RECT 431.000 232.200 432.600 232.800 ;
        RECT 426.800 231.000 430.600 231.600 ;
        RECT 423.600 230.300 424.400 230.400 ;
        RECT 426.800 230.300 427.600 230.400 ;
        RECT 423.600 229.700 427.600 230.300 ;
        RECT 423.600 229.600 424.400 229.700 ;
        RECT 426.800 228.800 427.600 229.700 ;
        RECT 428.400 228.800 429.200 230.400 ;
        RECT 430.000 229.000 430.600 231.000 ;
        RECT 432.000 230.400 432.600 232.200 ;
        RECT 431.600 229.600 432.600 230.400 ;
        RECT 433.200 230.300 434.000 231.200 ;
        RECT 438.000 230.300 438.800 239.800 ;
        RECT 441.200 231.200 442.000 239.800 ;
        RECT 444.400 231.200 445.200 239.800 ;
        RECT 447.600 231.200 448.400 239.800 ;
        RECT 450.800 231.200 451.600 239.800 ;
        RECT 455.600 236.400 456.400 239.800 ;
        RECT 455.400 235.800 456.400 236.400 ;
        RECT 455.400 235.200 456.000 235.800 ;
        RECT 458.800 235.200 459.600 239.800 ;
        RECT 462.000 237.000 462.800 239.800 ;
        RECT 463.600 237.000 464.400 239.800 ;
        RECT 454.000 234.600 456.000 235.200 ;
        RECT 441.200 230.400 443.000 231.200 ;
        RECT 444.400 230.400 446.600 231.200 ;
        RECT 447.600 230.400 449.800 231.200 ;
        RECT 450.800 230.400 453.200 231.200 ;
        RECT 433.200 229.700 438.800 230.300 ;
        RECT 433.200 229.600 434.000 229.700 ;
        RECT 430.000 228.200 431.400 229.000 ;
        RECT 432.000 228.400 432.600 229.600 ;
        RECT 430.000 227.800 431.000 228.200 ;
        RECT 418.800 226.300 419.800 226.800 ;
        RECT 426.800 227.200 431.000 227.800 ;
        RECT 432.000 227.600 434.000 228.400 ;
        RECT 425.200 226.300 426.000 226.400 ;
        RECT 418.800 225.700 426.000 226.300 ;
        RECT 418.800 222.200 419.600 225.700 ;
        RECT 425.200 225.600 426.000 225.700 ;
        RECT 426.800 225.000 427.400 227.200 ;
        RECT 432.000 227.000 432.600 227.600 ;
        RECT 431.800 226.600 432.600 227.000 ;
        RECT 431.000 226.000 432.600 226.600 ;
        RECT 426.800 223.000 427.600 225.000 ;
        RECT 431.000 223.000 431.800 226.000 ;
        RECT 436.400 224.800 437.200 226.400 ;
        RECT 438.000 222.200 438.800 229.700 ;
        RECT 442.200 229.000 443.000 230.400 ;
        RECT 445.800 229.000 446.600 230.400 ;
        RECT 449.000 229.000 449.800 230.400 ;
        RECT 439.600 228.200 441.400 229.000 ;
        RECT 442.200 228.200 444.800 229.000 ;
        RECT 445.800 228.200 448.200 229.000 ;
        RECT 449.000 228.200 451.600 229.000 ;
        RECT 439.600 227.600 440.400 228.200 ;
        RECT 442.200 227.600 443.000 228.200 ;
        RECT 445.800 227.600 446.600 228.200 ;
        RECT 449.000 227.600 449.800 228.200 ;
        RECT 452.400 227.600 453.200 230.400 ;
        RECT 441.200 226.800 443.000 227.600 ;
        RECT 444.400 226.800 446.600 227.600 ;
        RECT 447.600 226.800 449.800 227.600 ;
        RECT 450.800 226.800 453.200 227.600 ;
        RECT 454.000 229.000 454.800 234.600 ;
        RECT 456.600 234.400 460.800 235.200 ;
        RECT 465.200 235.000 466.000 239.800 ;
        RECT 468.400 235.000 469.200 239.800 ;
        RECT 456.600 234.000 457.200 234.400 ;
        RECT 455.600 233.200 457.200 234.000 ;
        RECT 460.200 233.800 466.000 234.400 ;
        RECT 458.200 233.200 459.600 233.800 ;
        RECT 458.200 233.000 464.400 233.200 ;
        RECT 459.000 232.600 464.400 233.000 ;
        RECT 463.600 232.400 464.400 232.600 ;
        RECT 465.400 233.000 466.000 233.800 ;
        RECT 466.600 233.600 469.200 234.400 ;
        RECT 471.600 233.600 472.400 239.800 ;
        RECT 473.200 237.000 474.000 239.800 ;
        RECT 474.800 237.000 475.600 239.800 ;
        RECT 476.400 237.000 477.200 239.800 ;
        RECT 474.800 234.400 479.000 235.200 ;
        RECT 479.600 234.400 480.400 239.800 ;
        RECT 482.800 235.200 483.600 239.800 ;
        RECT 482.800 234.600 485.400 235.200 ;
        RECT 479.600 233.600 482.200 234.400 ;
        RECT 473.200 233.000 474.000 233.200 ;
        RECT 465.400 232.400 474.000 233.000 ;
        RECT 476.400 233.000 477.200 233.200 ;
        RECT 484.800 233.000 485.400 234.600 ;
        RECT 476.400 232.400 485.400 233.000 ;
        RECT 484.800 230.600 485.400 232.400 ;
        RECT 486.000 232.000 486.800 239.800 ;
        RECT 489.200 235.000 490.000 239.000 ;
        RECT 486.000 231.200 487.000 232.000 ;
        RECT 455.400 230.000 478.800 230.600 ;
        RECT 484.800 230.000 485.600 230.600 ;
        RECT 455.400 229.800 456.200 230.000 ;
        RECT 457.200 229.600 458.000 230.000 ;
        RECT 460.400 229.600 461.200 230.000 ;
        RECT 478.000 229.400 478.800 230.000 ;
        RECT 454.000 228.200 462.800 229.000 ;
        RECT 463.400 228.600 465.400 229.400 ;
        RECT 469.200 228.600 472.400 229.400 ;
        RECT 441.200 222.200 442.000 226.800 ;
        RECT 444.400 222.200 445.200 226.800 ;
        RECT 447.600 222.200 448.400 226.800 ;
        RECT 450.800 222.200 451.600 226.800 ;
        RECT 454.000 222.200 454.800 228.200 ;
        RECT 456.400 226.800 459.400 227.600 ;
        RECT 458.600 226.200 459.400 226.800 ;
        RECT 464.600 226.200 465.400 228.600 ;
        RECT 466.800 226.800 467.600 228.400 ;
        RECT 472.000 227.800 472.800 228.000 ;
        RECT 468.400 227.200 472.800 227.800 ;
        RECT 468.400 227.000 469.200 227.200 ;
        RECT 474.800 226.400 475.600 229.200 ;
        RECT 480.600 228.600 484.400 229.400 ;
        RECT 480.600 227.400 481.400 228.600 ;
        RECT 485.000 228.000 485.600 230.000 ;
        RECT 468.400 226.200 469.200 226.400 ;
        RECT 458.600 225.400 461.200 226.200 ;
        RECT 464.600 225.600 469.200 226.200 ;
        RECT 470.000 225.600 471.600 226.400 ;
        RECT 474.600 225.600 475.600 226.400 ;
        RECT 479.600 226.800 481.400 227.400 ;
        RECT 484.400 227.400 485.600 228.000 ;
        RECT 479.600 226.200 480.400 226.800 ;
        RECT 460.400 222.200 461.200 225.400 ;
        RECT 478.000 225.400 480.400 226.200 ;
        RECT 462.000 222.200 462.800 225.000 ;
        RECT 463.600 222.200 464.400 225.000 ;
        RECT 465.200 222.200 466.000 225.000 ;
        RECT 468.400 222.200 469.200 225.000 ;
        RECT 471.600 222.200 472.400 225.000 ;
        RECT 473.200 222.200 474.000 225.000 ;
        RECT 474.800 222.200 475.600 225.000 ;
        RECT 476.400 222.200 477.200 225.000 ;
        RECT 478.000 222.200 478.800 225.400 ;
        RECT 484.400 222.200 485.200 227.400 ;
        RECT 486.200 226.800 487.000 231.200 ;
        RECT 489.200 231.600 489.800 235.000 ;
        RECT 493.400 232.800 494.200 239.800 ;
        RECT 493.400 232.200 495.000 232.800 ;
        RECT 489.200 231.000 493.000 231.600 ;
        RECT 489.200 228.800 490.000 230.400 ;
        RECT 490.800 228.800 491.600 230.400 ;
        RECT 492.400 229.000 493.000 231.000 ;
        RECT 492.400 228.200 493.800 229.000 ;
        RECT 494.400 228.400 495.000 232.200 ;
        RECT 495.600 230.300 496.400 231.200 ;
        RECT 498.800 230.300 499.600 239.800 ;
        RECT 503.600 236.400 504.400 239.800 ;
        RECT 503.400 235.800 504.400 236.400 ;
        RECT 503.400 235.200 504.000 235.800 ;
        RECT 506.800 235.200 507.600 239.800 ;
        RECT 510.000 237.000 510.800 239.800 ;
        RECT 511.600 237.000 512.400 239.800 ;
        RECT 495.600 229.700 499.600 230.300 ;
        RECT 495.600 229.600 496.400 229.700 ;
        RECT 492.400 227.800 493.400 228.200 ;
        RECT 486.000 226.000 487.000 226.800 ;
        RECT 489.200 227.200 493.400 227.800 ;
        RECT 494.400 227.600 496.400 228.400 ;
        RECT 486.000 222.200 486.800 226.000 ;
        RECT 489.200 225.000 489.800 227.200 ;
        RECT 494.400 227.000 495.000 227.600 ;
        RECT 494.200 226.600 495.000 227.000 ;
        RECT 493.400 226.400 495.000 226.600 ;
        RECT 492.400 226.000 495.000 226.400 ;
        RECT 492.400 225.600 494.200 226.000 ;
        RECT 489.200 223.000 490.000 225.000 ;
        RECT 493.400 223.000 494.200 225.600 ;
        RECT 498.800 222.200 499.600 229.700 ;
        RECT 502.000 234.600 504.000 235.200 ;
        RECT 502.000 229.000 502.800 234.600 ;
        RECT 504.600 234.400 508.800 235.200 ;
        RECT 513.200 235.000 514.000 239.800 ;
        RECT 516.400 235.000 517.200 239.800 ;
        RECT 504.600 234.000 505.200 234.400 ;
        RECT 503.600 233.200 505.200 234.000 ;
        RECT 508.200 233.800 514.000 234.400 ;
        RECT 506.200 233.200 507.600 233.800 ;
        RECT 506.200 233.000 512.400 233.200 ;
        RECT 507.000 232.600 512.400 233.000 ;
        RECT 511.600 232.400 512.400 232.600 ;
        RECT 513.400 233.000 514.000 233.800 ;
        RECT 514.600 233.600 517.200 234.400 ;
        RECT 519.600 233.600 520.400 239.800 ;
        RECT 521.200 237.000 522.000 239.800 ;
        RECT 522.800 237.000 523.600 239.800 ;
        RECT 524.400 237.000 525.200 239.800 ;
        RECT 522.800 234.400 527.000 235.200 ;
        RECT 527.600 234.400 528.400 239.800 ;
        RECT 530.800 235.200 531.600 239.800 ;
        RECT 530.800 234.600 533.400 235.200 ;
        RECT 527.600 233.600 530.200 234.400 ;
        RECT 521.200 233.000 522.000 233.200 ;
        RECT 513.400 232.400 522.000 233.000 ;
        RECT 524.400 233.000 525.200 233.200 ;
        RECT 532.800 233.000 533.400 234.600 ;
        RECT 524.400 232.400 533.400 233.000 ;
        RECT 532.800 230.600 533.400 232.400 ;
        RECT 534.000 232.000 534.800 239.800 ;
        RECT 534.000 231.200 535.000 232.000 ;
        RECT 503.400 230.000 526.800 230.600 ;
        RECT 532.800 230.000 533.600 230.600 ;
        RECT 503.400 229.800 504.200 230.000 ;
        RECT 506.800 229.600 507.600 230.000 ;
        RECT 508.400 229.600 509.200 230.000 ;
        RECT 526.000 229.400 526.800 230.000 ;
        RECT 502.000 228.200 510.800 229.000 ;
        RECT 511.400 228.600 513.400 229.400 ;
        RECT 517.200 228.600 520.400 229.400 ;
        RECT 500.400 224.800 501.200 226.400 ;
        RECT 502.000 222.200 502.800 228.200 ;
        RECT 504.400 226.800 507.400 227.600 ;
        RECT 506.600 226.200 507.400 226.800 ;
        RECT 512.600 226.200 513.400 228.600 ;
        RECT 514.800 226.800 515.600 228.400 ;
        RECT 520.000 227.800 520.800 228.000 ;
        RECT 516.400 227.200 520.800 227.800 ;
        RECT 516.400 227.000 517.200 227.200 ;
        RECT 522.800 226.400 523.600 229.200 ;
        RECT 528.600 228.600 532.400 229.400 ;
        RECT 528.600 227.400 529.400 228.600 ;
        RECT 533.000 228.000 533.600 230.000 ;
        RECT 516.400 226.200 517.200 226.400 ;
        RECT 506.600 225.400 509.200 226.200 ;
        RECT 512.600 225.600 517.200 226.200 ;
        RECT 518.000 225.600 519.600 226.400 ;
        RECT 522.600 225.600 523.600 226.400 ;
        RECT 527.600 226.800 529.400 227.400 ;
        RECT 532.400 227.400 533.600 228.000 ;
        RECT 527.600 226.200 528.400 226.800 ;
        RECT 508.400 222.200 509.200 225.400 ;
        RECT 526.000 225.400 528.400 226.200 ;
        RECT 510.000 222.200 510.800 225.000 ;
        RECT 511.600 222.200 512.400 225.000 ;
        RECT 513.200 222.200 514.000 225.000 ;
        RECT 516.400 222.200 517.200 225.000 ;
        RECT 519.600 222.200 520.400 225.000 ;
        RECT 521.200 222.200 522.000 225.000 ;
        RECT 522.800 222.200 523.600 225.000 ;
        RECT 524.400 222.200 525.200 225.000 ;
        RECT 526.000 222.200 526.800 225.400 ;
        RECT 532.400 222.200 533.200 227.400 ;
        RECT 534.200 226.800 535.000 231.200 ;
        RECT 534.000 226.000 535.000 226.800 ;
        RECT 534.000 222.200 534.800 226.000 ;
        RECT 537.200 222.200 538.000 239.800 ;
        RECT 542.000 235.800 542.800 239.800 ;
        RECT 542.200 231.600 542.800 235.800 ;
        RECT 545.200 231.800 546.000 239.800 ;
        RECT 542.200 231.000 544.600 231.600 ;
        RECT 542.000 229.600 542.800 230.400 ;
        RECT 540.400 227.600 541.200 229.200 ;
        RECT 542.200 228.800 542.800 229.600 ;
        RECT 542.200 228.200 543.200 228.800 ;
        RECT 542.400 228.000 543.200 228.200 ;
        RECT 544.000 227.600 544.600 231.000 ;
        RECT 545.400 230.400 546.000 231.800 ;
        RECT 545.200 229.600 546.000 230.400 ;
        RECT 544.000 227.400 544.800 227.600 ;
        RECT 541.800 227.000 544.800 227.400 ;
        RECT 540.600 226.800 544.800 227.000 ;
        RECT 540.600 226.400 542.400 226.800 ;
        RECT 538.800 224.800 539.600 226.400 ;
        RECT 540.600 226.200 541.200 226.400 ;
        RECT 545.400 226.200 546.000 229.600 ;
        RECT 540.400 222.200 541.200 226.200 ;
        RECT 544.600 225.200 546.000 226.200 ;
        RECT 544.600 224.400 545.400 225.200 ;
        RECT 546.800 224.800 547.600 226.400 ;
        RECT 544.600 223.600 546.000 224.400 ;
        RECT 544.600 222.200 545.400 223.600 ;
        RECT 548.400 222.200 549.200 239.800 ;
        RECT 553.200 232.400 554.000 239.800 ;
        RECT 555.600 233.600 556.400 234.400 ;
        RECT 555.600 232.400 556.200 233.600 ;
        RECT 557.000 232.400 557.800 239.800 ;
        RECT 551.800 231.800 554.000 232.400 ;
        RECT 554.800 231.800 556.200 232.400 ;
        RECT 556.800 231.800 557.800 232.400 ;
        RECT 551.800 231.200 552.400 231.800 ;
        RECT 554.800 231.600 555.600 231.800 ;
        RECT 551.200 230.400 552.400 231.200 ;
        RECT 556.800 230.400 557.400 231.800 ;
        RECT 551.800 227.400 552.400 230.400 ;
        RECT 553.200 228.800 554.000 230.400 ;
        RECT 556.400 229.600 557.400 230.400 ;
        RECT 556.800 228.400 557.400 229.600 ;
        RECT 558.000 228.800 558.800 230.400 ;
        RECT 554.800 227.600 557.400 228.400 ;
        RECT 559.600 228.200 560.400 228.400 ;
        RECT 558.800 227.600 560.400 228.200 ;
        RECT 551.800 226.800 554.000 227.400 ;
        RECT 553.200 222.200 554.000 226.800 ;
        RECT 555.000 226.200 555.600 227.600 ;
        RECT 558.800 227.200 559.600 227.600 ;
        RECT 561.200 226.800 562.000 228.400 ;
        RECT 556.600 226.200 560.200 226.600 ;
        RECT 562.800 226.200 563.600 239.800 ;
        RECT 564.400 231.600 565.200 233.200 ;
        RECT 566.000 231.600 566.800 233.200 ;
        RECT 564.500 230.300 565.100 231.600 ;
        RECT 567.600 230.300 568.400 239.800 ;
        RECT 577.200 232.000 578.000 239.800 ;
        RECT 580.400 235.200 581.200 239.800 ;
        RECT 577.000 231.200 578.000 232.000 ;
        RECT 578.600 234.600 581.200 235.200 ;
        RECT 578.600 233.000 579.200 234.600 ;
        RECT 583.600 234.400 584.400 239.800 ;
        RECT 586.800 237.000 587.600 239.800 ;
        RECT 588.400 237.000 589.200 239.800 ;
        RECT 590.000 237.000 590.800 239.800 ;
        RECT 585.000 234.400 589.200 235.200 ;
        RECT 581.800 233.600 584.400 234.400 ;
        RECT 591.600 233.600 592.400 239.800 ;
        RECT 594.800 235.000 595.600 239.800 ;
        RECT 598.000 235.000 598.800 239.800 ;
        RECT 599.600 237.000 600.400 239.800 ;
        RECT 601.200 237.000 602.000 239.800 ;
        RECT 604.400 235.200 605.200 239.800 ;
        RECT 607.600 236.400 608.400 239.800 ;
        RECT 607.600 235.800 608.600 236.400 ;
        RECT 608.000 235.200 608.600 235.800 ;
        RECT 603.200 234.400 607.400 235.200 ;
        RECT 608.000 234.600 610.000 235.200 ;
        RECT 594.800 233.600 597.400 234.400 ;
        RECT 598.000 233.800 603.800 234.400 ;
        RECT 606.800 234.000 607.400 234.400 ;
        RECT 586.800 233.000 587.600 233.200 ;
        RECT 578.600 232.400 587.600 233.000 ;
        RECT 590.000 233.000 590.800 233.200 ;
        RECT 598.000 233.000 598.600 233.800 ;
        RECT 604.400 233.200 605.800 233.800 ;
        RECT 606.800 233.200 608.400 234.000 ;
        RECT 590.000 232.400 598.600 233.000 ;
        RECT 599.600 233.000 605.800 233.200 ;
        RECT 599.600 232.600 605.000 233.000 ;
        RECT 599.600 232.400 600.400 232.600 ;
        RECT 564.500 229.700 568.400 230.300 ;
        RECT 567.600 226.200 568.400 229.700 ;
        RECT 572.400 230.300 573.200 230.400 ;
        RECT 577.000 230.300 577.800 231.200 ;
        RECT 578.600 230.600 579.200 232.400 ;
        RECT 572.400 229.700 577.800 230.300 ;
        RECT 572.400 229.600 573.200 229.700 ;
        RECT 569.200 226.800 570.000 228.400 ;
        RECT 577.000 226.800 577.800 229.700 ;
        RECT 578.400 230.000 579.200 230.600 ;
        RECT 585.200 230.000 608.600 230.600 ;
        RECT 578.400 228.000 579.000 230.000 ;
        RECT 585.200 229.400 586.000 230.000 ;
        RECT 602.800 229.600 603.600 230.000 ;
        RECT 607.600 229.800 608.600 230.000 ;
        RECT 607.600 229.600 608.400 229.800 ;
        RECT 579.600 228.600 583.400 229.400 ;
        RECT 578.400 227.400 579.600 228.000 ;
        RECT 554.800 222.200 555.600 226.200 ;
        RECT 556.400 226.000 560.400 226.200 ;
        RECT 556.400 222.200 557.200 226.000 ;
        RECT 559.600 222.200 560.400 226.000 ;
        RECT 562.800 225.600 564.600 226.200 ;
        RECT 563.800 224.400 564.600 225.600 ;
        RECT 562.800 223.600 564.600 224.400 ;
        RECT 563.800 222.200 564.600 223.600 ;
        RECT 566.600 225.600 568.400 226.200 ;
        RECT 577.000 226.000 578.000 226.800 ;
        RECT 566.600 222.200 567.400 225.600 ;
        RECT 577.200 222.200 578.000 226.000 ;
        RECT 578.800 222.200 579.600 227.400 ;
        RECT 582.600 227.400 583.400 228.600 ;
        RECT 582.600 226.800 584.400 227.400 ;
        RECT 583.600 226.200 584.400 226.800 ;
        RECT 588.400 226.400 589.200 229.200 ;
        RECT 591.600 228.600 594.800 229.400 ;
        RECT 598.600 228.600 600.600 229.400 ;
        RECT 609.200 229.000 610.000 234.600 ;
        RECT 591.200 227.800 592.000 228.000 ;
        RECT 591.200 227.200 595.600 227.800 ;
        RECT 594.800 227.000 595.600 227.200 ;
        RECT 596.400 226.800 597.200 228.400 ;
        RECT 583.600 225.400 586.000 226.200 ;
        RECT 588.400 225.600 589.400 226.400 ;
        RECT 592.400 225.600 594.000 226.400 ;
        RECT 594.800 226.200 595.600 226.400 ;
        RECT 598.600 226.200 599.400 228.600 ;
        RECT 601.200 228.200 610.000 229.000 ;
        RECT 604.600 226.800 607.600 227.600 ;
        RECT 604.600 226.200 605.400 226.800 ;
        RECT 594.800 225.600 599.400 226.200 ;
        RECT 585.200 222.200 586.000 225.400 ;
        RECT 602.800 225.400 605.400 226.200 ;
        RECT 586.800 222.200 587.600 225.000 ;
        RECT 588.400 222.200 589.200 225.000 ;
        RECT 590.000 222.200 590.800 225.000 ;
        RECT 591.600 222.200 592.400 225.000 ;
        RECT 594.800 222.200 595.600 225.000 ;
        RECT 598.000 222.200 598.800 225.000 ;
        RECT 599.600 222.200 600.400 225.000 ;
        RECT 601.200 222.200 602.000 225.000 ;
        RECT 602.800 222.200 603.600 225.400 ;
        RECT 609.200 222.200 610.000 228.200 ;
        RECT 610.800 231.200 611.600 239.800 ;
        RECT 615.000 235.800 616.200 239.800 ;
        RECT 619.600 235.800 620.400 239.800 ;
        RECT 624.000 236.400 624.800 239.800 ;
        RECT 624.000 235.800 626.000 236.400 ;
        RECT 615.600 235.000 616.400 235.800 ;
        RECT 619.800 235.200 620.400 235.800 ;
        RECT 619.000 234.600 622.600 235.200 ;
        RECT 625.200 235.000 626.000 235.800 ;
        RECT 619.000 234.400 619.800 234.600 ;
        RECT 621.800 234.400 622.600 234.600 ;
        RECT 614.800 233.200 616.200 234.000 ;
        RECT 615.600 232.200 616.200 233.200 ;
        RECT 617.800 233.000 620.000 233.600 ;
        RECT 617.800 232.800 618.600 233.000 ;
        RECT 615.600 231.600 618.000 232.200 ;
        RECT 610.800 230.600 615.000 231.200 ;
        RECT 610.800 227.200 611.600 230.600 ;
        RECT 614.200 230.400 615.000 230.600 ;
        RECT 617.400 230.300 618.000 231.600 ;
        RECT 619.400 231.800 620.000 233.000 ;
        RECT 620.600 233.000 621.400 233.200 ;
        RECT 625.200 233.000 626.000 233.200 ;
        RECT 620.600 232.400 626.000 233.000 ;
        RECT 619.400 231.400 624.200 231.800 ;
        RECT 628.400 231.400 629.200 239.800 ;
        RECT 631.600 236.400 632.400 239.800 ;
        RECT 631.400 235.800 632.400 236.400 ;
        RECT 631.400 235.200 632.000 235.800 ;
        RECT 634.800 235.200 635.600 239.800 ;
        RECT 638.000 237.000 638.800 239.800 ;
        RECT 639.600 237.000 640.400 239.800 ;
        RECT 619.400 231.200 629.200 231.400 ;
        RECT 623.400 231.000 629.200 231.200 ;
        RECT 623.600 230.800 629.200 231.000 ;
        RECT 630.000 234.600 632.000 235.200 ;
        RECT 618.800 230.300 619.600 230.400 ;
        RECT 612.600 229.800 613.400 230.000 ;
        RECT 612.600 229.200 616.400 229.800 ;
        RECT 617.300 229.700 619.600 230.300 ;
        RECT 615.600 229.000 616.400 229.200 ;
        RECT 617.400 228.400 618.000 229.700 ;
        RECT 618.800 229.600 619.600 229.700 ;
        RECT 622.000 230.200 622.800 230.400 ;
        RECT 622.000 229.600 627.000 230.200 ;
        RECT 623.600 229.400 624.400 229.600 ;
        RECT 626.200 229.400 627.000 229.600 ;
        RECT 630.000 229.000 630.800 234.600 ;
        RECT 632.600 234.400 636.800 235.200 ;
        RECT 641.200 235.000 642.000 239.800 ;
        RECT 644.400 235.000 645.200 239.800 ;
        RECT 632.600 234.000 633.200 234.400 ;
        RECT 631.600 233.200 633.200 234.000 ;
        RECT 636.200 233.800 642.000 234.400 ;
        RECT 634.200 233.200 635.600 233.800 ;
        RECT 634.200 233.000 640.400 233.200 ;
        RECT 635.000 232.600 640.400 233.000 ;
        RECT 639.600 232.400 640.400 232.600 ;
        RECT 641.400 233.000 642.000 233.800 ;
        RECT 642.600 233.600 645.200 234.400 ;
        RECT 647.600 233.600 648.400 239.800 ;
        RECT 649.200 237.000 650.000 239.800 ;
        RECT 650.800 237.000 651.600 239.800 ;
        RECT 652.400 237.000 653.200 239.800 ;
        RECT 650.800 234.400 655.000 235.200 ;
        RECT 655.600 234.400 656.400 239.800 ;
        RECT 658.800 235.200 659.600 239.800 ;
        RECT 658.800 234.600 661.400 235.200 ;
        RECT 655.600 233.600 658.200 234.400 ;
        RECT 649.200 233.000 650.000 233.200 ;
        RECT 641.400 232.400 650.000 233.000 ;
        RECT 652.400 233.000 653.200 233.200 ;
        RECT 660.800 233.000 661.400 234.600 ;
        RECT 652.400 232.400 661.400 233.000 ;
        RECT 660.800 230.600 661.400 232.400 ;
        RECT 662.000 232.000 662.800 239.800 ;
        RECT 662.000 231.200 663.000 232.000 ;
        RECT 631.400 230.000 654.800 230.600 ;
        RECT 660.800 230.000 661.600 230.600 ;
        RECT 631.400 229.800 632.200 230.000 ;
        RECT 633.200 229.600 634.000 230.000 ;
        RECT 636.400 229.600 637.200 230.000 ;
        RECT 654.000 229.400 654.800 230.000 ;
        RECT 624.600 228.400 625.400 228.600 ;
        RECT 617.400 227.800 628.400 228.400 ;
        RECT 617.800 227.600 618.600 227.800 ;
        RECT 610.800 226.600 614.600 227.200 ;
        RECT 610.800 222.200 611.600 226.600 ;
        RECT 613.800 226.400 614.600 226.600 ;
        RECT 623.600 225.600 624.200 227.800 ;
        RECT 626.800 227.600 628.400 227.800 ;
        RECT 630.000 228.200 638.800 229.000 ;
        RECT 639.400 228.600 641.400 229.400 ;
        RECT 645.200 228.600 648.400 229.400 ;
        RECT 621.800 225.400 622.600 225.600 ;
        RECT 615.600 224.200 616.400 225.000 ;
        RECT 619.800 224.800 622.600 225.400 ;
        RECT 623.600 224.800 624.400 225.600 ;
        RECT 619.800 224.200 620.400 224.800 ;
        RECT 625.200 224.200 626.000 225.000 ;
        RECT 615.000 223.600 616.400 224.200 ;
        RECT 615.000 222.200 616.200 223.600 ;
        RECT 619.600 222.200 620.400 224.200 ;
        RECT 624.000 223.600 626.000 224.200 ;
        RECT 624.000 222.200 624.800 223.600 ;
        RECT 628.400 222.200 629.200 227.000 ;
        RECT 630.000 222.200 630.800 228.200 ;
        RECT 632.400 226.800 635.400 227.600 ;
        RECT 634.600 226.200 635.400 226.800 ;
        RECT 640.600 226.200 641.400 228.600 ;
        RECT 642.800 226.800 643.600 228.400 ;
        RECT 648.000 227.800 648.800 228.000 ;
        RECT 644.400 227.200 648.800 227.800 ;
        RECT 644.400 227.000 645.200 227.200 ;
        RECT 650.800 226.400 651.600 229.200 ;
        RECT 656.600 228.600 660.400 229.400 ;
        RECT 656.600 227.400 657.400 228.600 ;
        RECT 661.000 228.000 661.600 230.000 ;
        RECT 644.400 226.200 645.200 226.400 ;
        RECT 634.600 225.400 637.200 226.200 ;
        RECT 640.600 225.600 645.200 226.200 ;
        RECT 646.000 225.600 647.600 226.400 ;
        RECT 650.600 225.600 651.600 226.400 ;
        RECT 655.600 226.800 657.400 227.400 ;
        RECT 660.400 227.400 661.600 228.000 ;
        RECT 655.600 226.200 656.400 226.800 ;
        RECT 636.400 222.200 637.200 225.400 ;
        RECT 654.000 225.400 656.400 226.200 ;
        RECT 638.000 222.200 638.800 225.000 ;
        RECT 639.600 222.200 640.400 225.000 ;
        RECT 641.200 222.200 642.000 225.000 ;
        RECT 644.400 222.200 645.200 225.000 ;
        RECT 647.600 222.200 648.400 225.000 ;
        RECT 649.200 222.200 650.000 225.000 ;
        RECT 650.800 222.200 651.600 225.000 ;
        RECT 652.400 222.200 653.200 225.000 ;
        RECT 654.000 222.200 654.800 225.400 ;
        RECT 660.400 222.200 661.200 227.400 ;
        RECT 662.200 226.800 663.000 231.200 ;
        RECT 662.000 226.000 663.000 226.800 ;
        RECT 663.600 226.300 664.400 226.400 ;
        RECT 665.200 226.300 666.000 226.400 ;
        RECT 662.000 222.200 662.800 226.000 ;
        RECT 663.600 225.700 666.000 226.300 ;
        RECT 663.600 225.600 664.400 225.700 ;
        RECT 665.200 224.800 666.000 225.700 ;
        RECT 666.800 222.200 667.600 239.800 ;
        RECT 668.400 231.400 669.200 239.800 ;
        RECT 672.800 236.400 673.600 239.800 ;
        RECT 671.600 235.800 673.600 236.400 ;
        RECT 677.200 235.800 678.000 239.800 ;
        RECT 681.400 235.800 682.600 239.800 ;
        RECT 671.600 235.000 672.400 235.800 ;
        RECT 677.200 235.200 677.800 235.800 ;
        RECT 675.000 234.600 678.600 235.200 ;
        RECT 681.200 235.000 682.000 235.800 ;
        RECT 675.000 234.400 675.800 234.600 ;
        RECT 677.800 234.400 678.600 234.600 ;
        RECT 671.600 233.000 672.400 233.200 ;
        RECT 676.200 233.000 677.000 233.200 ;
        RECT 671.600 232.400 677.000 233.000 ;
        RECT 677.600 233.000 679.800 233.600 ;
        RECT 677.600 231.800 678.200 233.000 ;
        RECT 679.000 232.800 679.800 233.000 ;
        RECT 681.400 233.200 682.800 234.000 ;
        RECT 681.400 232.200 682.000 233.200 ;
        RECT 673.400 231.400 678.200 231.800 ;
        RECT 668.400 231.200 678.200 231.400 ;
        RECT 679.600 231.600 682.000 232.200 ;
        RECT 668.400 231.000 674.200 231.200 ;
        RECT 668.400 230.800 674.000 231.000 ;
        RECT 674.800 230.200 675.600 230.400 ;
        RECT 670.600 229.600 675.600 230.200 ;
        RECT 670.600 229.400 671.400 229.600 ;
        RECT 672.200 228.400 673.000 228.600 ;
        RECT 679.600 228.400 680.200 231.600 ;
        RECT 686.000 231.200 686.800 239.800 ;
        RECT 682.600 230.600 686.800 231.200 ;
        RECT 682.600 230.400 683.400 230.600 ;
        RECT 684.200 229.800 685.000 230.000 ;
        RECT 681.200 229.200 685.000 229.800 ;
        RECT 681.200 229.000 682.000 229.200 ;
        RECT 669.200 227.800 680.200 228.400 ;
        RECT 669.200 227.600 670.800 227.800 ;
        RECT 668.400 222.200 669.200 227.000 ;
        RECT 673.400 225.600 674.000 227.800 ;
        RECT 674.800 227.600 675.600 227.800 ;
        RECT 679.000 227.600 679.800 227.800 ;
        RECT 686.000 227.200 686.800 230.600 ;
        RECT 683.000 226.600 686.800 227.200 ;
        RECT 683.000 226.400 683.800 226.600 ;
        RECT 671.600 224.200 672.400 225.000 ;
        RECT 673.200 224.800 674.000 225.600 ;
        RECT 675.000 225.400 675.800 225.600 ;
        RECT 675.000 224.800 677.800 225.400 ;
        RECT 677.200 224.200 677.800 224.800 ;
        RECT 681.200 224.200 682.000 225.000 ;
        RECT 671.600 223.600 673.600 224.200 ;
        RECT 672.800 222.200 673.600 223.600 ;
        RECT 677.200 222.200 678.000 224.200 ;
        RECT 681.200 223.600 682.600 224.200 ;
        RECT 681.400 222.200 682.600 223.600 ;
        RECT 686.000 222.200 686.800 226.600 ;
        RECT 2.800 214.300 3.600 219.800 ;
        RECT 4.400 216.000 5.200 219.800 ;
        RECT 7.600 216.000 8.400 219.800 ;
        RECT 4.400 215.800 8.400 216.000 ;
        RECT 9.200 215.800 10.000 219.800 ;
        RECT 4.600 215.400 8.200 215.800 ;
        RECT 5.200 214.400 6.000 214.800 ;
        RECT 9.200 214.400 9.800 215.800 ;
        RECT 4.400 214.300 6.000 214.400 ;
        RECT 2.800 213.800 6.000 214.300 ;
        RECT 2.800 213.700 5.200 213.800 ;
        RECT 2.800 202.200 3.600 213.700 ;
        RECT 4.400 213.600 5.200 213.700 ;
        RECT 7.400 213.600 10.000 214.400 ;
        RECT 10.800 213.800 11.600 219.800 ;
        RECT 17.200 216.600 18.000 219.800 ;
        RECT 18.800 217.000 19.600 219.800 ;
        RECT 20.400 217.000 21.200 219.800 ;
        RECT 22.000 217.000 22.800 219.800 ;
        RECT 25.200 217.000 26.000 219.800 ;
        RECT 28.400 217.000 29.200 219.800 ;
        RECT 30.000 217.000 30.800 219.800 ;
        RECT 31.600 217.000 32.400 219.800 ;
        RECT 33.200 217.000 34.000 219.800 ;
        RECT 15.400 215.800 18.000 216.600 ;
        RECT 34.800 216.600 35.600 219.800 ;
        RECT 21.400 215.800 26.000 216.400 ;
        RECT 15.400 215.200 16.200 215.800 ;
        RECT 13.200 214.400 16.200 215.200 ;
        RECT 6.000 211.600 6.800 213.200 ;
        RECT 7.400 210.200 8.000 213.600 ;
        RECT 10.800 213.000 19.600 213.800 ;
        RECT 21.400 213.400 22.200 215.800 ;
        RECT 25.200 215.600 26.000 215.800 ;
        RECT 26.800 215.600 28.400 216.400 ;
        RECT 31.400 215.600 32.400 216.400 ;
        RECT 34.800 215.800 37.200 216.600 ;
        RECT 23.600 213.600 24.400 215.200 ;
        RECT 25.200 214.800 26.000 215.000 ;
        RECT 25.200 214.200 29.600 214.800 ;
        RECT 28.800 214.000 29.600 214.200 ;
        RECT 9.200 210.200 10.000 210.400 ;
        RECT 7.000 209.600 8.000 210.200 ;
        RECT 8.600 209.600 10.000 210.200 ;
        RECT 7.000 202.200 7.800 209.600 ;
        RECT 8.600 208.400 9.200 209.600 ;
        RECT 8.400 207.600 9.200 208.400 ;
        RECT 10.800 207.400 11.600 213.000 ;
        RECT 20.200 212.600 22.200 213.400 ;
        RECT 26.000 212.600 29.200 213.400 ;
        RECT 31.600 212.800 32.400 215.600 ;
        RECT 36.400 215.200 37.200 215.800 ;
        RECT 36.400 214.600 38.200 215.200 ;
        RECT 37.400 213.400 38.200 214.600 ;
        RECT 41.200 214.600 42.000 219.800 ;
        RECT 42.800 216.000 43.600 219.800 ;
        RECT 42.800 215.200 43.800 216.000 ;
        RECT 47.600 215.200 48.400 219.800 ;
        RECT 50.800 215.200 51.600 219.800 ;
        RECT 54.000 215.200 54.800 219.800 ;
        RECT 57.200 215.200 58.000 219.800 ;
        RECT 62.000 216.000 62.800 219.800 ;
        RECT 41.200 214.000 42.400 214.600 ;
        RECT 37.400 212.600 41.200 213.400 ;
        RECT 12.200 212.000 13.000 212.200 ;
        RECT 17.200 212.000 18.000 212.400 ;
        RECT 23.600 212.000 24.400 212.400 ;
        RECT 34.800 212.000 35.600 212.600 ;
        RECT 41.800 212.000 42.400 214.000 ;
        RECT 12.200 211.400 35.600 212.000 ;
        RECT 41.600 211.400 42.400 212.000 ;
        RECT 41.600 209.600 42.200 211.400 ;
        RECT 43.000 210.800 43.800 215.200 ;
        RECT 46.000 214.400 48.400 215.200 ;
        RECT 49.400 214.400 51.600 215.200 ;
        RECT 52.600 214.400 54.800 215.200 ;
        RECT 56.200 214.400 58.000 215.200 ;
        RECT 61.800 215.200 62.800 216.000 ;
        RECT 46.000 211.600 46.800 214.400 ;
        RECT 49.400 213.800 50.200 214.400 ;
        RECT 52.600 213.800 53.400 214.400 ;
        RECT 56.200 213.800 57.000 214.400 ;
        RECT 58.800 213.800 59.600 214.400 ;
        RECT 47.600 213.000 50.200 213.800 ;
        RECT 51.000 213.000 53.400 213.800 ;
        RECT 54.400 213.000 57.000 213.800 ;
        RECT 57.800 213.000 59.600 213.800 ;
        RECT 49.400 211.600 50.200 213.000 ;
        RECT 52.600 211.600 53.400 213.000 ;
        RECT 56.200 211.600 57.000 213.000 ;
        RECT 46.000 210.800 48.400 211.600 ;
        RECT 49.400 210.800 51.600 211.600 ;
        RECT 52.600 210.800 54.800 211.600 ;
        RECT 56.200 210.800 58.000 211.600 ;
        RECT 20.400 209.400 21.200 209.600 ;
        RECT 15.800 209.000 21.200 209.400 ;
        RECT 15.000 208.800 21.200 209.000 ;
        RECT 22.200 209.000 30.800 209.600 ;
        RECT 12.400 208.000 14.000 208.800 ;
        RECT 15.000 208.200 16.400 208.800 ;
        RECT 22.200 208.200 22.800 209.000 ;
        RECT 30.000 208.800 30.800 209.000 ;
        RECT 33.200 209.000 42.200 209.600 ;
        RECT 33.200 208.800 34.000 209.000 ;
        RECT 13.400 207.600 14.000 208.000 ;
        RECT 17.000 207.600 22.800 208.200 ;
        RECT 23.400 207.600 26.000 208.400 ;
        RECT 10.800 206.800 12.800 207.400 ;
        RECT 13.400 206.800 17.600 207.600 ;
        RECT 12.200 206.200 12.800 206.800 ;
        RECT 12.200 205.600 13.200 206.200 ;
        RECT 12.400 202.200 13.200 205.600 ;
        RECT 15.600 202.200 16.400 206.800 ;
        RECT 18.800 202.200 19.600 205.000 ;
        RECT 20.400 202.200 21.200 205.000 ;
        RECT 22.000 202.200 22.800 207.000 ;
        RECT 25.200 202.200 26.000 207.000 ;
        RECT 28.400 202.200 29.200 208.400 ;
        RECT 36.400 207.600 39.000 208.400 ;
        RECT 31.600 206.800 35.800 207.600 ;
        RECT 30.000 202.200 30.800 205.000 ;
        RECT 31.600 202.200 32.400 205.000 ;
        RECT 33.200 202.200 34.000 205.000 ;
        RECT 36.400 202.200 37.200 207.600 ;
        RECT 41.600 207.400 42.200 209.000 ;
        RECT 39.600 206.800 42.200 207.400 ;
        RECT 42.800 210.000 43.800 210.800 ;
        RECT 39.600 202.200 40.400 206.800 ;
        RECT 42.800 202.200 43.600 210.000 ;
        RECT 47.600 202.200 48.400 210.800 ;
        RECT 50.800 202.200 51.600 210.800 ;
        RECT 54.000 202.200 54.800 210.800 ;
        RECT 57.200 202.200 58.000 210.800 ;
        RECT 61.800 210.800 62.600 215.200 ;
        RECT 63.600 214.600 64.400 219.800 ;
        RECT 70.000 216.600 70.800 219.800 ;
        RECT 71.600 217.000 72.400 219.800 ;
        RECT 73.200 217.000 74.000 219.800 ;
        RECT 74.800 217.000 75.600 219.800 ;
        RECT 76.400 217.000 77.200 219.800 ;
        RECT 79.600 217.000 80.400 219.800 ;
        RECT 82.800 217.000 83.600 219.800 ;
        RECT 84.400 217.000 85.200 219.800 ;
        RECT 86.000 217.000 86.800 219.800 ;
        RECT 68.400 215.800 70.800 216.600 ;
        RECT 87.600 216.600 88.400 219.800 ;
        RECT 68.400 215.200 69.200 215.800 ;
        RECT 63.200 214.000 64.400 214.600 ;
        RECT 67.400 214.600 69.200 215.200 ;
        RECT 73.200 215.600 74.200 216.400 ;
        RECT 77.200 215.600 78.800 216.400 ;
        RECT 79.600 215.800 84.200 216.400 ;
        RECT 87.600 215.800 90.200 216.600 ;
        RECT 79.600 215.600 80.400 215.800 ;
        RECT 63.200 212.000 63.800 214.000 ;
        RECT 67.400 213.400 68.200 214.600 ;
        RECT 64.400 212.600 68.200 213.400 ;
        RECT 73.200 212.800 74.000 215.600 ;
        RECT 79.600 214.800 80.400 215.000 ;
        RECT 76.000 214.200 80.400 214.800 ;
        RECT 76.000 214.000 76.800 214.200 ;
        RECT 81.200 213.600 82.000 215.200 ;
        RECT 83.400 213.400 84.200 215.800 ;
        RECT 89.400 215.200 90.200 215.800 ;
        RECT 89.400 214.400 92.400 215.200 ;
        RECT 94.000 213.800 94.800 219.800 ;
        RECT 97.200 215.200 98.000 219.800 ;
        RECT 100.400 215.200 101.200 219.800 ;
        RECT 103.600 215.200 104.400 219.800 ;
        RECT 106.800 215.200 107.600 219.800 ;
        RECT 97.200 214.400 99.000 215.200 ;
        RECT 100.400 214.400 102.600 215.200 ;
        RECT 103.600 214.400 105.800 215.200 ;
        RECT 106.800 214.400 109.200 215.200 ;
        RECT 76.400 212.600 79.600 213.400 ;
        RECT 83.400 212.600 85.400 213.400 ;
        RECT 86.000 213.000 94.800 213.800 ;
        RECT 95.600 213.800 96.400 214.400 ;
        RECT 98.200 213.800 99.000 214.400 ;
        RECT 101.800 213.800 102.600 214.400 ;
        RECT 105.000 213.800 105.800 214.400 ;
        RECT 95.600 213.000 97.400 213.800 ;
        RECT 98.200 213.000 100.800 213.800 ;
        RECT 101.800 213.000 104.200 213.800 ;
        RECT 105.000 213.000 107.600 213.800 ;
        RECT 70.000 212.000 70.800 212.600 ;
        RECT 87.600 212.000 88.400 212.400 ;
        RECT 90.800 212.000 91.600 212.400 ;
        RECT 92.600 212.000 93.400 212.200 ;
        RECT 63.200 211.400 64.000 212.000 ;
        RECT 70.000 211.400 93.400 212.000 ;
        RECT 61.800 210.000 62.800 210.800 ;
        RECT 62.000 202.200 62.800 210.000 ;
        RECT 63.400 209.600 64.000 211.400 ;
        RECT 63.400 209.000 72.400 209.600 ;
        RECT 63.400 207.400 64.000 209.000 ;
        RECT 71.600 208.800 72.400 209.000 ;
        RECT 74.800 209.000 83.400 209.600 ;
        RECT 74.800 208.800 75.600 209.000 ;
        RECT 66.600 207.600 69.200 208.400 ;
        RECT 63.400 206.800 66.000 207.400 ;
        RECT 65.200 202.200 66.000 206.800 ;
        RECT 68.400 202.200 69.200 207.600 ;
        RECT 69.800 206.800 74.000 207.600 ;
        RECT 71.600 202.200 72.400 205.000 ;
        RECT 73.200 202.200 74.000 205.000 ;
        RECT 74.800 202.200 75.600 205.000 ;
        RECT 76.400 202.200 77.200 208.400 ;
        RECT 79.600 207.600 82.200 208.400 ;
        RECT 82.800 208.200 83.400 209.000 ;
        RECT 84.400 209.400 85.200 209.600 ;
        RECT 84.400 209.000 89.800 209.400 ;
        RECT 84.400 208.800 90.600 209.000 ;
        RECT 89.200 208.200 90.600 208.800 ;
        RECT 82.800 207.600 88.600 208.200 ;
        RECT 91.600 208.000 93.200 208.800 ;
        RECT 91.600 207.600 92.200 208.000 ;
        RECT 79.600 202.200 80.400 207.000 ;
        RECT 82.800 202.200 83.600 207.000 ;
        RECT 88.000 206.800 92.200 207.600 ;
        RECT 94.000 207.400 94.800 213.000 ;
        RECT 98.200 211.600 99.000 213.000 ;
        RECT 101.800 211.600 102.600 213.000 ;
        RECT 105.000 211.600 105.800 213.000 ;
        RECT 108.400 211.600 109.200 214.400 ;
        RECT 92.800 206.800 94.800 207.400 ;
        RECT 97.200 210.800 99.000 211.600 ;
        RECT 100.400 210.800 102.600 211.600 ;
        RECT 103.600 210.800 105.800 211.600 ;
        RECT 106.800 210.800 109.200 211.600 ;
        RECT 84.400 202.200 85.200 205.000 ;
        RECT 86.000 202.200 86.800 205.000 ;
        RECT 89.200 202.200 90.000 206.800 ;
        RECT 92.800 206.200 93.400 206.800 ;
        RECT 92.400 205.600 93.400 206.200 ;
        RECT 92.400 202.200 93.200 205.600 ;
        RECT 97.200 202.200 98.000 210.800 ;
        RECT 100.400 202.200 101.200 210.800 ;
        RECT 103.600 202.200 104.400 210.800 ;
        RECT 106.800 202.200 107.600 210.800 ;
        RECT 114.800 208.300 115.600 219.800 ;
        RECT 116.400 216.300 117.200 217.200 ;
        RECT 119.600 216.300 120.400 219.800 ;
        RECT 116.400 215.700 120.400 216.300 ;
        RECT 116.400 215.600 117.200 215.700 ;
        RECT 119.400 215.200 120.400 215.700 ;
        RECT 119.400 210.800 120.200 215.200 ;
        RECT 121.200 214.600 122.000 219.800 ;
        RECT 127.600 216.600 128.400 219.800 ;
        RECT 129.200 217.000 130.000 219.800 ;
        RECT 130.800 217.000 131.600 219.800 ;
        RECT 132.400 217.000 133.200 219.800 ;
        RECT 134.000 217.000 134.800 219.800 ;
        RECT 137.200 217.000 138.000 219.800 ;
        RECT 140.400 217.000 141.200 219.800 ;
        RECT 142.000 217.000 142.800 219.800 ;
        RECT 143.600 217.000 144.400 219.800 ;
        RECT 126.000 215.800 128.400 216.600 ;
        RECT 145.200 216.600 146.000 219.800 ;
        RECT 126.000 215.200 126.800 215.800 ;
        RECT 120.800 214.000 122.000 214.600 ;
        RECT 125.000 214.600 126.800 215.200 ;
        RECT 130.800 215.600 131.800 216.400 ;
        RECT 134.800 215.600 136.400 216.400 ;
        RECT 137.200 215.800 141.800 216.400 ;
        RECT 145.200 215.800 147.800 216.600 ;
        RECT 137.200 215.600 138.000 215.800 ;
        RECT 120.800 212.000 121.400 214.000 ;
        RECT 125.000 213.400 125.800 214.600 ;
        RECT 122.000 212.600 125.800 213.400 ;
        RECT 130.800 212.800 131.600 215.600 ;
        RECT 137.200 214.800 138.000 215.000 ;
        RECT 133.600 214.200 138.000 214.800 ;
        RECT 133.600 214.000 134.400 214.200 ;
        RECT 138.800 213.600 139.600 215.200 ;
        RECT 141.000 213.400 141.800 215.800 ;
        RECT 147.000 215.200 147.800 215.800 ;
        RECT 147.000 214.400 150.000 215.200 ;
        RECT 151.600 213.800 152.400 219.800 ;
        RECT 154.800 216.000 155.600 219.800 ;
        RECT 134.000 212.600 137.200 213.400 ;
        RECT 141.000 212.600 143.000 213.400 ;
        RECT 143.600 213.000 152.400 213.800 ;
        RECT 127.600 212.000 128.400 212.600 ;
        RECT 145.200 212.000 146.000 212.400 ;
        RECT 148.400 212.000 149.200 212.400 ;
        RECT 150.200 212.000 151.000 212.200 ;
        RECT 120.800 211.400 121.600 212.000 ;
        RECT 127.600 211.400 151.000 212.000 ;
        RECT 119.400 210.000 120.400 210.800 ;
        RECT 118.000 208.300 118.800 208.400 ;
        RECT 114.800 207.700 118.800 208.300 ;
        RECT 114.800 202.200 115.600 207.700 ;
        RECT 118.000 207.600 118.800 207.700 ;
        RECT 119.600 202.200 120.400 210.000 ;
        RECT 121.000 209.600 121.600 211.400 ;
        RECT 121.000 209.000 130.000 209.600 ;
        RECT 121.000 207.400 121.600 209.000 ;
        RECT 129.200 208.800 130.000 209.000 ;
        RECT 132.400 209.000 141.000 209.600 ;
        RECT 132.400 208.800 133.200 209.000 ;
        RECT 124.200 207.600 126.800 208.400 ;
        RECT 121.000 206.800 123.600 207.400 ;
        RECT 122.800 202.200 123.600 206.800 ;
        RECT 126.000 202.200 126.800 207.600 ;
        RECT 127.400 206.800 131.600 207.600 ;
        RECT 129.200 202.200 130.000 205.000 ;
        RECT 130.800 202.200 131.600 205.000 ;
        RECT 132.400 202.200 133.200 205.000 ;
        RECT 134.000 202.200 134.800 208.400 ;
        RECT 137.200 207.600 139.800 208.400 ;
        RECT 140.400 208.200 141.000 209.000 ;
        RECT 142.000 209.400 142.800 209.600 ;
        RECT 142.000 209.000 147.400 209.400 ;
        RECT 142.000 208.800 148.200 209.000 ;
        RECT 146.800 208.200 148.200 208.800 ;
        RECT 140.400 207.600 146.200 208.200 ;
        RECT 149.200 208.000 150.800 208.800 ;
        RECT 149.200 207.600 149.800 208.000 ;
        RECT 137.200 202.200 138.000 207.000 ;
        RECT 140.400 202.200 141.200 207.000 ;
        RECT 145.600 206.800 149.800 207.600 ;
        RECT 151.600 207.400 152.400 213.000 ;
        RECT 154.600 215.200 155.600 216.000 ;
        RECT 154.600 210.800 155.400 215.200 ;
        RECT 156.400 214.600 157.200 219.800 ;
        RECT 162.800 216.600 163.600 219.800 ;
        RECT 164.400 217.000 165.200 219.800 ;
        RECT 166.000 217.000 166.800 219.800 ;
        RECT 167.600 217.000 168.400 219.800 ;
        RECT 169.200 217.000 170.000 219.800 ;
        RECT 172.400 217.000 173.200 219.800 ;
        RECT 175.600 217.000 176.400 219.800 ;
        RECT 177.200 217.000 178.000 219.800 ;
        RECT 178.800 217.000 179.600 219.800 ;
        RECT 161.200 215.800 163.600 216.600 ;
        RECT 180.400 216.600 181.200 219.800 ;
        RECT 161.200 215.200 162.000 215.800 ;
        RECT 156.000 214.000 157.200 214.600 ;
        RECT 160.200 214.600 162.000 215.200 ;
        RECT 166.000 215.600 167.000 216.400 ;
        RECT 170.000 215.600 171.600 216.400 ;
        RECT 172.400 215.800 177.000 216.400 ;
        RECT 180.400 215.800 183.000 216.600 ;
        RECT 172.400 215.600 173.200 215.800 ;
        RECT 156.000 212.000 156.600 214.000 ;
        RECT 160.200 213.400 161.000 214.600 ;
        RECT 157.200 212.600 161.000 213.400 ;
        RECT 166.000 212.800 166.800 215.600 ;
        RECT 172.400 214.800 173.200 215.000 ;
        RECT 168.800 214.200 173.200 214.800 ;
        RECT 168.800 214.000 169.600 214.200 ;
        RECT 174.000 213.600 174.800 215.200 ;
        RECT 176.200 213.400 177.000 215.800 ;
        RECT 182.200 215.200 183.000 215.800 ;
        RECT 182.200 214.400 185.200 215.200 ;
        RECT 186.800 213.800 187.600 219.800 ;
        RECT 169.200 212.600 172.400 213.400 ;
        RECT 176.200 212.600 178.200 213.400 ;
        RECT 178.800 213.000 187.600 213.800 ;
        RECT 162.800 212.000 163.600 212.600 ;
        RECT 180.400 212.000 181.200 212.400 ;
        RECT 183.600 212.000 184.400 212.400 ;
        RECT 185.400 212.000 186.200 212.200 ;
        RECT 156.000 211.400 156.800 212.000 ;
        RECT 162.800 211.400 186.200 212.000 ;
        RECT 154.600 210.000 155.600 210.800 ;
        RECT 150.400 206.800 152.400 207.400 ;
        RECT 142.000 202.200 142.800 205.000 ;
        RECT 143.600 202.200 144.400 205.000 ;
        RECT 146.800 202.200 147.600 206.800 ;
        RECT 150.400 206.200 151.000 206.800 ;
        RECT 150.000 205.600 151.000 206.200 ;
        RECT 150.000 202.200 150.800 205.600 ;
        RECT 154.800 202.200 155.600 210.000 ;
        RECT 156.200 209.600 156.800 211.400 ;
        RECT 156.200 209.000 165.200 209.600 ;
        RECT 156.200 207.400 156.800 209.000 ;
        RECT 164.400 208.800 165.200 209.000 ;
        RECT 167.600 209.000 176.200 209.600 ;
        RECT 167.600 208.800 168.400 209.000 ;
        RECT 159.400 207.600 162.000 208.400 ;
        RECT 156.200 206.800 158.800 207.400 ;
        RECT 158.000 202.200 158.800 206.800 ;
        RECT 161.200 202.200 162.000 207.600 ;
        RECT 162.600 206.800 166.800 207.600 ;
        RECT 164.400 202.200 165.200 205.000 ;
        RECT 166.000 202.200 166.800 205.000 ;
        RECT 167.600 202.200 168.400 205.000 ;
        RECT 169.200 202.200 170.000 208.400 ;
        RECT 172.400 207.600 175.000 208.400 ;
        RECT 175.600 208.200 176.200 209.000 ;
        RECT 177.200 209.400 178.000 209.600 ;
        RECT 177.200 209.000 182.600 209.400 ;
        RECT 177.200 208.800 183.400 209.000 ;
        RECT 182.000 208.200 183.400 208.800 ;
        RECT 175.600 207.600 181.400 208.200 ;
        RECT 184.400 208.000 186.000 208.800 ;
        RECT 184.400 207.600 185.000 208.000 ;
        RECT 172.400 202.200 173.200 207.000 ;
        RECT 175.600 202.200 176.400 207.000 ;
        RECT 180.800 206.800 185.000 207.600 ;
        RECT 186.800 207.400 187.600 213.000 ;
        RECT 185.600 206.800 187.600 207.400 ;
        RECT 188.400 213.800 189.200 219.800 ;
        RECT 194.800 216.600 195.600 219.800 ;
        RECT 196.400 217.000 197.200 219.800 ;
        RECT 198.000 217.000 198.800 219.800 ;
        RECT 199.600 217.000 200.400 219.800 ;
        RECT 202.800 217.000 203.600 219.800 ;
        RECT 206.000 217.000 206.800 219.800 ;
        RECT 207.600 217.000 208.400 219.800 ;
        RECT 209.200 217.000 210.000 219.800 ;
        RECT 210.800 217.000 211.600 219.800 ;
        RECT 193.000 215.800 195.600 216.600 ;
        RECT 212.400 216.600 213.200 219.800 ;
        RECT 199.000 215.800 203.600 216.400 ;
        RECT 193.000 215.200 193.800 215.800 ;
        RECT 190.800 214.400 193.800 215.200 ;
        RECT 188.400 213.000 197.200 213.800 ;
        RECT 199.000 213.400 199.800 215.800 ;
        RECT 202.800 215.600 203.600 215.800 ;
        RECT 204.400 215.600 206.000 216.400 ;
        RECT 209.000 215.600 210.000 216.400 ;
        RECT 212.400 215.800 214.800 216.600 ;
        RECT 201.200 213.600 202.000 215.200 ;
        RECT 202.800 214.800 203.600 215.000 ;
        RECT 202.800 214.200 207.200 214.800 ;
        RECT 206.400 214.000 207.200 214.200 ;
        RECT 188.400 207.400 189.200 213.000 ;
        RECT 197.800 212.600 199.800 213.400 ;
        RECT 203.600 212.600 206.800 213.400 ;
        RECT 209.200 212.800 210.000 215.600 ;
        RECT 214.000 215.200 214.800 215.800 ;
        RECT 214.000 214.600 215.800 215.200 ;
        RECT 215.000 213.400 215.800 214.600 ;
        RECT 218.800 214.600 219.600 219.800 ;
        RECT 220.400 216.300 221.200 219.800 ;
        RECT 225.200 217.800 226.000 219.800 ;
        RECT 223.600 216.300 224.400 217.200 ;
        RECT 225.400 216.300 226.000 217.800 ;
        RECT 228.600 216.400 229.400 217.200 ;
        RECT 228.400 216.300 229.200 216.400 ;
        RECT 220.400 215.700 224.400 216.300 ;
        RECT 225.300 215.700 229.200 216.300 ;
        RECT 230.000 215.800 230.800 219.800 ;
        RECT 237.400 218.400 238.200 219.800 ;
        RECT 236.400 217.600 238.200 218.400 ;
        RECT 241.200 217.800 242.000 219.800 ;
        RECT 237.400 216.400 238.200 217.600 ;
        RECT 220.400 215.200 221.400 215.700 ;
        RECT 223.600 215.600 224.400 215.700 ;
        RECT 218.800 214.000 220.000 214.600 ;
        RECT 215.000 212.600 218.800 213.400 ;
        RECT 190.000 212.200 190.800 212.400 ;
        RECT 189.800 212.000 190.800 212.200 ;
        RECT 194.800 212.000 195.600 212.400 ;
        RECT 212.400 212.000 213.200 212.600 ;
        RECT 219.400 212.000 220.000 214.000 ;
        RECT 189.800 211.400 213.200 212.000 ;
        RECT 219.200 211.400 220.000 212.000 ;
        RECT 219.200 209.600 219.800 211.400 ;
        RECT 220.600 210.800 221.400 215.200 ;
        RECT 225.400 214.400 226.000 215.700 ;
        RECT 228.400 215.600 229.200 215.700 ;
        RECT 225.200 213.600 226.000 214.400 ;
        RECT 226.800 214.300 227.600 214.400 ;
        RECT 230.200 214.300 230.800 215.800 ;
        RECT 236.400 215.800 238.200 216.400 ;
        RECT 226.800 213.700 230.800 214.300 ;
        RECT 226.800 213.600 227.600 213.700 ;
        RECT 198.000 209.400 198.800 209.600 ;
        RECT 193.400 209.000 198.800 209.400 ;
        RECT 192.600 208.800 198.800 209.000 ;
        RECT 199.800 209.000 208.400 209.600 ;
        RECT 190.000 208.000 191.600 208.800 ;
        RECT 192.600 208.200 194.000 208.800 ;
        RECT 199.800 208.200 200.400 209.000 ;
        RECT 207.600 208.800 208.400 209.000 ;
        RECT 210.800 209.000 219.800 209.600 ;
        RECT 210.800 208.800 211.600 209.000 ;
        RECT 191.000 207.600 191.600 208.000 ;
        RECT 194.600 207.600 200.400 208.200 ;
        RECT 201.000 207.600 203.600 208.400 ;
        RECT 188.400 206.800 190.400 207.400 ;
        RECT 191.000 206.800 195.200 207.600 ;
        RECT 177.200 202.200 178.000 205.000 ;
        RECT 178.800 202.200 179.600 205.000 ;
        RECT 182.000 202.200 182.800 206.800 ;
        RECT 185.600 206.200 186.200 206.800 ;
        RECT 185.200 205.600 186.200 206.200 ;
        RECT 189.800 206.200 190.400 206.800 ;
        RECT 189.800 205.600 190.800 206.200 ;
        RECT 185.200 202.200 186.000 205.600 ;
        RECT 190.000 202.200 190.800 205.600 ;
        RECT 193.200 202.200 194.000 206.800 ;
        RECT 196.400 202.200 197.200 205.000 ;
        RECT 198.000 202.200 198.800 205.000 ;
        RECT 199.600 202.200 200.400 207.000 ;
        RECT 202.800 202.200 203.600 207.000 ;
        RECT 206.000 202.200 206.800 208.400 ;
        RECT 214.000 207.600 216.600 208.400 ;
        RECT 209.200 206.800 213.400 207.600 ;
        RECT 207.600 202.200 208.400 205.000 ;
        RECT 209.200 202.200 210.000 205.000 ;
        RECT 210.800 202.200 211.600 205.000 ;
        RECT 214.000 202.200 214.800 207.600 ;
        RECT 219.200 207.400 219.800 209.000 ;
        RECT 217.200 206.800 219.800 207.400 ;
        RECT 220.400 210.000 221.400 210.800 ;
        RECT 225.400 210.200 226.000 213.600 ;
        RECT 226.800 210.800 227.600 212.400 ;
        RECT 228.400 212.200 229.200 212.400 ;
        RECT 230.200 212.200 230.800 213.700 ;
        RECT 231.600 212.800 232.400 214.400 ;
        RECT 234.800 213.600 235.600 215.200 ;
        RECT 233.200 212.200 234.000 212.400 ;
        RECT 228.400 211.600 230.800 212.200 ;
        RECT 232.400 211.600 234.000 212.200 ;
        RECT 228.600 210.200 229.200 211.600 ;
        RECT 232.400 211.200 233.200 211.600 ;
        RECT 217.200 202.200 218.000 206.800 ;
        RECT 220.400 202.200 221.200 210.000 ;
        RECT 225.200 209.400 227.000 210.200 ;
        RECT 226.200 202.200 227.000 209.400 ;
        RECT 228.400 202.200 229.200 210.200 ;
        RECT 230.000 209.600 234.000 210.200 ;
        RECT 230.000 202.200 230.800 209.600 ;
        RECT 233.200 202.200 234.000 209.600 ;
        RECT 236.400 202.200 237.200 215.800 ;
        RECT 239.600 215.600 240.400 217.200 ;
        RECT 241.400 214.400 242.000 217.800 ;
        RECT 246.000 216.400 246.800 219.800 ;
        RECT 245.800 215.800 246.800 216.400 ;
        RECT 245.800 214.400 246.400 215.800 ;
        RECT 249.200 215.200 250.000 219.800 ;
        RECT 252.400 216.400 253.200 219.800 ;
        RECT 247.400 214.600 250.000 215.200 ;
        RECT 252.200 215.800 253.200 216.400 ;
        RECT 238.000 214.300 238.800 214.400 ;
        RECT 241.200 214.300 242.000 214.400 ;
        RECT 238.000 213.700 242.000 214.300 ;
        RECT 238.000 213.600 238.800 213.700 ;
        RECT 241.200 213.600 242.000 213.700 ;
        RECT 244.400 214.300 245.200 214.400 ;
        RECT 245.800 214.300 246.800 214.400 ;
        RECT 244.400 213.700 246.800 214.300 ;
        RECT 244.400 213.600 245.200 213.700 ;
        RECT 245.800 213.600 246.800 213.700 ;
        RECT 238.000 208.800 238.800 210.400 ;
        RECT 241.400 210.200 242.000 213.600 ;
        RECT 242.800 210.800 243.600 212.400 ;
        RECT 245.800 210.200 246.400 213.600 ;
        RECT 247.400 213.000 248.000 214.600 ;
        RECT 252.200 214.400 252.800 215.800 ;
        RECT 255.600 215.200 256.400 219.800 ;
        RECT 253.800 214.600 256.400 215.200 ;
        RECT 252.200 213.600 253.200 214.400 ;
        RECT 247.000 212.200 248.000 213.000 ;
        RECT 247.400 210.200 248.000 212.200 ;
        RECT 249.000 212.400 249.800 213.200 ;
        RECT 249.000 211.600 250.000 212.400 ;
        RECT 252.200 210.200 252.800 213.600 ;
        RECT 253.800 213.000 254.400 214.600 ;
        RECT 253.400 212.200 254.400 213.000 ;
        RECT 253.800 210.200 254.400 212.200 ;
        RECT 255.400 212.400 256.200 213.200 ;
        RECT 255.400 211.600 256.400 212.400 ;
        RECT 241.200 209.400 243.000 210.200 ;
        RECT 242.200 202.200 243.000 209.400 ;
        RECT 245.800 209.200 246.800 210.200 ;
        RECT 247.400 209.600 250.000 210.200 ;
        RECT 246.000 202.200 246.800 209.200 ;
        RECT 249.200 202.200 250.000 209.600 ;
        RECT 252.200 209.200 253.200 210.200 ;
        RECT 253.800 209.600 256.400 210.200 ;
        RECT 252.400 202.200 253.200 209.200 ;
        RECT 255.600 202.200 256.400 209.600 ;
        RECT 257.200 202.200 258.000 219.800 ;
        RECT 258.800 215.600 259.600 217.200 ;
        RECT 265.200 213.800 266.000 219.800 ;
        RECT 271.600 216.600 272.400 219.800 ;
        RECT 273.200 217.000 274.000 219.800 ;
        RECT 274.800 217.000 275.600 219.800 ;
        RECT 276.400 217.000 277.200 219.800 ;
        RECT 279.600 217.000 280.400 219.800 ;
        RECT 282.800 217.000 283.600 219.800 ;
        RECT 284.400 217.000 285.200 219.800 ;
        RECT 286.000 217.000 286.800 219.800 ;
        RECT 287.600 217.000 288.400 219.800 ;
        RECT 269.800 215.800 272.400 216.600 ;
        RECT 289.200 216.600 290.000 219.800 ;
        RECT 275.800 215.800 280.400 216.400 ;
        RECT 269.800 215.200 270.600 215.800 ;
        RECT 267.600 214.400 270.600 215.200 ;
        RECT 265.200 213.000 274.000 213.800 ;
        RECT 275.800 213.400 276.600 215.800 ;
        RECT 279.600 215.600 280.400 215.800 ;
        RECT 281.200 215.600 282.800 216.400 ;
        RECT 285.800 215.600 286.800 216.400 ;
        RECT 289.200 215.800 291.600 216.600 ;
        RECT 278.000 213.600 278.800 215.200 ;
        RECT 279.600 214.800 280.400 215.000 ;
        RECT 279.600 214.200 284.000 214.800 ;
        RECT 283.200 214.000 284.000 214.200 ;
        RECT 265.200 207.400 266.000 213.000 ;
        RECT 274.600 212.600 276.600 213.400 ;
        RECT 280.400 212.600 283.600 213.400 ;
        RECT 286.000 212.800 286.800 215.600 ;
        RECT 290.800 215.200 291.600 215.800 ;
        RECT 290.800 214.600 292.600 215.200 ;
        RECT 291.800 213.400 292.600 214.600 ;
        RECT 295.600 214.600 296.400 219.800 ;
        RECT 297.200 216.000 298.000 219.800 ;
        RECT 303.000 218.400 303.800 219.800 ;
        RECT 302.000 217.600 303.800 218.400 ;
        RECT 303.000 216.400 303.800 217.600 ;
        RECT 297.200 215.200 298.200 216.000 ;
        RECT 302.000 215.800 303.800 216.400 ;
        RECT 305.200 216.000 306.000 219.800 ;
        RECT 308.400 216.000 309.200 219.800 ;
        RECT 305.200 215.800 309.200 216.000 ;
        RECT 310.000 215.800 310.800 219.800 ;
        RECT 295.600 214.000 296.800 214.600 ;
        RECT 291.800 212.600 295.600 213.400 ;
        RECT 266.600 212.000 267.400 212.200 ;
        RECT 270.000 212.000 270.800 212.400 ;
        RECT 271.600 212.000 272.400 212.400 ;
        RECT 289.200 212.000 290.000 212.600 ;
        RECT 296.200 212.000 296.800 214.000 ;
        RECT 266.600 211.400 290.000 212.000 ;
        RECT 296.000 211.400 296.800 212.000 ;
        RECT 297.400 212.300 298.200 215.200 ;
        RECT 298.800 214.300 299.600 214.400 ;
        RECT 300.400 214.300 301.200 215.200 ;
        RECT 298.800 213.700 301.200 214.300 ;
        RECT 298.800 213.600 299.600 213.700 ;
        RECT 300.400 213.600 301.200 213.700 ;
        RECT 298.800 212.300 299.600 212.400 ;
        RECT 297.400 211.700 299.600 212.300 ;
        RECT 296.000 209.600 296.600 211.400 ;
        RECT 297.400 210.800 298.200 211.700 ;
        RECT 298.800 211.600 299.600 211.700 ;
        RECT 274.800 209.400 275.600 209.600 ;
        RECT 270.200 209.000 275.600 209.400 ;
        RECT 269.400 208.800 275.600 209.000 ;
        RECT 276.600 209.000 285.200 209.600 ;
        RECT 266.800 208.000 268.400 208.800 ;
        RECT 269.400 208.200 270.800 208.800 ;
        RECT 276.600 208.200 277.200 209.000 ;
        RECT 284.400 208.800 285.200 209.000 ;
        RECT 287.600 209.000 296.600 209.600 ;
        RECT 287.600 208.800 288.400 209.000 ;
        RECT 267.800 207.600 268.400 208.000 ;
        RECT 271.400 207.600 277.200 208.200 ;
        RECT 277.800 207.600 280.400 208.400 ;
        RECT 265.200 206.800 267.200 207.400 ;
        RECT 267.800 206.800 272.000 207.600 ;
        RECT 266.600 206.200 267.200 206.800 ;
        RECT 266.600 205.600 267.600 206.200 ;
        RECT 266.800 202.200 267.600 205.600 ;
        RECT 270.000 202.200 270.800 206.800 ;
        RECT 273.200 202.200 274.000 205.000 ;
        RECT 274.800 202.200 275.600 205.000 ;
        RECT 276.400 202.200 277.200 207.000 ;
        RECT 279.600 202.200 280.400 207.000 ;
        RECT 282.800 202.200 283.600 208.400 ;
        RECT 290.800 207.600 293.400 208.400 ;
        RECT 286.000 206.800 290.200 207.600 ;
        RECT 284.400 202.200 285.200 205.000 ;
        RECT 286.000 202.200 286.800 205.000 ;
        RECT 287.600 202.200 288.400 205.000 ;
        RECT 290.800 202.200 291.600 207.600 ;
        RECT 296.000 207.400 296.600 209.000 ;
        RECT 294.000 206.800 296.600 207.400 ;
        RECT 297.200 210.000 298.200 210.800 ;
        RECT 294.000 202.200 294.800 206.800 ;
        RECT 297.200 202.200 298.000 210.000 ;
        RECT 302.000 202.200 302.800 215.800 ;
        RECT 305.400 215.400 309.000 215.800 ;
        RECT 306.000 214.400 306.800 214.800 ;
        RECT 310.000 214.400 310.600 215.800 ;
        RECT 305.200 213.800 306.800 214.400 ;
        RECT 305.200 213.600 306.000 213.800 ;
        RECT 308.200 213.600 310.800 214.400 ;
        RECT 311.600 213.600 312.400 215.200 ;
        RECT 303.600 212.300 304.400 212.400 ;
        RECT 306.800 212.300 307.600 213.200 ;
        RECT 303.600 211.700 307.600 212.300 ;
        RECT 303.600 211.600 304.400 211.700 ;
        RECT 306.800 211.600 307.600 211.700 ;
        RECT 308.200 210.400 308.800 213.600 ;
        RECT 310.000 212.300 310.800 212.400 ;
        RECT 311.700 212.300 312.300 213.600 ;
        RECT 310.000 211.700 312.300 212.300 ;
        RECT 310.000 211.600 310.800 211.700 ;
        RECT 310.100 210.400 310.700 211.600 ;
        RECT 303.600 208.800 304.400 210.400 ;
        RECT 306.800 209.600 308.800 210.400 ;
        RECT 310.000 210.200 310.800 210.400 ;
        RECT 309.400 209.600 310.800 210.200 ;
        RECT 307.800 202.200 308.600 209.600 ;
        RECT 309.400 208.400 310.000 209.600 ;
        RECT 309.200 207.600 310.000 208.400 ;
        RECT 313.200 202.200 314.000 219.800 ;
        RECT 318.000 202.200 318.800 219.800 ;
        RECT 321.200 215.200 322.000 219.800 ;
        RECT 324.400 216.400 325.200 219.800 ;
        RECT 324.400 215.800 325.400 216.400 ;
        RECT 327.600 215.800 328.400 219.800 ;
        RECT 329.200 216.000 330.000 219.800 ;
        RECT 332.400 216.000 333.200 219.800 ;
        RECT 334.600 216.400 335.400 219.800 ;
        RECT 339.400 216.400 340.200 219.800 ;
        RECT 329.200 215.800 333.200 216.000 ;
        RECT 321.200 214.600 323.800 215.200 ;
        RECT 321.400 212.400 322.200 213.200 ;
        RECT 321.200 211.600 322.200 212.400 ;
        RECT 323.200 213.000 323.800 214.600 ;
        RECT 324.800 214.400 325.400 215.800 ;
        RECT 327.800 214.400 328.400 215.800 ;
        RECT 329.400 215.400 333.000 215.800 ;
        RECT 334.000 215.600 336.400 216.400 ;
        RECT 339.400 215.800 341.200 216.400 ;
        RECT 343.600 216.000 344.400 219.800 ;
        RECT 346.800 216.000 347.600 219.800 ;
        RECT 343.600 215.800 347.600 216.000 ;
        RECT 348.400 215.800 349.200 219.800 ;
        RECT 350.600 218.400 351.400 219.800 ;
        RECT 350.000 217.600 351.400 218.400 ;
        RECT 350.600 216.400 351.400 217.600 ;
        RECT 350.600 215.800 352.400 216.400 ;
        RECT 356.400 216.000 357.200 219.800 ;
        RECT 331.600 214.400 332.400 214.800 ;
        RECT 324.400 213.600 325.400 214.400 ;
        RECT 327.600 213.600 330.200 214.400 ;
        RECT 331.600 213.800 333.200 214.400 ;
        RECT 332.400 213.600 333.200 213.800 ;
        RECT 323.200 212.200 324.200 213.000 ;
        RECT 323.200 210.200 323.800 212.200 ;
        RECT 324.800 210.200 325.400 213.600 ;
        RECT 321.200 209.600 323.800 210.200 ;
        RECT 321.200 202.200 322.000 209.600 ;
        RECT 324.400 209.200 325.400 210.200 ;
        RECT 327.600 210.200 328.400 210.400 ;
        RECT 329.600 210.200 330.200 213.600 ;
        RECT 330.800 211.600 331.600 213.200 ;
        RECT 327.600 209.600 329.000 210.200 ;
        RECT 329.600 209.600 330.600 210.200 ;
        RECT 324.400 202.200 325.200 209.200 ;
        RECT 328.400 208.400 329.000 209.600 ;
        RECT 328.400 207.600 329.200 208.400 ;
        RECT 329.800 204.400 330.600 209.600 ;
        RECT 334.000 208.800 334.800 210.400 ;
        RECT 329.800 203.600 331.600 204.400 ;
        RECT 329.800 202.200 330.600 203.600 ;
        RECT 335.600 202.200 336.400 215.600 ;
        RECT 337.200 213.600 338.000 215.200 ;
        RECT 337.200 212.300 338.000 212.400 ;
        RECT 340.400 212.300 341.200 215.800 ;
        RECT 343.800 215.400 347.400 215.800 ;
        RECT 342.000 213.600 342.800 215.200 ;
        RECT 348.400 214.400 349.000 215.800 ;
        RECT 346.600 213.600 349.200 214.400 ;
        RECT 337.200 211.700 341.200 212.300 ;
        RECT 337.200 211.600 338.000 211.700 ;
        RECT 338.800 208.800 339.600 210.400 ;
        RECT 340.400 202.200 341.200 211.700 ;
        RECT 345.200 211.600 346.000 213.200 ;
        RECT 346.600 210.200 347.200 213.600 ;
        RECT 348.400 210.200 349.200 210.400 ;
        RECT 346.200 209.600 347.200 210.200 ;
        RECT 347.800 209.600 349.200 210.200 ;
        RECT 346.200 204.400 347.000 209.600 ;
        RECT 347.800 208.400 348.400 209.600 ;
        RECT 350.000 208.800 350.800 210.400 ;
        RECT 347.600 207.600 348.400 208.400 ;
        RECT 345.200 203.600 347.000 204.400 ;
        RECT 346.200 202.200 347.000 203.600 ;
        RECT 351.600 202.200 352.400 215.800 ;
        RECT 356.200 215.200 357.200 216.000 ;
        RECT 353.200 214.300 354.000 215.200 ;
        RECT 356.200 214.300 357.000 215.200 ;
        RECT 358.000 214.600 358.800 219.800 ;
        RECT 364.400 216.600 365.200 219.800 ;
        RECT 366.000 217.000 366.800 219.800 ;
        RECT 367.600 217.000 368.400 219.800 ;
        RECT 369.200 217.000 370.000 219.800 ;
        RECT 370.800 217.000 371.600 219.800 ;
        RECT 374.000 217.000 374.800 219.800 ;
        RECT 377.200 217.000 378.000 219.800 ;
        RECT 378.800 217.000 379.600 219.800 ;
        RECT 380.400 217.000 381.200 219.800 ;
        RECT 362.800 215.800 365.200 216.600 ;
        RECT 382.000 216.600 382.800 219.800 ;
        RECT 362.800 215.200 363.600 215.800 ;
        RECT 353.200 213.700 357.000 214.300 ;
        RECT 353.200 213.600 354.000 213.700 ;
        RECT 356.200 210.800 357.000 213.700 ;
        RECT 357.600 214.000 358.800 214.600 ;
        RECT 361.800 214.600 363.600 215.200 ;
        RECT 367.600 215.600 368.600 216.400 ;
        RECT 371.600 215.600 373.200 216.400 ;
        RECT 374.000 215.800 378.600 216.400 ;
        RECT 382.000 215.800 384.600 216.600 ;
        RECT 374.000 215.600 374.800 215.800 ;
        RECT 357.600 212.000 358.200 214.000 ;
        RECT 361.800 213.400 362.600 214.600 ;
        RECT 358.800 212.600 362.600 213.400 ;
        RECT 367.600 212.800 368.400 215.600 ;
        RECT 374.000 214.800 374.800 215.000 ;
        RECT 370.400 214.200 374.800 214.800 ;
        RECT 370.400 214.000 371.200 214.200 ;
        RECT 375.600 213.600 376.400 215.200 ;
        RECT 377.800 213.400 378.600 215.800 ;
        RECT 383.800 215.200 384.600 215.800 ;
        RECT 383.800 214.400 386.800 215.200 ;
        RECT 388.400 213.800 389.200 219.800 ;
        RECT 391.600 216.400 392.400 219.800 ;
        RECT 370.800 212.600 374.000 213.400 ;
        RECT 377.800 212.600 379.800 213.400 ;
        RECT 380.400 213.000 389.200 213.800 ;
        RECT 364.400 212.000 365.200 212.600 ;
        RECT 382.000 212.000 382.800 212.400 ;
        RECT 385.200 212.000 386.000 212.400 ;
        RECT 387.000 212.000 387.800 212.200 ;
        RECT 357.600 211.400 358.400 212.000 ;
        RECT 364.400 211.400 387.800 212.000 ;
        RECT 356.200 210.000 357.200 210.800 ;
        RECT 356.400 202.200 357.200 210.000 ;
        RECT 357.800 209.600 358.400 211.400 ;
        RECT 357.800 209.000 366.800 209.600 ;
        RECT 357.800 207.400 358.400 209.000 ;
        RECT 366.000 208.800 366.800 209.000 ;
        RECT 369.200 209.000 377.800 209.600 ;
        RECT 369.200 208.800 370.000 209.000 ;
        RECT 361.000 207.600 363.600 208.400 ;
        RECT 357.800 206.800 360.400 207.400 ;
        RECT 359.600 202.200 360.400 206.800 ;
        RECT 362.800 202.200 363.600 207.600 ;
        RECT 364.200 206.800 368.400 207.600 ;
        RECT 366.000 202.200 366.800 205.000 ;
        RECT 367.600 202.200 368.400 205.000 ;
        RECT 369.200 202.200 370.000 205.000 ;
        RECT 370.800 202.200 371.600 208.400 ;
        RECT 374.000 207.600 376.600 208.400 ;
        RECT 377.200 208.200 377.800 209.000 ;
        RECT 378.800 209.400 379.600 209.600 ;
        RECT 378.800 209.000 384.200 209.400 ;
        RECT 378.800 208.800 385.000 209.000 ;
        RECT 383.600 208.200 385.000 208.800 ;
        RECT 377.200 207.600 383.000 208.200 ;
        RECT 386.000 208.000 387.600 208.800 ;
        RECT 386.000 207.600 386.600 208.000 ;
        RECT 374.000 202.200 374.800 207.000 ;
        RECT 377.200 202.200 378.000 207.000 ;
        RECT 382.400 206.800 386.600 207.600 ;
        RECT 388.400 207.400 389.200 213.000 ;
        RECT 391.400 215.800 392.400 216.400 ;
        RECT 391.400 214.400 392.000 215.800 ;
        RECT 394.800 215.200 395.600 219.800 ;
        RECT 396.400 216.000 397.200 219.800 ;
        RECT 399.600 216.000 400.400 219.800 ;
        RECT 396.400 215.800 400.400 216.000 ;
        RECT 401.200 215.800 402.000 219.800 ;
        RECT 396.600 215.400 400.200 215.800 ;
        RECT 393.000 214.600 395.600 215.200 ;
        RECT 391.400 213.600 392.400 214.400 ;
        RECT 391.400 210.200 392.000 213.600 ;
        RECT 393.000 213.000 393.600 214.600 ;
        RECT 397.200 214.400 398.000 214.800 ;
        RECT 401.200 214.400 401.800 215.800 ;
        RECT 396.400 213.800 398.000 214.400 ;
        RECT 396.400 213.600 397.200 213.800 ;
        RECT 399.400 213.600 402.000 214.400 ;
        RECT 407.600 213.800 408.400 219.800 ;
        RECT 414.000 216.600 414.800 219.800 ;
        RECT 415.600 217.000 416.400 219.800 ;
        RECT 417.200 217.000 418.000 219.800 ;
        RECT 418.800 217.000 419.600 219.800 ;
        RECT 422.000 217.000 422.800 219.800 ;
        RECT 425.200 217.000 426.000 219.800 ;
        RECT 426.800 217.000 427.600 219.800 ;
        RECT 428.400 217.000 429.200 219.800 ;
        RECT 430.000 217.000 430.800 219.800 ;
        RECT 412.200 215.800 414.800 216.600 ;
        RECT 431.600 216.600 432.400 219.800 ;
        RECT 418.200 215.800 422.800 216.400 ;
        RECT 412.200 215.200 413.000 215.800 ;
        RECT 410.000 214.400 413.000 215.200 ;
        RECT 392.600 212.200 393.600 213.000 ;
        RECT 393.000 210.200 393.600 212.200 ;
        RECT 394.600 212.400 395.400 213.200 ;
        RECT 394.600 212.300 395.600 212.400 ;
        RECT 396.400 212.300 397.200 212.400 ;
        RECT 394.600 211.700 397.200 212.300 ;
        RECT 394.600 211.600 395.600 211.700 ;
        RECT 396.400 211.600 397.200 211.700 ;
        RECT 398.000 211.600 398.800 213.200 ;
        RECT 399.400 212.300 400.000 213.600 ;
        RECT 407.600 213.000 416.400 213.800 ;
        RECT 418.200 213.400 419.000 215.800 ;
        RECT 422.000 215.600 422.800 215.800 ;
        RECT 423.600 215.600 425.200 216.400 ;
        RECT 428.200 215.600 429.200 216.400 ;
        RECT 431.600 215.800 434.000 216.600 ;
        RECT 420.400 213.600 421.200 215.200 ;
        RECT 422.000 214.800 422.800 215.000 ;
        RECT 422.000 214.200 426.400 214.800 ;
        RECT 425.600 214.000 426.400 214.200 ;
        RECT 406.000 212.300 406.800 212.400 ;
        RECT 399.400 211.700 406.800 212.300 ;
        RECT 399.400 210.200 400.000 211.700 ;
        RECT 406.000 211.600 406.800 211.700 ;
        RECT 401.200 210.200 402.000 210.400 ;
        RECT 391.400 209.200 392.400 210.200 ;
        RECT 393.000 209.600 395.600 210.200 ;
        RECT 387.200 206.800 389.200 207.400 ;
        RECT 378.800 202.200 379.600 205.000 ;
        RECT 380.400 202.200 381.200 205.000 ;
        RECT 383.600 202.200 384.400 206.800 ;
        RECT 387.200 206.200 387.800 206.800 ;
        RECT 386.800 205.600 387.800 206.200 ;
        RECT 386.800 202.200 387.600 205.600 ;
        RECT 391.600 202.200 392.400 209.200 ;
        RECT 394.800 202.200 395.600 209.600 ;
        RECT 399.000 209.600 400.000 210.200 ;
        RECT 400.600 209.600 402.000 210.200 ;
        RECT 399.000 202.200 399.800 209.600 ;
        RECT 400.600 208.400 401.200 209.600 ;
        RECT 400.400 207.600 401.200 208.400 ;
        RECT 407.600 207.400 408.400 213.000 ;
        RECT 417.000 212.600 419.000 213.400 ;
        RECT 422.800 212.600 426.000 213.400 ;
        RECT 428.400 212.800 429.200 215.600 ;
        RECT 433.200 215.200 434.000 215.800 ;
        RECT 433.200 214.600 435.000 215.200 ;
        RECT 434.200 213.400 435.000 214.600 ;
        RECT 438.000 214.600 438.800 219.800 ;
        RECT 439.600 216.000 440.400 219.800 ;
        RECT 439.600 215.200 440.600 216.000 ;
        RECT 438.000 214.000 439.200 214.600 ;
        RECT 434.200 212.600 438.000 213.400 ;
        RECT 409.000 212.000 409.800 212.200 ;
        RECT 410.800 212.000 411.600 212.400 ;
        RECT 414.000 212.000 414.800 212.400 ;
        RECT 431.600 212.000 432.400 212.600 ;
        RECT 438.600 212.000 439.200 214.000 ;
        RECT 409.000 211.400 432.400 212.000 ;
        RECT 438.400 211.400 439.200 212.000 ;
        RECT 438.400 209.600 439.000 211.400 ;
        RECT 439.800 210.800 440.600 215.200 ;
        RECT 442.800 215.200 443.600 219.800 ;
        RECT 446.000 216.400 446.800 219.800 ;
        RECT 446.000 215.800 447.000 216.400 ;
        RECT 450.800 216.000 451.600 219.800 ;
        RECT 442.800 214.600 445.400 215.200 ;
        RECT 443.000 212.400 443.800 213.200 ;
        RECT 442.800 211.600 443.800 212.400 ;
        RECT 444.800 213.000 445.400 214.600 ;
        RECT 446.400 214.400 447.000 215.800 ;
        RECT 446.000 213.600 447.000 214.400 ;
        RECT 444.800 212.200 445.800 213.000 ;
        RECT 417.200 209.400 418.000 209.600 ;
        RECT 412.600 209.000 418.000 209.400 ;
        RECT 411.800 208.800 418.000 209.000 ;
        RECT 419.000 209.000 427.600 209.600 ;
        RECT 409.200 208.000 410.800 208.800 ;
        RECT 411.800 208.200 413.200 208.800 ;
        RECT 419.000 208.200 419.600 209.000 ;
        RECT 426.800 208.800 427.600 209.000 ;
        RECT 430.000 209.000 439.000 209.600 ;
        RECT 430.000 208.800 430.800 209.000 ;
        RECT 410.200 207.600 410.800 208.000 ;
        RECT 413.800 207.600 419.600 208.200 ;
        RECT 420.200 207.600 422.800 208.400 ;
        RECT 407.600 206.800 409.600 207.400 ;
        RECT 410.200 206.800 414.400 207.600 ;
        RECT 409.000 206.200 409.600 206.800 ;
        RECT 409.000 205.600 410.000 206.200 ;
        RECT 409.200 202.200 410.000 205.600 ;
        RECT 412.400 202.200 413.200 206.800 ;
        RECT 415.600 202.200 416.400 205.000 ;
        RECT 417.200 202.200 418.000 205.000 ;
        RECT 418.800 202.200 419.600 207.000 ;
        RECT 422.000 202.200 422.800 207.000 ;
        RECT 425.200 202.200 426.000 208.400 ;
        RECT 433.200 207.600 435.800 208.400 ;
        RECT 428.400 206.800 432.600 207.600 ;
        RECT 426.800 202.200 427.600 205.000 ;
        RECT 428.400 202.200 429.200 205.000 ;
        RECT 430.000 202.200 430.800 205.000 ;
        RECT 433.200 202.200 434.000 207.600 ;
        RECT 438.400 207.400 439.000 209.000 ;
        RECT 436.400 206.800 439.000 207.400 ;
        RECT 439.600 210.000 440.600 210.800 ;
        RECT 444.800 210.200 445.400 212.200 ;
        RECT 446.400 210.200 447.000 213.600 ;
        RECT 436.400 202.200 437.200 206.800 ;
        RECT 439.600 202.200 440.400 210.000 ;
        RECT 442.800 209.600 445.400 210.200 ;
        RECT 442.800 202.200 443.600 209.600 ;
        RECT 446.000 209.200 447.000 210.200 ;
        RECT 450.600 215.200 451.600 216.000 ;
        RECT 450.600 210.800 451.400 215.200 ;
        RECT 452.400 214.600 453.200 219.800 ;
        RECT 458.800 216.600 459.600 219.800 ;
        RECT 460.400 217.000 461.200 219.800 ;
        RECT 462.000 217.000 462.800 219.800 ;
        RECT 463.600 217.000 464.400 219.800 ;
        RECT 465.200 217.000 466.000 219.800 ;
        RECT 468.400 217.000 469.200 219.800 ;
        RECT 471.600 217.000 472.400 219.800 ;
        RECT 473.200 217.000 474.000 219.800 ;
        RECT 474.800 217.000 475.600 219.800 ;
        RECT 457.200 215.800 459.600 216.600 ;
        RECT 476.400 216.600 477.200 219.800 ;
        RECT 457.200 215.200 458.000 215.800 ;
        RECT 452.000 214.000 453.200 214.600 ;
        RECT 456.200 214.600 458.000 215.200 ;
        RECT 462.000 215.600 463.000 216.400 ;
        RECT 466.000 215.600 467.600 216.400 ;
        RECT 468.400 215.800 473.000 216.400 ;
        RECT 476.400 215.800 479.000 216.600 ;
        RECT 468.400 215.600 469.200 215.800 ;
        RECT 452.000 212.000 452.600 214.000 ;
        RECT 456.200 213.400 457.000 214.600 ;
        RECT 453.200 212.600 457.000 213.400 ;
        RECT 462.000 212.800 462.800 215.600 ;
        RECT 468.400 214.800 469.200 215.000 ;
        RECT 464.800 214.200 469.200 214.800 ;
        RECT 464.800 214.000 465.600 214.200 ;
        RECT 470.000 213.600 470.800 215.200 ;
        RECT 472.200 213.400 473.000 215.800 ;
        RECT 478.200 215.200 479.000 215.800 ;
        RECT 478.200 214.400 481.200 215.200 ;
        RECT 482.800 213.800 483.600 219.800 ;
        RECT 484.400 215.600 485.200 217.200 ;
        RECT 465.200 212.600 468.400 213.400 ;
        RECT 472.200 212.600 474.200 213.400 ;
        RECT 474.800 213.000 483.600 213.800 ;
        RECT 452.000 211.400 452.800 212.000 ;
        RECT 450.600 210.000 451.600 210.800 ;
        RECT 446.000 202.200 446.800 209.200 ;
        RECT 450.800 202.200 451.600 210.000 ;
        RECT 452.200 209.600 452.800 211.400 ;
        RECT 453.400 210.800 454.200 211.000 ;
        RECT 453.400 210.200 480.400 210.800 ;
        RECT 476.200 210.000 477.000 210.200 ;
        RECT 479.600 209.600 480.400 210.200 ;
        RECT 452.200 209.000 461.200 209.600 ;
        RECT 452.200 207.400 452.800 209.000 ;
        RECT 460.400 208.800 461.200 209.000 ;
        RECT 463.600 209.000 472.200 209.600 ;
        RECT 463.600 208.800 464.400 209.000 ;
        RECT 455.400 207.600 458.000 208.400 ;
        RECT 452.200 206.800 454.800 207.400 ;
        RECT 454.000 202.200 454.800 206.800 ;
        RECT 457.200 202.200 458.000 207.600 ;
        RECT 458.600 206.800 462.800 207.600 ;
        RECT 460.400 202.200 461.200 205.000 ;
        RECT 462.000 202.200 462.800 205.000 ;
        RECT 463.600 202.200 464.400 205.000 ;
        RECT 465.200 202.200 466.000 208.400 ;
        RECT 468.400 207.600 471.000 208.400 ;
        RECT 471.600 208.200 472.200 209.000 ;
        RECT 473.200 209.400 474.000 209.600 ;
        RECT 473.200 209.000 478.600 209.400 ;
        RECT 473.200 208.800 479.400 209.000 ;
        RECT 478.000 208.200 479.400 208.800 ;
        RECT 471.600 207.600 477.400 208.200 ;
        RECT 480.400 208.000 482.000 208.800 ;
        RECT 480.400 207.600 481.000 208.000 ;
        RECT 468.400 202.200 469.200 207.000 ;
        RECT 471.600 202.200 472.400 207.000 ;
        RECT 476.800 206.800 481.000 207.600 ;
        RECT 482.800 207.400 483.600 213.000 ;
        RECT 481.600 206.800 483.600 207.400 ;
        RECT 473.200 202.200 474.000 205.000 ;
        RECT 474.800 202.200 475.600 205.000 ;
        RECT 478.000 202.200 478.800 206.800 ;
        RECT 481.600 206.200 482.200 206.800 ;
        RECT 481.200 205.600 482.200 206.200 ;
        RECT 481.200 202.200 482.000 205.600 ;
        RECT 486.000 202.200 486.800 219.800 ;
        RECT 487.600 213.800 488.400 219.800 ;
        RECT 494.000 216.600 494.800 219.800 ;
        RECT 495.600 217.000 496.400 219.800 ;
        RECT 497.200 217.000 498.000 219.800 ;
        RECT 498.800 217.000 499.600 219.800 ;
        RECT 502.000 217.000 502.800 219.800 ;
        RECT 505.200 217.000 506.000 219.800 ;
        RECT 506.800 217.000 507.600 219.800 ;
        RECT 508.400 217.000 509.200 219.800 ;
        RECT 510.000 217.000 510.800 219.800 ;
        RECT 492.200 215.800 494.800 216.600 ;
        RECT 511.600 216.600 512.400 219.800 ;
        RECT 498.200 215.800 502.800 216.400 ;
        RECT 492.200 215.200 493.000 215.800 ;
        RECT 490.000 214.400 493.000 215.200 ;
        RECT 487.600 213.000 496.400 213.800 ;
        RECT 498.200 213.400 499.000 215.800 ;
        RECT 502.000 215.600 502.800 215.800 ;
        RECT 503.600 215.600 505.200 216.400 ;
        RECT 508.200 215.600 509.200 216.400 ;
        RECT 511.600 215.800 514.000 216.600 ;
        RECT 500.400 213.600 501.200 215.200 ;
        RECT 502.000 214.800 502.800 215.000 ;
        RECT 502.000 214.200 506.400 214.800 ;
        RECT 505.600 214.000 506.400 214.200 ;
        RECT 487.600 207.400 488.400 213.000 ;
        RECT 497.000 212.600 499.000 213.400 ;
        RECT 502.800 212.600 506.000 213.400 ;
        RECT 508.400 212.800 509.200 215.600 ;
        RECT 513.200 215.200 514.000 215.800 ;
        RECT 513.200 214.600 515.000 215.200 ;
        RECT 514.200 213.400 515.000 214.600 ;
        RECT 518.000 214.600 518.800 219.800 ;
        RECT 519.600 216.000 520.400 219.800 ;
        RECT 522.800 216.000 523.600 219.800 ;
        RECT 526.000 216.000 526.800 219.800 ;
        RECT 519.600 215.200 520.600 216.000 ;
        RECT 522.800 215.800 526.800 216.000 ;
        RECT 527.600 215.800 528.400 219.800 ;
        RECT 529.800 218.400 530.600 219.800 ;
        RECT 529.200 217.600 530.600 218.400 ;
        RECT 529.800 216.400 530.600 217.600 ;
        RECT 529.800 215.800 531.600 216.400 ;
        RECT 534.000 215.800 534.800 219.800 ;
        RECT 535.600 216.000 536.400 219.800 ;
        RECT 538.800 216.000 539.600 219.800 ;
        RECT 542.000 217.800 542.800 219.800 ;
        RECT 535.600 215.800 539.600 216.000 ;
        RECT 523.000 215.400 526.600 215.800 ;
        RECT 518.000 214.000 519.200 214.600 ;
        RECT 514.200 212.600 518.000 213.400 ;
        RECT 489.200 212.200 490.000 212.400 ;
        RECT 489.000 212.000 490.000 212.200 ;
        RECT 494.000 212.000 494.800 212.400 ;
        RECT 500.400 212.000 501.200 212.400 ;
        RECT 511.600 212.000 512.400 212.600 ;
        RECT 518.600 212.000 519.200 214.000 ;
        RECT 489.000 211.400 512.400 212.000 ;
        RECT 518.400 211.400 519.200 212.000 ;
        RECT 518.400 209.600 519.000 211.400 ;
        RECT 519.800 210.800 520.600 215.200 ;
        RECT 523.600 214.400 524.400 214.800 ;
        RECT 527.600 214.400 528.200 215.800 ;
        RECT 522.800 213.800 524.400 214.400 ;
        RECT 522.800 213.600 523.600 213.800 ;
        RECT 525.800 213.600 528.400 214.400 ;
        RECT 524.400 211.600 525.200 213.200 ;
        RECT 497.200 209.400 498.000 209.600 ;
        RECT 492.600 209.000 498.000 209.400 ;
        RECT 491.800 208.800 498.000 209.000 ;
        RECT 499.000 209.000 507.600 209.600 ;
        RECT 489.200 208.000 490.800 208.800 ;
        RECT 491.800 208.200 493.200 208.800 ;
        RECT 499.000 208.200 499.600 209.000 ;
        RECT 506.800 208.800 507.600 209.000 ;
        RECT 510.000 209.000 519.000 209.600 ;
        RECT 510.000 208.800 510.800 209.000 ;
        RECT 490.200 207.600 490.800 208.000 ;
        RECT 493.800 207.600 499.600 208.200 ;
        RECT 500.200 207.600 502.800 208.400 ;
        RECT 487.600 206.800 489.600 207.400 ;
        RECT 490.200 206.800 494.400 207.600 ;
        RECT 489.000 206.200 489.600 206.800 ;
        RECT 489.000 205.600 490.000 206.200 ;
        RECT 489.200 202.200 490.000 205.600 ;
        RECT 492.400 202.200 493.200 206.800 ;
        RECT 495.600 202.200 496.400 205.000 ;
        RECT 497.200 202.200 498.000 205.000 ;
        RECT 498.800 202.200 499.600 207.000 ;
        RECT 502.000 202.200 502.800 207.000 ;
        RECT 505.200 202.200 506.000 208.400 ;
        RECT 513.200 207.600 515.800 208.400 ;
        RECT 508.400 206.800 512.600 207.600 ;
        RECT 506.800 202.200 507.600 205.000 ;
        RECT 508.400 202.200 509.200 205.000 ;
        RECT 510.000 202.200 510.800 205.000 ;
        RECT 513.200 202.200 514.000 207.600 ;
        RECT 518.400 207.400 519.000 209.000 ;
        RECT 516.400 206.800 519.000 207.400 ;
        RECT 519.600 210.000 520.600 210.800 ;
        RECT 525.800 210.200 526.400 213.600 ;
        RECT 527.600 210.200 528.400 210.400 ;
        RECT 516.400 202.200 517.200 206.800 ;
        RECT 519.600 202.200 520.400 210.000 ;
        RECT 525.400 209.600 526.400 210.200 ;
        RECT 527.000 209.600 528.400 210.200 ;
        RECT 525.400 202.200 526.200 209.600 ;
        RECT 527.000 208.400 527.600 209.600 ;
        RECT 529.200 208.800 530.000 210.400 ;
        RECT 526.800 207.600 527.600 208.400 ;
        RECT 530.800 202.200 531.600 215.800 ;
        RECT 532.400 214.300 533.200 215.200 ;
        RECT 534.200 214.400 534.800 215.800 ;
        RECT 535.800 215.400 539.400 215.800 ;
        RECT 540.400 215.600 541.200 217.200 ;
        RECT 538.000 214.400 538.800 214.800 ;
        RECT 542.200 214.400 542.800 217.800 ;
        RECT 546.800 217.800 547.600 219.800 ;
        RECT 546.800 214.400 547.400 217.800 ;
        RECT 548.400 215.600 549.200 217.200 ;
        RECT 550.000 216.000 550.800 219.800 ;
        RECT 553.200 216.000 554.000 219.800 ;
        RECT 550.000 215.800 554.000 216.000 ;
        RECT 554.800 215.800 555.600 219.800 ;
        RECT 556.600 216.400 557.400 217.200 ;
        RECT 550.200 215.400 553.800 215.800 ;
        RECT 550.800 214.400 551.600 214.800 ;
        RECT 554.800 214.400 555.400 215.800 ;
        RECT 556.400 215.600 557.200 216.400 ;
        RECT 558.000 215.800 558.800 219.800 ;
        RECT 534.000 214.300 536.600 214.400 ;
        RECT 532.400 213.700 536.600 214.300 ;
        RECT 538.000 213.800 539.600 214.400 ;
        RECT 532.400 213.600 533.200 213.700 ;
        RECT 534.000 213.600 536.600 213.700 ;
        RECT 538.800 213.600 539.600 213.800 ;
        RECT 542.000 213.600 542.800 214.400 ;
        RECT 543.600 214.300 544.400 214.400 ;
        RECT 546.800 214.300 547.600 214.400 ;
        RECT 543.600 213.700 547.600 214.300 ;
        RECT 543.600 213.600 544.400 213.700 ;
        RECT 546.800 213.600 547.600 213.700 ;
        RECT 548.400 214.300 549.200 214.400 ;
        RECT 550.000 214.300 551.600 214.400 ;
        RECT 548.400 213.800 551.600 214.300 ;
        RECT 548.400 213.700 550.800 213.800 ;
        RECT 548.400 213.600 549.200 213.700 ;
        RECT 550.000 213.600 550.800 213.700 ;
        RECT 553.000 213.600 555.600 214.400 ;
        RECT 534.000 210.200 534.800 210.400 ;
        RECT 536.000 210.200 536.600 213.600 ;
        RECT 537.200 212.300 538.000 213.200 ;
        RECT 542.200 212.300 542.800 213.600 ;
        RECT 537.200 211.700 542.800 212.300 ;
        RECT 537.200 211.600 538.000 211.700 ;
        RECT 542.200 210.200 542.800 211.700 ;
        RECT 543.600 212.300 544.400 212.400 ;
        RECT 545.200 212.300 546.000 212.400 ;
        RECT 543.600 211.700 546.000 212.300 ;
        RECT 543.600 210.800 544.400 211.700 ;
        RECT 545.200 210.800 546.000 211.700 ;
        RECT 546.800 210.200 547.400 213.600 ;
        RECT 551.600 211.600 552.400 213.200 ;
        RECT 553.000 210.200 553.600 213.600 ;
        RECT 554.800 212.300 555.600 212.400 ;
        RECT 556.400 212.300 557.200 212.400 ;
        RECT 554.800 212.200 557.200 212.300 ;
        RECT 558.200 212.200 558.800 215.800 ;
        RECT 559.600 214.300 560.400 214.400 ;
        RECT 564.000 214.300 564.800 219.800 ;
        RECT 559.600 213.800 564.800 214.300 ;
        RECT 574.000 215.800 574.800 219.800 ;
        RECT 577.200 217.800 578.000 219.800 ;
        RECT 559.600 213.700 564.600 213.800 ;
        RECT 559.600 212.800 560.400 213.700 ;
        RECT 563.000 213.600 564.600 213.700 ;
        RECT 561.200 212.200 562.000 212.400 ;
        RECT 554.800 211.700 558.800 212.200 ;
        RECT 554.800 211.600 555.600 211.700 ;
        RECT 556.400 211.600 558.800 211.700 ;
        RECT 560.400 211.600 562.000 212.200 ;
        RECT 554.800 210.200 555.600 210.400 ;
        RECT 556.600 210.200 557.200 211.600 ;
        RECT 560.400 211.200 561.200 211.600 ;
        RECT 563.000 210.400 563.600 213.600 ;
        RECT 574.000 212.400 574.600 215.800 ;
        RECT 577.200 215.600 577.800 217.800 ;
        RECT 578.800 215.600 579.600 217.200 ;
        RECT 580.400 215.800 581.200 219.800 ;
        RECT 584.800 218.400 586.400 219.800 ;
        RECT 584.800 217.600 587.600 218.400 ;
        RECT 584.800 216.200 586.400 217.600 ;
        RECT 575.400 215.000 577.800 215.600 ;
        RECT 580.400 215.200 583.000 215.800 ;
        RECT 582.200 215.000 583.000 215.200 ;
        RECT 565.200 211.600 566.800 212.400 ;
        RECT 569.200 212.300 570.000 212.400 ;
        RECT 574.000 212.300 574.800 212.400 ;
        RECT 569.200 211.700 574.800 212.300 ;
        RECT 569.200 211.600 570.000 211.700 ;
        RECT 574.000 211.600 574.800 211.700 ;
        RECT 575.400 212.000 576.000 215.000 ;
        RECT 583.600 214.800 585.200 215.600 ;
        RECT 577.000 213.600 578.000 214.400 ;
        RECT 580.400 214.200 582.000 214.400 ;
        RECT 585.800 214.200 586.400 216.200 ;
        RECT 590.000 215.800 590.800 219.800 ;
        RECT 587.000 214.800 587.800 215.600 ;
        RECT 588.400 215.200 590.800 215.800 ;
        RECT 591.600 217.000 592.400 219.000 ;
        RECT 588.400 215.000 589.200 215.200 ;
        RECT 580.400 214.000 582.600 214.200 ;
        RECT 580.400 213.600 584.800 214.000 ;
        RECT 576.800 212.800 577.600 213.600 ;
        RECT 582.000 213.400 584.800 213.600 ;
        RECT 584.000 213.200 584.800 213.400 ;
        RECT 585.400 213.600 586.400 214.200 ;
        RECT 587.200 214.400 587.800 214.800 ;
        RECT 591.600 214.800 592.200 217.000 ;
        RECT 595.800 216.000 596.600 219.000 ;
        RECT 601.200 217.000 602.000 219.000 ;
        RECT 595.800 215.400 597.400 216.000 ;
        RECT 596.600 215.000 597.400 215.400 ;
        RECT 587.200 213.600 588.000 214.400 ;
        RECT 589.200 213.600 590.800 214.400 ;
        RECT 591.600 214.200 595.800 214.800 ;
        RECT 594.800 213.800 595.800 214.200 ;
        RECT 596.800 214.400 597.400 215.000 ;
        RECT 601.200 214.800 601.800 217.000 ;
        RECT 605.400 216.000 606.200 219.000 ;
        RECT 612.400 216.000 613.200 219.800 ;
        RECT 605.400 215.400 607.000 216.000 ;
        RECT 606.200 215.000 607.000 215.400 ;
        RECT 596.800 214.300 598.800 214.400 ;
        RECT 599.600 214.300 600.400 214.400 ;
        RECT 585.400 212.400 586.000 213.600 ;
        RECT 582.600 212.200 583.400 212.400 ;
        RECT 534.000 209.600 535.400 210.200 ;
        RECT 536.000 209.600 537.000 210.200 ;
        RECT 534.800 208.400 535.400 209.600 ;
        RECT 534.800 207.600 535.600 208.400 ;
        RECT 536.200 202.200 537.000 209.600 ;
        RECT 542.000 209.400 543.800 210.200 ;
        RECT 543.000 202.200 543.800 209.400 ;
        RECT 545.800 209.400 547.600 210.200 ;
        RECT 552.600 209.600 553.600 210.200 ;
        RECT 554.200 209.600 555.600 210.200 ;
        RECT 545.800 202.200 546.600 209.400 ;
        RECT 552.600 208.400 553.400 209.600 ;
        RECT 554.200 208.400 554.800 209.600 ;
        RECT 551.600 207.600 553.400 208.400 ;
        RECT 554.000 207.600 554.800 208.400 ;
        RECT 552.600 202.200 553.400 207.600 ;
        RECT 556.400 202.200 557.200 210.200 ;
        RECT 558.000 209.600 562.000 210.200 ;
        RECT 562.800 209.600 563.600 210.400 ;
        RECT 567.600 209.600 568.400 211.200 ;
        RECT 574.000 210.200 574.600 211.600 ;
        RECT 575.400 211.400 576.200 212.000 ;
        RECT 582.600 211.600 584.200 212.200 ;
        RECT 585.200 211.600 586.000 212.400 ;
        RECT 590.000 212.300 590.800 212.400 ;
        RECT 591.600 212.300 592.400 213.200 ;
        RECT 590.000 211.700 592.400 212.300 ;
        RECT 590.000 211.600 590.800 211.700 ;
        RECT 591.600 211.600 592.400 211.700 ;
        RECT 593.200 211.600 594.000 213.200 ;
        RECT 594.800 213.000 596.200 213.800 ;
        RECT 596.800 213.700 600.400 214.300 ;
        RECT 601.200 214.200 605.400 214.800 ;
        RECT 596.800 213.600 598.800 213.700 ;
        RECT 599.600 213.600 600.400 213.700 ;
        RECT 604.400 213.800 605.400 214.200 ;
        RECT 606.400 214.400 607.000 215.000 ;
        RECT 612.200 215.200 613.200 216.000 ;
        RECT 606.400 214.300 608.400 214.400 ;
        RECT 610.800 214.300 611.600 214.400 ;
        RECT 583.400 211.400 584.200 211.600 ;
        RECT 575.400 211.200 579.600 211.400 ;
        RECT 575.600 210.800 579.600 211.200 ;
        RECT 574.000 209.600 575.400 210.200 ;
        RECT 558.000 202.200 558.800 209.600 ;
        RECT 561.200 202.200 562.000 209.600 ;
        RECT 563.000 207.000 563.600 209.600 ;
        RECT 564.400 207.600 565.200 209.200 ;
        RECT 563.000 206.400 566.600 207.000 ;
        RECT 563.000 206.200 563.600 206.400 ;
        RECT 562.800 202.200 563.600 206.200 ;
        RECT 566.000 206.200 566.600 206.400 ;
        RECT 566.000 202.200 566.800 206.200 ;
        RECT 574.600 202.200 575.400 209.600 ;
        RECT 578.800 202.200 579.600 210.800 ;
        RECT 585.400 210.200 586.000 211.600 ;
        RECT 594.800 211.000 595.400 213.000 ;
        RECT 591.600 210.400 595.400 211.000 ;
        RECT 580.400 209.600 583.000 210.200 ;
        RECT 580.400 202.200 581.200 209.600 ;
        RECT 582.200 209.400 583.000 209.600 ;
        RECT 584.800 202.200 586.400 210.200 ;
        RECT 588.400 209.600 590.800 210.200 ;
        RECT 588.400 209.400 589.200 209.600 ;
        RECT 590.000 202.200 590.800 209.600 ;
        RECT 591.600 207.000 592.200 210.400 ;
        RECT 596.800 209.800 597.400 213.600 ;
        RECT 598.000 210.800 598.800 212.400 ;
        RECT 601.200 211.600 602.000 213.200 ;
        RECT 602.800 211.600 603.600 213.200 ;
        RECT 604.400 213.000 605.800 213.800 ;
        RECT 606.400 213.700 611.600 214.300 ;
        RECT 606.400 213.600 608.400 213.700 ;
        RECT 610.800 213.600 611.600 213.700 ;
        RECT 604.400 211.000 605.000 213.000 ;
        RECT 595.800 209.200 597.400 209.800 ;
        RECT 601.200 210.400 605.000 211.000 ;
        RECT 591.600 203.000 592.400 207.000 ;
        RECT 595.800 202.200 596.600 209.200 ;
        RECT 601.200 207.000 601.800 210.400 ;
        RECT 606.400 209.800 607.000 213.600 ;
        RECT 607.600 210.800 608.400 212.400 ;
        RECT 612.200 210.800 613.000 215.200 ;
        RECT 614.000 214.600 614.800 219.800 ;
        RECT 620.400 216.600 621.200 219.800 ;
        RECT 622.000 217.000 622.800 219.800 ;
        RECT 623.600 217.000 624.400 219.800 ;
        RECT 625.200 217.000 626.000 219.800 ;
        RECT 626.800 217.000 627.600 219.800 ;
        RECT 630.000 217.000 630.800 219.800 ;
        RECT 633.200 217.000 634.000 219.800 ;
        RECT 634.800 217.000 635.600 219.800 ;
        RECT 636.400 217.000 637.200 219.800 ;
        RECT 618.800 215.800 621.200 216.600 ;
        RECT 638.000 216.600 638.800 219.800 ;
        RECT 618.800 215.200 619.600 215.800 ;
        RECT 613.600 214.000 614.800 214.600 ;
        RECT 617.800 214.600 619.600 215.200 ;
        RECT 623.600 215.600 624.600 216.400 ;
        RECT 627.600 215.600 629.200 216.400 ;
        RECT 630.000 215.800 634.600 216.400 ;
        RECT 638.000 215.800 640.600 216.600 ;
        RECT 630.000 215.600 630.800 215.800 ;
        RECT 613.600 212.000 614.200 214.000 ;
        RECT 617.800 213.400 618.600 214.600 ;
        RECT 614.800 212.600 618.600 213.400 ;
        RECT 623.600 212.800 624.400 215.600 ;
        RECT 630.000 214.800 630.800 215.000 ;
        RECT 626.400 214.200 630.800 214.800 ;
        RECT 626.400 214.000 627.200 214.200 ;
        RECT 631.600 213.600 632.400 215.200 ;
        RECT 633.800 213.400 634.600 215.800 ;
        RECT 639.800 215.200 640.600 215.800 ;
        RECT 639.800 214.400 642.800 215.200 ;
        RECT 644.400 213.800 645.200 219.800 ;
        RECT 646.000 215.800 646.800 219.800 ;
        RECT 650.400 218.400 652.000 219.800 ;
        RECT 649.200 217.600 652.000 218.400 ;
        RECT 650.400 216.200 652.000 217.600 ;
        RECT 646.000 215.200 648.200 215.800 ;
        RECT 649.200 215.400 650.800 215.600 ;
        RECT 647.400 215.000 648.200 215.200 ;
        RECT 648.800 214.800 650.800 215.400 ;
        RECT 648.800 214.400 649.400 214.800 ;
        RECT 626.800 212.600 630.000 213.400 ;
        RECT 633.800 212.600 635.800 213.400 ;
        RECT 636.400 213.000 645.200 213.800 ;
        RECT 646.000 213.800 649.400 214.400 ;
        RECT 646.000 213.600 647.600 213.800 ;
        RECT 620.400 212.000 621.200 212.600 ;
        RECT 638.000 212.000 638.800 212.400 ;
        RECT 642.800 212.200 643.600 212.400 ;
        RECT 642.800 212.000 643.800 212.200 ;
        RECT 613.600 211.400 614.400 212.000 ;
        RECT 620.400 211.400 643.800 212.000 ;
        RECT 612.200 210.000 613.200 210.800 ;
        RECT 605.400 209.200 607.000 209.800 ;
        RECT 601.200 203.000 602.000 207.000 ;
        RECT 605.400 202.200 606.200 209.200 ;
        RECT 612.400 202.200 613.200 210.000 ;
        RECT 613.800 209.600 614.400 211.400 ;
        RECT 613.800 209.000 622.800 209.600 ;
        RECT 613.800 207.400 614.400 209.000 ;
        RECT 622.000 208.800 622.800 209.000 ;
        RECT 625.200 209.000 633.800 209.600 ;
        RECT 625.200 208.800 626.000 209.000 ;
        RECT 617.000 207.600 619.600 208.400 ;
        RECT 613.800 206.800 616.400 207.400 ;
        RECT 615.600 202.200 616.400 206.800 ;
        RECT 618.800 202.200 619.600 207.600 ;
        RECT 620.200 206.800 624.400 207.600 ;
        RECT 622.000 202.200 622.800 205.000 ;
        RECT 623.600 202.200 624.400 205.000 ;
        RECT 625.200 202.200 626.000 205.000 ;
        RECT 626.800 202.200 627.600 208.400 ;
        RECT 630.000 207.600 632.600 208.400 ;
        RECT 633.200 208.200 633.800 209.000 ;
        RECT 634.800 209.400 635.600 209.600 ;
        RECT 634.800 209.000 640.200 209.400 ;
        RECT 634.800 208.800 641.000 209.000 ;
        RECT 639.600 208.200 641.000 208.800 ;
        RECT 633.200 207.600 639.000 208.200 ;
        RECT 642.000 208.000 643.600 208.800 ;
        RECT 642.000 207.600 642.600 208.000 ;
        RECT 630.000 202.200 630.800 207.000 ;
        RECT 633.200 202.200 634.000 207.000 ;
        RECT 638.400 206.800 642.600 207.600 ;
        RECT 644.400 207.400 645.200 213.000 ;
        RECT 650.000 213.400 650.800 214.200 ;
        RECT 650.000 212.800 650.600 213.400 ;
        RECT 648.000 212.200 650.600 212.800 ;
        RECT 651.400 212.800 652.000 216.200 ;
        RECT 655.600 215.800 656.400 219.800 ;
        RECT 652.600 214.800 653.400 215.600 ;
        RECT 654.000 215.200 656.400 215.800 ;
        RECT 658.800 215.200 659.600 219.800 ;
        RECT 662.000 215.200 662.800 219.800 ;
        RECT 665.200 215.200 666.000 219.800 ;
        RECT 668.400 215.200 669.200 219.800 ;
        RECT 673.200 215.200 674.000 219.800 ;
        RECT 676.400 215.200 677.200 219.800 ;
        RECT 679.600 215.200 680.400 219.800 ;
        RECT 682.800 215.200 683.600 219.800 ;
        RECT 654.000 215.000 654.800 215.200 ;
        RECT 652.800 214.400 653.400 214.800 ;
        RECT 658.800 214.400 660.600 215.200 ;
        RECT 662.000 214.400 664.200 215.200 ;
        RECT 665.200 214.400 667.400 215.200 ;
        RECT 668.400 214.400 670.800 215.200 ;
        RECT 673.200 214.400 675.000 215.200 ;
        RECT 676.400 214.400 678.600 215.200 ;
        RECT 679.600 214.400 681.800 215.200 ;
        RECT 682.800 214.400 685.200 215.200 ;
        RECT 652.800 213.600 653.600 214.400 ;
        RECT 654.800 213.600 656.400 214.400 ;
        RECT 657.200 213.800 658.000 214.400 ;
        RECT 659.800 213.800 660.600 214.400 ;
        RECT 663.400 213.800 664.200 214.400 ;
        RECT 666.600 213.800 667.400 214.400 ;
        RECT 657.200 213.000 659.000 213.800 ;
        RECT 659.800 213.000 662.400 213.800 ;
        RECT 663.400 213.000 665.800 213.800 ;
        RECT 666.600 213.000 669.200 213.800 ;
        RECT 651.400 212.400 652.400 212.800 ;
        RECT 651.400 212.200 653.200 212.400 ;
        RECT 648.000 212.000 648.800 212.200 ;
        RECT 651.800 211.600 653.200 212.200 ;
        RECT 655.600 212.300 656.400 212.400 ;
        RECT 657.300 212.300 657.900 213.000 ;
        RECT 655.600 211.700 657.900 212.300 ;
        RECT 655.600 211.600 656.400 211.700 ;
        RECT 659.800 211.600 660.600 213.000 ;
        RECT 663.400 211.600 664.200 213.000 ;
        RECT 666.600 211.600 667.400 213.000 ;
        RECT 670.000 211.600 670.800 214.400 ;
        RECT 671.600 213.800 672.400 214.400 ;
        RECT 674.200 213.800 675.000 214.400 ;
        RECT 677.800 213.800 678.600 214.400 ;
        RECT 681.000 213.800 681.800 214.400 ;
        RECT 671.600 213.000 673.400 213.800 ;
        RECT 674.200 213.000 676.800 213.800 ;
        RECT 677.800 213.000 680.200 213.800 ;
        RECT 681.000 213.000 683.600 213.800 ;
        RECT 674.200 211.600 675.000 213.000 ;
        RECT 677.800 211.600 678.600 213.000 ;
        RECT 681.000 211.600 681.800 213.000 ;
        RECT 684.400 211.600 685.200 214.400 ;
        RECT 650.200 211.400 651.000 211.600 ;
        RECT 647.600 210.800 651.000 211.400 ;
        RECT 647.600 210.200 648.200 210.800 ;
        RECT 651.800 210.200 652.400 211.600 ;
        RECT 658.800 210.800 660.600 211.600 ;
        RECT 662.000 210.800 664.200 211.600 ;
        RECT 665.200 210.800 667.400 211.600 ;
        RECT 668.400 210.800 670.800 211.600 ;
        RECT 673.200 210.800 675.000 211.600 ;
        RECT 676.400 210.800 678.600 211.600 ;
        RECT 679.600 210.800 681.800 211.600 ;
        RECT 682.800 210.800 685.200 211.600 ;
        RECT 643.200 206.800 645.200 207.400 ;
        RECT 646.000 209.600 648.200 210.200 ;
        RECT 634.800 202.200 635.600 205.000 ;
        RECT 636.400 202.200 637.200 205.000 ;
        RECT 639.600 202.200 640.400 206.800 ;
        RECT 643.200 206.200 643.800 206.800 ;
        RECT 642.800 205.600 643.800 206.200 ;
        RECT 642.800 202.200 643.600 205.600 ;
        RECT 646.000 202.200 646.800 209.600 ;
        RECT 647.400 209.400 648.200 209.600 ;
        RECT 650.400 209.600 652.400 210.200 ;
        RECT 654.000 209.600 656.400 210.200 ;
        RECT 650.400 202.200 652.000 209.600 ;
        RECT 654.000 209.400 654.800 209.600 ;
        RECT 655.600 202.200 656.400 209.600 ;
        RECT 658.800 202.200 659.600 210.800 ;
        RECT 662.000 202.200 662.800 210.800 ;
        RECT 665.200 202.200 666.000 210.800 ;
        RECT 668.400 202.200 669.200 210.800 ;
        RECT 673.200 202.200 674.000 210.800 ;
        RECT 676.400 202.200 677.200 210.800 ;
        RECT 679.600 202.200 680.400 210.800 ;
        RECT 682.800 202.200 683.600 210.800 ;
        RECT 2.800 188.300 3.600 199.800 ;
        RECT 7.000 192.400 7.800 199.800 ;
        RECT 13.000 198.400 13.800 199.800 ;
        RECT 13.000 197.600 14.800 198.400 ;
        RECT 8.400 193.600 9.200 194.400 ;
        RECT 8.600 192.400 9.200 193.600 ;
        RECT 11.600 193.600 12.400 194.400 ;
        RECT 11.600 192.400 12.200 193.600 ;
        RECT 13.000 192.400 13.800 197.600 ;
        RECT 18.800 196.400 19.600 199.800 ;
        RECT 18.600 195.800 19.600 196.400 ;
        RECT 18.600 195.200 19.200 195.800 ;
        RECT 22.000 195.200 22.800 199.800 ;
        RECT 25.200 197.000 26.000 199.800 ;
        RECT 26.800 197.000 27.600 199.800 ;
        RECT 7.000 191.800 8.000 192.400 ;
        RECT 8.600 191.800 10.000 192.400 ;
        RECT 6.000 188.800 6.800 190.400 ;
        RECT 7.400 188.400 8.000 191.800 ;
        RECT 9.200 191.600 10.000 191.800 ;
        RECT 10.800 191.800 12.200 192.400 ;
        RECT 12.800 191.800 13.800 192.400 ;
        RECT 17.200 194.600 19.200 195.200 ;
        RECT 10.800 191.600 11.600 191.800 ;
        RECT 12.800 188.400 13.400 191.800 ;
        RECT 14.000 188.800 14.800 190.400 ;
        RECT 17.200 189.000 18.000 194.600 ;
        RECT 19.800 194.400 24.000 195.200 ;
        RECT 28.400 195.000 29.200 199.800 ;
        RECT 31.600 195.000 32.400 199.800 ;
        RECT 19.800 194.000 20.400 194.400 ;
        RECT 18.800 193.200 20.400 194.000 ;
        RECT 23.400 193.800 29.200 194.400 ;
        RECT 21.400 193.200 22.800 193.800 ;
        RECT 21.400 193.000 27.600 193.200 ;
        RECT 22.200 192.600 27.600 193.000 ;
        RECT 26.800 192.400 27.600 192.600 ;
        RECT 28.600 193.000 29.200 193.800 ;
        RECT 29.800 193.600 32.400 194.400 ;
        RECT 34.800 193.600 35.600 199.800 ;
        RECT 36.400 197.000 37.200 199.800 ;
        RECT 38.000 197.000 38.800 199.800 ;
        RECT 39.600 197.000 40.400 199.800 ;
        RECT 38.000 194.400 42.200 195.200 ;
        RECT 42.800 194.400 43.600 199.800 ;
        RECT 46.000 195.200 46.800 199.800 ;
        RECT 46.000 194.600 48.600 195.200 ;
        RECT 42.800 193.600 45.400 194.400 ;
        RECT 36.400 193.000 37.200 193.200 ;
        RECT 28.600 192.400 37.200 193.000 ;
        RECT 39.600 193.000 40.400 193.200 ;
        RECT 48.000 193.000 48.600 194.600 ;
        RECT 39.600 192.400 48.600 193.000 ;
        RECT 48.000 190.600 48.600 192.400 ;
        RECT 49.200 192.300 50.000 199.800 ;
        RECT 53.200 193.600 54.000 194.400 ;
        RECT 53.200 192.400 53.800 193.600 ;
        RECT 54.600 192.400 55.400 199.800 ;
        RECT 52.400 192.300 53.800 192.400 ;
        RECT 49.200 191.800 53.800 192.300 ;
        RECT 54.400 191.800 55.400 192.400 ;
        RECT 49.200 191.700 53.200 191.800 ;
        RECT 49.200 191.200 50.200 191.700 ;
        RECT 52.400 191.600 53.200 191.700 ;
        RECT 18.600 190.000 42.000 190.600 ;
        RECT 48.000 190.000 48.800 190.600 ;
        RECT 18.600 189.800 19.400 190.000 ;
        RECT 23.600 189.600 24.400 190.000 ;
        RECT 41.200 189.400 42.000 190.000 ;
        RECT 4.400 188.300 5.200 188.400 ;
        RECT 2.800 188.200 5.200 188.300 ;
        RECT 2.800 187.700 6.000 188.200 ;
        RECT 2.800 182.200 3.600 187.700 ;
        RECT 4.400 187.600 6.000 187.700 ;
        RECT 7.400 187.600 10.000 188.400 ;
        RECT 10.800 187.600 13.400 188.400 ;
        RECT 15.600 188.200 16.400 188.400 ;
        RECT 14.800 187.600 16.400 188.200 ;
        RECT 17.200 188.200 26.000 189.000 ;
        RECT 26.600 188.600 28.600 189.400 ;
        RECT 32.400 188.600 35.600 189.400 ;
        RECT 5.200 187.200 6.000 187.600 ;
        RECT 4.600 186.200 8.200 186.600 ;
        RECT 9.200 186.400 9.800 187.600 ;
        RECT 4.400 186.000 8.400 186.200 ;
        RECT 4.400 182.200 5.200 186.000 ;
        RECT 7.600 182.200 8.400 186.000 ;
        RECT 9.200 182.200 10.000 186.400 ;
        RECT 11.000 186.200 11.600 187.600 ;
        RECT 14.800 187.200 15.600 187.600 ;
        RECT 12.600 186.200 16.200 186.600 ;
        RECT 10.800 182.200 11.600 186.200 ;
        RECT 12.400 186.000 16.400 186.200 ;
        RECT 12.400 182.200 13.200 186.000 ;
        RECT 15.600 182.200 16.400 186.000 ;
        RECT 17.200 182.200 18.000 188.200 ;
        RECT 19.600 186.800 22.600 187.600 ;
        RECT 21.800 186.200 22.600 186.800 ;
        RECT 27.800 186.200 28.600 188.600 ;
        RECT 30.000 186.800 30.800 188.400 ;
        RECT 35.200 187.800 36.000 188.000 ;
        RECT 31.600 187.200 36.000 187.800 ;
        RECT 31.600 187.000 32.400 187.200 ;
        RECT 38.000 186.400 38.800 189.200 ;
        RECT 43.800 188.600 47.600 189.400 ;
        RECT 43.800 187.400 44.600 188.600 ;
        RECT 48.200 188.000 48.800 190.000 ;
        RECT 31.600 186.200 32.400 186.400 ;
        RECT 21.800 185.400 24.400 186.200 ;
        RECT 27.800 185.600 32.400 186.200 ;
        RECT 33.200 185.600 34.800 186.400 ;
        RECT 37.800 185.600 38.800 186.400 ;
        RECT 42.800 186.800 44.600 187.400 ;
        RECT 47.600 187.400 48.800 188.000 ;
        RECT 42.800 186.200 43.600 186.800 ;
        RECT 23.600 182.200 24.400 185.400 ;
        RECT 41.200 185.400 43.600 186.200 ;
        RECT 25.200 182.200 26.000 185.000 ;
        RECT 26.800 182.200 27.600 185.000 ;
        RECT 28.400 182.200 29.200 185.000 ;
        RECT 31.600 182.200 32.400 185.000 ;
        RECT 34.800 182.200 35.600 185.000 ;
        RECT 36.400 182.200 37.200 185.000 ;
        RECT 38.000 182.200 38.800 185.000 ;
        RECT 39.600 182.200 40.400 185.000 ;
        RECT 41.200 182.200 42.000 185.400 ;
        RECT 47.600 182.200 48.400 187.400 ;
        RECT 49.400 186.800 50.200 191.200 ;
        RECT 50.800 190.300 51.600 190.400 ;
        RECT 54.400 190.300 55.000 191.800 ;
        RECT 58.800 191.200 59.600 199.800 ;
        RECT 63.000 192.400 63.800 199.800 ;
        RECT 63.000 191.800 64.400 192.400 ;
        RECT 58.800 190.800 62.800 191.200 ;
        RECT 58.800 190.600 63.000 190.800 ;
        RECT 50.800 189.700 55.000 190.300 ;
        RECT 50.800 189.600 51.600 189.700 ;
        RECT 54.400 188.400 55.000 189.700 ;
        RECT 55.600 188.800 56.400 190.400 ;
        RECT 62.200 190.000 63.000 190.600 ;
        RECT 63.800 190.400 64.400 191.800 ;
        RECT 60.800 188.400 61.600 189.200 ;
        RECT 52.400 187.600 55.000 188.400 ;
        RECT 57.200 188.300 58.000 188.400 ;
        RECT 57.200 188.200 59.500 188.300 ;
        RECT 56.400 187.700 59.500 188.200 ;
        RECT 56.400 187.600 58.000 187.700 ;
        RECT 49.200 186.000 50.200 186.800 ;
        RECT 52.600 186.200 53.200 187.600 ;
        RECT 56.400 187.200 57.200 187.600 ;
        RECT 54.200 186.200 57.800 186.600 ;
        RECT 58.900 186.400 59.500 187.700 ;
        RECT 60.400 187.600 61.400 188.400 ;
        RECT 62.400 187.000 63.000 190.000 ;
        RECT 63.600 189.600 64.400 190.400 ;
        RECT 60.600 186.400 63.000 187.000 ;
        RECT 49.200 182.200 50.000 186.000 ;
        RECT 52.400 182.200 53.200 186.200 ;
        RECT 54.000 186.000 58.000 186.200 ;
        RECT 54.000 182.200 54.800 186.000 ;
        RECT 57.200 182.200 58.000 186.000 ;
        RECT 58.800 184.800 59.600 186.400 ;
        RECT 60.600 184.200 61.200 186.400 ;
        RECT 63.800 186.200 64.400 189.600 ;
        RECT 66.800 190.300 67.600 199.800 ;
        RECT 68.400 191.600 69.200 194.400 ;
        RECT 70.000 190.300 70.800 190.400 ;
        RECT 66.800 189.700 70.800 190.300 ;
        RECT 65.200 186.800 66.000 188.400 ;
        RECT 60.400 182.200 61.200 184.200 ;
        RECT 63.600 182.200 64.400 186.200 ;
        RECT 66.800 186.200 67.600 189.700 ;
        RECT 70.000 189.600 70.800 189.700 ;
        RECT 66.800 185.600 68.600 186.200 ;
        RECT 67.800 182.200 68.600 185.600 ;
        RECT 70.000 184.800 70.800 186.400 ;
        RECT 71.600 182.200 72.400 199.800 ;
        RECT 74.000 193.600 74.800 194.400 ;
        RECT 74.000 192.400 74.600 193.600 ;
        RECT 75.400 192.400 76.200 199.800 ;
        RECT 80.400 193.600 81.200 194.400 ;
        RECT 80.400 192.400 81.000 193.600 ;
        RECT 81.800 192.400 82.600 199.800 ;
        RECT 73.200 191.800 74.600 192.400 ;
        RECT 75.200 191.800 76.200 192.400 ;
        RECT 79.600 191.800 81.000 192.400 ;
        RECT 81.600 191.800 82.600 192.400 ;
        RECT 73.200 191.600 74.000 191.800 ;
        RECT 75.200 188.400 75.800 191.800 ;
        RECT 79.600 191.600 80.400 191.800 ;
        RECT 76.400 188.800 77.200 190.400 ;
        RECT 81.600 188.400 82.200 191.800 ;
        RECT 86.000 191.400 86.800 199.800 ;
        RECT 90.400 196.400 91.200 199.800 ;
        RECT 89.200 195.800 91.200 196.400 ;
        RECT 94.800 195.800 95.600 199.800 ;
        RECT 99.000 195.800 100.200 199.800 ;
        RECT 89.200 195.000 90.000 195.800 ;
        RECT 94.800 195.200 95.400 195.800 ;
        RECT 92.600 194.600 96.200 195.200 ;
        RECT 98.800 195.000 99.600 195.800 ;
        RECT 92.600 194.400 93.400 194.600 ;
        RECT 95.400 194.400 96.200 194.600 ;
        RECT 89.200 193.000 90.000 193.200 ;
        RECT 93.800 193.000 94.600 193.200 ;
        RECT 89.200 192.400 94.600 193.000 ;
        RECT 95.200 193.000 97.400 193.600 ;
        RECT 95.200 191.800 95.800 193.000 ;
        RECT 96.600 192.800 97.400 193.000 ;
        RECT 99.000 193.200 100.400 194.000 ;
        RECT 99.000 192.200 99.600 193.200 ;
        RECT 91.000 191.400 95.800 191.800 ;
        RECT 86.000 191.200 95.800 191.400 ;
        RECT 97.200 191.600 99.600 192.200 ;
        RECT 86.000 191.000 91.800 191.200 ;
        RECT 86.000 190.800 91.600 191.000 ;
        RECT 82.800 188.800 83.600 190.400 ;
        RECT 92.400 190.200 93.200 190.400 ;
        RECT 88.200 189.600 93.200 190.200 ;
        RECT 88.200 189.400 89.000 189.600 ;
        RECT 90.800 189.400 91.600 189.600 ;
        RECT 89.800 188.400 90.600 188.600 ;
        RECT 97.200 188.400 97.800 191.600 ;
        RECT 103.600 191.200 104.400 199.800 ;
        RECT 105.200 191.600 106.000 194.400 ;
        RECT 106.800 192.300 107.600 199.800 ;
        RECT 115.600 193.600 116.400 194.400 ;
        RECT 115.600 192.400 116.200 193.600 ;
        RECT 117.000 192.400 117.800 199.800 ;
        RECT 114.800 192.300 116.200 192.400 ;
        RECT 106.800 191.800 116.200 192.300 ;
        RECT 116.800 191.800 117.800 192.400 ;
        RECT 106.800 191.700 115.600 191.800 ;
        RECT 100.200 190.600 104.400 191.200 ;
        RECT 100.200 190.400 101.000 190.600 ;
        RECT 101.800 189.800 102.600 190.000 ;
        RECT 98.800 189.200 102.600 189.800 ;
        RECT 98.800 189.000 99.600 189.200 ;
        RECT 73.200 187.600 75.800 188.400 ;
        RECT 78.000 188.200 78.800 188.400 ;
        RECT 77.200 187.600 78.800 188.200 ;
        RECT 79.600 187.600 82.200 188.400 ;
        RECT 84.400 188.200 85.200 188.400 ;
        RECT 83.600 187.600 85.200 188.200 ;
        RECT 86.800 187.800 97.800 188.400 ;
        RECT 86.800 187.600 88.400 187.800 ;
        RECT 73.400 186.200 74.000 187.600 ;
        RECT 77.200 187.200 78.000 187.600 ;
        RECT 75.000 186.200 78.600 186.600 ;
        RECT 79.800 186.200 80.400 187.600 ;
        RECT 83.600 187.200 84.400 187.600 ;
        RECT 81.400 186.200 85.000 186.600 ;
        RECT 73.200 182.200 74.000 186.200 ;
        RECT 74.800 186.000 78.800 186.200 ;
        RECT 74.800 182.200 75.600 186.000 ;
        RECT 78.000 182.200 78.800 186.000 ;
        RECT 79.600 182.200 80.400 186.200 ;
        RECT 81.200 186.000 85.200 186.200 ;
        RECT 81.200 182.200 82.000 186.000 ;
        RECT 84.400 182.200 85.200 186.000 ;
        RECT 86.000 182.200 86.800 187.000 ;
        RECT 91.000 185.600 91.600 187.800 ;
        RECT 92.400 187.600 93.200 187.800 ;
        RECT 96.600 187.600 97.400 187.800 ;
        RECT 103.600 187.200 104.400 190.600 ;
        RECT 100.600 186.600 104.400 187.200 ;
        RECT 100.600 186.400 101.400 186.600 ;
        RECT 89.200 184.200 90.000 185.000 ;
        RECT 90.800 184.800 91.600 185.600 ;
        RECT 92.600 185.400 93.400 185.600 ;
        RECT 92.600 184.800 95.400 185.400 ;
        RECT 94.800 184.200 95.400 184.800 ;
        RECT 98.800 184.200 99.600 185.000 ;
        RECT 89.200 183.600 91.200 184.200 ;
        RECT 90.400 182.200 91.200 183.600 ;
        RECT 94.800 182.200 95.600 184.200 ;
        RECT 98.800 183.600 100.200 184.200 ;
        RECT 99.000 182.200 100.200 183.600 ;
        RECT 103.600 182.200 104.400 186.600 ;
        RECT 106.800 186.200 107.600 191.700 ;
        RECT 114.800 191.600 115.600 191.700 ;
        RECT 116.800 188.400 117.400 191.800 ;
        RECT 121.200 191.400 122.000 199.800 ;
        RECT 125.600 196.400 126.400 199.800 ;
        RECT 124.400 195.800 126.400 196.400 ;
        RECT 130.000 195.800 130.800 199.800 ;
        RECT 134.200 195.800 135.400 199.800 ;
        RECT 124.400 195.000 125.200 195.800 ;
        RECT 130.000 195.200 130.600 195.800 ;
        RECT 127.800 194.600 131.400 195.200 ;
        RECT 134.000 195.000 134.800 195.800 ;
        RECT 127.800 194.400 128.600 194.600 ;
        RECT 130.600 194.400 131.400 194.600 ;
        RECT 124.400 193.000 125.200 193.200 ;
        RECT 129.000 193.000 129.800 193.200 ;
        RECT 124.400 192.400 129.800 193.000 ;
        RECT 130.400 193.000 132.600 193.600 ;
        RECT 130.400 191.800 131.000 193.000 ;
        RECT 131.800 192.800 132.600 193.000 ;
        RECT 134.200 193.200 135.600 194.000 ;
        RECT 134.200 192.200 134.800 193.200 ;
        RECT 126.200 191.400 131.000 191.800 ;
        RECT 121.200 191.200 131.000 191.400 ;
        RECT 132.400 191.600 134.800 192.200 ;
        RECT 121.200 191.000 127.000 191.200 ;
        RECT 121.200 190.800 126.800 191.000 ;
        RECT 118.000 188.800 118.800 190.400 ;
        RECT 127.600 190.300 128.400 190.400 ;
        RECT 130.800 190.300 131.600 190.400 ;
        RECT 127.600 190.200 131.600 190.300 ;
        RECT 123.400 189.700 131.600 190.200 ;
        RECT 123.400 189.600 128.400 189.700 ;
        RECT 130.800 189.600 131.600 189.700 ;
        RECT 123.400 189.400 124.200 189.600 ;
        RECT 125.000 188.400 125.800 188.600 ;
        RECT 132.400 188.400 133.000 191.600 ;
        RECT 138.800 191.200 139.600 199.800 ;
        RECT 135.400 190.600 139.600 191.200 ;
        RECT 135.400 190.400 136.200 190.600 ;
        RECT 137.000 189.800 137.800 190.000 ;
        RECT 134.000 189.200 137.800 189.800 ;
        RECT 134.000 189.000 134.800 189.200 ;
        RECT 108.400 186.800 109.200 188.400 ;
        RECT 114.800 187.600 117.400 188.400 ;
        RECT 119.600 188.200 120.400 188.400 ;
        RECT 118.800 187.600 120.400 188.200 ;
        RECT 122.000 187.800 133.000 188.400 ;
        RECT 122.000 187.600 123.600 187.800 ;
        RECT 115.000 186.200 115.600 187.600 ;
        RECT 118.800 187.200 119.600 187.600 ;
        RECT 116.600 186.200 120.200 186.600 ;
        RECT 105.800 185.600 107.600 186.200 ;
        RECT 105.800 182.200 106.600 185.600 ;
        RECT 114.800 182.200 115.600 186.200 ;
        RECT 116.400 186.000 120.400 186.200 ;
        RECT 116.400 182.200 117.200 186.000 ;
        RECT 119.600 182.200 120.400 186.000 ;
        RECT 121.200 182.200 122.000 187.000 ;
        RECT 126.200 185.600 126.800 187.800 ;
        RECT 131.800 187.600 132.600 187.800 ;
        RECT 138.800 187.200 139.600 190.600 ;
        RECT 135.800 186.600 139.600 187.200 ;
        RECT 135.800 186.400 136.600 186.600 ;
        RECT 124.400 184.200 125.200 185.000 ;
        RECT 126.000 184.800 126.800 185.600 ;
        RECT 127.800 185.400 128.600 185.600 ;
        RECT 127.800 184.800 130.600 185.400 ;
        RECT 130.000 184.200 130.600 184.800 ;
        RECT 134.000 184.200 134.800 185.000 ;
        RECT 124.400 183.600 126.400 184.200 ;
        RECT 125.600 182.200 126.400 183.600 ;
        RECT 130.000 182.200 130.800 184.200 ;
        RECT 134.000 183.600 135.400 184.200 ;
        RECT 134.200 182.200 135.400 183.600 ;
        RECT 138.800 182.200 139.600 186.600 ;
        RECT 140.400 182.200 141.200 199.800 ;
        RECT 143.600 191.400 144.400 199.800 ;
        RECT 148.000 196.400 148.800 199.800 ;
        RECT 146.800 195.800 148.800 196.400 ;
        RECT 152.400 195.800 153.200 199.800 ;
        RECT 156.600 195.800 157.800 199.800 ;
        RECT 146.800 195.000 147.600 195.800 ;
        RECT 152.400 195.200 153.000 195.800 ;
        RECT 150.200 194.600 153.800 195.200 ;
        RECT 156.400 195.000 157.200 195.800 ;
        RECT 150.200 194.400 151.000 194.600 ;
        RECT 153.000 194.400 153.800 194.600 ;
        RECT 146.800 193.000 147.600 193.200 ;
        RECT 151.400 193.000 152.200 193.200 ;
        RECT 146.800 192.400 152.200 193.000 ;
        RECT 152.800 193.000 155.000 193.600 ;
        RECT 152.800 191.800 153.400 193.000 ;
        RECT 154.200 192.800 155.000 193.000 ;
        RECT 156.600 193.200 158.000 194.000 ;
        RECT 156.600 192.200 157.200 193.200 ;
        RECT 148.600 191.400 153.400 191.800 ;
        RECT 143.600 191.200 153.400 191.400 ;
        RECT 154.800 191.600 157.200 192.200 ;
        RECT 143.600 191.000 149.400 191.200 ;
        RECT 143.600 190.800 149.200 191.000 ;
        RECT 150.000 190.300 150.800 190.400 ;
        RECT 153.200 190.300 154.000 190.400 ;
        RECT 150.000 190.200 154.000 190.300 ;
        RECT 145.800 189.700 154.000 190.200 ;
        RECT 145.800 189.600 150.800 189.700 ;
        RECT 153.200 189.600 154.000 189.700 ;
        RECT 145.800 189.400 146.600 189.600 ;
        RECT 147.400 188.400 148.200 188.600 ;
        RECT 154.800 188.400 155.400 191.600 ;
        RECT 161.200 191.200 162.000 199.800 ;
        RECT 157.800 190.600 162.000 191.200 ;
        RECT 162.800 191.400 163.600 199.800 ;
        RECT 167.200 196.400 168.000 199.800 ;
        RECT 166.000 195.800 168.000 196.400 ;
        RECT 171.600 195.800 172.400 199.800 ;
        RECT 175.800 195.800 177.000 199.800 ;
        RECT 166.000 195.000 166.800 195.800 ;
        RECT 171.600 195.200 172.200 195.800 ;
        RECT 169.400 194.600 173.000 195.200 ;
        RECT 175.600 195.000 176.400 195.800 ;
        RECT 169.400 194.400 170.200 194.600 ;
        RECT 172.200 194.400 173.000 194.600 ;
        RECT 166.000 193.000 166.800 193.200 ;
        RECT 170.600 193.000 171.400 193.200 ;
        RECT 166.000 192.400 171.400 193.000 ;
        RECT 172.000 193.000 174.200 193.600 ;
        RECT 172.000 191.800 172.600 193.000 ;
        RECT 173.400 192.800 174.200 193.000 ;
        RECT 175.800 193.200 177.200 194.000 ;
        RECT 175.800 192.200 176.400 193.200 ;
        RECT 167.800 191.400 172.600 191.800 ;
        RECT 162.800 191.200 172.600 191.400 ;
        RECT 174.000 191.600 176.400 192.200 ;
        RECT 162.800 191.000 168.600 191.200 ;
        RECT 162.800 190.800 168.400 191.000 ;
        RECT 157.800 190.400 158.600 190.600 ;
        RECT 159.400 189.800 160.200 190.000 ;
        RECT 156.400 189.200 160.200 189.800 ;
        RECT 156.400 189.000 157.200 189.200 ;
        RECT 144.400 187.800 155.400 188.400 ;
        RECT 144.400 187.600 146.000 187.800 ;
        RECT 142.000 184.800 142.800 186.400 ;
        RECT 143.600 182.200 144.400 187.000 ;
        RECT 148.600 185.600 149.200 187.800 ;
        RECT 150.000 187.600 150.800 187.800 ;
        RECT 154.200 187.600 155.000 187.800 ;
        RECT 161.200 187.200 162.000 190.600 ;
        RECT 169.200 190.200 170.000 190.400 ;
        RECT 165.000 189.600 170.000 190.200 ;
        RECT 165.000 189.400 165.800 189.600 ;
        RECT 166.600 188.400 167.400 188.600 ;
        RECT 174.000 188.400 174.600 191.600 ;
        RECT 180.400 191.200 181.200 199.800 ;
        RECT 183.600 192.000 184.400 199.800 ;
        RECT 186.800 195.200 187.600 199.800 ;
        RECT 177.000 190.600 181.200 191.200 ;
        RECT 177.000 190.400 177.800 190.600 ;
        RECT 178.600 189.800 179.400 190.000 ;
        RECT 175.600 189.200 179.400 189.800 ;
        RECT 175.600 189.000 176.400 189.200 ;
        RECT 163.600 187.800 174.600 188.400 ;
        RECT 163.600 187.600 165.200 187.800 ;
        RECT 158.200 186.600 162.000 187.200 ;
        RECT 158.200 186.400 159.000 186.600 ;
        RECT 146.800 184.200 147.600 185.000 ;
        RECT 148.400 184.800 149.200 185.600 ;
        RECT 150.200 185.400 151.000 185.600 ;
        RECT 150.200 184.800 153.000 185.400 ;
        RECT 152.400 184.200 153.000 184.800 ;
        RECT 156.400 184.200 157.200 185.000 ;
        RECT 146.800 183.600 148.800 184.200 ;
        RECT 148.000 182.200 148.800 183.600 ;
        RECT 152.400 182.200 153.200 184.200 ;
        RECT 156.400 183.600 157.800 184.200 ;
        RECT 156.600 182.200 157.800 183.600 ;
        RECT 161.200 182.200 162.000 186.600 ;
        RECT 162.800 182.200 163.600 187.000 ;
        RECT 167.800 185.600 168.400 187.800 ;
        RECT 173.400 187.600 174.200 187.800 ;
        RECT 180.400 187.200 181.200 190.600 ;
        RECT 177.400 186.600 181.200 187.200 ;
        RECT 177.400 186.400 178.200 186.600 ;
        RECT 166.000 184.200 166.800 185.000 ;
        RECT 167.600 184.800 168.400 185.600 ;
        RECT 169.400 185.400 170.200 185.600 ;
        RECT 169.400 184.800 172.200 185.400 ;
        RECT 171.600 184.200 172.200 184.800 ;
        RECT 175.600 184.200 176.400 185.000 ;
        RECT 166.000 183.600 168.000 184.200 ;
        RECT 167.200 182.200 168.000 183.600 ;
        RECT 171.600 182.200 172.400 184.200 ;
        RECT 175.600 183.600 177.000 184.200 ;
        RECT 175.800 182.200 177.000 183.600 ;
        RECT 180.400 182.200 181.200 186.600 ;
        RECT 183.400 191.200 184.400 192.000 ;
        RECT 185.000 194.600 187.600 195.200 ;
        RECT 185.000 193.000 185.600 194.600 ;
        RECT 190.000 194.400 190.800 199.800 ;
        RECT 193.200 197.000 194.000 199.800 ;
        RECT 194.800 197.000 195.600 199.800 ;
        RECT 196.400 197.000 197.200 199.800 ;
        RECT 191.400 194.400 195.600 195.200 ;
        RECT 188.200 193.600 190.800 194.400 ;
        RECT 198.000 193.600 198.800 199.800 ;
        RECT 201.200 195.000 202.000 199.800 ;
        RECT 204.400 195.000 205.200 199.800 ;
        RECT 206.000 197.000 206.800 199.800 ;
        RECT 207.600 197.000 208.400 199.800 ;
        RECT 210.800 195.200 211.600 199.800 ;
        RECT 214.000 196.400 214.800 199.800 ;
        RECT 214.000 195.800 215.000 196.400 ;
        RECT 214.400 195.200 215.000 195.800 ;
        RECT 209.600 194.400 213.800 195.200 ;
        RECT 214.400 194.600 216.400 195.200 ;
        RECT 201.200 193.600 203.800 194.400 ;
        RECT 204.400 193.800 210.200 194.400 ;
        RECT 213.200 194.000 213.800 194.400 ;
        RECT 193.200 193.000 194.000 193.200 ;
        RECT 185.000 192.400 194.000 193.000 ;
        RECT 196.400 193.000 197.200 193.200 ;
        RECT 204.400 193.000 205.000 193.800 ;
        RECT 210.800 193.200 212.200 193.800 ;
        RECT 213.200 193.200 214.800 194.000 ;
        RECT 196.400 192.400 205.000 193.000 ;
        RECT 206.000 193.000 212.200 193.200 ;
        RECT 206.000 192.600 211.400 193.000 ;
        RECT 206.000 192.400 206.800 192.600 ;
        RECT 183.400 186.800 184.200 191.200 ;
        RECT 185.000 190.600 185.600 192.400 ;
        RECT 184.800 190.000 185.600 190.600 ;
        RECT 191.600 190.000 215.000 190.600 ;
        RECT 184.800 188.000 185.400 190.000 ;
        RECT 191.600 189.400 192.400 190.000 ;
        RECT 209.200 189.600 210.000 190.000 ;
        RECT 210.800 189.600 211.600 190.000 ;
        RECT 214.200 189.800 215.000 190.000 ;
        RECT 186.000 188.600 189.800 189.400 ;
        RECT 184.800 187.400 186.000 188.000 ;
        RECT 183.400 186.000 184.400 186.800 ;
        RECT 183.600 182.200 184.400 186.000 ;
        RECT 185.200 182.200 186.000 187.400 ;
        RECT 189.000 187.400 189.800 188.600 ;
        RECT 189.000 186.800 190.800 187.400 ;
        RECT 190.000 186.200 190.800 186.800 ;
        RECT 194.800 186.400 195.600 189.200 ;
        RECT 198.000 188.600 201.200 189.400 ;
        RECT 205.000 188.600 207.000 189.400 ;
        RECT 215.600 189.000 216.400 194.600 ;
        RECT 217.800 192.600 218.600 199.800 ;
        RECT 217.800 191.800 219.600 192.600 ;
        RECT 222.000 191.800 222.800 199.800 ;
        RECT 223.600 192.400 224.400 199.800 ;
        RECT 226.800 192.400 227.600 199.800 ;
        RECT 223.600 191.800 227.600 192.400 ;
        RECT 230.000 192.000 230.800 199.800 ;
        RECT 233.200 195.200 234.000 199.800 ;
        RECT 217.200 189.600 218.000 191.200 ;
        RECT 197.600 187.800 198.400 188.000 ;
        RECT 197.600 187.200 202.000 187.800 ;
        RECT 201.200 187.000 202.000 187.200 ;
        RECT 202.800 186.800 203.600 188.400 ;
        RECT 190.000 185.400 192.400 186.200 ;
        RECT 194.800 185.600 195.800 186.400 ;
        RECT 198.800 185.600 200.400 186.400 ;
        RECT 201.200 186.200 202.000 186.400 ;
        RECT 205.000 186.200 205.800 188.600 ;
        RECT 207.600 188.200 216.400 189.000 ;
        RECT 211.000 186.800 214.000 187.600 ;
        RECT 211.000 186.200 211.800 186.800 ;
        RECT 201.200 185.600 205.800 186.200 ;
        RECT 191.600 182.200 192.400 185.400 ;
        RECT 209.200 185.400 211.800 186.200 ;
        RECT 193.200 182.200 194.000 185.000 ;
        RECT 194.800 182.200 195.600 185.000 ;
        RECT 196.400 182.200 197.200 185.000 ;
        RECT 198.000 182.200 198.800 185.000 ;
        RECT 201.200 182.200 202.000 185.000 ;
        RECT 204.400 182.200 205.200 185.000 ;
        RECT 206.000 182.200 206.800 185.000 ;
        RECT 207.600 182.200 208.400 185.000 ;
        RECT 209.200 182.200 210.000 185.400 ;
        RECT 215.600 182.200 216.400 188.200 ;
        RECT 218.800 188.400 219.400 191.800 ;
        RECT 222.200 190.400 222.800 191.800 ;
        RECT 229.800 191.200 230.800 192.000 ;
        RECT 231.400 194.600 234.000 195.200 ;
        RECT 231.400 193.000 232.000 194.600 ;
        RECT 236.400 194.400 237.200 199.800 ;
        RECT 239.600 197.000 240.400 199.800 ;
        RECT 241.200 197.000 242.000 199.800 ;
        RECT 242.800 197.000 243.600 199.800 ;
        RECT 237.800 194.400 242.000 195.200 ;
        RECT 234.600 193.600 237.200 194.400 ;
        RECT 244.400 193.600 245.200 199.800 ;
        RECT 247.600 195.000 248.400 199.800 ;
        RECT 250.800 195.000 251.600 199.800 ;
        RECT 252.400 197.000 253.200 199.800 ;
        RECT 254.000 197.000 254.800 199.800 ;
        RECT 257.200 195.200 258.000 199.800 ;
        RECT 260.400 196.400 261.200 199.800 ;
        RECT 260.400 195.800 261.400 196.400 ;
        RECT 260.800 195.200 261.400 195.800 ;
        RECT 256.000 194.400 260.200 195.200 ;
        RECT 260.800 194.600 262.800 195.200 ;
        RECT 247.600 193.600 250.200 194.400 ;
        RECT 250.800 193.800 256.600 194.400 ;
        RECT 259.600 194.000 260.200 194.400 ;
        RECT 239.600 193.000 240.400 193.200 ;
        RECT 231.400 192.400 240.400 193.000 ;
        RECT 242.800 193.000 243.600 193.200 ;
        RECT 250.800 193.000 251.400 193.800 ;
        RECT 257.200 193.200 258.600 193.800 ;
        RECT 259.600 193.200 261.200 194.000 ;
        RECT 242.800 192.400 251.400 193.000 ;
        RECT 252.400 193.000 258.600 193.200 ;
        RECT 252.400 192.600 257.800 193.000 ;
        RECT 252.400 192.400 253.200 192.600 ;
        RECT 226.000 190.400 226.800 190.800 ;
        RECT 222.000 189.800 224.400 190.400 ;
        RECT 226.000 189.800 227.600 190.400 ;
        RECT 222.000 189.600 222.800 189.800 ;
        RECT 218.800 188.300 219.600 188.400 ;
        RECT 218.800 187.700 222.700 188.300 ;
        RECT 218.800 187.600 219.600 187.700 ;
        RECT 218.800 184.200 219.400 187.600 ;
        RECT 222.100 186.400 222.700 187.700 ;
        RECT 223.800 186.400 224.400 189.800 ;
        RECT 226.800 189.600 227.600 189.800 ;
        RECT 225.200 187.600 226.000 189.200 ;
        RECT 220.400 184.800 221.200 186.400 ;
        RECT 222.000 185.600 222.800 186.400 ;
        RECT 222.200 184.800 223.000 185.600 ;
        RECT 218.800 182.200 219.600 184.200 ;
        RECT 223.600 182.200 224.400 186.400 ;
        RECT 229.800 186.800 230.600 191.200 ;
        RECT 231.400 190.600 232.000 192.400 ;
        RECT 231.200 190.000 232.000 190.600 ;
        RECT 238.000 190.000 261.400 190.600 ;
        RECT 231.200 188.000 231.800 190.000 ;
        RECT 238.000 189.400 238.800 190.000 ;
        RECT 255.600 189.600 256.400 190.000 ;
        RECT 260.600 189.800 261.400 190.000 ;
        RECT 232.400 188.600 236.200 189.400 ;
        RECT 231.200 187.400 232.400 188.000 ;
        RECT 229.800 186.000 230.800 186.800 ;
        RECT 230.000 182.200 230.800 186.000 ;
        RECT 231.600 182.200 232.400 187.400 ;
        RECT 235.400 187.400 236.200 188.600 ;
        RECT 235.400 186.800 237.200 187.400 ;
        RECT 236.400 186.200 237.200 186.800 ;
        RECT 241.200 186.400 242.000 189.200 ;
        RECT 244.400 188.600 247.600 189.400 ;
        RECT 251.400 188.600 253.400 189.400 ;
        RECT 262.000 189.000 262.800 194.600 ;
        RECT 270.000 192.000 270.800 199.800 ;
        RECT 273.200 195.200 274.000 199.800 ;
        RECT 244.000 187.800 244.800 188.000 ;
        RECT 244.000 187.200 248.400 187.800 ;
        RECT 247.600 187.000 248.400 187.200 ;
        RECT 249.200 186.800 250.000 188.400 ;
        RECT 236.400 185.400 238.800 186.200 ;
        RECT 241.200 185.600 242.200 186.400 ;
        RECT 245.200 185.600 246.800 186.400 ;
        RECT 247.600 186.200 248.400 186.400 ;
        RECT 251.400 186.200 252.200 188.600 ;
        RECT 254.000 188.200 262.800 189.000 ;
        RECT 257.400 186.800 260.400 187.600 ;
        RECT 257.400 186.200 258.200 186.800 ;
        RECT 247.600 185.600 252.200 186.200 ;
        RECT 238.000 182.200 238.800 185.400 ;
        RECT 255.600 185.400 258.200 186.200 ;
        RECT 239.600 182.200 240.400 185.000 ;
        RECT 241.200 182.200 242.000 185.000 ;
        RECT 242.800 182.200 243.600 185.000 ;
        RECT 244.400 182.200 245.200 185.000 ;
        RECT 247.600 182.200 248.400 185.000 ;
        RECT 250.800 182.200 251.600 185.000 ;
        RECT 252.400 182.200 253.200 185.000 ;
        RECT 254.000 182.200 254.800 185.000 ;
        RECT 255.600 182.200 256.400 185.400 ;
        RECT 262.000 182.200 262.800 188.200 ;
        RECT 269.800 191.200 270.800 192.000 ;
        RECT 271.400 194.600 274.000 195.200 ;
        RECT 271.400 193.000 272.000 194.600 ;
        RECT 276.400 194.400 277.200 199.800 ;
        RECT 279.600 197.000 280.400 199.800 ;
        RECT 281.200 197.000 282.000 199.800 ;
        RECT 282.800 197.000 283.600 199.800 ;
        RECT 277.800 194.400 282.000 195.200 ;
        RECT 274.600 193.600 277.200 194.400 ;
        RECT 284.400 193.600 285.200 199.800 ;
        RECT 287.600 195.000 288.400 199.800 ;
        RECT 290.800 195.000 291.600 199.800 ;
        RECT 292.400 197.000 293.200 199.800 ;
        RECT 294.000 197.000 294.800 199.800 ;
        RECT 297.200 195.200 298.000 199.800 ;
        RECT 300.400 196.400 301.200 199.800 ;
        RECT 300.400 195.800 301.400 196.400 ;
        RECT 300.800 195.200 301.400 195.800 ;
        RECT 296.000 194.400 300.200 195.200 ;
        RECT 300.800 194.600 302.800 195.200 ;
        RECT 287.600 193.600 290.200 194.400 ;
        RECT 290.800 193.800 296.600 194.400 ;
        RECT 299.600 194.000 300.200 194.400 ;
        RECT 279.600 193.000 280.400 193.200 ;
        RECT 271.400 192.400 280.400 193.000 ;
        RECT 282.800 193.000 283.600 193.200 ;
        RECT 290.800 193.000 291.400 193.800 ;
        RECT 297.200 193.200 298.600 193.800 ;
        RECT 299.600 193.200 301.200 194.000 ;
        RECT 282.800 192.400 291.400 193.000 ;
        RECT 292.400 193.000 298.600 193.200 ;
        RECT 292.400 192.600 297.800 193.000 ;
        RECT 292.400 192.400 293.200 192.600 ;
        RECT 269.800 186.800 270.600 191.200 ;
        RECT 271.400 190.600 272.000 192.400 ;
        RECT 271.200 190.000 272.000 190.600 ;
        RECT 278.000 190.000 301.400 190.600 ;
        RECT 271.200 188.000 271.800 190.000 ;
        RECT 278.000 189.400 278.800 190.000 ;
        RECT 295.600 189.600 296.400 190.000 ;
        RECT 300.400 189.800 301.400 190.000 ;
        RECT 300.400 189.600 301.200 189.800 ;
        RECT 272.400 188.600 276.200 189.400 ;
        RECT 271.200 187.400 272.400 188.000 ;
        RECT 269.800 186.000 270.800 186.800 ;
        RECT 270.000 182.200 270.800 186.000 ;
        RECT 271.600 182.200 272.400 187.400 ;
        RECT 275.400 187.400 276.200 188.600 ;
        RECT 275.400 186.800 277.200 187.400 ;
        RECT 276.400 186.200 277.200 186.800 ;
        RECT 281.200 186.400 282.000 189.200 ;
        RECT 284.400 188.600 287.600 189.400 ;
        RECT 291.400 188.600 293.400 189.400 ;
        RECT 302.000 189.000 302.800 194.600 ;
        RECT 284.000 187.800 284.800 188.000 ;
        RECT 284.000 187.200 288.400 187.800 ;
        RECT 287.600 187.000 288.400 187.200 ;
        RECT 289.200 186.800 290.000 188.400 ;
        RECT 276.400 185.400 278.800 186.200 ;
        RECT 281.200 185.600 282.200 186.400 ;
        RECT 285.200 185.600 286.800 186.400 ;
        RECT 287.600 186.200 288.400 186.400 ;
        RECT 291.400 186.200 292.200 188.600 ;
        RECT 294.000 188.200 302.800 189.000 ;
        RECT 297.400 186.800 300.400 187.600 ;
        RECT 297.400 186.200 298.200 186.800 ;
        RECT 287.600 185.600 292.200 186.200 ;
        RECT 278.000 182.200 278.800 185.400 ;
        RECT 295.600 185.400 298.200 186.200 ;
        RECT 279.600 182.200 280.400 185.000 ;
        RECT 281.200 182.200 282.000 185.000 ;
        RECT 282.800 182.200 283.600 185.000 ;
        RECT 284.400 182.200 285.200 185.000 ;
        RECT 287.600 182.200 288.400 185.000 ;
        RECT 290.800 182.200 291.600 185.000 ;
        RECT 292.400 182.200 293.200 185.000 ;
        RECT 294.000 182.200 294.800 185.000 ;
        RECT 295.600 182.200 296.400 185.400 ;
        RECT 302.000 182.200 302.800 188.200 ;
        RECT 303.600 182.200 304.400 199.800 ;
        RECT 308.400 196.400 309.200 199.800 ;
        RECT 308.200 195.800 309.200 196.400 ;
        RECT 308.200 195.200 308.800 195.800 ;
        RECT 311.600 195.200 312.400 199.800 ;
        RECT 314.800 197.000 315.600 199.800 ;
        RECT 316.400 197.000 317.200 199.800 ;
        RECT 306.800 194.600 308.800 195.200 ;
        RECT 306.800 189.000 307.600 194.600 ;
        RECT 309.400 194.400 313.600 195.200 ;
        RECT 318.000 195.000 318.800 199.800 ;
        RECT 321.200 195.000 322.000 199.800 ;
        RECT 309.400 194.000 310.000 194.400 ;
        RECT 308.400 193.200 310.000 194.000 ;
        RECT 313.000 193.800 318.800 194.400 ;
        RECT 311.000 193.200 312.400 193.800 ;
        RECT 311.000 193.000 317.200 193.200 ;
        RECT 311.800 192.600 317.200 193.000 ;
        RECT 316.400 192.400 317.200 192.600 ;
        RECT 318.200 193.000 318.800 193.800 ;
        RECT 319.400 193.600 322.000 194.400 ;
        RECT 324.400 193.600 325.200 199.800 ;
        RECT 326.000 197.000 326.800 199.800 ;
        RECT 327.600 197.000 328.400 199.800 ;
        RECT 329.200 197.000 330.000 199.800 ;
        RECT 327.600 194.400 331.800 195.200 ;
        RECT 332.400 194.400 333.200 199.800 ;
        RECT 335.600 195.200 336.400 199.800 ;
        RECT 335.600 194.600 338.200 195.200 ;
        RECT 332.400 193.600 335.000 194.400 ;
        RECT 326.000 193.000 326.800 193.200 ;
        RECT 318.200 192.400 326.800 193.000 ;
        RECT 329.200 193.000 330.000 193.200 ;
        RECT 337.600 193.000 338.200 194.600 ;
        RECT 329.200 192.400 338.200 193.000 ;
        RECT 337.600 190.600 338.200 192.400 ;
        RECT 338.800 192.000 339.600 199.800 ;
        RECT 340.400 192.300 341.200 192.400 ;
        RECT 342.000 192.300 342.800 193.200 ;
        RECT 338.800 191.200 339.800 192.000 ;
        RECT 340.400 191.700 342.800 192.300 ;
        RECT 340.400 191.600 341.200 191.700 ;
        RECT 342.000 191.600 342.800 191.700 ;
        RECT 308.200 190.000 331.600 190.600 ;
        RECT 337.600 190.000 338.400 190.600 ;
        RECT 308.200 189.800 309.000 190.000 ;
        RECT 310.000 189.600 310.800 190.000 ;
        RECT 313.200 189.600 314.000 190.000 ;
        RECT 330.800 189.400 331.600 190.000 ;
        RECT 306.800 188.200 315.600 189.000 ;
        RECT 316.200 188.600 318.200 189.400 ;
        RECT 322.000 188.600 325.200 189.400 ;
        RECT 305.200 184.800 306.000 186.400 ;
        RECT 306.800 182.200 307.600 188.200 ;
        RECT 309.200 186.800 312.200 187.600 ;
        RECT 311.400 186.200 312.200 186.800 ;
        RECT 317.400 186.200 318.200 188.600 ;
        RECT 319.600 186.800 320.400 188.400 ;
        RECT 324.800 187.800 325.600 188.000 ;
        RECT 321.200 187.200 325.600 187.800 ;
        RECT 321.200 187.000 322.000 187.200 ;
        RECT 327.600 186.400 328.400 189.200 ;
        RECT 333.400 188.600 337.200 189.400 ;
        RECT 333.400 187.400 334.200 188.600 ;
        RECT 337.800 188.000 338.400 190.000 ;
        RECT 321.200 186.200 322.000 186.400 ;
        RECT 311.400 185.400 314.000 186.200 ;
        RECT 317.400 185.600 322.000 186.200 ;
        RECT 322.800 185.600 324.400 186.400 ;
        RECT 327.400 185.600 328.400 186.400 ;
        RECT 332.400 186.800 334.200 187.400 ;
        RECT 337.200 187.400 338.400 188.000 ;
        RECT 332.400 186.200 333.200 186.800 ;
        RECT 313.200 182.200 314.000 185.400 ;
        RECT 330.800 185.400 333.200 186.200 ;
        RECT 314.800 182.200 315.600 185.000 ;
        RECT 316.400 182.200 317.200 185.000 ;
        RECT 318.000 182.200 318.800 185.000 ;
        RECT 321.200 182.200 322.000 185.000 ;
        RECT 324.400 182.200 325.200 185.000 ;
        RECT 326.000 182.200 326.800 185.000 ;
        RECT 327.600 182.200 328.400 185.000 ;
        RECT 329.200 182.200 330.000 185.000 ;
        RECT 330.800 182.200 331.600 185.400 ;
        RECT 337.200 182.200 338.000 187.400 ;
        RECT 339.000 186.800 339.800 191.200 ;
        RECT 340.400 190.300 341.200 190.400 ;
        RECT 343.600 190.300 344.400 199.800 ;
        RECT 346.800 191.600 347.600 193.200 ;
        RECT 340.400 189.700 344.400 190.300 ;
        RECT 340.400 189.600 341.200 189.700 ;
        RECT 338.800 186.000 339.800 186.800 ;
        RECT 343.600 186.200 344.400 189.700 ;
        RECT 345.200 188.300 346.000 188.400 ;
        RECT 348.400 188.300 349.200 199.800 ;
        RECT 345.200 187.700 349.200 188.300 ;
        RECT 345.200 186.800 346.000 187.700 ;
        RECT 348.400 186.200 349.200 187.700 ;
        RECT 350.000 188.300 350.800 188.400 ;
        RECT 351.600 188.300 352.400 188.400 ;
        RECT 350.000 187.700 352.400 188.300 ;
        RECT 350.000 186.800 350.800 187.700 ;
        RECT 351.600 186.800 352.400 187.700 ;
        RECT 338.800 182.200 339.600 186.000 ;
        RECT 342.600 185.600 344.400 186.200 ;
        RECT 347.400 185.600 349.200 186.200 ;
        RECT 342.600 182.200 343.400 185.600 ;
        RECT 347.400 182.200 348.200 185.600 ;
        RECT 353.200 182.200 354.000 199.800 ;
        RECT 356.400 191.200 357.200 199.800 ;
        RECT 359.600 191.200 360.400 199.800 ;
        RECT 362.800 191.200 363.600 199.800 ;
        RECT 366.000 191.200 366.800 199.800 ;
        RECT 354.800 190.400 357.200 191.200 ;
        RECT 358.200 190.400 360.400 191.200 ;
        RECT 361.400 190.400 363.600 191.200 ;
        RECT 365.000 190.400 366.800 191.200 ;
        RECT 354.800 187.600 355.600 190.400 ;
        RECT 358.200 189.000 359.000 190.400 ;
        RECT 361.400 189.000 362.200 190.400 ;
        RECT 365.000 189.000 365.800 190.400 ;
        RECT 356.400 188.200 359.000 189.000 ;
        RECT 359.800 188.200 362.200 189.000 ;
        RECT 363.200 188.200 365.800 189.000 ;
        RECT 366.600 188.200 368.400 189.000 ;
        RECT 358.200 187.600 359.000 188.200 ;
        RECT 361.400 187.600 362.200 188.200 ;
        RECT 365.000 187.600 365.800 188.200 ;
        RECT 367.600 187.600 368.400 188.200 ;
        RECT 354.800 186.800 357.200 187.600 ;
        RECT 358.200 186.800 360.400 187.600 ;
        RECT 361.400 186.800 363.600 187.600 ;
        RECT 365.000 186.800 366.800 187.600 ;
        RECT 369.200 186.800 370.000 188.400 ;
        RECT 356.400 182.200 357.200 186.800 ;
        RECT 359.600 182.200 360.400 186.800 ;
        RECT 362.800 182.200 363.600 186.800 ;
        RECT 366.000 182.200 366.800 186.800 ;
        RECT 370.800 182.200 371.600 199.800 ;
        RECT 372.400 186.800 373.200 188.400 ;
        RECT 374.000 188.300 374.800 199.800 ;
        RECT 375.600 191.600 376.400 193.200 ;
        RECT 377.200 188.300 378.000 188.400 ;
        RECT 374.000 187.700 378.000 188.300 ;
        RECT 374.000 186.200 374.800 187.700 ;
        RECT 377.200 186.800 378.000 187.700 ;
        RECT 378.800 186.200 379.600 199.800 ;
        RECT 380.400 191.600 381.200 193.200 ;
        RECT 384.600 191.800 386.600 199.800 ;
        RECT 382.000 187.600 382.800 189.200 ;
        RECT 383.600 188.800 384.400 190.400 ;
        RECT 385.400 188.400 386.000 191.800 ;
        RECT 390.000 191.600 390.800 193.200 ;
        RECT 386.800 190.300 387.600 190.400 ;
        RECT 391.600 190.300 392.400 199.800 ;
        RECT 396.400 195.800 397.200 199.800 ;
        RECT 396.600 195.600 397.200 195.800 ;
        RECT 399.600 195.800 400.400 199.800 ;
        RECT 402.800 195.800 403.600 199.800 ;
        RECT 399.600 195.600 400.200 195.800 ;
        RECT 396.600 195.000 400.200 195.600 ;
        RECT 403.000 195.600 403.600 195.800 ;
        RECT 406.000 195.800 406.800 199.800 ;
        RECT 406.000 195.600 406.600 195.800 ;
        RECT 403.000 195.000 406.600 195.600 ;
        RECT 398.000 192.800 398.800 194.400 ;
        RECT 399.600 192.400 400.200 195.000 ;
        RECT 404.400 192.800 405.200 194.400 ;
        RECT 406.000 192.400 406.600 195.000 ;
        RECT 393.200 192.300 394.000 192.400 ;
        RECT 394.800 192.300 395.600 192.400 ;
        RECT 393.200 191.700 395.600 192.300 ;
        RECT 393.200 191.600 394.000 191.700 ;
        RECT 394.800 190.800 395.600 191.700 ;
        RECT 399.600 191.600 400.400 192.400 ;
        RECT 386.800 189.700 392.400 190.300 ;
        RECT 386.800 188.800 387.600 189.700 ;
        RECT 385.200 188.200 386.000 188.400 ;
        RECT 388.400 188.200 389.200 188.400 ;
        RECT 383.600 187.600 386.000 188.200 ;
        RECT 387.600 187.600 389.200 188.200 ;
        RECT 383.600 186.200 384.200 187.600 ;
        RECT 387.600 187.200 388.400 187.600 ;
        RECT 385.400 186.200 389.000 186.600 ;
        RECT 391.600 186.200 392.400 189.700 ;
        RECT 396.400 189.600 398.000 190.400 ;
        RECT 399.600 188.400 400.200 191.600 ;
        RECT 401.200 190.800 402.000 192.400 ;
        RECT 406.000 191.600 406.800 192.400 ;
        RECT 402.800 189.600 404.400 190.400 ;
        RECT 406.000 188.400 406.600 191.600 ;
        RECT 409.200 191.200 410.000 199.800 ;
        RECT 412.400 191.200 413.200 199.800 ;
        RECT 415.600 191.200 416.400 199.800 ;
        RECT 418.800 191.200 419.600 199.800 ;
        RECT 428.400 192.000 429.200 199.800 ;
        RECT 431.600 195.200 432.400 199.800 ;
        RECT 393.200 186.800 394.000 188.400 ;
        RECT 398.600 188.200 400.200 188.400 ;
        RECT 405.000 188.200 406.600 188.400 ;
        RECT 398.400 187.800 400.200 188.200 ;
        RECT 404.800 187.800 406.600 188.200 ;
        RECT 407.600 190.400 410.000 191.200 ;
        RECT 411.000 190.400 413.200 191.200 ;
        RECT 414.200 190.400 416.400 191.200 ;
        RECT 417.800 190.400 419.600 191.200 ;
        RECT 428.200 191.200 429.200 192.000 ;
        RECT 429.800 194.600 432.400 195.200 ;
        RECT 429.800 193.000 430.400 194.600 ;
        RECT 434.800 194.400 435.600 199.800 ;
        RECT 438.000 197.000 438.800 199.800 ;
        RECT 439.600 197.000 440.400 199.800 ;
        RECT 441.200 197.000 442.000 199.800 ;
        RECT 436.200 194.400 440.400 195.200 ;
        RECT 433.000 193.600 435.600 194.400 ;
        RECT 442.800 193.600 443.600 199.800 ;
        RECT 446.000 195.000 446.800 199.800 ;
        RECT 449.200 195.000 450.000 199.800 ;
        RECT 450.800 197.000 451.600 199.800 ;
        RECT 452.400 197.000 453.200 199.800 ;
        RECT 455.600 195.200 456.400 199.800 ;
        RECT 458.800 196.400 459.600 199.800 ;
        RECT 458.800 195.800 459.800 196.400 ;
        RECT 459.200 195.200 459.800 195.800 ;
        RECT 454.400 194.400 458.600 195.200 ;
        RECT 459.200 194.600 461.200 195.200 ;
        RECT 446.000 193.600 448.600 194.400 ;
        RECT 449.200 193.800 455.000 194.400 ;
        RECT 458.000 194.000 458.600 194.400 ;
        RECT 438.000 193.000 438.800 193.200 ;
        RECT 429.800 192.400 438.800 193.000 ;
        RECT 441.200 193.000 442.000 193.200 ;
        RECT 449.200 193.000 449.800 193.800 ;
        RECT 455.600 193.200 457.000 193.800 ;
        RECT 458.000 193.200 459.600 194.000 ;
        RECT 441.200 192.400 449.800 193.000 ;
        RECT 450.800 193.000 457.000 193.200 ;
        RECT 450.800 192.600 456.200 193.000 ;
        RECT 450.800 192.400 451.600 192.600 ;
        RECT 374.000 185.600 375.800 186.200 ;
        RECT 378.800 185.600 380.600 186.200 ;
        RECT 375.000 182.200 375.800 185.600 ;
        RECT 379.800 184.400 380.600 185.600 ;
        RECT 379.800 183.600 381.200 184.400 ;
        RECT 379.800 182.200 380.600 183.600 ;
        RECT 382.000 182.800 382.800 186.200 ;
        RECT 383.600 183.400 384.400 186.200 ;
        RECT 385.200 186.000 389.200 186.200 ;
        RECT 385.200 182.800 386.000 186.000 ;
        RECT 382.000 182.200 386.000 182.800 ;
        RECT 388.400 182.200 389.200 186.000 ;
        RECT 390.600 185.600 392.400 186.200 ;
        RECT 390.600 182.200 391.400 185.600 ;
        RECT 398.400 182.200 399.200 187.800 ;
        RECT 404.800 182.200 405.600 187.800 ;
        RECT 407.600 187.600 408.400 190.400 ;
        RECT 411.000 189.000 411.800 190.400 ;
        RECT 414.200 189.000 415.000 190.400 ;
        RECT 417.800 189.000 418.600 190.400 ;
        RECT 409.200 188.200 411.800 189.000 ;
        RECT 412.600 188.200 415.000 189.000 ;
        RECT 416.000 188.200 418.600 189.000 ;
        RECT 419.400 188.200 421.200 189.000 ;
        RECT 411.000 187.600 411.800 188.200 ;
        RECT 414.200 187.600 415.000 188.200 ;
        RECT 417.800 187.600 418.600 188.200 ;
        RECT 420.400 187.600 421.200 188.200 ;
        RECT 407.600 186.800 410.000 187.600 ;
        RECT 411.000 186.800 413.200 187.600 ;
        RECT 414.200 186.800 416.400 187.600 ;
        RECT 417.800 186.800 419.600 187.600 ;
        RECT 409.200 182.200 410.000 186.800 ;
        RECT 412.400 182.200 413.200 186.800 ;
        RECT 415.600 182.200 416.400 186.800 ;
        RECT 418.800 182.200 419.600 186.800 ;
        RECT 428.200 186.800 429.000 191.200 ;
        RECT 429.800 190.600 430.400 192.400 ;
        RECT 429.600 190.000 430.400 190.600 ;
        RECT 436.400 190.000 459.800 190.600 ;
        RECT 429.600 188.000 430.200 190.000 ;
        RECT 436.400 189.400 437.200 190.000 ;
        RECT 454.000 189.600 454.800 190.000 ;
        RECT 457.200 189.600 458.000 190.000 ;
        RECT 459.000 189.800 459.800 190.000 ;
        RECT 430.800 188.600 434.600 189.400 ;
        RECT 429.600 187.400 430.800 188.000 ;
        RECT 428.200 186.000 429.200 186.800 ;
        RECT 428.400 182.200 429.200 186.000 ;
        RECT 430.000 182.200 430.800 187.400 ;
        RECT 433.800 187.400 434.600 188.600 ;
        RECT 433.800 186.800 435.600 187.400 ;
        RECT 434.800 186.200 435.600 186.800 ;
        RECT 439.600 186.400 440.400 189.200 ;
        RECT 442.800 188.600 446.000 189.400 ;
        RECT 449.800 188.600 451.800 189.400 ;
        RECT 460.400 189.000 461.200 194.600 ;
        RECT 462.800 193.600 463.600 194.400 ;
        RECT 462.800 192.400 463.400 193.600 ;
        RECT 464.200 192.400 465.000 199.800 ;
        RECT 462.000 191.800 463.400 192.400 ;
        RECT 464.000 191.800 465.000 192.400 ;
        RECT 462.000 191.600 462.800 191.800 ;
        RECT 442.400 187.800 443.200 188.000 ;
        RECT 442.400 187.200 446.800 187.800 ;
        RECT 446.000 187.000 446.800 187.200 ;
        RECT 447.600 186.800 448.400 188.400 ;
        RECT 434.800 185.400 437.200 186.200 ;
        RECT 439.600 185.600 440.600 186.400 ;
        RECT 443.600 185.600 445.200 186.400 ;
        RECT 446.000 186.200 446.800 186.400 ;
        RECT 449.800 186.200 450.600 188.600 ;
        RECT 452.400 188.200 461.200 189.000 ;
        RECT 464.000 188.400 464.600 191.800 ;
        RECT 470.000 191.200 470.800 199.800 ;
        RECT 473.200 191.200 474.000 199.800 ;
        RECT 476.400 191.200 477.200 199.800 ;
        RECT 479.600 191.200 480.400 199.800 ;
        RECT 468.400 190.400 470.800 191.200 ;
        RECT 471.800 190.400 474.000 191.200 ;
        RECT 475.000 190.400 477.200 191.200 ;
        RECT 478.600 190.400 480.400 191.200 ;
        RECT 482.800 195.000 483.600 199.000 ;
        RECT 482.800 191.600 483.400 195.000 ;
        RECT 487.000 192.800 487.800 199.800 ;
        RECT 487.000 192.200 488.600 192.800 ;
        RECT 482.800 191.000 486.600 191.600 ;
        RECT 465.200 188.800 466.000 190.400 ;
        RECT 455.800 186.800 458.800 187.600 ;
        RECT 455.800 186.200 456.600 186.800 ;
        RECT 446.000 185.600 450.600 186.200 ;
        RECT 436.400 182.200 437.200 185.400 ;
        RECT 454.000 185.400 456.600 186.200 ;
        RECT 438.000 182.200 438.800 185.000 ;
        RECT 439.600 182.200 440.400 185.000 ;
        RECT 441.200 182.200 442.000 185.000 ;
        RECT 442.800 182.200 443.600 185.000 ;
        RECT 446.000 182.200 446.800 185.000 ;
        RECT 449.200 182.200 450.000 185.000 ;
        RECT 450.800 182.200 451.600 185.000 ;
        RECT 452.400 182.200 453.200 185.000 ;
        RECT 454.000 182.200 454.800 185.400 ;
        RECT 460.400 182.200 461.200 188.200 ;
        RECT 462.000 187.600 464.600 188.400 ;
        RECT 466.800 188.200 467.600 188.400 ;
        RECT 466.000 187.600 467.600 188.200 ;
        RECT 468.400 187.600 469.200 190.400 ;
        RECT 471.800 189.000 472.600 190.400 ;
        RECT 475.000 189.000 475.800 190.400 ;
        RECT 478.600 189.000 479.400 190.400 ;
        RECT 470.000 188.200 472.600 189.000 ;
        RECT 473.400 188.200 475.800 189.000 ;
        RECT 476.800 188.200 479.400 189.000 ;
        RECT 480.200 188.200 482.000 189.000 ;
        RECT 482.800 188.800 483.600 190.400 ;
        RECT 484.400 188.800 485.200 190.400 ;
        RECT 486.000 189.000 486.600 191.000 ;
        RECT 488.000 190.400 488.600 192.200 ;
        RECT 487.600 189.600 488.600 190.400 ;
        RECT 489.200 190.300 490.000 191.200 ;
        RECT 492.400 190.300 493.200 199.800 ;
        RECT 497.200 191.200 498.000 199.800 ;
        RECT 500.400 191.200 501.200 199.800 ;
        RECT 503.600 191.200 504.400 199.800 ;
        RECT 506.800 191.200 507.600 199.800 ;
        RECT 510.000 192.400 510.800 199.800 ;
        RECT 513.200 192.800 514.000 199.800 ;
        RECT 510.000 191.800 512.600 192.400 ;
        RECT 513.200 191.800 514.200 192.800 ;
        RECT 497.200 190.400 499.000 191.200 ;
        RECT 500.400 190.400 502.600 191.200 ;
        RECT 503.600 190.400 505.800 191.200 ;
        RECT 506.800 190.400 509.200 191.200 ;
        RECT 489.200 189.700 493.200 190.300 ;
        RECT 489.200 189.600 490.000 189.700 ;
        RECT 471.800 187.600 472.600 188.200 ;
        RECT 475.000 187.600 475.800 188.200 ;
        RECT 478.600 187.600 479.400 188.200 ;
        RECT 481.200 187.600 482.000 188.200 ;
        RECT 486.000 188.200 487.400 189.000 ;
        RECT 488.000 188.400 488.600 189.600 ;
        RECT 486.000 187.800 487.000 188.200 ;
        RECT 462.200 186.200 462.800 187.600 ;
        RECT 466.000 187.200 466.800 187.600 ;
        RECT 468.400 186.800 470.800 187.600 ;
        RECT 471.800 186.800 474.000 187.600 ;
        RECT 475.000 186.800 477.200 187.600 ;
        RECT 478.600 186.800 480.400 187.600 ;
        RECT 463.800 186.200 467.400 186.600 ;
        RECT 462.000 182.200 462.800 186.200 ;
        RECT 463.600 186.000 467.600 186.200 ;
        RECT 463.600 182.200 464.400 186.000 ;
        RECT 466.800 182.200 467.600 186.000 ;
        RECT 470.000 182.200 470.800 186.800 ;
        RECT 473.200 182.200 474.000 186.800 ;
        RECT 476.400 182.200 477.200 186.800 ;
        RECT 479.600 182.200 480.400 186.800 ;
        RECT 482.800 187.200 487.000 187.800 ;
        RECT 488.000 187.600 490.000 188.400 ;
        RECT 482.800 185.000 483.400 187.200 ;
        RECT 488.000 187.000 488.600 187.600 ;
        RECT 487.800 186.600 488.600 187.000 ;
        RECT 487.000 186.000 488.600 186.600 ;
        RECT 482.800 183.000 483.600 185.000 ;
        RECT 487.000 183.000 487.800 186.000 ;
        RECT 492.400 182.200 493.200 189.700 ;
        RECT 498.200 189.000 499.000 190.400 ;
        RECT 501.800 189.000 502.600 190.400 ;
        RECT 505.000 189.000 505.800 190.400 ;
        RECT 495.600 188.200 497.400 189.000 ;
        RECT 498.200 188.200 500.800 189.000 ;
        RECT 501.800 188.200 504.200 189.000 ;
        RECT 505.000 188.200 507.600 189.000 ;
        RECT 495.600 187.600 496.400 188.200 ;
        RECT 498.200 187.600 499.000 188.200 ;
        RECT 501.800 187.600 502.600 188.200 ;
        RECT 505.000 187.600 505.800 188.200 ;
        RECT 508.400 187.600 509.200 190.400 ;
        RECT 497.200 186.800 499.000 187.600 ;
        RECT 500.400 186.800 502.600 187.600 ;
        RECT 503.600 186.800 505.800 187.600 ;
        RECT 506.800 186.800 509.200 187.600 ;
        RECT 512.000 189.800 512.600 191.800 ;
        RECT 512.000 189.000 513.000 189.800 ;
        RECT 512.000 187.400 512.600 189.000 ;
        RECT 513.600 188.400 514.200 191.800 ;
        RECT 516.400 191.200 517.200 199.800 ;
        RECT 520.600 192.400 521.400 199.800 ;
        RECT 525.400 198.400 526.200 199.800 ;
        RECT 525.400 197.600 526.800 198.400 ;
        RECT 525.400 192.600 526.200 197.600 ;
        RECT 520.600 191.800 522.000 192.400 ;
        RECT 524.400 191.800 526.200 192.600 ;
        RECT 527.600 192.400 528.400 199.800 ;
        RECT 529.000 192.400 529.800 192.600 ;
        RECT 527.600 191.800 529.800 192.400 ;
        RECT 532.000 192.400 533.600 199.800 ;
        RECT 535.600 192.400 536.400 192.600 ;
        RECT 537.200 192.400 538.000 199.800 ;
        RECT 532.000 191.800 534.000 192.400 ;
        RECT 535.600 191.800 538.000 192.400 ;
        RECT 516.400 190.800 520.400 191.200 ;
        RECT 516.400 190.600 520.600 190.800 ;
        RECT 519.800 190.000 520.600 190.600 ;
        RECT 521.400 190.400 522.000 191.800 ;
        RECT 518.400 188.400 519.200 189.200 ;
        RECT 513.200 187.600 514.200 188.400 ;
        RECT 518.000 187.600 519.000 188.400 ;
        RECT 510.000 186.800 512.600 187.400 ;
        RECT 494.000 184.800 494.800 186.400 ;
        RECT 497.200 182.200 498.000 186.800 ;
        RECT 500.400 182.200 501.200 186.800 ;
        RECT 503.600 182.200 504.400 186.800 ;
        RECT 506.800 182.200 507.600 186.800 ;
        RECT 510.000 182.200 510.800 186.800 ;
        RECT 513.600 186.200 514.200 187.600 ;
        RECT 520.000 187.000 520.600 190.000 ;
        RECT 521.200 189.600 522.000 190.400 ;
        RECT 518.200 186.400 520.600 187.000 ;
        RECT 513.200 185.600 514.200 186.200 ;
        RECT 513.200 182.200 514.000 185.600 ;
        RECT 516.400 184.800 517.200 186.400 ;
        RECT 518.200 184.200 518.800 186.400 ;
        RECT 521.400 186.200 522.000 189.600 ;
        RECT 524.600 188.400 525.200 191.800 ;
        RECT 529.200 191.200 529.800 191.800 ;
        RECT 526.000 189.600 526.800 191.200 ;
        RECT 529.200 190.600 532.600 191.200 ;
        RECT 531.800 190.400 532.600 190.600 ;
        RECT 533.400 190.400 534.000 191.800 ;
        RECT 538.800 191.400 539.600 199.800 ;
        RECT 543.200 196.400 544.000 199.800 ;
        RECT 542.000 195.800 544.000 196.400 ;
        RECT 547.600 195.800 548.400 199.800 ;
        RECT 551.800 195.800 553.000 199.800 ;
        RECT 542.000 195.000 542.800 195.800 ;
        RECT 547.600 195.200 548.200 195.800 ;
        RECT 545.400 194.600 549.000 195.200 ;
        RECT 551.600 195.000 552.400 195.800 ;
        RECT 545.400 194.400 546.200 194.600 ;
        RECT 548.200 194.400 549.000 194.600 ;
        RECT 542.000 193.000 542.800 193.200 ;
        RECT 546.600 193.000 547.400 193.200 ;
        RECT 542.000 192.400 547.400 193.000 ;
        RECT 548.000 193.000 550.200 193.600 ;
        RECT 548.000 191.800 548.600 193.000 ;
        RECT 549.400 192.800 550.200 193.000 ;
        RECT 551.800 193.200 553.200 194.000 ;
        RECT 551.800 192.200 552.400 193.200 ;
        RECT 543.800 191.400 548.600 191.800 ;
        RECT 538.800 191.200 548.600 191.400 ;
        RECT 550.000 191.600 552.400 192.200 ;
        RECT 538.800 191.000 544.600 191.200 ;
        RECT 538.800 190.800 544.400 191.000 ;
        RECT 529.600 189.800 530.400 190.000 ;
        RECT 533.400 189.800 534.800 190.400 ;
        RECT 545.200 190.200 546.000 190.400 ;
        RECT 529.600 189.200 532.200 189.800 ;
        RECT 531.600 188.600 532.200 189.200 ;
        RECT 533.000 189.600 534.800 189.800 ;
        RECT 541.000 189.600 546.000 190.200 ;
        RECT 533.000 189.200 534.000 189.600 ;
        RECT 541.000 189.400 541.800 189.600 ;
        RECT 524.400 188.300 525.200 188.400 ;
        RECT 527.600 188.300 529.200 188.400 ;
        RECT 524.400 188.200 529.200 188.300 ;
        RECT 524.400 187.700 531.000 188.200 ;
        RECT 531.600 187.800 532.400 188.600 ;
        RECT 524.400 187.600 525.200 187.700 ;
        RECT 527.600 187.600 531.000 187.700 ;
        RECT 518.000 182.200 518.800 184.200 ;
        RECT 521.200 182.200 522.000 186.200 ;
        RECT 522.800 184.800 523.600 186.400 ;
        RECT 524.600 184.200 525.200 187.600 ;
        RECT 530.400 187.200 531.000 187.600 ;
        RECT 529.000 186.800 529.800 187.000 ;
        RECT 524.400 182.200 525.200 184.200 ;
        RECT 527.600 186.200 529.800 186.800 ;
        RECT 530.400 186.600 532.400 187.200 ;
        RECT 530.800 186.400 532.400 186.600 ;
        RECT 527.600 182.200 528.400 186.200 ;
        RECT 533.000 185.800 533.600 189.200 ;
        RECT 542.600 188.400 543.400 188.600 ;
        RECT 550.000 188.400 550.600 191.600 ;
        RECT 556.400 191.200 557.200 199.800 ;
        RECT 560.600 192.400 561.400 199.800 ;
        RECT 562.000 193.600 562.800 194.400 ;
        RECT 562.200 192.400 562.800 193.600 ;
        RECT 565.200 193.600 566.000 194.400 ;
        RECT 565.200 192.400 565.800 193.600 ;
        RECT 566.600 192.400 567.400 199.800 ;
        RECT 560.600 191.800 561.600 192.400 ;
        RECT 562.200 191.800 563.600 192.400 ;
        RECT 553.000 190.600 557.200 191.200 ;
        RECT 553.000 190.400 553.800 190.600 ;
        RECT 554.600 189.800 555.400 190.000 ;
        RECT 551.600 189.200 555.400 189.800 ;
        RECT 551.600 189.000 552.400 189.200 ;
        RECT 534.400 187.600 535.200 188.400 ;
        RECT 536.400 187.600 538.000 188.400 ;
        RECT 539.600 187.800 550.600 188.400 ;
        RECT 539.600 187.600 541.200 187.800 ;
        RECT 534.400 187.200 535.000 187.600 ;
        RECT 534.200 186.400 535.000 187.200 ;
        RECT 535.600 186.800 536.400 187.000 ;
        RECT 535.600 186.200 538.000 186.800 ;
        RECT 532.000 184.400 533.600 185.800 ;
        RECT 530.800 183.600 533.600 184.400 ;
        RECT 532.000 182.200 533.600 183.600 ;
        RECT 537.200 182.200 538.000 186.200 ;
        RECT 538.800 182.200 539.600 187.000 ;
        RECT 543.800 185.600 544.400 187.800 ;
        RECT 549.400 187.600 550.200 187.800 ;
        RECT 556.400 187.200 557.200 190.600 ;
        RECT 561.000 190.400 561.600 191.800 ;
        RECT 562.800 191.600 563.600 191.800 ;
        RECT 564.400 191.800 565.800 192.400 ;
        RECT 566.400 191.800 567.400 192.400 ;
        RECT 575.600 195.000 576.400 199.000 ;
        RECT 564.400 191.600 565.200 191.800 ;
        RECT 559.600 188.800 560.400 190.400 ;
        RECT 561.000 189.600 562.000 190.400 ;
        RECT 562.900 190.300 563.500 191.600 ;
        RECT 566.400 190.300 567.000 191.800 ;
        RECT 575.600 191.600 576.200 195.000 ;
        RECT 579.800 194.400 580.600 199.800 ;
        RECT 578.800 193.600 580.600 194.400 ;
        RECT 579.800 192.800 580.600 193.600 ;
        RECT 579.800 192.200 581.400 192.800 ;
        RECT 575.600 191.000 579.400 191.600 ;
        RECT 562.900 189.700 567.000 190.300 ;
        RECT 561.000 188.400 561.600 189.600 ;
        RECT 566.400 188.400 567.000 189.700 ;
        RECT 567.600 188.800 568.400 190.400 ;
        RECT 575.600 188.800 576.400 190.400 ;
        RECT 577.200 188.800 578.000 190.400 ;
        RECT 578.800 189.000 579.400 191.000 ;
        RECT 558.000 188.200 558.800 188.400 ;
        RECT 558.000 187.600 559.600 188.200 ;
        RECT 561.000 187.600 563.600 188.400 ;
        RECT 564.400 187.600 567.000 188.400 ;
        RECT 569.200 188.200 570.000 188.400 ;
        RECT 568.400 187.600 570.000 188.200 ;
        RECT 578.800 188.200 580.200 189.000 ;
        RECT 580.800 188.400 581.400 192.200 ;
        RECT 587.800 192.400 588.600 199.800 ;
        RECT 589.200 193.600 590.000 194.400 ;
        RECT 589.400 192.400 590.000 193.600 ;
        RECT 592.400 193.600 593.200 194.400 ;
        RECT 592.400 192.400 593.000 193.600 ;
        RECT 593.800 192.400 594.600 199.800 ;
        RECT 587.800 191.800 588.800 192.400 ;
        RECT 589.400 191.800 590.800 192.400 ;
        RECT 582.000 189.600 582.800 191.200 ;
        RECT 588.200 190.400 588.800 191.800 ;
        RECT 590.000 191.600 590.800 191.800 ;
        RECT 591.600 191.800 593.000 192.400 ;
        RECT 593.600 191.800 594.600 192.400 ;
        RECT 591.600 191.600 592.400 191.800 ;
        RECT 586.800 188.800 587.600 190.400 ;
        RECT 588.200 189.600 589.200 190.400 ;
        RECT 590.100 190.300 590.700 191.600 ;
        RECT 593.600 190.300 594.200 191.800 ;
        RECT 598.000 191.200 598.800 199.800 ;
        RECT 602.200 195.800 603.400 199.800 ;
        RECT 606.800 195.800 607.600 199.800 ;
        RECT 611.200 196.400 612.000 199.800 ;
        RECT 611.200 195.800 613.200 196.400 ;
        RECT 602.800 195.000 603.600 195.800 ;
        RECT 607.000 195.200 607.600 195.800 ;
        RECT 606.200 194.600 609.800 195.200 ;
        RECT 612.400 195.000 613.200 195.800 ;
        RECT 606.200 194.400 607.000 194.600 ;
        RECT 609.000 194.400 609.800 194.600 ;
        RECT 602.000 193.200 603.400 194.000 ;
        RECT 602.800 192.200 603.400 193.200 ;
        RECT 605.000 193.000 607.200 193.600 ;
        RECT 605.000 192.800 605.800 193.000 ;
        RECT 602.800 191.600 605.200 192.200 ;
        RECT 598.000 190.600 602.200 191.200 ;
        RECT 590.100 189.700 594.200 190.300 ;
        RECT 588.200 188.400 588.800 189.600 ;
        RECT 593.600 188.400 594.200 189.700 ;
        RECT 594.800 188.800 595.600 190.400 ;
        RECT 578.800 187.800 579.800 188.200 ;
        RECT 558.800 187.200 559.600 187.600 ;
        RECT 553.400 186.600 557.200 187.200 ;
        RECT 553.400 186.400 554.200 186.600 ;
        RECT 542.000 184.200 542.800 185.000 ;
        RECT 543.600 184.800 544.400 185.600 ;
        RECT 545.400 185.400 546.200 185.600 ;
        RECT 545.400 184.800 548.200 185.400 ;
        RECT 547.600 184.200 548.200 184.800 ;
        RECT 551.600 184.200 552.400 185.000 ;
        RECT 542.000 183.600 544.000 184.200 ;
        RECT 543.200 182.200 544.000 183.600 ;
        RECT 547.600 182.200 548.400 184.200 ;
        RECT 551.600 183.600 553.000 184.200 ;
        RECT 551.800 182.200 553.000 183.600 ;
        RECT 556.400 182.200 557.200 186.600 ;
        RECT 558.200 186.200 561.800 186.600 ;
        RECT 562.800 186.200 563.400 187.600 ;
        RECT 564.600 186.200 565.200 187.600 ;
        RECT 568.400 187.200 569.200 187.600 ;
        RECT 575.600 187.200 579.800 187.800 ;
        RECT 580.800 187.600 582.800 188.400 ;
        RECT 585.200 188.200 586.000 188.400 ;
        RECT 585.200 187.600 586.800 188.200 ;
        RECT 588.200 187.600 590.800 188.400 ;
        RECT 591.600 187.600 594.200 188.400 ;
        RECT 596.400 188.200 597.200 188.400 ;
        RECT 595.600 187.600 597.200 188.200 ;
        RECT 566.200 186.200 569.800 186.600 ;
        RECT 558.000 186.000 562.000 186.200 ;
        RECT 558.000 182.200 558.800 186.000 ;
        RECT 561.200 182.200 562.000 186.000 ;
        RECT 562.800 182.200 563.600 186.200 ;
        RECT 564.400 182.200 565.200 186.200 ;
        RECT 566.000 186.000 570.000 186.200 ;
        RECT 566.000 182.200 566.800 186.000 ;
        RECT 569.200 182.200 570.000 186.000 ;
        RECT 575.600 185.000 576.200 187.200 ;
        RECT 580.800 187.000 581.400 187.600 ;
        RECT 586.000 187.200 586.800 187.600 ;
        RECT 580.600 186.600 581.400 187.000 ;
        RECT 579.800 186.000 581.400 186.600 ;
        RECT 585.400 186.200 589.000 186.600 ;
        RECT 590.000 186.200 590.600 187.600 ;
        RECT 591.800 186.200 592.400 187.600 ;
        RECT 595.600 187.200 596.400 187.600 ;
        RECT 598.000 187.200 598.800 190.600 ;
        RECT 601.400 190.400 602.200 190.600 ;
        RECT 599.800 189.800 600.600 190.000 ;
        RECT 599.800 189.200 603.600 189.800 ;
        RECT 602.800 189.000 603.600 189.200 ;
        RECT 604.600 188.400 605.200 191.600 ;
        RECT 606.600 191.800 607.200 193.000 ;
        RECT 607.800 193.000 608.600 193.200 ;
        RECT 612.400 193.000 613.200 193.200 ;
        RECT 607.800 192.400 613.200 193.000 ;
        RECT 606.600 191.400 611.400 191.800 ;
        RECT 615.600 191.400 616.400 199.800 ;
        RECT 619.800 192.400 620.600 199.800 ;
        RECT 621.200 193.600 622.000 194.400 ;
        RECT 621.400 192.400 622.000 193.600 ;
        RECT 626.200 192.400 627.000 199.800 ;
        RECT 627.600 193.600 628.400 194.400 ;
        RECT 627.800 192.400 628.400 193.600 ;
        RECT 633.800 192.800 634.600 199.800 ;
        RECT 638.000 195.000 638.800 199.000 ;
        RECT 619.800 191.800 620.800 192.400 ;
        RECT 621.400 191.800 622.800 192.400 ;
        RECT 626.200 191.800 627.200 192.400 ;
        RECT 627.800 191.800 629.200 192.400 ;
        RECT 606.600 191.200 616.400 191.400 ;
        RECT 610.600 191.000 616.400 191.200 ;
        RECT 610.800 190.800 616.400 191.000 ;
        RECT 620.200 190.400 620.800 191.800 ;
        RECT 622.000 191.600 622.800 191.800 ;
        RECT 609.200 190.200 610.000 190.400 ;
        RECT 609.200 189.600 614.200 190.200 ;
        RECT 613.400 189.400 614.200 189.600 ;
        RECT 618.800 188.800 619.600 190.400 ;
        RECT 620.200 189.600 621.200 190.400 ;
        RECT 611.800 188.400 612.600 188.600 ;
        RECT 620.200 188.400 620.800 189.600 ;
        RECT 625.200 188.800 626.000 190.400 ;
        RECT 626.600 190.300 627.200 191.800 ;
        RECT 628.400 191.600 629.200 191.800 ;
        RECT 633.000 192.200 634.600 192.800 ;
        RECT 630.000 190.300 630.800 190.400 ;
        RECT 626.600 189.700 630.800 190.300 ;
        RECT 626.600 188.400 627.200 189.700 ;
        RECT 630.000 189.600 630.800 189.700 ;
        RECT 631.600 189.600 632.400 191.200 ;
        RECT 633.000 188.400 633.600 192.200 ;
        RECT 638.200 191.600 638.800 195.000 ;
        RECT 635.000 191.000 638.800 191.600 ;
        RECT 639.600 191.200 640.400 199.800 ;
        RECT 643.800 195.800 645.000 199.800 ;
        RECT 648.400 195.800 649.200 199.800 ;
        RECT 652.800 196.400 653.600 199.800 ;
        RECT 652.800 195.800 654.800 196.400 ;
        RECT 644.400 195.000 645.200 195.800 ;
        RECT 648.600 195.200 649.200 195.800 ;
        RECT 647.800 194.600 651.400 195.200 ;
        RECT 654.000 195.000 654.800 195.800 ;
        RECT 647.800 194.400 648.600 194.600 ;
        RECT 650.600 194.400 651.400 194.600 ;
        RECT 643.600 193.200 645.000 194.000 ;
        RECT 644.400 192.200 645.000 193.200 ;
        RECT 646.600 193.000 648.800 193.600 ;
        RECT 646.600 192.800 647.400 193.000 ;
        RECT 644.400 191.600 646.800 192.200 ;
        RECT 635.000 189.000 635.600 191.000 ;
        RECT 639.600 190.600 643.800 191.200 ;
        RECT 604.600 187.800 615.600 188.400 ;
        RECT 605.000 187.600 605.800 187.800 ;
        RECT 607.600 187.600 608.400 187.800 ;
        RECT 598.000 186.600 601.800 187.200 ;
        RECT 593.400 186.200 597.000 186.600 ;
        RECT 585.200 186.000 589.200 186.200 ;
        RECT 575.600 183.000 576.400 185.000 ;
        RECT 579.800 183.000 580.600 186.000 ;
        RECT 585.200 182.200 586.000 186.000 ;
        RECT 588.400 182.200 589.200 186.000 ;
        RECT 590.000 182.200 590.800 186.200 ;
        RECT 591.600 182.200 592.400 186.200 ;
        RECT 593.200 186.000 597.200 186.200 ;
        RECT 593.200 182.200 594.000 186.000 ;
        RECT 596.400 182.200 597.200 186.000 ;
        RECT 598.000 182.200 598.800 186.600 ;
        RECT 601.000 186.400 601.800 186.600 ;
        RECT 610.800 185.600 611.400 187.800 ;
        RECT 614.000 187.600 615.600 187.800 ;
        RECT 617.200 188.200 618.000 188.400 ;
        RECT 617.200 187.600 618.800 188.200 ;
        RECT 620.200 187.600 622.800 188.400 ;
        RECT 623.600 188.200 624.400 188.400 ;
        RECT 623.600 187.600 625.200 188.200 ;
        RECT 626.600 187.600 629.200 188.400 ;
        RECT 630.000 188.300 630.800 188.400 ;
        RECT 631.600 188.300 633.600 188.400 ;
        RECT 630.000 187.700 633.600 188.300 ;
        RECT 634.200 188.200 635.600 189.000 ;
        RECT 636.400 188.800 637.200 190.400 ;
        RECT 638.000 188.800 638.800 190.400 ;
        RECT 630.000 187.600 630.800 187.700 ;
        RECT 631.600 187.600 633.600 187.700 ;
        RECT 618.000 187.200 618.800 187.600 ;
        RECT 609.000 185.400 609.800 185.600 ;
        RECT 602.800 184.200 603.600 185.000 ;
        RECT 607.000 184.800 609.800 185.400 ;
        RECT 610.800 184.800 611.600 185.600 ;
        RECT 607.000 184.200 607.600 184.800 ;
        RECT 612.400 184.200 613.200 185.000 ;
        RECT 602.200 183.600 603.600 184.200 ;
        RECT 602.200 182.200 603.400 183.600 ;
        RECT 606.800 182.200 607.600 184.200 ;
        RECT 611.200 183.600 613.200 184.200 ;
        RECT 611.200 182.200 612.000 183.600 ;
        RECT 615.600 182.200 616.400 187.000 ;
        RECT 617.400 186.200 621.000 186.600 ;
        RECT 622.000 186.200 622.600 187.600 ;
        RECT 624.400 187.200 625.200 187.600 ;
        RECT 623.800 186.200 627.400 186.600 ;
        RECT 628.400 186.200 629.000 187.600 ;
        RECT 633.000 187.000 633.600 187.600 ;
        RECT 634.600 187.800 635.600 188.200 ;
        RECT 634.600 187.200 638.800 187.800 ;
        RECT 633.000 186.600 633.800 187.000 ;
        RECT 617.200 186.000 621.200 186.200 ;
        RECT 617.200 182.200 618.000 186.000 ;
        RECT 620.400 182.200 621.200 186.000 ;
        RECT 622.000 182.200 622.800 186.200 ;
        RECT 623.600 186.000 627.600 186.200 ;
        RECT 623.600 182.200 624.400 186.000 ;
        RECT 626.800 182.200 627.600 186.000 ;
        RECT 628.400 182.200 629.200 186.200 ;
        RECT 633.000 186.000 634.600 186.600 ;
        RECT 633.800 183.000 634.600 186.000 ;
        RECT 638.200 185.000 638.800 187.200 ;
        RECT 638.000 183.000 638.800 185.000 ;
        RECT 639.600 187.200 640.400 190.600 ;
        RECT 643.000 190.400 643.800 190.600 ;
        RECT 641.400 189.800 642.200 190.000 ;
        RECT 641.400 189.200 645.200 189.800 ;
        RECT 644.400 189.000 645.200 189.200 ;
        RECT 646.200 188.400 646.800 191.600 ;
        RECT 648.200 191.800 648.800 193.000 ;
        RECT 649.400 193.000 650.200 193.200 ;
        RECT 654.000 193.000 654.800 193.200 ;
        RECT 649.400 192.400 654.800 193.000 ;
        RECT 648.200 191.400 653.000 191.800 ;
        RECT 657.200 191.400 658.000 199.800 ;
        RECT 661.400 192.600 662.200 199.800 ;
        RECT 660.400 191.800 662.200 192.600 ;
        RECT 648.200 191.200 658.000 191.400 ;
        RECT 652.200 191.000 658.000 191.200 ;
        RECT 652.400 190.800 658.000 191.000 ;
        RECT 650.800 190.200 651.600 190.400 ;
        RECT 650.800 189.600 655.800 190.200 ;
        RECT 655.000 189.400 655.800 189.600 ;
        RECT 653.400 188.400 654.200 188.600 ;
        RECT 660.600 188.400 661.200 191.800 ;
        RECT 662.000 189.600 662.800 191.200 ;
        RECT 646.200 187.800 657.200 188.400 ;
        RECT 646.600 187.600 647.400 187.800 ;
        RECT 652.400 187.600 653.200 187.800 ;
        RECT 655.600 187.600 657.200 187.800 ;
        RECT 660.400 187.600 661.200 188.400 ;
        RECT 639.600 186.600 643.400 187.200 ;
        RECT 639.600 182.200 640.400 186.600 ;
        RECT 642.600 186.400 643.400 186.600 ;
        RECT 652.400 185.600 653.000 187.600 ;
        RECT 650.600 185.400 651.400 185.600 ;
        RECT 644.400 184.200 645.200 185.000 ;
        RECT 648.600 184.800 651.400 185.400 ;
        RECT 652.400 184.800 653.200 185.600 ;
        RECT 648.600 184.200 649.200 184.800 ;
        RECT 654.000 184.200 654.800 185.000 ;
        RECT 643.800 183.600 645.200 184.200 ;
        RECT 643.800 182.200 645.000 183.600 ;
        RECT 648.400 182.200 649.200 184.200 ;
        RECT 652.800 183.600 654.800 184.200 ;
        RECT 652.800 182.200 653.600 183.600 ;
        RECT 657.200 182.200 658.000 187.000 ;
        RECT 660.600 186.400 661.200 187.600 ;
        RECT 658.800 184.800 659.600 186.400 ;
        RECT 660.400 185.600 661.200 186.400 ;
        RECT 662.000 186.300 662.800 186.400 ;
        RECT 663.600 186.300 664.400 186.400 ;
        RECT 662.000 185.700 664.400 186.300 ;
        RECT 662.000 185.600 662.800 185.700 ;
        RECT 660.600 184.200 661.200 185.600 ;
        RECT 663.600 184.800 664.400 185.700 ;
        RECT 665.200 186.300 666.000 199.800 ;
        RECT 667.400 192.600 668.200 199.800 ;
        RECT 672.400 193.600 673.200 194.400 ;
        RECT 667.400 191.800 669.200 192.600 ;
        RECT 672.400 192.400 673.000 193.600 ;
        RECT 673.800 192.400 674.600 199.800 ;
        RECT 671.600 191.800 673.000 192.400 ;
        RECT 673.600 191.800 674.600 192.400 ;
        RECT 678.000 192.400 678.800 199.800 ;
        RECT 679.600 192.400 680.400 192.600 ;
        RECT 682.400 192.400 684.000 199.800 ;
        RECT 678.000 191.800 680.400 192.400 ;
        RECT 682.000 191.800 684.000 192.400 ;
        RECT 686.200 192.400 687.000 192.600 ;
        RECT 687.600 192.400 688.400 199.800 ;
        RECT 686.200 191.800 688.400 192.400 ;
        RECT 666.800 189.600 667.600 191.200 ;
        RECT 668.400 190.300 669.000 191.800 ;
        RECT 671.600 191.600 672.400 191.800 ;
        RECT 671.600 190.300 672.400 190.400 ;
        RECT 668.400 189.700 672.400 190.300 ;
        RECT 668.400 188.400 669.000 189.700 ;
        RECT 671.600 189.600 672.400 189.700 ;
        RECT 673.600 188.400 674.200 191.800 ;
        RECT 682.000 190.400 682.600 191.800 ;
        RECT 686.200 191.200 686.800 191.800 ;
        RECT 683.400 190.600 686.800 191.200 ;
        RECT 683.400 190.400 684.200 190.600 ;
        RECT 674.800 190.300 675.600 190.400 ;
        RECT 676.400 190.300 677.200 190.400 ;
        RECT 674.800 189.700 677.200 190.300 ;
        RECT 674.800 188.800 675.600 189.700 ;
        RECT 676.400 189.600 677.200 189.700 ;
        RECT 681.200 189.800 682.600 190.400 ;
        RECT 685.600 189.800 686.400 190.000 ;
        RECT 681.200 189.600 683.000 189.800 ;
        RECT 682.000 189.200 683.000 189.600 ;
        RECT 668.400 187.600 669.200 188.400 ;
        RECT 671.600 187.600 674.200 188.400 ;
        RECT 676.400 188.200 677.200 188.400 ;
        RECT 675.600 187.600 677.200 188.200 ;
        RECT 678.000 187.600 679.600 188.400 ;
        RECT 680.800 187.600 681.600 188.400 ;
        RECT 666.800 186.300 667.600 186.400 ;
        RECT 665.200 185.700 667.600 186.300 ;
        RECT 660.400 182.200 661.200 184.200 ;
        RECT 665.200 182.200 666.000 185.700 ;
        RECT 666.800 185.600 667.600 185.700 ;
        RECT 668.400 184.200 669.000 187.600 ;
        RECT 670.000 184.800 670.800 186.400 ;
        RECT 671.800 186.200 672.400 187.600 ;
        RECT 675.600 187.200 676.400 187.600 ;
        RECT 681.000 187.200 681.600 187.600 ;
        RECT 679.600 186.800 680.400 187.000 ;
        RECT 673.400 186.200 677.000 186.600 ;
        RECT 678.000 186.200 680.400 186.800 ;
        RECT 681.000 186.400 681.800 187.200 ;
        RECT 668.400 182.200 669.200 184.200 ;
        RECT 671.600 182.200 672.400 186.200 ;
        RECT 673.200 186.000 677.200 186.200 ;
        RECT 673.200 182.200 674.000 186.000 ;
        RECT 676.400 182.200 677.200 186.000 ;
        RECT 678.000 182.200 678.800 186.200 ;
        RECT 682.400 185.800 683.000 189.200 ;
        RECT 683.800 189.200 686.400 189.800 ;
        RECT 683.800 188.600 684.400 189.200 ;
        RECT 683.600 187.800 684.400 188.600 ;
        RECT 686.800 188.200 688.400 188.400 ;
        RECT 685.000 187.600 688.400 188.200 ;
        RECT 685.000 187.200 685.600 187.600 ;
        RECT 683.600 186.600 685.600 187.200 ;
        RECT 686.200 186.800 687.000 187.000 ;
        RECT 683.600 186.400 685.200 186.600 ;
        RECT 686.200 186.200 688.400 186.800 ;
        RECT 682.400 184.400 684.000 185.800 ;
        RECT 681.200 183.600 684.000 184.400 ;
        RECT 682.400 182.200 684.000 183.600 ;
        RECT 687.600 182.200 688.400 186.200 ;
        RECT 1.200 173.800 2.000 179.800 ;
        RECT 7.600 176.600 8.400 179.800 ;
        RECT 9.200 177.000 10.000 179.800 ;
        RECT 10.800 177.000 11.600 179.800 ;
        RECT 12.400 177.000 13.200 179.800 ;
        RECT 15.600 177.000 16.400 179.800 ;
        RECT 18.800 177.000 19.600 179.800 ;
        RECT 20.400 177.000 21.200 179.800 ;
        RECT 22.000 177.000 22.800 179.800 ;
        RECT 23.600 177.000 24.400 179.800 ;
        RECT 5.800 175.800 8.400 176.600 ;
        RECT 25.200 176.600 26.000 179.800 ;
        RECT 11.800 175.800 16.400 176.400 ;
        RECT 5.800 175.200 6.600 175.800 ;
        RECT 3.600 174.400 6.600 175.200 ;
        RECT 1.200 173.000 10.000 173.800 ;
        RECT 11.800 173.400 12.600 175.800 ;
        RECT 15.600 175.600 16.400 175.800 ;
        RECT 17.200 175.600 18.800 176.400 ;
        RECT 21.800 175.600 22.800 176.400 ;
        RECT 25.200 175.800 27.600 176.600 ;
        RECT 14.000 173.600 14.800 175.200 ;
        RECT 15.600 174.800 16.400 175.000 ;
        RECT 15.600 174.200 20.000 174.800 ;
        RECT 19.200 174.000 20.000 174.200 ;
        RECT 1.200 167.400 2.000 173.000 ;
        RECT 10.600 172.600 12.600 173.400 ;
        RECT 16.400 172.600 19.600 173.400 ;
        RECT 22.000 172.800 22.800 175.600 ;
        RECT 26.800 175.200 27.600 175.800 ;
        RECT 26.800 174.600 28.600 175.200 ;
        RECT 27.800 173.400 28.600 174.600 ;
        RECT 31.600 174.600 32.400 179.800 ;
        RECT 33.200 176.000 34.000 179.800 ;
        RECT 33.200 175.200 34.200 176.000 ;
        RECT 31.600 174.000 32.800 174.600 ;
        RECT 27.800 172.600 31.600 173.400 ;
        RECT 2.600 172.000 3.400 172.200 ;
        RECT 7.600 172.000 8.400 172.400 ;
        RECT 14.000 172.000 14.800 172.400 ;
        RECT 25.200 172.000 26.000 172.600 ;
        RECT 32.200 172.000 32.800 174.000 ;
        RECT 2.600 171.400 26.000 172.000 ;
        RECT 32.000 171.400 32.800 172.000 ;
        RECT 32.000 169.600 32.600 171.400 ;
        RECT 33.400 170.800 34.200 175.200 ;
        RECT 36.400 175.000 37.200 179.800 ;
        RECT 40.800 178.400 41.600 179.800 ;
        RECT 39.600 177.800 41.600 178.400 ;
        RECT 45.200 177.800 46.000 179.800 ;
        RECT 49.400 178.400 50.600 179.800 ;
        RECT 49.200 177.800 50.600 178.400 ;
        RECT 39.600 177.000 40.400 177.800 ;
        RECT 45.200 177.200 45.800 177.800 ;
        RECT 41.200 175.600 42.000 177.200 ;
        RECT 43.000 176.600 45.800 177.200 ;
        RECT 49.200 177.000 50.000 177.800 ;
        RECT 43.000 176.400 43.800 176.600 ;
        RECT 37.200 174.200 38.800 174.400 ;
        RECT 41.400 174.200 42.000 175.600 ;
        RECT 51.000 175.400 51.800 175.600 ;
        RECT 54.000 175.400 54.800 179.800 ;
        RECT 56.200 178.400 57.000 179.800 ;
        RECT 56.200 177.600 58.000 178.400 ;
        RECT 56.200 176.400 57.000 177.600 ;
        RECT 56.200 175.800 58.000 176.400 ;
        RECT 60.400 176.000 61.200 179.800 ;
        RECT 63.600 176.000 64.400 179.800 ;
        RECT 60.400 175.800 64.400 176.000 ;
        RECT 65.200 175.800 66.000 179.800 ;
        RECT 66.800 175.800 67.600 179.800 ;
        RECT 68.400 176.000 69.200 179.800 ;
        RECT 71.600 176.000 72.400 179.800 ;
        RECT 68.400 175.800 72.400 176.000 ;
        RECT 51.000 174.800 54.800 175.400 ;
        RECT 47.000 174.200 47.800 174.400 ;
        RECT 37.200 173.600 48.200 174.200 ;
        RECT 40.200 173.400 41.000 173.600 ;
        RECT 38.600 172.400 39.400 172.600 ;
        RECT 41.200 172.400 42.000 172.600 ;
        RECT 38.600 171.800 43.600 172.400 ;
        RECT 42.800 171.600 43.600 171.800 ;
        RECT 10.800 169.400 11.600 169.600 ;
        RECT 6.200 169.000 11.600 169.400 ;
        RECT 5.400 168.800 11.600 169.000 ;
        RECT 12.600 169.000 21.200 169.600 ;
        RECT 2.800 168.000 4.400 168.800 ;
        RECT 5.400 168.200 6.800 168.800 ;
        RECT 12.600 168.200 13.200 169.000 ;
        RECT 20.400 168.800 21.200 169.000 ;
        RECT 23.600 169.000 32.600 169.600 ;
        RECT 23.600 168.800 24.400 169.000 ;
        RECT 3.800 167.600 4.400 168.000 ;
        RECT 7.400 167.600 13.200 168.200 ;
        RECT 13.800 167.600 16.400 168.400 ;
        RECT 1.200 166.800 3.200 167.400 ;
        RECT 3.800 166.800 8.000 167.600 ;
        RECT 2.600 166.200 3.200 166.800 ;
        RECT 2.600 165.600 3.600 166.200 ;
        RECT 2.800 162.200 3.600 165.600 ;
        RECT 6.000 162.200 6.800 166.800 ;
        RECT 9.200 162.200 10.000 165.000 ;
        RECT 10.800 162.200 11.600 165.000 ;
        RECT 12.400 162.200 13.200 167.000 ;
        RECT 15.600 162.200 16.400 167.000 ;
        RECT 18.800 162.200 19.600 168.400 ;
        RECT 26.800 167.600 29.400 168.400 ;
        RECT 22.000 166.800 26.200 167.600 ;
        RECT 20.400 162.200 21.200 165.000 ;
        RECT 22.000 162.200 22.800 165.000 ;
        RECT 23.600 162.200 24.400 165.000 ;
        RECT 26.800 162.200 27.600 167.600 ;
        RECT 32.000 167.400 32.600 169.000 ;
        RECT 30.000 166.800 32.600 167.400 ;
        RECT 33.200 170.000 34.200 170.800 ;
        RECT 36.400 171.000 42.000 171.200 ;
        RECT 36.400 170.800 42.200 171.000 ;
        RECT 36.400 170.600 46.200 170.800 ;
        RECT 30.000 162.200 30.800 166.800 ;
        RECT 33.200 162.200 34.000 170.000 ;
        RECT 36.400 162.200 37.200 170.600 ;
        RECT 41.400 170.200 46.200 170.600 ;
        RECT 39.600 169.000 45.000 169.600 ;
        RECT 39.600 168.800 40.400 169.000 ;
        RECT 44.200 168.800 45.000 169.000 ;
        RECT 45.600 169.000 46.200 170.200 ;
        RECT 47.600 170.400 48.200 173.600 ;
        RECT 49.200 172.800 50.000 173.000 ;
        RECT 49.200 172.200 53.000 172.800 ;
        RECT 52.200 172.000 53.000 172.200 ;
        RECT 50.600 171.400 51.400 171.600 ;
        RECT 54.000 171.400 54.800 174.800 ;
        RECT 50.600 170.800 54.800 171.400 ;
        RECT 47.600 169.800 50.000 170.400 ;
        RECT 47.000 169.000 47.800 169.200 ;
        RECT 45.600 168.400 47.800 169.000 ;
        RECT 49.400 168.800 50.000 169.800 ;
        RECT 49.400 168.000 50.800 168.800 ;
        RECT 43.000 167.400 43.800 167.600 ;
        RECT 45.800 167.400 46.600 167.600 ;
        RECT 39.600 166.200 40.400 167.000 ;
        RECT 43.000 166.800 46.600 167.400 ;
        RECT 45.200 166.200 45.800 166.800 ;
        RECT 49.200 166.200 50.000 167.000 ;
        RECT 39.600 165.600 41.600 166.200 ;
        RECT 40.800 162.200 41.600 165.600 ;
        RECT 45.200 162.200 46.000 166.200 ;
        RECT 49.400 162.200 50.600 166.200 ;
        RECT 54.000 162.200 54.800 170.800 ;
        RECT 55.600 167.600 56.400 170.400 ;
        RECT 57.200 162.200 58.000 175.800 ;
        RECT 60.600 175.400 64.200 175.800 ;
        RECT 58.800 173.600 59.600 175.200 ;
        RECT 61.200 174.400 62.000 174.800 ;
        RECT 65.200 174.400 65.800 175.800 ;
        RECT 67.000 174.400 67.600 175.800 ;
        RECT 68.600 175.400 72.200 175.800 ;
        RECT 70.800 174.400 71.600 174.800 ;
        RECT 60.400 173.800 62.000 174.400 ;
        RECT 60.400 173.600 61.200 173.800 ;
        RECT 63.400 173.600 66.000 174.400 ;
        RECT 66.800 173.600 69.400 174.400 ;
        RECT 70.800 174.300 72.400 174.400 ;
        RECT 73.200 174.300 74.000 179.800 ;
        RECT 74.800 175.600 75.600 177.200 ;
        RECT 70.800 173.800 74.000 174.300 ;
        RECT 71.600 173.700 74.000 173.800 ;
        RECT 71.600 173.600 72.400 173.700 ;
        RECT 62.000 171.600 62.800 173.200 ;
        RECT 63.400 172.300 64.000 173.600 ;
        RECT 63.400 171.700 67.500 172.300 ;
        RECT 63.400 170.200 64.000 171.700 ;
        RECT 66.900 170.400 67.500 171.700 ;
        RECT 65.200 170.200 66.000 170.400 ;
        RECT 63.000 169.600 64.000 170.200 ;
        RECT 64.600 169.600 66.000 170.200 ;
        RECT 66.800 170.200 67.600 170.400 ;
        RECT 68.800 170.200 69.400 173.600 ;
        RECT 70.000 171.600 70.800 173.200 ;
        RECT 66.800 169.600 68.200 170.200 ;
        RECT 68.800 169.600 69.800 170.200 ;
        RECT 63.000 162.200 63.800 169.600 ;
        RECT 64.600 168.400 65.200 169.600 ;
        RECT 64.400 167.600 65.200 168.400 ;
        RECT 67.600 168.400 68.200 169.600 ;
        RECT 67.600 167.600 68.400 168.400 ;
        RECT 69.000 162.200 69.800 169.600 ;
        RECT 73.200 162.200 74.000 173.700 ;
        RECT 76.400 173.800 77.200 179.800 ;
        RECT 82.800 176.600 83.600 179.800 ;
        RECT 84.400 177.000 85.200 179.800 ;
        RECT 86.000 177.000 86.800 179.800 ;
        RECT 87.600 177.000 88.400 179.800 ;
        RECT 90.800 177.000 91.600 179.800 ;
        RECT 94.000 177.000 94.800 179.800 ;
        RECT 95.600 177.000 96.400 179.800 ;
        RECT 97.200 177.000 98.000 179.800 ;
        RECT 98.800 177.000 99.600 179.800 ;
        RECT 81.000 175.800 83.600 176.600 ;
        RECT 100.400 176.600 101.200 179.800 ;
        RECT 87.000 175.800 91.600 176.400 ;
        RECT 81.000 175.200 81.800 175.800 ;
        RECT 78.800 174.400 81.800 175.200 ;
        RECT 76.400 173.000 85.200 173.800 ;
        RECT 87.000 173.400 87.800 175.800 ;
        RECT 90.800 175.600 91.600 175.800 ;
        RECT 92.400 175.600 94.000 176.400 ;
        RECT 97.000 175.600 98.000 176.400 ;
        RECT 100.400 175.800 102.800 176.600 ;
        RECT 89.200 173.600 90.000 175.200 ;
        RECT 90.800 174.800 91.600 175.000 ;
        RECT 90.800 174.200 95.200 174.800 ;
        RECT 94.400 174.000 95.200 174.200 ;
        RECT 76.400 167.400 77.200 173.000 ;
        RECT 85.800 172.600 87.800 173.400 ;
        RECT 91.600 172.600 94.800 173.400 ;
        RECT 97.200 172.800 98.000 175.600 ;
        RECT 102.000 175.200 102.800 175.800 ;
        RECT 102.000 174.600 103.800 175.200 ;
        RECT 103.000 173.400 103.800 174.600 ;
        RECT 106.800 174.600 107.600 179.800 ;
        RECT 108.400 176.000 109.200 179.800 ;
        RECT 108.400 175.200 109.400 176.000 ;
        RECT 106.800 174.000 108.000 174.600 ;
        RECT 103.000 172.600 106.800 173.400 ;
        RECT 77.800 172.000 78.600 172.200 ;
        RECT 79.600 172.000 80.400 172.400 ;
        RECT 82.800 172.000 83.600 172.400 ;
        RECT 100.400 172.000 101.200 172.600 ;
        RECT 107.400 172.000 108.000 174.000 ;
        RECT 77.800 171.400 101.200 172.000 ;
        RECT 107.200 171.400 108.000 172.000 ;
        RECT 107.200 169.600 107.800 171.400 ;
        RECT 108.600 170.800 109.400 175.200 ;
        RECT 86.000 169.400 86.800 169.600 ;
        RECT 81.400 169.000 86.800 169.400 ;
        RECT 80.600 168.800 86.800 169.000 ;
        RECT 87.800 169.000 96.400 169.600 ;
        RECT 78.000 168.000 79.600 168.800 ;
        RECT 80.600 168.200 82.000 168.800 ;
        RECT 87.800 168.200 88.400 169.000 ;
        RECT 95.600 168.800 96.400 169.000 ;
        RECT 98.800 169.000 107.800 169.600 ;
        RECT 98.800 168.800 99.600 169.000 ;
        RECT 79.000 167.600 79.600 168.000 ;
        RECT 82.600 167.600 88.400 168.200 ;
        RECT 89.000 167.600 91.600 168.400 ;
        RECT 76.400 166.800 78.400 167.400 ;
        RECT 79.000 166.800 83.200 167.600 ;
        RECT 77.800 166.200 78.400 166.800 ;
        RECT 77.800 165.600 78.800 166.200 ;
        RECT 78.000 162.200 78.800 165.600 ;
        RECT 81.200 162.200 82.000 166.800 ;
        RECT 84.400 162.200 85.200 165.000 ;
        RECT 86.000 162.200 86.800 165.000 ;
        RECT 87.600 162.200 88.400 167.000 ;
        RECT 90.800 162.200 91.600 167.000 ;
        RECT 94.000 162.200 94.800 168.400 ;
        RECT 102.000 167.600 104.600 168.400 ;
        RECT 97.200 166.800 101.400 167.600 ;
        RECT 95.600 162.200 96.400 165.000 ;
        RECT 97.200 162.200 98.000 165.000 ;
        RECT 98.800 162.200 99.600 165.000 ;
        RECT 102.000 162.200 102.800 167.600 ;
        RECT 107.200 167.400 107.800 169.000 ;
        RECT 105.200 166.800 107.800 167.400 ;
        RECT 108.400 170.000 109.400 170.800 ;
        RECT 105.200 162.200 106.000 166.800 ;
        RECT 108.400 162.200 109.200 170.000 ;
        RECT 111.600 166.300 112.400 166.400 ;
        RECT 116.400 166.300 117.200 179.800 ;
        RECT 118.000 175.600 118.800 177.200 ;
        RECT 120.200 176.400 121.000 179.800 ;
        RECT 120.200 175.800 122.000 176.400 ;
        RECT 118.000 170.300 118.800 170.400 ;
        RECT 119.600 170.300 120.400 170.400 ;
        RECT 118.000 169.700 120.400 170.300 ;
        RECT 118.000 169.600 118.800 169.700 ;
        RECT 119.600 168.800 120.400 169.700 ;
        RECT 111.600 165.700 117.200 166.300 ;
        RECT 111.600 165.600 112.400 165.700 ;
        RECT 116.400 162.200 117.200 165.700 ;
        RECT 121.200 162.200 122.000 175.800 ;
        RECT 124.400 175.200 125.200 179.800 ;
        RECT 127.600 176.400 128.400 179.800 ;
        RECT 127.600 175.800 128.600 176.400 ;
        RECT 130.800 175.800 131.600 179.800 ;
        RECT 132.400 176.000 133.200 179.800 ;
        RECT 135.600 176.000 136.400 179.800 ;
        RECT 132.400 175.800 136.400 176.000 ;
        RECT 137.200 177.000 138.000 179.000 ;
        RECT 122.800 173.600 123.600 175.200 ;
        RECT 124.400 174.600 127.000 175.200 ;
        RECT 124.600 172.400 125.400 173.200 ;
        RECT 124.400 171.600 125.400 172.400 ;
        RECT 126.400 173.000 127.000 174.600 ;
        RECT 128.000 174.400 128.600 175.800 ;
        RECT 131.000 174.400 131.600 175.800 ;
        RECT 132.600 175.400 136.200 175.800 ;
        RECT 137.200 174.800 137.800 177.000 ;
        RECT 141.400 176.400 142.200 179.000 ;
        RECT 140.400 176.000 142.200 176.400 ;
        RECT 148.400 177.800 149.200 179.800 ;
        RECT 140.400 175.600 143.000 176.000 ;
        RECT 141.400 175.400 143.000 175.600 ;
        RECT 142.200 175.000 143.000 175.400 ;
        RECT 134.800 174.400 135.600 174.800 ;
        RECT 127.600 173.600 128.600 174.400 ;
        RECT 130.800 173.600 133.400 174.400 ;
        RECT 134.800 173.800 136.400 174.400 ;
        RECT 137.200 174.200 141.400 174.800 ;
        RECT 135.600 173.600 136.400 173.800 ;
        RECT 140.400 173.800 141.400 174.200 ;
        RECT 142.400 174.400 143.000 175.000 ;
        RECT 148.400 174.400 149.000 177.800 ;
        RECT 150.000 175.600 150.800 177.200 ;
        RECT 151.600 175.800 152.400 179.800 ;
        RECT 153.200 176.000 154.000 179.800 ;
        RECT 156.400 176.000 157.200 179.800 ;
        RECT 153.200 175.800 157.200 176.000 ;
        RECT 158.000 176.000 158.800 179.800 ;
        RECT 161.200 176.000 162.000 179.800 ;
        RECT 158.000 175.800 162.000 176.000 ;
        RECT 162.800 175.800 163.600 179.800 ;
        RECT 151.800 174.400 152.400 175.800 ;
        RECT 153.400 175.400 157.000 175.800 ;
        RECT 158.200 175.400 161.800 175.800 ;
        RECT 155.600 174.400 156.400 174.800 ;
        RECT 158.800 174.400 159.600 174.800 ;
        RECT 162.800 174.400 163.400 175.800 ;
        RECT 126.400 172.200 127.400 173.000 ;
        RECT 126.400 170.200 127.000 172.200 ;
        RECT 128.000 170.200 128.600 173.600 ;
        RECT 124.400 169.600 127.000 170.200 ;
        RECT 124.400 162.200 125.200 169.600 ;
        RECT 127.600 169.200 128.600 170.200 ;
        RECT 130.800 170.200 131.600 170.400 ;
        RECT 132.800 170.200 133.400 173.600 ;
        RECT 134.000 171.600 134.800 173.200 ;
        RECT 137.200 171.600 138.000 173.200 ;
        RECT 138.800 171.600 139.600 173.200 ;
        RECT 140.400 173.000 141.800 173.800 ;
        RECT 142.400 173.600 144.400 174.400 ;
        RECT 148.400 173.600 149.200 174.400 ;
        RECT 151.600 173.600 154.200 174.400 ;
        RECT 155.600 173.800 157.200 174.400 ;
        RECT 156.400 173.600 157.200 173.800 ;
        RECT 158.000 173.800 159.600 174.400 ;
        RECT 158.000 173.600 158.800 173.800 ;
        RECT 161.000 173.600 163.600 174.400 ;
        RECT 140.400 171.000 141.000 173.000 ;
        RECT 137.200 170.400 141.000 171.000 ;
        RECT 130.800 169.600 132.200 170.200 ;
        RECT 132.800 169.600 133.800 170.200 ;
        RECT 127.600 162.200 128.400 169.200 ;
        RECT 131.600 168.400 132.200 169.600 ;
        RECT 131.600 167.600 132.400 168.400 ;
        RECT 133.000 162.200 133.800 169.600 ;
        RECT 137.200 167.000 137.800 170.400 ;
        RECT 142.400 169.800 143.000 173.600 ;
        RECT 143.600 170.800 144.400 172.400 ;
        RECT 146.800 170.800 147.600 172.400 ;
        RECT 148.400 170.400 149.000 173.600 ;
        RECT 148.400 170.200 149.200 170.400 ;
        RECT 141.400 169.200 143.000 169.800 ;
        RECT 147.400 169.400 149.200 170.200 ;
        RECT 151.600 170.200 152.400 170.400 ;
        RECT 153.600 170.200 154.200 173.600 ;
        RECT 154.800 171.600 155.600 173.200 ;
        RECT 156.500 172.400 157.100 173.600 ;
        RECT 156.400 172.300 157.200 172.400 ;
        RECT 159.600 172.300 160.400 173.200 ;
        RECT 156.400 171.700 160.400 172.300 ;
        RECT 156.400 171.600 157.200 171.700 ;
        RECT 159.600 171.600 160.400 171.700 ;
        RECT 161.000 170.200 161.600 173.600 ;
        RECT 162.800 170.300 163.600 170.400 ;
        RECT 164.400 170.300 165.200 179.800 ;
        RECT 166.000 175.600 166.800 177.200 ;
        RECT 167.600 177.000 168.400 179.000 ;
        RECT 167.600 174.800 168.200 177.000 ;
        RECT 171.800 176.000 172.600 179.000 ;
        RECT 177.200 176.000 178.000 179.800 ;
        RECT 180.400 176.000 181.200 179.800 ;
        RECT 171.800 175.400 173.400 176.000 ;
        RECT 177.200 175.800 181.200 176.000 ;
        RECT 182.000 175.800 182.800 179.800 ;
        RECT 183.600 176.000 184.400 179.800 ;
        RECT 186.800 176.000 187.600 179.800 ;
        RECT 183.600 175.800 187.600 176.000 ;
        RECT 188.400 175.800 189.200 179.800 ;
        RECT 190.000 175.800 190.800 179.800 ;
        RECT 191.600 176.000 192.400 179.800 ;
        RECT 194.800 176.000 195.600 179.800 ;
        RECT 191.600 175.800 195.600 176.000 ;
        RECT 177.400 175.400 181.000 175.800 ;
        RECT 172.600 175.000 173.400 175.400 ;
        RECT 167.600 174.200 171.800 174.800 ;
        RECT 170.800 173.800 171.800 174.200 ;
        RECT 172.800 174.400 173.400 175.000 ;
        RECT 178.000 174.400 178.800 174.800 ;
        RECT 182.000 174.400 182.600 175.800 ;
        RECT 183.800 175.400 187.400 175.800 ;
        RECT 184.400 174.400 185.200 174.800 ;
        RECT 188.400 174.400 189.000 175.800 ;
        RECT 190.200 174.400 190.800 175.800 ;
        RECT 191.800 175.400 195.400 175.800 ;
        RECT 194.000 174.400 194.800 174.800 ;
        RECT 172.800 174.300 174.800 174.400 ;
        RECT 167.600 171.600 168.400 173.200 ;
        RECT 169.200 171.600 170.000 173.200 ;
        RECT 170.800 173.000 172.200 173.800 ;
        RECT 172.800 173.700 176.300 174.300 ;
        RECT 172.800 173.600 174.800 173.700 ;
        RECT 170.800 171.000 171.400 173.000 ;
        RECT 162.800 170.200 165.200 170.300 ;
        RECT 151.600 169.600 153.000 170.200 ;
        RECT 153.600 169.600 154.600 170.200 ;
        RECT 137.200 163.000 138.000 167.000 ;
        RECT 141.400 162.200 142.200 169.200 ;
        RECT 147.400 162.200 148.200 169.400 ;
        RECT 152.400 168.400 153.000 169.600 ;
        RECT 153.800 168.400 154.600 169.600 ;
        RECT 160.600 169.600 161.600 170.200 ;
        RECT 162.200 169.700 165.200 170.200 ;
        RECT 162.200 169.600 163.600 169.700 ;
        RECT 152.400 167.600 153.200 168.400 ;
        RECT 153.800 167.600 155.600 168.400 ;
        RECT 153.800 162.200 154.600 167.600 ;
        RECT 160.600 162.200 161.400 169.600 ;
        RECT 162.200 168.400 162.800 169.600 ;
        RECT 162.000 167.600 162.800 168.400 ;
        RECT 164.400 162.200 165.200 169.700 ;
        RECT 167.600 170.400 171.400 171.000 ;
        RECT 167.600 167.000 168.200 170.400 ;
        RECT 172.800 169.800 173.400 173.600 ;
        RECT 174.000 170.800 174.800 172.400 ;
        RECT 175.700 172.300 176.300 173.700 ;
        RECT 177.200 173.800 178.800 174.400 ;
        RECT 177.200 173.600 178.000 173.800 ;
        RECT 180.200 173.600 182.800 174.400 ;
        RECT 183.600 173.800 185.200 174.400 ;
        RECT 183.600 173.600 184.400 173.800 ;
        RECT 186.600 173.600 189.200 174.400 ;
        RECT 190.000 173.600 192.600 174.400 ;
        RECT 194.000 173.800 195.600 174.400 ;
        RECT 194.800 173.600 195.600 173.800 ;
        RECT 178.800 172.300 179.600 173.200 ;
        RECT 175.700 171.700 179.600 172.300 ;
        RECT 178.800 171.600 179.600 171.700 ;
        RECT 180.200 170.400 180.800 173.600 ;
        RECT 185.200 171.600 186.000 173.200 ;
        RECT 171.800 169.200 173.400 169.800 ;
        RECT 178.800 169.600 180.800 170.400 ;
        RECT 182.000 170.200 182.800 170.400 ;
        RECT 186.600 170.200 187.200 173.600 ;
        RECT 192.000 172.300 192.600 173.600 ;
        RECT 188.500 171.700 192.600 172.300 ;
        RECT 188.500 170.400 189.100 171.700 ;
        RECT 188.400 170.200 189.200 170.400 ;
        RECT 181.400 169.600 182.800 170.200 ;
        RECT 186.200 169.600 187.200 170.200 ;
        RECT 187.800 169.600 189.200 170.200 ;
        RECT 190.000 170.200 190.800 170.400 ;
        RECT 192.000 170.200 192.600 171.700 ;
        RECT 193.200 172.300 194.000 173.200 ;
        RECT 194.800 172.300 195.600 172.400 ;
        RECT 193.200 171.700 195.600 172.300 ;
        RECT 193.200 171.600 194.000 171.700 ;
        RECT 194.800 171.600 195.600 171.700 ;
        RECT 190.000 169.600 191.400 170.200 ;
        RECT 192.000 169.600 193.000 170.200 ;
        RECT 167.600 163.000 168.400 167.000 ;
        RECT 171.800 162.200 172.600 169.200 ;
        RECT 179.800 162.200 180.600 169.600 ;
        RECT 181.400 168.400 182.000 169.600 ;
        RECT 181.200 167.600 182.000 168.400 ;
        RECT 186.200 162.200 187.000 169.600 ;
        RECT 187.800 168.400 188.400 169.600 ;
        RECT 187.600 167.600 188.400 168.400 ;
        RECT 190.800 168.400 191.400 169.600 ;
        RECT 190.800 167.600 191.600 168.400 ;
        RECT 192.200 162.200 193.000 169.600 ;
        RECT 196.400 162.200 197.200 179.800 ;
        RECT 198.000 175.600 198.800 177.200 ;
        RECT 199.600 175.800 200.400 179.800 ;
        RECT 201.200 176.000 202.000 179.800 ;
        RECT 204.400 176.000 205.200 179.800 ;
        RECT 207.600 177.800 208.400 179.800 ;
        RECT 201.200 175.800 205.200 176.000 ;
        RECT 199.800 174.400 200.400 175.800 ;
        RECT 201.400 175.400 205.000 175.800 ;
        RECT 206.000 175.600 206.800 177.200 ;
        RECT 207.800 176.300 208.400 177.800 ;
        RECT 211.000 176.400 211.800 177.200 ;
        RECT 210.800 176.300 211.600 176.400 ;
        RECT 207.700 175.700 211.600 176.300 ;
        RECT 212.400 175.800 213.200 179.800 ;
        RECT 203.600 174.400 204.400 174.800 ;
        RECT 207.800 174.400 208.400 175.700 ;
        RECT 210.800 175.600 211.600 175.700 ;
        RECT 199.600 173.600 202.200 174.400 ;
        RECT 203.600 173.800 205.200 174.400 ;
        RECT 204.400 173.600 205.200 173.800 ;
        RECT 207.600 173.600 208.400 174.400 ;
        RECT 198.000 170.300 198.800 170.400 ;
        RECT 199.600 170.300 200.400 170.400 ;
        RECT 198.000 170.200 200.400 170.300 ;
        RECT 201.600 170.200 202.200 173.600 ;
        RECT 202.800 172.300 203.600 173.200 ;
        RECT 206.000 172.300 206.800 172.400 ;
        RECT 202.800 171.700 206.800 172.300 ;
        RECT 202.800 171.600 203.600 171.700 ;
        RECT 206.000 171.600 206.800 171.700 ;
        RECT 207.800 170.200 208.400 173.600 ;
        RECT 209.200 170.800 210.000 172.400 ;
        RECT 210.800 172.200 211.600 172.400 ;
        RECT 212.600 172.200 213.200 175.800 ;
        RECT 214.000 172.800 214.800 174.400 ;
        RECT 215.600 172.200 216.400 172.400 ;
        RECT 210.800 171.600 213.200 172.200 ;
        RECT 214.800 171.600 216.400 172.200 ;
        RECT 211.000 170.200 211.600 171.600 ;
        RECT 214.800 171.200 215.600 171.600 ;
        RECT 198.000 169.700 201.000 170.200 ;
        RECT 198.000 169.600 198.800 169.700 ;
        RECT 199.600 169.600 201.000 169.700 ;
        RECT 201.600 169.600 202.600 170.200 ;
        RECT 200.400 168.400 201.000 169.600 ;
        RECT 201.800 168.400 202.600 169.600 ;
        RECT 207.600 169.400 209.400 170.200 ;
        RECT 200.400 167.600 201.200 168.400 ;
        RECT 201.800 167.600 203.600 168.400 ;
        RECT 201.800 162.200 202.600 167.600 ;
        RECT 208.600 162.200 209.400 169.400 ;
        RECT 210.800 162.200 211.600 170.200 ;
        RECT 212.400 169.600 216.400 170.200 ;
        RECT 212.400 162.200 213.200 169.600 ;
        RECT 215.600 162.200 216.400 169.600 ;
        RECT 217.200 162.200 218.000 179.800 ;
        RECT 218.800 175.600 219.600 177.200 ;
        RECT 222.000 176.000 222.800 179.800 ;
        RECT 221.800 175.200 222.800 176.000 ;
        RECT 221.800 170.800 222.600 175.200 ;
        RECT 223.600 174.600 224.400 179.800 ;
        RECT 230.000 176.600 230.800 179.800 ;
        RECT 231.600 177.000 232.400 179.800 ;
        RECT 233.200 177.000 234.000 179.800 ;
        RECT 234.800 177.000 235.600 179.800 ;
        RECT 236.400 177.000 237.200 179.800 ;
        RECT 239.600 177.000 240.400 179.800 ;
        RECT 242.800 177.000 243.600 179.800 ;
        RECT 244.400 177.000 245.200 179.800 ;
        RECT 246.000 177.000 246.800 179.800 ;
        RECT 228.400 175.800 230.800 176.600 ;
        RECT 247.600 176.600 248.400 179.800 ;
        RECT 228.400 175.200 229.200 175.800 ;
        RECT 223.200 174.000 224.400 174.600 ;
        RECT 227.400 174.600 229.200 175.200 ;
        RECT 233.200 175.600 234.200 176.400 ;
        RECT 237.200 175.600 238.800 176.400 ;
        RECT 239.600 175.800 244.200 176.400 ;
        RECT 247.600 175.800 250.200 176.600 ;
        RECT 239.600 175.600 240.400 175.800 ;
        RECT 223.200 172.000 223.800 174.000 ;
        RECT 227.400 173.400 228.200 174.600 ;
        RECT 224.400 172.600 228.200 173.400 ;
        RECT 233.200 172.800 234.000 175.600 ;
        RECT 239.600 174.800 240.400 175.000 ;
        RECT 236.000 174.200 240.400 174.800 ;
        RECT 236.000 174.000 236.800 174.200 ;
        RECT 241.200 173.600 242.000 175.200 ;
        RECT 243.400 173.400 244.200 175.800 ;
        RECT 249.400 175.200 250.200 175.800 ;
        RECT 249.400 174.400 252.400 175.200 ;
        RECT 254.000 173.800 254.800 179.800 ;
        RECT 236.400 172.600 239.600 173.400 ;
        RECT 243.400 172.600 245.400 173.400 ;
        RECT 246.000 173.000 254.800 173.800 ;
        RECT 230.000 172.000 230.800 172.600 ;
        RECT 247.600 172.000 248.400 172.400 ;
        RECT 250.800 172.000 251.600 172.400 ;
        RECT 252.600 172.000 253.400 172.200 ;
        RECT 223.200 171.400 224.000 172.000 ;
        RECT 230.000 171.400 253.400 172.000 ;
        RECT 221.800 170.000 222.800 170.800 ;
        RECT 220.400 168.300 221.200 168.400 ;
        RECT 222.000 168.300 222.800 170.000 ;
        RECT 220.400 167.700 222.800 168.300 ;
        RECT 220.400 167.600 221.200 167.700 ;
        RECT 222.000 162.200 222.800 167.700 ;
        RECT 223.400 169.600 224.000 171.400 ;
        RECT 223.400 169.000 232.400 169.600 ;
        RECT 223.400 167.400 224.000 169.000 ;
        RECT 231.600 168.800 232.400 169.000 ;
        RECT 234.800 169.000 243.400 169.600 ;
        RECT 234.800 168.800 235.600 169.000 ;
        RECT 226.600 167.600 229.200 168.400 ;
        RECT 223.400 166.800 226.000 167.400 ;
        RECT 225.200 162.200 226.000 166.800 ;
        RECT 228.400 162.200 229.200 167.600 ;
        RECT 229.800 166.800 234.000 167.600 ;
        RECT 231.600 162.200 232.400 165.000 ;
        RECT 233.200 162.200 234.000 165.000 ;
        RECT 234.800 162.200 235.600 165.000 ;
        RECT 236.400 162.200 237.200 168.400 ;
        RECT 239.600 167.600 242.200 168.400 ;
        RECT 242.800 168.200 243.400 169.000 ;
        RECT 244.400 169.400 245.200 169.600 ;
        RECT 244.400 169.000 249.800 169.400 ;
        RECT 244.400 168.800 250.600 169.000 ;
        RECT 249.200 168.200 250.600 168.800 ;
        RECT 242.800 167.600 248.600 168.200 ;
        RECT 251.600 168.000 253.200 168.800 ;
        RECT 251.600 167.600 252.200 168.000 ;
        RECT 239.600 162.200 240.400 167.000 ;
        RECT 242.800 162.200 243.600 167.000 ;
        RECT 248.000 166.800 252.200 167.600 ;
        RECT 254.000 167.400 254.800 173.000 ;
        RECT 257.200 177.800 258.000 179.800 ;
        RECT 257.200 174.400 257.800 177.800 ;
        RECT 258.800 175.600 259.600 177.200 ;
        RECT 260.600 176.400 261.400 177.200 ;
        RECT 260.400 175.600 261.200 176.400 ;
        RECT 262.000 175.800 262.800 179.800 ;
        RECT 257.200 174.300 258.000 174.400 ;
        RECT 260.500 174.300 261.100 175.600 ;
        RECT 257.200 173.700 261.100 174.300 ;
        RECT 257.200 173.600 258.000 173.700 ;
        RECT 255.600 170.800 256.400 172.400 ;
        RECT 257.200 170.200 257.800 173.600 ;
        RECT 260.400 172.200 261.200 172.400 ;
        RECT 262.200 172.200 262.800 175.800 ;
        RECT 263.600 172.800 264.400 174.400 ;
        RECT 271.600 173.800 272.400 179.800 ;
        RECT 278.000 176.600 278.800 179.800 ;
        RECT 279.600 177.000 280.400 179.800 ;
        RECT 281.200 177.000 282.000 179.800 ;
        RECT 282.800 177.000 283.600 179.800 ;
        RECT 286.000 177.000 286.800 179.800 ;
        RECT 289.200 177.000 290.000 179.800 ;
        RECT 290.800 177.000 291.600 179.800 ;
        RECT 292.400 177.000 293.200 179.800 ;
        RECT 294.000 177.000 294.800 179.800 ;
        RECT 276.200 175.800 278.800 176.600 ;
        RECT 295.600 176.600 296.400 179.800 ;
        RECT 282.200 175.800 286.800 176.400 ;
        RECT 276.200 175.200 277.000 175.800 ;
        RECT 274.000 174.400 277.000 175.200 ;
        RECT 271.600 173.000 280.400 173.800 ;
        RECT 282.200 173.400 283.000 175.800 ;
        RECT 286.000 175.600 286.800 175.800 ;
        RECT 287.600 175.600 289.200 176.400 ;
        RECT 292.200 175.600 293.200 176.400 ;
        RECT 295.600 175.800 298.000 176.600 ;
        RECT 284.400 173.600 285.200 175.200 ;
        RECT 286.000 174.800 286.800 175.000 ;
        RECT 286.000 174.200 290.400 174.800 ;
        RECT 289.600 174.000 290.400 174.200 ;
        RECT 265.200 172.200 266.000 172.400 ;
        RECT 260.400 171.600 262.800 172.200 ;
        RECT 264.400 171.600 266.000 172.200 ;
        RECT 260.600 170.200 261.200 171.600 ;
        RECT 264.400 171.200 265.200 171.600 ;
        RECT 252.800 166.800 254.800 167.400 ;
        RECT 256.200 169.400 258.000 170.200 ;
        RECT 244.400 162.200 245.200 165.000 ;
        RECT 246.000 162.200 246.800 165.000 ;
        RECT 249.200 162.200 250.000 166.800 ;
        RECT 252.800 166.200 253.400 166.800 ;
        RECT 252.400 165.600 253.400 166.200 ;
        RECT 252.400 162.200 253.200 165.600 ;
        RECT 256.200 162.200 257.000 169.400 ;
        RECT 260.400 162.200 261.200 170.200 ;
        RECT 262.000 169.600 266.000 170.200 ;
        RECT 262.000 162.200 262.800 169.600 ;
        RECT 265.200 162.200 266.000 169.600 ;
        RECT 271.600 167.400 272.400 173.000 ;
        RECT 281.000 172.600 283.000 173.400 ;
        RECT 286.800 172.600 290.000 173.400 ;
        RECT 292.400 172.800 293.200 175.600 ;
        RECT 297.200 175.200 298.000 175.800 ;
        RECT 297.200 174.600 299.000 175.200 ;
        RECT 298.200 173.400 299.000 174.600 ;
        RECT 302.000 174.600 302.800 179.800 ;
        RECT 303.600 176.000 304.400 179.800 ;
        RECT 303.600 175.200 304.600 176.000 ;
        RECT 302.000 174.000 303.200 174.600 ;
        RECT 298.200 172.600 302.000 173.400 ;
        RECT 273.000 172.000 273.800 172.200 ;
        RECT 274.800 172.000 275.600 172.400 ;
        RECT 278.000 172.000 278.800 172.400 ;
        RECT 295.600 172.000 296.400 172.600 ;
        RECT 302.600 172.000 303.200 174.000 ;
        RECT 273.000 171.400 296.400 172.000 ;
        RECT 302.400 171.400 303.200 172.000 ;
        RECT 302.400 169.600 303.000 171.400 ;
        RECT 303.800 170.800 304.600 175.200 ;
        RECT 306.800 175.200 307.600 179.800 ;
        RECT 310.000 176.400 310.800 179.800 ;
        RECT 313.800 176.400 314.600 179.800 ;
        RECT 310.000 175.800 311.000 176.400 ;
        RECT 313.800 175.800 315.600 176.400 ;
        RECT 318.000 176.000 318.800 179.800 ;
        RECT 321.200 176.000 322.000 179.800 ;
        RECT 318.000 175.800 322.000 176.000 ;
        RECT 322.800 175.800 323.600 179.800 ;
        RECT 306.800 174.600 309.400 175.200 ;
        RECT 307.000 172.400 307.800 173.200 ;
        RECT 305.200 172.300 306.000 172.400 ;
        RECT 306.800 172.300 307.800 172.400 ;
        RECT 305.200 171.700 307.800 172.300 ;
        RECT 305.200 171.600 306.000 171.700 ;
        RECT 306.800 171.600 307.800 171.700 ;
        RECT 308.800 173.000 309.400 174.600 ;
        RECT 310.400 174.400 311.000 175.800 ;
        RECT 310.000 174.300 311.000 174.400 ;
        RECT 313.200 174.300 314.000 174.400 ;
        RECT 310.000 173.700 314.000 174.300 ;
        RECT 310.000 173.600 311.000 173.700 ;
        RECT 313.200 173.600 314.000 173.700 ;
        RECT 308.800 172.200 309.800 173.000 ;
        RECT 281.200 169.400 282.000 169.600 ;
        RECT 276.600 169.000 282.000 169.400 ;
        RECT 275.800 168.800 282.000 169.000 ;
        RECT 283.000 169.000 291.600 169.600 ;
        RECT 273.200 168.000 274.800 168.800 ;
        RECT 275.800 168.200 277.200 168.800 ;
        RECT 283.000 168.200 283.600 169.000 ;
        RECT 290.800 168.800 291.600 169.000 ;
        RECT 294.000 169.000 303.000 169.600 ;
        RECT 294.000 168.800 294.800 169.000 ;
        RECT 274.200 167.600 274.800 168.000 ;
        RECT 277.800 167.600 283.600 168.200 ;
        RECT 284.200 167.600 286.800 168.400 ;
        RECT 271.600 166.800 273.600 167.400 ;
        RECT 274.200 166.800 278.400 167.600 ;
        RECT 273.000 166.200 273.600 166.800 ;
        RECT 273.000 165.600 274.000 166.200 ;
        RECT 273.200 162.200 274.000 165.600 ;
        RECT 276.400 162.200 277.200 166.800 ;
        RECT 279.600 162.200 280.400 165.000 ;
        RECT 281.200 162.200 282.000 165.000 ;
        RECT 282.800 162.200 283.600 167.000 ;
        RECT 286.000 162.200 286.800 167.000 ;
        RECT 289.200 162.200 290.000 168.400 ;
        RECT 297.200 167.600 299.800 168.400 ;
        RECT 292.400 166.800 296.600 167.600 ;
        RECT 290.800 162.200 291.600 165.000 ;
        RECT 292.400 162.200 293.200 165.000 ;
        RECT 294.000 162.200 294.800 165.000 ;
        RECT 297.200 162.200 298.000 167.600 ;
        RECT 302.400 167.400 303.000 169.000 ;
        RECT 300.400 166.800 303.000 167.400 ;
        RECT 303.600 170.000 304.600 170.800 ;
        RECT 308.800 170.200 309.400 172.200 ;
        RECT 310.400 170.200 311.000 173.600 ;
        RECT 300.400 162.200 301.200 166.800 ;
        RECT 303.600 162.200 304.400 170.000 ;
        RECT 306.800 169.600 309.400 170.200 ;
        RECT 306.800 162.200 307.600 169.600 ;
        RECT 310.000 169.200 311.000 170.200 ;
        RECT 310.000 162.200 310.800 169.200 ;
        RECT 313.200 168.800 314.000 170.400 ;
        RECT 314.800 162.200 315.600 175.800 ;
        RECT 318.200 175.400 321.800 175.800 ;
        RECT 316.400 173.600 317.200 175.200 ;
        RECT 318.800 174.400 319.600 174.800 ;
        RECT 322.800 174.400 323.400 175.800 ;
        RECT 318.000 173.800 319.600 174.400 ;
        RECT 318.000 173.600 318.800 173.800 ;
        RECT 321.000 173.600 323.600 174.400 ;
        RECT 324.400 173.800 325.200 179.800 ;
        RECT 330.800 176.600 331.600 179.800 ;
        RECT 332.400 177.000 333.200 179.800 ;
        RECT 334.000 177.000 334.800 179.800 ;
        RECT 335.600 177.000 336.400 179.800 ;
        RECT 338.800 177.000 339.600 179.800 ;
        RECT 342.000 177.000 342.800 179.800 ;
        RECT 343.600 177.000 344.400 179.800 ;
        RECT 345.200 177.000 346.000 179.800 ;
        RECT 346.800 177.000 347.600 179.800 ;
        RECT 329.000 175.800 331.600 176.600 ;
        RECT 348.400 176.600 349.200 179.800 ;
        RECT 335.000 175.800 339.600 176.400 ;
        RECT 329.000 175.200 329.800 175.800 ;
        RECT 326.800 174.400 329.800 175.200 ;
        RECT 319.600 171.600 320.400 173.200 ;
        RECT 321.000 172.400 321.600 173.600 ;
        RECT 324.400 173.000 333.200 173.800 ;
        RECT 335.000 173.400 335.800 175.800 ;
        RECT 338.800 175.600 339.600 175.800 ;
        RECT 340.400 175.600 342.000 176.400 ;
        RECT 345.000 175.600 346.000 176.400 ;
        RECT 348.400 175.800 350.800 176.600 ;
        RECT 337.200 173.600 338.000 175.200 ;
        RECT 338.800 174.800 339.600 175.000 ;
        RECT 338.800 174.200 343.200 174.800 ;
        RECT 342.400 174.000 343.200 174.200 ;
        RECT 321.000 171.600 322.000 172.400 ;
        RECT 321.000 170.200 321.600 171.600 ;
        RECT 322.800 170.200 323.600 170.400 ;
        RECT 320.600 169.600 321.600 170.200 ;
        RECT 322.200 169.600 323.600 170.200 ;
        RECT 320.600 162.200 321.400 169.600 ;
        RECT 322.200 168.400 322.800 169.600 ;
        RECT 322.000 167.600 322.800 168.400 ;
        RECT 324.400 167.400 325.200 173.000 ;
        RECT 333.800 172.600 335.800 173.400 ;
        RECT 339.600 172.600 342.800 173.400 ;
        RECT 345.200 172.800 346.000 175.600 ;
        RECT 350.000 175.200 350.800 175.800 ;
        RECT 350.000 174.600 351.800 175.200 ;
        RECT 351.000 173.400 351.800 174.600 ;
        RECT 354.800 174.600 355.600 179.800 ;
        RECT 356.400 176.000 357.200 179.800 ;
        RECT 361.200 176.000 362.000 179.800 ;
        RECT 356.400 175.200 357.400 176.000 ;
        RECT 354.800 174.000 356.000 174.600 ;
        RECT 351.000 172.600 354.800 173.400 ;
        RECT 325.800 172.000 326.600 172.200 ;
        RECT 329.200 172.000 330.000 172.400 ;
        RECT 330.800 172.000 331.600 172.400 ;
        RECT 348.400 172.000 349.200 172.600 ;
        RECT 355.400 172.000 356.000 174.000 ;
        RECT 325.800 171.400 349.200 172.000 ;
        RECT 355.200 171.400 356.000 172.000 ;
        RECT 355.200 169.600 355.800 171.400 ;
        RECT 356.600 170.800 357.400 175.200 ;
        RECT 334.000 169.400 334.800 169.600 ;
        RECT 329.400 169.000 334.800 169.400 ;
        RECT 328.600 168.800 334.800 169.000 ;
        RECT 335.800 169.000 344.400 169.600 ;
        RECT 326.000 168.000 327.600 168.800 ;
        RECT 328.600 168.200 330.000 168.800 ;
        RECT 335.800 168.200 336.400 169.000 ;
        RECT 343.600 168.800 344.400 169.000 ;
        RECT 346.800 169.000 355.800 169.600 ;
        RECT 346.800 168.800 347.600 169.000 ;
        RECT 327.000 167.600 327.600 168.000 ;
        RECT 330.600 167.600 336.400 168.200 ;
        RECT 337.000 167.600 339.600 168.400 ;
        RECT 324.400 166.800 326.400 167.400 ;
        RECT 327.000 166.800 331.200 167.600 ;
        RECT 325.800 166.200 326.400 166.800 ;
        RECT 325.800 165.600 326.800 166.200 ;
        RECT 326.000 162.200 326.800 165.600 ;
        RECT 329.200 162.200 330.000 166.800 ;
        RECT 332.400 162.200 333.200 165.000 ;
        RECT 334.000 162.200 334.800 165.000 ;
        RECT 335.600 162.200 336.400 167.000 ;
        RECT 338.800 162.200 339.600 167.000 ;
        RECT 342.000 162.200 342.800 168.400 ;
        RECT 350.000 167.600 352.600 168.400 ;
        RECT 345.200 166.800 349.400 167.600 ;
        RECT 343.600 162.200 344.400 165.000 ;
        RECT 345.200 162.200 346.000 165.000 ;
        RECT 346.800 162.200 347.600 165.000 ;
        RECT 350.000 162.200 350.800 167.600 ;
        RECT 355.200 167.400 355.800 169.000 ;
        RECT 353.200 166.800 355.800 167.400 ;
        RECT 356.400 170.000 357.400 170.800 ;
        RECT 361.000 175.200 362.000 176.000 ;
        RECT 361.000 170.800 361.800 175.200 ;
        RECT 362.800 174.600 363.600 179.800 ;
        RECT 369.200 176.600 370.000 179.800 ;
        RECT 370.800 177.000 371.600 179.800 ;
        RECT 372.400 177.000 373.200 179.800 ;
        RECT 374.000 177.000 374.800 179.800 ;
        RECT 375.600 177.000 376.400 179.800 ;
        RECT 378.800 177.000 379.600 179.800 ;
        RECT 382.000 177.000 382.800 179.800 ;
        RECT 383.600 177.000 384.400 179.800 ;
        RECT 385.200 177.000 386.000 179.800 ;
        RECT 367.600 175.800 370.000 176.600 ;
        RECT 386.800 176.600 387.600 179.800 ;
        RECT 367.600 175.200 368.400 175.800 ;
        RECT 362.400 174.000 363.600 174.600 ;
        RECT 366.600 174.600 368.400 175.200 ;
        RECT 372.400 175.600 373.400 176.400 ;
        RECT 376.400 175.600 378.000 176.400 ;
        RECT 378.800 175.800 383.400 176.400 ;
        RECT 386.800 175.800 389.400 176.600 ;
        RECT 378.800 175.600 379.600 175.800 ;
        RECT 362.400 172.000 363.000 174.000 ;
        RECT 366.600 173.400 367.400 174.600 ;
        RECT 363.600 172.600 367.400 173.400 ;
        RECT 372.400 172.800 373.200 175.600 ;
        RECT 378.800 174.800 379.600 175.000 ;
        RECT 375.200 174.200 379.600 174.800 ;
        RECT 375.200 174.000 376.000 174.200 ;
        RECT 380.400 173.600 381.200 175.200 ;
        RECT 382.600 173.400 383.400 175.800 ;
        RECT 388.600 175.200 389.400 175.800 ;
        RECT 388.600 174.400 391.600 175.200 ;
        RECT 393.200 173.800 394.000 179.800 ;
        RECT 394.800 177.000 395.600 179.000 ;
        RECT 394.800 174.800 395.400 177.000 ;
        RECT 399.000 176.000 399.800 179.000 ;
        RECT 399.000 175.400 400.600 176.000 ;
        RECT 399.800 175.000 400.600 175.400 ;
        RECT 394.800 174.200 399.000 174.800 ;
        RECT 375.600 172.600 378.800 173.400 ;
        RECT 382.600 172.600 384.600 173.400 ;
        RECT 385.200 173.000 394.000 173.800 ;
        RECT 398.000 173.800 399.000 174.200 ;
        RECT 400.000 174.400 400.600 175.000 ;
        RECT 404.400 175.200 405.200 179.800 ;
        RECT 407.600 176.400 408.400 179.800 ;
        RECT 407.600 175.800 408.600 176.400 ;
        RECT 417.200 176.000 418.000 179.800 ;
        RECT 404.400 174.600 407.000 175.200 ;
        RECT 369.200 172.000 370.000 172.600 ;
        RECT 380.400 172.000 381.200 172.400 ;
        RECT 386.800 172.000 387.600 172.400 ;
        RECT 391.800 172.000 392.600 172.200 ;
        RECT 362.400 171.400 363.200 172.000 ;
        RECT 369.200 171.400 392.600 172.000 ;
        RECT 361.000 170.000 362.000 170.800 ;
        RECT 353.200 162.200 354.000 166.800 ;
        RECT 356.400 162.200 357.200 170.000 ;
        RECT 361.200 162.200 362.000 170.000 ;
        RECT 362.600 169.600 363.200 171.400 ;
        RECT 362.600 169.000 371.600 169.600 ;
        RECT 362.600 167.400 363.200 169.000 ;
        RECT 370.800 168.800 371.600 169.000 ;
        RECT 374.000 169.000 382.600 169.600 ;
        RECT 374.000 168.800 374.800 169.000 ;
        RECT 365.800 167.600 368.400 168.400 ;
        RECT 362.600 166.800 365.200 167.400 ;
        RECT 364.400 162.200 365.200 166.800 ;
        RECT 367.600 162.200 368.400 167.600 ;
        RECT 369.000 166.800 373.200 167.600 ;
        RECT 370.800 162.200 371.600 165.000 ;
        RECT 372.400 162.200 373.200 165.000 ;
        RECT 374.000 162.200 374.800 165.000 ;
        RECT 375.600 162.200 376.400 168.400 ;
        RECT 378.800 167.600 381.400 168.400 ;
        RECT 382.000 168.200 382.600 169.000 ;
        RECT 383.600 169.400 384.400 169.600 ;
        RECT 383.600 169.000 389.000 169.400 ;
        RECT 383.600 168.800 389.800 169.000 ;
        RECT 388.400 168.200 389.800 168.800 ;
        RECT 382.000 167.600 387.800 168.200 ;
        RECT 390.800 168.000 392.400 168.800 ;
        RECT 390.800 167.600 391.400 168.000 ;
        RECT 378.800 162.200 379.600 167.000 ;
        RECT 382.000 162.200 382.800 167.000 ;
        RECT 387.200 166.800 391.400 167.600 ;
        RECT 393.200 167.400 394.000 173.000 ;
        RECT 394.800 171.600 395.600 173.200 ;
        RECT 396.400 171.600 397.200 173.200 ;
        RECT 398.000 173.000 399.400 173.800 ;
        RECT 400.000 173.600 402.000 174.400 ;
        RECT 398.000 171.000 398.600 173.000 ;
        RECT 392.000 166.800 394.000 167.400 ;
        RECT 394.800 170.400 398.600 171.000 ;
        RECT 394.800 167.000 395.400 170.400 ;
        RECT 400.000 169.800 400.600 173.600 ;
        RECT 406.400 173.000 407.000 174.600 ;
        RECT 408.000 174.400 408.600 175.800 ;
        RECT 407.600 173.600 408.600 174.400 ;
        RECT 401.200 170.800 402.000 172.400 ;
        RECT 406.400 172.200 407.400 173.000 ;
        RECT 406.400 170.200 407.000 172.200 ;
        RECT 408.000 170.200 408.600 173.600 ;
        RECT 399.000 169.200 400.600 169.800 ;
        RECT 404.400 169.600 407.000 170.200 ;
        RECT 383.600 162.200 384.400 165.000 ;
        RECT 385.200 162.200 386.000 165.000 ;
        RECT 388.400 162.200 389.200 166.800 ;
        RECT 392.000 166.200 392.600 166.800 ;
        RECT 391.600 165.600 392.600 166.200 ;
        RECT 391.600 162.200 392.400 165.600 ;
        RECT 394.800 163.000 395.600 167.000 ;
        RECT 399.000 164.400 399.800 169.200 ;
        RECT 398.000 163.600 399.800 164.400 ;
        RECT 399.000 162.200 399.800 163.600 ;
        RECT 404.400 162.200 405.200 169.600 ;
        RECT 407.600 169.200 408.600 170.200 ;
        RECT 417.000 175.200 418.000 176.000 ;
        RECT 417.000 170.800 417.800 175.200 ;
        RECT 418.800 174.600 419.600 179.800 ;
        RECT 425.200 176.600 426.000 179.800 ;
        RECT 426.800 177.000 427.600 179.800 ;
        RECT 428.400 177.000 429.200 179.800 ;
        RECT 430.000 177.000 430.800 179.800 ;
        RECT 431.600 177.000 432.400 179.800 ;
        RECT 434.800 177.000 435.600 179.800 ;
        RECT 438.000 177.000 438.800 179.800 ;
        RECT 439.600 177.000 440.400 179.800 ;
        RECT 441.200 177.000 442.000 179.800 ;
        RECT 423.600 175.800 426.000 176.600 ;
        RECT 442.800 176.600 443.600 179.800 ;
        RECT 423.600 175.200 424.400 175.800 ;
        RECT 418.400 174.000 419.600 174.600 ;
        RECT 422.600 174.600 424.400 175.200 ;
        RECT 428.400 175.600 429.400 176.400 ;
        RECT 432.400 175.600 434.000 176.400 ;
        RECT 434.800 175.800 439.400 176.400 ;
        RECT 442.800 175.800 445.400 176.600 ;
        RECT 434.800 175.600 435.600 175.800 ;
        RECT 418.400 172.000 419.000 174.000 ;
        RECT 422.600 173.400 423.400 174.600 ;
        RECT 419.600 172.600 423.400 173.400 ;
        RECT 428.400 172.800 429.200 175.600 ;
        RECT 434.800 174.800 435.600 175.000 ;
        RECT 431.200 174.200 435.600 174.800 ;
        RECT 431.200 174.000 432.000 174.200 ;
        RECT 436.400 173.600 437.200 175.200 ;
        RECT 438.600 173.400 439.400 175.800 ;
        RECT 444.600 175.200 445.400 175.800 ;
        RECT 444.600 174.400 447.600 175.200 ;
        RECT 449.200 173.800 450.000 179.800 ;
        RECT 453.400 178.400 454.200 179.800 ;
        RECT 452.400 177.600 454.200 178.400 ;
        RECT 453.400 176.400 454.200 177.600 ;
        RECT 452.400 175.800 454.200 176.400 ;
        RECT 431.600 172.600 434.800 173.400 ;
        RECT 438.600 172.600 440.600 173.400 ;
        RECT 441.200 173.000 450.000 173.800 ;
        RECT 450.800 173.600 451.600 175.200 ;
        RECT 425.200 172.000 426.000 172.600 ;
        RECT 442.800 172.000 443.600 172.400 ;
        RECT 447.600 172.200 448.400 172.400 ;
        RECT 447.600 172.000 448.600 172.200 ;
        RECT 418.400 171.400 419.200 172.000 ;
        RECT 425.200 171.400 448.600 172.000 ;
        RECT 417.000 170.000 418.000 170.800 ;
        RECT 407.600 162.200 408.400 169.200 ;
        RECT 417.200 162.200 418.000 170.000 ;
        RECT 418.600 169.600 419.200 171.400 ;
        RECT 418.600 169.000 427.600 169.600 ;
        RECT 418.600 167.400 419.200 169.000 ;
        RECT 426.800 168.800 427.600 169.000 ;
        RECT 430.000 169.000 438.600 169.600 ;
        RECT 430.000 168.800 430.800 169.000 ;
        RECT 421.800 167.600 424.400 168.400 ;
        RECT 418.600 166.800 421.200 167.400 ;
        RECT 420.400 162.200 421.200 166.800 ;
        RECT 423.600 162.200 424.400 167.600 ;
        RECT 425.000 166.800 429.200 167.600 ;
        RECT 426.800 162.200 427.600 165.000 ;
        RECT 428.400 162.200 429.200 165.000 ;
        RECT 430.000 162.200 430.800 165.000 ;
        RECT 431.600 162.200 432.400 168.400 ;
        RECT 434.800 167.600 437.400 168.400 ;
        RECT 438.000 168.200 438.600 169.000 ;
        RECT 439.600 169.400 440.400 169.600 ;
        RECT 439.600 169.000 445.000 169.400 ;
        RECT 439.600 168.800 445.800 169.000 ;
        RECT 444.400 168.200 445.800 168.800 ;
        RECT 438.000 167.600 443.800 168.200 ;
        RECT 446.800 168.000 448.400 168.800 ;
        RECT 446.800 167.600 447.400 168.000 ;
        RECT 434.800 162.200 435.600 167.000 ;
        RECT 438.000 162.200 438.800 167.000 ;
        RECT 443.200 166.800 447.400 167.600 ;
        RECT 449.200 167.400 450.000 173.000 ;
        RECT 448.000 166.800 450.000 167.400 ;
        RECT 439.600 162.200 440.400 165.000 ;
        RECT 441.200 162.200 442.000 165.000 ;
        RECT 444.400 162.200 445.200 166.800 ;
        RECT 448.000 166.200 448.600 166.800 ;
        RECT 447.600 165.600 448.600 166.200 ;
        RECT 447.600 162.200 448.400 165.600 ;
        RECT 452.400 162.200 453.200 175.800 ;
        RECT 455.600 175.600 456.400 177.200 ;
        RECT 454.000 168.800 454.800 170.400 ;
        RECT 457.200 162.200 458.000 179.800 ;
        RECT 459.400 178.400 460.200 179.800 ;
        RECT 458.800 177.600 460.200 178.400 ;
        RECT 459.400 176.400 460.200 177.600 ;
        RECT 463.600 177.000 464.400 179.000 ;
        RECT 459.400 175.800 461.200 176.400 ;
        RECT 458.800 168.800 459.600 170.400 ;
        RECT 460.400 162.200 461.200 175.800 ;
        RECT 462.000 173.600 462.800 175.200 ;
        RECT 463.600 174.800 464.200 177.000 ;
        RECT 467.800 176.000 468.600 179.000 ;
        RECT 473.200 177.000 474.000 179.000 ;
        RECT 467.800 175.400 469.400 176.000 ;
        RECT 468.600 175.000 469.400 175.400 ;
        RECT 463.600 174.200 467.800 174.800 ;
        RECT 466.800 173.800 467.800 174.200 ;
        RECT 468.800 174.400 469.400 175.000 ;
        RECT 473.200 174.800 473.800 177.000 ;
        RECT 477.400 176.000 478.200 179.000 ;
        RECT 477.400 175.400 479.000 176.000 ;
        RECT 478.200 175.000 479.000 175.400 ;
        RECT 463.600 171.600 464.400 173.200 ;
        RECT 465.200 171.600 466.000 173.200 ;
        RECT 466.800 173.000 468.200 173.800 ;
        RECT 468.800 173.600 470.800 174.400 ;
        RECT 473.200 174.200 477.400 174.800 ;
        RECT 476.400 173.800 477.400 174.200 ;
        RECT 478.400 174.400 479.000 175.000 ;
        RECT 466.800 171.000 467.400 173.000 ;
        RECT 463.600 170.400 467.400 171.000 ;
        RECT 463.600 167.000 464.200 170.400 ;
        RECT 468.800 169.800 469.400 173.600 ;
        RECT 470.000 172.300 470.800 172.400 ;
        RECT 471.600 172.300 472.400 172.400 ;
        RECT 470.000 171.700 472.400 172.300 ;
        RECT 470.000 170.800 470.800 171.700 ;
        RECT 471.600 171.600 472.400 171.700 ;
        RECT 473.200 171.600 474.000 173.200 ;
        RECT 474.800 171.600 475.600 173.200 ;
        RECT 476.400 173.000 477.800 173.800 ;
        RECT 478.400 173.600 480.400 174.400 ;
        RECT 476.400 171.000 477.000 173.000 ;
        RECT 467.800 169.200 469.400 169.800 ;
        RECT 473.200 170.400 477.000 171.000 ;
        RECT 463.600 163.000 464.400 167.000 ;
        RECT 467.800 164.400 468.600 169.200 ;
        RECT 466.800 163.600 468.600 164.400 ;
        RECT 467.800 162.200 468.600 163.600 ;
        RECT 473.200 167.000 473.800 170.400 ;
        RECT 478.400 169.800 479.000 173.600 ;
        RECT 479.600 172.300 480.400 172.400 ;
        RECT 482.800 172.300 483.600 179.800 ;
        RECT 484.400 175.600 485.200 177.200 ;
        RECT 486.000 175.800 486.800 179.800 ;
        RECT 487.600 176.000 488.400 179.800 ;
        RECT 490.800 176.000 491.600 179.800 ;
        RECT 487.600 175.800 491.600 176.000 ;
        RECT 486.200 174.400 486.800 175.800 ;
        RECT 487.800 175.400 491.400 175.800 ;
        RECT 490.000 174.400 490.800 174.800 ;
        RECT 486.000 173.600 488.600 174.400 ;
        RECT 490.000 174.300 491.600 174.400 ;
        RECT 492.400 174.300 493.200 179.800 ;
        RECT 494.000 175.600 494.800 177.200 ;
        RECT 495.600 175.600 496.400 177.200 ;
        RECT 490.000 173.800 493.200 174.300 ;
        RECT 490.800 173.700 493.200 173.800 ;
        RECT 490.800 173.600 491.600 173.700 ;
        RECT 479.600 171.700 483.600 172.300 ;
        RECT 479.600 170.800 480.400 171.700 ;
        RECT 477.400 169.200 479.000 169.800 ;
        RECT 473.200 163.000 474.000 167.000 ;
        RECT 477.400 164.400 478.200 169.200 ;
        RECT 476.400 163.600 478.200 164.400 ;
        RECT 477.400 162.200 478.200 163.600 ;
        RECT 482.800 162.200 483.600 171.700 ;
        RECT 484.400 170.300 485.200 170.400 ;
        RECT 486.000 170.300 486.800 170.400 ;
        RECT 484.400 170.200 486.800 170.300 ;
        RECT 488.000 170.200 488.600 173.600 ;
        RECT 489.200 171.600 490.000 173.200 ;
        RECT 484.400 169.700 487.400 170.200 ;
        RECT 484.400 169.600 485.200 169.700 ;
        RECT 486.000 169.600 487.400 169.700 ;
        RECT 488.000 169.600 489.000 170.200 ;
        RECT 486.800 168.400 487.400 169.600 ;
        RECT 486.800 167.600 487.600 168.400 ;
        RECT 488.200 164.400 489.000 169.600 ;
        RECT 488.200 163.600 490.000 164.400 ;
        RECT 488.200 162.200 489.000 163.600 ;
        RECT 492.400 162.200 493.200 173.700 ;
        RECT 497.200 162.200 498.000 179.800 ;
        RECT 500.400 176.400 501.200 179.800 ;
        RECT 500.200 175.800 501.200 176.400 ;
        RECT 500.200 174.400 500.800 175.800 ;
        RECT 503.600 175.200 504.400 179.800 ;
        RECT 501.800 174.600 504.400 175.200 ;
        RECT 500.200 173.600 501.200 174.400 ;
        RECT 500.200 170.200 500.800 173.600 ;
        RECT 501.800 173.000 502.400 174.600 ;
        RECT 505.200 173.800 506.000 179.800 ;
        RECT 511.600 176.600 512.400 179.800 ;
        RECT 513.200 177.000 514.000 179.800 ;
        RECT 514.800 177.000 515.600 179.800 ;
        RECT 516.400 177.000 517.200 179.800 ;
        RECT 519.600 177.000 520.400 179.800 ;
        RECT 522.800 177.000 523.600 179.800 ;
        RECT 524.400 177.000 525.200 179.800 ;
        RECT 526.000 177.000 526.800 179.800 ;
        RECT 527.600 177.000 528.400 179.800 ;
        RECT 509.800 175.800 512.400 176.600 ;
        RECT 529.200 176.600 530.000 179.800 ;
        RECT 515.800 175.800 520.400 176.400 ;
        RECT 509.800 175.200 510.600 175.800 ;
        RECT 507.600 174.400 510.600 175.200 ;
        RECT 501.400 172.200 502.400 173.000 ;
        RECT 501.800 170.200 502.400 172.200 ;
        RECT 503.400 172.400 504.200 173.200 ;
        RECT 505.200 173.000 514.000 173.800 ;
        RECT 515.800 173.400 516.600 175.800 ;
        RECT 519.600 175.600 520.400 175.800 ;
        RECT 521.200 175.600 522.800 176.400 ;
        RECT 525.800 175.600 526.800 176.400 ;
        RECT 529.200 175.800 531.600 176.600 ;
        RECT 518.000 173.600 518.800 175.200 ;
        RECT 519.600 174.800 520.400 175.000 ;
        RECT 519.600 174.200 524.000 174.800 ;
        RECT 523.200 174.000 524.000 174.200 ;
        RECT 503.400 171.600 504.400 172.400 ;
        RECT 500.200 169.200 501.200 170.200 ;
        RECT 501.800 169.600 504.400 170.200 ;
        RECT 500.400 162.200 501.200 169.200 ;
        RECT 503.600 162.200 504.400 169.600 ;
        RECT 505.200 167.400 506.000 173.000 ;
        RECT 514.600 172.600 516.600 173.400 ;
        RECT 520.400 172.600 523.600 173.400 ;
        RECT 526.000 172.800 526.800 175.600 ;
        RECT 530.800 175.200 531.600 175.800 ;
        RECT 530.800 174.600 532.600 175.200 ;
        RECT 531.800 173.400 532.600 174.600 ;
        RECT 535.600 174.600 536.400 179.800 ;
        RECT 537.200 176.000 538.000 179.800 ;
        RECT 542.000 176.400 542.800 179.800 ;
        RECT 537.200 175.200 538.200 176.000 ;
        RECT 535.600 174.000 536.800 174.600 ;
        RECT 531.800 172.600 535.600 173.400 ;
        RECT 506.600 172.000 507.400 172.200 ;
        RECT 508.400 172.000 509.200 172.400 ;
        RECT 511.600 172.000 512.400 172.400 ;
        RECT 529.200 172.000 530.000 172.600 ;
        RECT 536.200 172.000 536.800 174.000 ;
        RECT 506.600 171.400 530.000 172.000 ;
        RECT 536.000 171.400 536.800 172.000 ;
        RECT 536.000 169.600 536.600 171.400 ;
        RECT 537.400 170.800 538.200 175.200 ;
        RECT 514.800 169.400 515.600 169.600 ;
        RECT 510.200 169.000 515.600 169.400 ;
        RECT 509.400 168.800 515.600 169.000 ;
        RECT 516.600 169.000 525.200 169.600 ;
        RECT 506.800 168.000 508.400 168.800 ;
        RECT 509.400 168.200 510.800 168.800 ;
        RECT 516.600 168.200 517.200 169.000 ;
        RECT 524.400 168.800 525.200 169.000 ;
        RECT 527.600 169.000 536.600 169.600 ;
        RECT 527.600 168.800 528.400 169.000 ;
        RECT 507.800 167.600 508.400 168.000 ;
        RECT 511.400 167.600 517.200 168.200 ;
        RECT 517.800 167.600 520.400 168.400 ;
        RECT 505.200 166.800 507.200 167.400 ;
        RECT 507.800 166.800 512.000 167.600 ;
        RECT 506.600 166.200 507.200 166.800 ;
        RECT 506.600 165.600 507.600 166.200 ;
        RECT 506.800 162.200 507.600 165.600 ;
        RECT 510.000 162.200 510.800 166.800 ;
        RECT 513.200 162.200 514.000 165.000 ;
        RECT 514.800 162.200 515.600 165.000 ;
        RECT 516.400 162.200 517.200 167.000 ;
        RECT 519.600 162.200 520.400 167.000 ;
        RECT 522.800 162.200 523.600 168.400 ;
        RECT 530.800 167.600 533.400 168.400 ;
        RECT 526.000 166.800 530.200 167.600 ;
        RECT 524.400 162.200 525.200 165.000 ;
        RECT 526.000 162.200 526.800 165.000 ;
        RECT 527.600 162.200 528.400 165.000 ;
        RECT 530.800 162.200 531.600 167.600 ;
        RECT 536.000 167.400 536.600 169.000 ;
        RECT 534.000 166.800 536.600 167.400 ;
        RECT 537.200 170.000 538.200 170.800 ;
        RECT 541.800 175.600 542.800 176.400 ;
        RECT 541.800 174.400 542.400 175.600 ;
        RECT 545.200 175.200 546.000 179.800 ;
        RECT 543.400 174.600 546.000 175.200 ;
        RECT 546.800 175.200 547.600 179.800 ;
        RECT 550.000 176.400 550.800 179.800 ;
        RECT 550.000 175.800 551.000 176.400 ;
        RECT 546.800 174.600 549.400 175.200 ;
        RECT 541.800 173.600 542.800 174.400 ;
        RECT 541.800 170.200 542.400 173.600 ;
        RECT 543.400 173.000 544.000 174.600 ;
        RECT 543.000 172.200 544.000 173.000 ;
        RECT 543.400 170.200 544.000 172.200 ;
        RECT 545.000 172.400 545.800 173.200 ;
        RECT 547.000 172.400 547.800 173.200 ;
        RECT 545.000 171.600 546.000 172.400 ;
        RECT 546.800 171.600 547.800 172.400 ;
        RECT 548.800 173.000 549.400 174.600 ;
        RECT 550.400 174.400 551.000 175.800 ;
        RECT 550.000 173.600 551.000 174.400 ;
        RECT 548.800 172.200 549.800 173.000 ;
        RECT 548.800 170.200 549.400 172.200 ;
        RECT 550.400 170.200 551.000 173.600 ;
        RECT 534.000 162.200 534.800 166.800 ;
        RECT 537.200 162.200 538.000 170.000 ;
        RECT 541.800 169.200 542.800 170.200 ;
        RECT 543.400 169.600 546.000 170.200 ;
        RECT 542.000 162.200 542.800 169.200 ;
        RECT 545.200 162.200 546.000 169.600 ;
        RECT 546.800 169.600 549.400 170.200 ;
        RECT 546.800 162.200 547.600 169.600 ;
        RECT 550.000 169.200 551.000 170.200 ;
        RECT 550.000 162.200 550.800 169.200 ;
        RECT 553.200 162.200 554.000 179.800 ;
        RECT 554.800 175.600 555.600 177.200 ;
        RECT 556.400 175.800 557.200 179.800 ;
        RECT 558.000 176.000 558.800 179.800 ;
        RECT 561.200 176.000 562.000 179.800 ;
        RECT 565.400 176.400 566.200 179.800 ;
        RECT 558.000 175.800 562.000 176.000 ;
        RECT 564.400 175.800 566.200 176.400 ;
        RECT 576.200 178.400 577.000 179.000 ;
        RECT 576.200 177.600 578.000 178.400 ;
        RECT 576.200 176.000 577.000 177.600 ;
        RECT 580.400 177.000 581.200 179.000 ;
        RECT 556.600 174.400 557.200 175.800 ;
        RECT 558.200 175.400 561.800 175.800 ;
        RECT 560.400 174.400 561.200 174.800 ;
        RECT 554.800 174.300 555.600 174.400 ;
        RECT 556.400 174.300 559.000 174.400 ;
        RECT 554.800 173.700 559.000 174.300 ;
        RECT 560.400 173.800 562.000 174.400 ;
        RECT 554.800 173.600 555.600 173.700 ;
        RECT 556.400 173.600 559.000 173.700 ;
        RECT 561.200 173.600 562.000 173.800 ;
        RECT 562.800 173.600 563.600 175.200 ;
        RECT 556.400 170.200 557.200 170.400 ;
        RECT 558.400 170.200 559.000 173.600 ;
        RECT 559.600 171.600 560.400 173.200 ;
        RECT 556.400 169.600 557.800 170.200 ;
        RECT 558.400 169.600 559.400 170.200 ;
        RECT 557.200 168.400 557.800 169.600 ;
        RECT 557.200 167.600 558.000 168.400 ;
        RECT 558.600 162.200 559.400 169.600 ;
        RECT 564.400 162.200 565.200 175.800 ;
        RECT 575.400 175.400 577.000 176.000 ;
        RECT 575.400 175.000 576.200 175.400 ;
        RECT 575.400 174.400 576.000 175.000 ;
        RECT 580.600 174.800 581.200 177.000 ;
        RECT 582.000 175.800 582.800 179.800 ;
        RECT 583.600 176.000 584.400 179.800 ;
        RECT 586.800 176.000 587.600 179.800 ;
        RECT 583.600 175.800 587.600 176.000 ;
        RECT 574.000 173.600 576.000 174.400 ;
        RECT 577.000 174.200 581.200 174.800 ;
        RECT 582.200 174.400 582.800 175.800 ;
        RECT 583.800 175.400 587.400 175.800 ;
        RECT 586.000 174.400 586.800 174.800 ;
        RECT 577.000 173.800 578.000 174.200 ;
        RECT 566.000 172.300 566.800 172.400 ;
        RECT 570.800 172.300 571.600 172.400 ;
        RECT 566.000 171.700 571.600 172.300 ;
        RECT 566.000 171.600 566.800 171.700 ;
        RECT 570.800 171.600 571.600 171.700 ;
        RECT 574.000 170.800 574.800 172.400 ;
        RECT 566.000 168.800 566.800 170.400 ;
        RECT 575.400 169.800 576.000 173.600 ;
        RECT 576.600 173.000 578.000 173.800 ;
        RECT 582.000 173.600 584.600 174.400 ;
        RECT 586.000 174.300 587.600 174.400 ;
        RECT 588.400 174.300 589.200 179.800 ;
        RECT 590.000 176.300 590.800 177.200 ;
        RECT 591.600 176.300 592.400 179.800 ;
        RECT 595.800 178.400 597.000 179.800 ;
        RECT 595.800 177.800 597.200 178.400 ;
        RECT 600.400 177.800 601.200 179.800 ;
        RECT 604.800 178.400 605.600 179.800 ;
        RECT 604.800 177.800 606.800 178.400 ;
        RECT 596.400 177.000 597.200 177.800 ;
        RECT 600.600 177.200 601.200 177.800 ;
        RECT 600.600 176.600 603.400 177.200 ;
        RECT 602.600 176.400 603.400 176.600 ;
        RECT 604.400 176.400 605.200 177.200 ;
        RECT 606.000 177.000 606.800 177.800 ;
        RECT 590.000 175.700 592.400 176.300 ;
        RECT 590.000 175.600 590.800 175.700 ;
        RECT 586.000 173.800 589.200 174.300 ;
        RECT 586.800 173.700 589.200 173.800 ;
        RECT 586.800 173.600 587.600 173.700 ;
        RECT 577.400 171.000 578.000 173.000 ;
        RECT 578.800 171.600 579.600 173.200 ;
        RECT 580.400 171.600 581.200 173.200 ;
        RECT 582.000 172.300 582.800 172.400 ;
        RECT 584.000 172.300 584.600 173.600 ;
        RECT 582.000 171.700 584.600 172.300 ;
        RECT 582.000 171.600 582.800 171.700 ;
        RECT 577.400 170.400 581.200 171.000 ;
        RECT 575.400 169.200 577.000 169.800 ;
        RECT 576.200 162.200 577.000 169.200 ;
        RECT 580.600 167.000 581.200 170.400 ;
        RECT 582.000 170.200 582.800 170.400 ;
        RECT 584.000 170.200 584.600 171.700 ;
        RECT 585.200 171.600 586.000 173.200 ;
        RECT 582.000 169.600 583.400 170.200 ;
        RECT 584.000 169.600 585.000 170.200 ;
        RECT 582.800 168.400 583.400 169.600 ;
        RECT 582.800 167.600 583.600 168.400 ;
        RECT 580.400 163.000 581.200 167.000 ;
        RECT 584.200 162.200 585.000 169.600 ;
        RECT 588.400 162.200 589.200 173.700 ;
        RECT 591.600 175.400 592.400 175.700 ;
        RECT 594.600 175.400 595.400 175.600 ;
        RECT 591.600 174.800 595.400 175.400 ;
        RECT 591.600 171.400 592.400 174.800 ;
        RECT 598.600 174.200 599.400 174.400 ;
        RECT 604.400 174.200 605.000 176.400 ;
        RECT 609.200 175.000 610.000 179.800 ;
        RECT 607.600 174.200 609.200 174.400 ;
        RECT 598.200 173.600 609.200 174.200 ;
        RECT 596.400 172.800 597.200 173.000 ;
        RECT 593.400 172.200 597.200 172.800 ;
        RECT 593.400 172.000 594.200 172.200 ;
        RECT 595.000 171.400 595.800 171.600 ;
        RECT 591.600 170.800 595.800 171.400 ;
        RECT 591.600 162.200 592.400 170.800 ;
        RECT 598.200 170.400 598.800 173.600 ;
        RECT 605.400 173.400 606.200 173.600 ;
        RECT 604.400 172.400 605.200 172.600 ;
        RECT 607.000 172.400 607.800 172.600 ;
        RECT 602.800 171.800 607.800 172.400 ;
        RECT 602.800 171.600 603.600 171.800 ;
        RECT 604.400 171.000 610.000 171.200 ;
        RECT 604.200 170.800 610.000 171.000 ;
        RECT 596.400 169.800 598.800 170.400 ;
        RECT 600.200 170.600 610.000 170.800 ;
        RECT 600.200 170.200 605.000 170.600 ;
        RECT 596.400 168.800 597.000 169.800 ;
        RECT 595.600 168.000 597.000 168.800 ;
        RECT 598.600 169.000 599.400 169.200 ;
        RECT 600.200 169.000 600.800 170.200 ;
        RECT 598.600 168.400 600.800 169.000 ;
        RECT 601.400 169.000 606.800 169.600 ;
        RECT 601.400 168.800 602.200 169.000 ;
        RECT 606.000 168.800 606.800 169.000 ;
        RECT 599.800 167.400 600.600 167.600 ;
        RECT 602.600 167.400 603.400 167.600 ;
        RECT 596.400 166.200 597.200 167.000 ;
        RECT 599.800 166.800 603.400 167.400 ;
        RECT 600.600 166.200 601.200 166.800 ;
        RECT 606.000 166.200 606.800 167.000 ;
        RECT 595.800 162.200 597.000 166.200 ;
        RECT 600.400 162.200 601.200 166.200 ;
        RECT 604.800 165.600 606.800 166.200 ;
        RECT 604.800 162.200 605.600 165.600 ;
        RECT 609.200 162.200 610.000 170.600 ;
        RECT 610.800 162.200 611.600 179.800 ;
        RECT 612.400 175.600 613.200 177.200 ;
        RECT 614.000 176.000 614.800 179.800 ;
        RECT 617.200 176.000 618.000 179.800 ;
        RECT 614.000 175.800 618.000 176.000 ;
        RECT 618.800 175.800 619.600 179.800 ;
        RECT 620.400 175.800 621.200 179.800 ;
        RECT 622.000 176.000 622.800 179.800 ;
        RECT 625.200 176.000 626.000 179.800 ;
        RECT 622.000 175.800 626.000 176.000 ;
        RECT 626.800 177.000 627.600 179.000 ;
        RECT 614.200 175.400 617.800 175.800 ;
        RECT 614.800 174.400 615.600 174.800 ;
        RECT 618.800 174.400 619.400 175.800 ;
        RECT 620.600 174.400 621.200 175.800 ;
        RECT 622.200 175.400 625.800 175.800 ;
        RECT 626.800 174.800 627.400 177.000 ;
        RECT 631.000 176.400 631.800 179.000 ;
        RECT 637.000 178.400 637.800 179.800 ;
        RECT 636.400 177.600 637.800 178.400 ;
        RECT 642.800 177.800 643.600 179.800 ;
        RECT 630.000 176.000 631.800 176.400 ;
        RECT 637.000 176.400 637.800 177.600 ;
        RECT 630.000 175.600 632.600 176.000 ;
        RECT 637.000 175.800 638.800 176.400 ;
        RECT 631.000 175.400 632.600 175.600 ;
        RECT 631.800 175.000 632.600 175.400 ;
        RECT 624.400 174.400 625.200 174.800 ;
        RECT 614.000 173.800 615.600 174.400 ;
        RECT 614.000 173.600 614.800 173.800 ;
        RECT 617.000 173.600 619.600 174.400 ;
        RECT 620.400 173.600 623.000 174.400 ;
        RECT 624.400 173.800 626.000 174.400 ;
        RECT 626.800 174.200 631.000 174.800 ;
        RECT 625.200 173.600 626.000 173.800 ;
        RECT 630.000 173.800 631.000 174.200 ;
        RECT 632.000 174.400 632.600 175.000 ;
        RECT 615.600 171.600 616.400 173.200 ;
        RECT 617.000 172.300 617.600 173.600 ;
        RECT 617.000 171.700 621.100 172.300 ;
        RECT 617.000 170.200 617.600 171.700 ;
        RECT 620.500 170.400 621.100 171.700 ;
        RECT 618.800 170.200 619.600 170.400 ;
        RECT 616.600 169.600 617.600 170.200 ;
        RECT 618.200 169.600 619.600 170.200 ;
        RECT 620.400 170.200 621.200 170.400 ;
        RECT 622.400 170.200 623.000 173.600 ;
        RECT 623.600 171.600 624.400 173.200 ;
        RECT 626.800 171.600 627.600 173.200 ;
        RECT 628.400 171.600 629.200 173.200 ;
        RECT 630.000 173.000 631.400 173.800 ;
        RECT 632.000 173.600 634.000 174.400 ;
        RECT 630.000 171.000 630.600 173.000 ;
        RECT 626.800 170.400 630.600 171.000 ;
        RECT 620.400 169.600 621.800 170.200 ;
        RECT 622.400 169.600 623.400 170.200 ;
        RECT 616.600 162.200 617.400 169.600 ;
        RECT 618.200 168.400 618.800 169.600 ;
        RECT 618.000 167.600 618.800 168.400 ;
        RECT 621.200 168.400 621.800 169.600 ;
        RECT 622.600 168.400 623.400 169.600 ;
        RECT 621.200 167.600 622.000 168.400 ;
        RECT 622.600 167.600 624.400 168.400 ;
        RECT 622.600 162.200 623.400 167.600 ;
        RECT 626.800 167.000 627.400 170.400 ;
        RECT 632.000 169.800 632.600 173.600 ;
        RECT 633.200 170.800 634.000 172.400 ;
        RECT 631.000 169.200 632.600 169.800 ;
        RECT 626.800 163.000 627.600 167.000 ;
        RECT 631.000 162.200 631.800 169.200 ;
        RECT 636.400 168.800 637.200 170.400 ;
        RECT 638.000 168.300 638.800 175.800 ;
        RECT 641.200 175.600 642.000 177.200 ;
        RECT 639.600 174.300 640.400 175.200 ;
        RECT 641.300 174.300 641.900 175.600 ;
        RECT 643.000 174.400 643.600 177.800 ;
        RECT 639.600 173.700 641.900 174.300 ;
        RECT 639.600 173.600 640.400 173.700 ;
        RECT 642.800 173.600 643.600 174.400 ;
        RECT 639.600 172.300 640.400 172.400 ;
        RECT 643.000 172.300 643.600 173.600 ;
        RECT 647.600 177.800 648.400 179.800 ;
        RECT 647.600 174.400 648.200 177.800 ;
        RECT 649.200 176.300 650.000 177.200 ;
        RECT 650.800 176.300 651.600 179.800 ;
        RECT 649.200 175.700 651.600 176.300 ;
        RECT 649.200 175.600 650.000 175.700 ;
        RECT 647.600 173.600 648.400 174.400 ;
        RECT 639.600 171.700 643.600 172.300 ;
        RECT 639.600 171.600 640.400 171.700 ;
        RECT 643.000 170.200 643.600 171.700 ;
        RECT 644.400 172.300 645.200 172.400 ;
        RECT 646.000 172.300 646.800 172.400 ;
        RECT 644.400 171.700 646.800 172.300 ;
        RECT 644.400 170.800 645.200 171.700 ;
        RECT 646.000 170.800 646.800 171.700 ;
        RECT 647.600 170.200 648.200 173.600 ;
        RECT 642.800 169.400 644.600 170.200 ;
        RECT 639.600 168.300 640.400 168.400 ;
        RECT 638.000 167.700 640.400 168.300 ;
        RECT 638.000 162.200 638.800 167.700 ;
        RECT 639.600 167.600 640.400 167.700 ;
        RECT 643.800 164.400 644.600 169.400 ;
        RECT 646.600 169.400 648.400 170.200 ;
        RECT 646.600 164.400 647.400 169.400 ;
        RECT 643.800 163.600 645.200 164.400 ;
        RECT 646.000 163.600 647.400 164.400 ;
        RECT 643.800 162.200 644.600 163.600 ;
        RECT 646.600 162.200 647.400 163.600 ;
        RECT 650.800 162.200 651.600 175.700 ;
        RECT 652.400 176.300 653.200 177.200 ;
        RECT 655.600 176.300 656.400 179.800 ;
        RECT 652.400 175.700 656.400 176.300 ;
        RECT 652.400 175.600 653.200 175.700 ;
        RECT 655.400 175.200 656.400 175.700 ;
        RECT 655.400 170.800 656.200 175.200 ;
        RECT 657.200 174.600 658.000 179.800 ;
        RECT 663.600 176.600 664.400 179.800 ;
        RECT 665.200 177.000 666.000 179.800 ;
        RECT 666.800 177.000 667.600 179.800 ;
        RECT 668.400 177.000 669.200 179.800 ;
        RECT 670.000 177.000 670.800 179.800 ;
        RECT 673.200 177.000 674.000 179.800 ;
        RECT 676.400 177.000 677.200 179.800 ;
        RECT 678.000 177.000 678.800 179.800 ;
        RECT 679.600 177.000 680.400 179.800 ;
        RECT 662.000 175.800 664.400 176.600 ;
        RECT 681.200 176.600 682.000 179.800 ;
        RECT 662.000 175.200 662.800 175.800 ;
        RECT 656.800 174.000 658.000 174.600 ;
        RECT 661.000 174.600 662.800 175.200 ;
        RECT 666.800 175.600 667.800 176.400 ;
        RECT 670.800 175.600 672.400 176.400 ;
        RECT 673.200 175.800 677.800 176.400 ;
        RECT 681.200 175.800 683.800 176.600 ;
        RECT 673.200 175.600 674.000 175.800 ;
        RECT 656.800 172.000 657.400 174.000 ;
        RECT 661.000 173.400 661.800 174.600 ;
        RECT 658.000 172.600 661.800 173.400 ;
        RECT 666.800 172.800 667.600 175.600 ;
        RECT 673.200 174.800 674.000 175.000 ;
        RECT 669.600 174.200 674.000 174.800 ;
        RECT 669.600 174.000 670.400 174.200 ;
        RECT 674.800 173.600 675.600 175.200 ;
        RECT 677.000 173.400 677.800 175.800 ;
        RECT 683.000 175.200 683.800 175.800 ;
        RECT 683.000 174.400 686.000 175.200 ;
        RECT 687.600 173.800 688.400 179.800 ;
        RECT 670.000 172.600 673.200 173.400 ;
        RECT 677.000 172.600 679.000 173.400 ;
        RECT 679.600 173.000 688.400 173.800 ;
        RECT 663.600 172.000 664.400 172.600 ;
        RECT 674.800 172.000 675.600 172.400 ;
        RECT 681.200 172.000 682.000 172.400 ;
        RECT 686.200 172.000 687.000 172.200 ;
        RECT 656.800 171.400 657.600 172.000 ;
        RECT 663.600 171.400 687.000 172.000 ;
        RECT 655.400 170.000 656.400 170.800 ;
        RECT 655.600 162.200 656.400 170.000 ;
        RECT 657.000 169.600 657.600 171.400 ;
        RECT 657.000 169.000 666.000 169.600 ;
        RECT 657.000 167.400 657.600 169.000 ;
        RECT 665.200 168.800 666.000 169.000 ;
        RECT 668.400 169.000 677.000 169.600 ;
        RECT 668.400 168.800 669.200 169.000 ;
        RECT 660.200 167.600 662.800 168.400 ;
        RECT 657.000 166.800 659.600 167.400 ;
        RECT 658.800 162.200 659.600 166.800 ;
        RECT 662.000 162.200 662.800 167.600 ;
        RECT 663.400 166.800 667.600 167.600 ;
        RECT 665.200 162.200 666.000 165.000 ;
        RECT 666.800 162.200 667.600 165.000 ;
        RECT 668.400 162.200 669.200 165.000 ;
        RECT 670.000 162.200 670.800 168.400 ;
        RECT 673.200 167.600 675.800 168.400 ;
        RECT 676.400 168.200 677.000 169.000 ;
        RECT 678.000 169.400 678.800 169.600 ;
        RECT 678.000 169.000 683.400 169.400 ;
        RECT 678.000 168.800 684.200 169.000 ;
        RECT 682.800 168.200 684.200 168.800 ;
        RECT 676.400 167.600 682.200 168.200 ;
        RECT 685.200 168.000 686.800 168.800 ;
        RECT 685.200 167.600 685.800 168.000 ;
        RECT 673.200 162.200 674.000 167.000 ;
        RECT 676.400 162.200 677.200 167.000 ;
        RECT 681.600 166.800 685.800 167.600 ;
        RECT 687.600 167.400 688.400 173.000 ;
        RECT 686.400 166.800 688.400 167.400 ;
        RECT 678.000 162.200 678.800 165.000 ;
        RECT 679.600 162.200 680.400 165.000 ;
        RECT 682.800 162.200 683.600 166.800 ;
        RECT 686.400 166.200 687.000 166.800 ;
        RECT 686.000 165.600 687.000 166.200 ;
        RECT 686.000 162.200 686.800 165.600 ;
        RECT 1.200 148.300 2.000 159.800 ;
        RECT 7.000 158.400 7.800 159.800 ;
        RECT 6.000 157.600 7.800 158.400 ;
        RECT 7.000 152.400 7.800 157.600 ;
        RECT 8.400 153.600 9.200 154.400 ;
        RECT 8.600 152.400 9.200 153.600 ;
        RECT 11.600 153.600 12.400 154.400 ;
        RECT 11.600 152.400 12.200 153.600 ;
        RECT 13.000 152.400 13.800 159.800 ;
        RECT 18.800 152.800 19.600 159.800 ;
        RECT 7.000 151.800 8.000 152.400 ;
        RECT 8.600 151.800 10.000 152.400 ;
        RECT 6.000 148.800 6.800 150.400 ;
        RECT 7.400 148.400 8.000 151.800 ;
        RECT 9.200 151.600 10.000 151.800 ;
        RECT 10.800 151.800 12.200 152.400 ;
        RECT 12.800 151.800 13.800 152.400 ;
        RECT 18.600 151.800 19.600 152.800 ;
        RECT 22.000 152.400 22.800 159.800 ;
        RECT 25.200 152.800 26.000 159.800 ;
        RECT 20.200 151.800 22.800 152.400 ;
        RECT 25.000 151.800 26.000 152.800 ;
        RECT 28.400 152.400 29.200 159.800 ;
        RECT 26.600 151.800 29.200 152.400 ;
        RECT 32.600 152.400 33.400 159.800 ;
        RECT 38.600 158.400 39.400 159.800 ;
        RECT 38.600 157.600 40.400 158.400 ;
        RECT 34.000 153.600 34.800 154.400 ;
        RECT 34.200 152.400 34.800 153.600 ;
        RECT 37.200 153.600 38.000 154.400 ;
        RECT 37.200 152.400 37.800 153.600 ;
        RECT 38.600 152.400 39.400 157.600 ;
        RECT 46.600 152.800 47.400 159.800 ;
        RECT 50.800 155.000 51.600 159.000 ;
        RECT 32.600 151.800 33.600 152.400 ;
        RECT 34.200 151.800 35.600 152.400 ;
        RECT 10.800 151.600 11.600 151.800 ;
        RECT 9.300 150.300 9.900 151.600 ;
        RECT 12.800 150.300 13.400 151.800 ;
        RECT 9.300 149.700 13.400 150.300 ;
        RECT 12.800 148.400 13.400 149.700 ;
        RECT 14.000 148.800 14.800 150.400 ;
        RECT 18.600 148.400 19.200 151.800 ;
        RECT 20.200 149.800 20.800 151.800 ;
        RECT 19.800 149.000 20.800 149.800 ;
        RECT 4.400 148.300 5.200 148.400 ;
        RECT 1.200 148.200 5.200 148.300 ;
        RECT 1.200 147.700 6.000 148.200 ;
        RECT 1.200 142.200 2.000 147.700 ;
        RECT 4.400 147.600 6.000 147.700 ;
        RECT 7.400 147.600 10.000 148.400 ;
        RECT 10.800 147.600 13.400 148.400 ;
        RECT 15.600 148.300 16.400 148.400 ;
        RECT 18.600 148.300 19.600 148.400 ;
        RECT 15.600 148.200 19.600 148.300 ;
        RECT 14.800 147.700 19.600 148.200 ;
        RECT 14.800 147.600 16.400 147.700 ;
        RECT 18.600 147.600 19.600 147.700 ;
        RECT 5.200 147.200 6.000 147.600 ;
        RECT 2.800 144.800 3.600 146.400 ;
        RECT 4.600 146.200 8.200 146.600 ;
        RECT 9.200 146.200 9.800 147.600 ;
        RECT 11.000 146.200 11.600 147.600 ;
        RECT 14.800 147.200 15.600 147.600 ;
        RECT 12.600 146.200 16.200 146.600 ;
        RECT 18.600 146.200 19.200 147.600 ;
        RECT 20.200 147.400 20.800 149.000 ;
        RECT 21.800 149.600 22.800 150.400 ;
        RECT 21.800 148.800 22.600 149.600 ;
        RECT 25.000 148.400 25.600 151.800 ;
        RECT 26.600 149.800 27.200 151.800 ;
        RECT 26.200 149.000 27.200 149.800 ;
        RECT 25.000 147.600 26.000 148.400 ;
        RECT 20.200 146.800 22.800 147.400 ;
        RECT 4.400 146.000 8.400 146.200 ;
        RECT 4.400 142.200 5.200 146.000 ;
        RECT 7.600 142.200 8.400 146.000 ;
        RECT 9.200 142.200 10.000 146.200 ;
        RECT 10.800 142.200 11.600 146.200 ;
        RECT 12.400 146.000 16.400 146.200 ;
        RECT 12.400 142.200 13.200 146.000 ;
        RECT 15.600 142.200 16.400 146.000 ;
        RECT 18.600 145.600 19.600 146.200 ;
        RECT 18.800 142.200 19.600 145.600 ;
        RECT 22.000 142.200 22.800 146.800 ;
        RECT 25.000 146.200 25.600 147.600 ;
        RECT 26.600 147.400 27.200 149.000 ;
        RECT 28.200 149.600 29.200 150.400 ;
        RECT 28.200 148.800 29.000 149.600 ;
        RECT 31.600 148.800 32.400 150.400 ;
        RECT 33.000 150.300 33.600 151.800 ;
        RECT 34.800 151.600 35.600 151.800 ;
        RECT 36.400 151.800 37.800 152.400 ;
        RECT 38.400 151.800 39.400 152.400 ;
        RECT 45.800 152.200 47.400 152.800 ;
        RECT 36.400 151.600 37.200 151.800 ;
        RECT 36.500 150.300 37.100 151.600 ;
        RECT 33.000 149.700 37.100 150.300 ;
        RECT 33.000 148.400 33.600 149.700 ;
        RECT 38.400 148.400 39.000 151.800 ;
        RECT 39.600 148.800 40.400 150.400 ;
        RECT 41.200 150.300 42.000 150.400 ;
        RECT 44.400 150.300 45.200 151.200 ;
        RECT 41.200 149.700 45.200 150.300 ;
        RECT 41.200 149.600 42.000 149.700 ;
        RECT 44.400 149.600 45.200 149.700 ;
        RECT 45.800 148.400 46.400 152.200 ;
        RECT 51.000 151.600 51.600 155.000 ;
        RECT 56.200 152.800 57.000 159.800 ;
        RECT 60.400 155.000 61.200 159.000 ;
        RECT 47.800 151.000 51.600 151.600 ;
        RECT 55.400 152.200 57.000 152.800 ;
        RECT 47.800 149.000 48.400 151.000 ;
        RECT 30.000 148.200 30.800 148.400 ;
        RECT 30.000 147.600 31.600 148.200 ;
        RECT 33.000 147.600 35.600 148.400 ;
        RECT 36.400 147.600 39.000 148.400 ;
        RECT 41.200 148.200 42.000 148.400 ;
        RECT 40.400 147.600 42.000 148.200 ;
        RECT 42.800 148.300 43.600 148.400 ;
        RECT 44.400 148.300 46.400 148.400 ;
        RECT 42.800 147.700 46.400 148.300 ;
        RECT 47.000 148.200 48.400 149.000 ;
        RECT 49.200 148.800 50.000 150.400 ;
        RECT 50.800 148.800 51.600 150.400 ;
        RECT 52.400 150.300 53.200 150.400 ;
        RECT 54.000 150.300 54.800 151.200 ;
        RECT 52.400 149.700 54.800 150.300 ;
        RECT 52.400 149.600 53.200 149.700 ;
        RECT 54.000 149.600 54.800 149.700 ;
        RECT 55.400 150.400 56.000 152.200 ;
        RECT 60.600 151.600 61.200 155.000 ;
        RECT 64.600 152.400 65.400 159.800 ;
        RECT 66.000 153.600 66.800 154.400 ;
        RECT 66.200 152.400 66.800 153.600 ;
        RECT 69.200 153.600 70.000 154.400 ;
        RECT 69.200 152.400 69.800 153.600 ;
        RECT 70.600 152.400 71.400 159.800 ;
        RECT 76.400 152.800 77.200 159.800 ;
        RECT 64.600 151.800 65.600 152.400 ;
        RECT 66.200 151.800 67.600 152.400 ;
        RECT 57.400 151.000 61.200 151.600 ;
        RECT 55.400 149.600 56.400 150.400 ;
        RECT 55.400 148.400 56.000 149.600 ;
        RECT 57.400 149.000 58.000 151.000 ;
        RECT 42.800 147.600 43.600 147.700 ;
        RECT 44.400 147.600 46.400 147.700 ;
        RECT 26.600 146.800 29.200 147.400 ;
        RECT 30.800 147.200 31.600 147.600 ;
        RECT 25.000 145.600 26.000 146.200 ;
        RECT 25.200 142.200 26.000 145.600 ;
        RECT 28.400 142.200 29.200 146.800 ;
        RECT 30.200 146.200 33.800 146.600 ;
        RECT 34.800 146.200 35.400 147.600 ;
        RECT 36.600 146.200 37.200 147.600 ;
        RECT 40.400 147.200 41.200 147.600 ;
        RECT 45.800 147.000 46.400 147.600 ;
        RECT 47.400 147.800 48.400 148.200 ;
        RECT 47.400 147.200 51.600 147.800 ;
        RECT 54.000 147.600 56.000 148.400 ;
        RECT 56.600 148.200 58.000 149.000 ;
        RECT 58.800 148.800 59.600 150.400 ;
        RECT 60.400 148.800 61.200 150.400 ;
        RECT 63.600 148.800 64.400 150.400 ;
        RECT 65.000 148.400 65.600 151.800 ;
        RECT 66.800 151.600 67.600 151.800 ;
        RECT 68.400 151.800 69.800 152.400 ;
        RECT 70.400 151.800 71.400 152.400 ;
        RECT 76.200 151.800 77.200 152.800 ;
        RECT 79.600 152.400 80.400 159.800 ;
        RECT 77.800 151.800 80.400 152.400 ;
        RECT 83.800 152.400 84.600 159.800 ;
        RECT 89.800 158.400 90.600 159.800 ;
        RECT 89.800 157.600 91.600 158.400 ;
        RECT 85.200 153.600 86.000 154.400 ;
        RECT 85.400 152.400 86.000 153.600 ;
        RECT 88.400 153.600 89.200 154.400 ;
        RECT 88.400 152.400 89.000 153.600 ;
        RECT 89.800 152.400 90.600 157.600 ;
        RECT 83.800 151.800 84.800 152.400 ;
        RECT 85.400 151.800 86.800 152.400 ;
        RECT 68.400 151.600 69.200 151.800 ;
        RECT 66.900 150.300 67.500 151.600 ;
        RECT 70.400 150.300 71.000 151.800 ;
        RECT 66.900 149.700 71.000 150.300 ;
        RECT 70.400 148.400 71.000 149.700 ;
        RECT 71.600 148.800 72.400 150.400 ;
        RECT 76.200 148.400 76.800 151.800 ;
        RECT 77.800 149.800 78.400 151.800 ;
        RECT 77.400 149.000 78.400 149.800 ;
        RECT 45.800 146.600 46.600 147.000 ;
        RECT 38.200 146.200 41.800 146.600 ;
        RECT 30.000 146.000 34.000 146.200 ;
        RECT 30.000 142.200 30.800 146.000 ;
        RECT 33.200 142.200 34.000 146.000 ;
        RECT 34.800 142.200 35.600 146.200 ;
        RECT 36.400 142.200 37.200 146.200 ;
        RECT 38.000 146.000 42.000 146.200 ;
        RECT 45.800 146.000 47.400 146.600 ;
        RECT 38.000 142.200 38.800 146.000 ;
        RECT 41.200 142.200 42.000 146.000 ;
        RECT 46.600 143.000 47.400 146.000 ;
        RECT 51.000 145.000 51.600 147.200 ;
        RECT 55.400 147.000 56.000 147.600 ;
        RECT 57.000 147.800 58.000 148.200 ;
        RECT 62.000 148.200 62.800 148.400 ;
        RECT 57.000 147.200 61.200 147.800 ;
        RECT 62.000 147.600 63.600 148.200 ;
        RECT 65.000 147.600 67.600 148.400 ;
        RECT 68.400 147.600 71.000 148.400 ;
        RECT 73.200 148.200 74.000 148.400 ;
        RECT 72.400 147.600 74.000 148.200 ;
        RECT 74.800 148.300 75.600 148.400 ;
        RECT 76.200 148.300 77.200 148.400 ;
        RECT 74.800 147.700 77.200 148.300 ;
        RECT 74.800 147.600 75.600 147.700 ;
        RECT 76.200 147.600 77.200 147.700 ;
        RECT 62.800 147.200 63.600 147.600 ;
        RECT 55.400 146.600 56.200 147.000 ;
        RECT 55.400 146.000 57.000 146.600 ;
        RECT 50.800 143.000 51.600 145.000 ;
        RECT 56.200 143.000 57.000 146.000 ;
        RECT 60.600 145.000 61.200 147.200 ;
        RECT 62.200 146.200 65.800 146.600 ;
        RECT 66.800 146.200 67.400 147.600 ;
        RECT 68.600 146.200 69.200 147.600 ;
        RECT 72.400 147.200 73.200 147.600 ;
        RECT 70.200 146.200 73.800 146.600 ;
        RECT 76.200 146.200 76.800 147.600 ;
        RECT 77.800 147.400 78.400 149.000 ;
        RECT 79.400 149.600 80.400 150.400 ;
        RECT 79.400 148.800 80.200 149.600 ;
        RECT 82.800 148.800 83.600 150.400 ;
        RECT 84.200 150.300 84.800 151.800 ;
        RECT 86.000 151.600 86.800 151.800 ;
        RECT 87.600 151.800 89.000 152.400 ;
        RECT 89.600 151.800 90.600 152.400 ;
        RECT 87.600 151.600 88.400 151.800 ;
        RECT 87.700 150.300 88.300 151.600 ;
        RECT 84.200 149.700 88.300 150.300 ;
        RECT 84.200 148.400 84.800 149.700 ;
        RECT 89.600 148.400 90.200 151.800 ;
        RECT 94.000 151.200 94.800 159.800 ;
        RECT 98.200 155.800 99.400 159.800 ;
        RECT 102.800 155.800 103.600 159.800 ;
        RECT 107.200 156.400 108.000 159.800 ;
        RECT 107.200 155.800 109.200 156.400 ;
        RECT 98.800 155.000 99.600 155.800 ;
        RECT 103.000 155.200 103.600 155.800 ;
        RECT 102.200 154.600 105.800 155.200 ;
        RECT 108.400 155.000 109.200 155.800 ;
        RECT 102.200 154.400 103.000 154.600 ;
        RECT 105.000 154.400 105.800 154.600 ;
        RECT 98.000 153.200 99.400 154.000 ;
        RECT 98.800 152.200 99.400 153.200 ;
        RECT 101.000 153.000 103.200 153.600 ;
        RECT 101.000 152.800 101.800 153.000 ;
        RECT 98.800 151.600 101.200 152.200 ;
        RECT 94.000 150.600 98.200 151.200 ;
        RECT 90.800 148.800 91.600 150.400 ;
        RECT 81.200 148.200 82.000 148.400 ;
        RECT 81.200 147.600 82.800 148.200 ;
        RECT 84.200 147.600 86.800 148.400 ;
        RECT 87.600 147.600 90.200 148.400 ;
        RECT 92.400 148.200 93.200 148.400 ;
        RECT 91.600 147.600 93.200 148.200 ;
        RECT 77.800 146.800 80.400 147.400 ;
        RECT 82.000 147.200 82.800 147.600 ;
        RECT 60.400 143.000 61.200 145.000 ;
        RECT 62.000 146.000 66.000 146.200 ;
        RECT 62.000 142.200 62.800 146.000 ;
        RECT 65.200 142.200 66.000 146.000 ;
        RECT 66.800 142.200 67.600 146.200 ;
        RECT 68.400 142.200 69.200 146.200 ;
        RECT 70.000 146.000 74.000 146.200 ;
        RECT 70.000 142.200 70.800 146.000 ;
        RECT 73.200 142.200 74.000 146.000 ;
        RECT 76.200 145.600 77.200 146.200 ;
        RECT 76.400 142.200 77.200 145.600 ;
        RECT 79.600 142.200 80.400 146.800 ;
        RECT 81.400 146.200 85.000 146.600 ;
        RECT 86.000 146.200 86.600 147.600 ;
        RECT 87.800 146.200 88.400 147.600 ;
        RECT 91.600 147.200 92.400 147.600 ;
        RECT 94.000 147.200 94.800 150.600 ;
        RECT 97.400 150.400 98.200 150.600 ;
        RECT 95.800 149.800 96.600 150.000 ;
        RECT 95.800 149.200 99.600 149.800 ;
        RECT 98.800 149.000 99.600 149.200 ;
        RECT 100.600 148.400 101.200 151.600 ;
        RECT 102.600 151.800 103.200 153.000 ;
        RECT 103.800 153.000 104.600 153.200 ;
        RECT 108.400 153.000 109.200 153.200 ;
        RECT 103.800 152.400 109.200 153.000 ;
        RECT 102.600 151.400 107.400 151.800 ;
        RECT 111.600 151.400 112.400 159.800 ;
        RECT 102.600 151.200 112.400 151.400 ;
        RECT 106.600 151.000 112.400 151.200 ;
        RECT 118.000 155.000 118.800 159.000 ;
        RECT 118.000 151.600 118.600 155.000 ;
        RECT 122.200 152.800 123.000 159.800 ;
        RECT 122.200 152.200 123.800 152.800 ;
        RECT 118.000 151.000 121.800 151.600 ;
        RECT 106.800 150.800 112.400 151.000 ;
        RECT 105.200 150.200 106.000 150.400 ;
        RECT 105.200 149.600 110.200 150.200 ;
        RECT 109.400 149.400 110.200 149.600 ;
        RECT 118.000 148.800 118.800 150.400 ;
        RECT 119.600 148.800 120.400 150.400 ;
        RECT 121.200 149.000 121.800 151.000 ;
        RECT 107.800 148.400 108.600 148.600 ;
        RECT 100.600 147.800 111.600 148.400 ;
        RECT 121.200 148.200 122.600 149.000 ;
        RECT 123.200 148.400 123.800 152.200 ;
        RECT 130.200 152.400 131.000 159.800 ;
        RECT 131.600 153.600 132.400 154.400 ;
        RECT 131.800 152.400 132.400 153.600 ;
        RECT 134.000 152.400 134.800 159.800 ;
        RECT 137.200 152.800 138.000 159.800 ;
        RECT 140.400 155.000 141.200 159.000 ;
        RECT 130.200 151.800 131.200 152.400 ;
        RECT 131.800 151.800 133.200 152.400 ;
        RECT 134.000 151.800 136.600 152.400 ;
        RECT 137.200 151.800 138.200 152.800 ;
        RECT 124.400 149.600 125.200 151.200 ;
        RECT 130.600 150.400 131.200 151.800 ;
        RECT 132.400 151.600 133.200 151.800 ;
        RECT 127.600 150.300 128.400 150.400 ;
        RECT 129.200 150.300 130.000 150.400 ;
        RECT 127.600 149.700 130.000 150.300 ;
        RECT 127.600 149.600 128.400 149.700 ;
        RECT 129.200 148.800 130.000 149.700 ;
        RECT 130.600 149.600 131.600 150.400 ;
        RECT 134.000 149.600 135.000 150.400 ;
        RECT 130.600 148.400 131.200 149.600 ;
        RECT 134.200 148.800 135.000 149.600 ;
        RECT 136.000 149.800 136.600 151.800 ;
        RECT 136.000 149.000 137.000 149.800 ;
        RECT 121.200 147.800 122.200 148.200 ;
        RECT 101.000 147.600 101.800 147.800 ;
        RECT 106.800 147.600 107.600 147.800 ;
        RECT 110.000 147.600 111.600 147.800 ;
        RECT 94.000 146.600 98.000 147.200 ;
        RECT 89.400 146.200 93.000 146.600 ;
        RECT 81.200 146.000 85.200 146.200 ;
        RECT 81.200 142.200 82.000 146.000 ;
        RECT 84.400 142.200 85.200 146.000 ;
        RECT 86.000 142.200 86.800 146.200 ;
        RECT 87.600 142.200 88.400 146.200 ;
        RECT 89.200 146.000 93.200 146.200 ;
        RECT 89.200 142.200 90.000 146.000 ;
        RECT 92.400 142.200 93.200 146.000 ;
        RECT 94.000 142.200 94.800 146.600 ;
        RECT 97.000 146.400 98.000 146.600 ;
        RECT 97.200 146.300 98.000 146.400 ;
        RECT 100.400 146.300 101.200 146.400 ;
        RECT 97.200 145.700 101.200 146.300 ;
        RECT 100.400 145.600 101.200 145.700 ;
        RECT 106.800 145.600 107.400 147.600 ;
        RECT 118.000 147.200 122.200 147.800 ;
        RECT 123.200 147.600 125.200 148.400 ;
        RECT 127.600 148.200 128.400 148.400 ;
        RECT 127.600 147.600 129.200 148.200 ;
        RECT 130.600 147.600 133.200 148.400 ;
        RECT 105.000 145.400 105.800 145.600 ;
        RECT 98.800 144.200 99.600 145.000 ;
        RECT 103.000 144.800 105.800 145.400 ;
        RECT 106.800 144.800 107.600 145.600 ;
        RECT 103.000 144.200 103.600 144.800 ;
        RECT 108.400 144.200 109.200 145.000 ;
        RECT 98.200 143.600 99.600 144.200 ;
        RECT 98.200 142.200 99.400 143.600 ;
        RECT 102.800 142.200 103.600 144.200 ;
        RECT 107.200 143.600 109.200 144.200 ;
        RECT 107.200 142.200 108.000 143.600 ;
        RECT 111.600 142.200 112.400 147.000 ;
        RECT 118.000 145.000 118.600 147.200 ;
        RECT 123.200 147.000 123.800 147.600 ;
        RECT 128.400 147.200 129.200 147.600 ;
        RECT 123.000 146.600 123.800 147.000 ;
        RECT 122.200 146.400 123.800 146.600 ;
        RECT 121.200 146.000 123.800 146.400 ;
        RECT 127.800 146.200 131.400 146.600 ;
        RECT 132.400 146.200 133.000 147.600 ;
        RECT 136.000 147.400 136.600 149.000 ;
        RECT 137.600 148.400 138.200 151.800 ;
        RECT 140.400 151.600 141.000 155.000 ;
        RECT 144.600 152.800 145.400 159.800 ;
        RECT 144.600 152.200 146.200 152.800 ;
        RECT 140.400 151.000 144.200 151.600 ;
        RECT 140.400 148.800 141.200 150.400 ;
        RECT 142.000 148.800 142.800 150.400 ;
        RECT 143.600 149.000 144.200 151.000 ;
        RECT 137.200 148.300 138.200 148.400 ;
        RECT 138.800 148.300 139.600 148.400 ;
        RECT 137.200 147.700 139.600 148.300 ;
        RECT 143.600 148.200 145.000 149.000 ;
        RECT 145.600 148.400 146.200 152.200 ;
        RECT 152.600 152.400 153.400 159.800 ;
        RECT 154.000 153.600 154.800 154.400 ;
        RECT 154.200 152.400 154.800 153.600 ;
        RECT 157.200 153.600 158.000 154.400 ;
        RECT 157.200 152.400 157.800 153.600 ;
        RECT 158.600 152.400 159.400 159.800 ;
        RECT 152.600 151.800 153.600 152.400 ;
        RECT 154.200 151.800 155.600 152.400 ;
        RECT 146.800 150.300 147.600 151.200 ;
        RECT 148.400 150.300 149.200 150.400 ;
        RECT 146.800 149.700 149.200 150.300 ;
        RECT 146.800 149.600 147.600 149.700 ;
        RECT 148.400 149.600 149.200 149.700 ;
        RECT 151.600 148.800 152.400 150.400 ;
        RECT 153.000 148.400 153.600 151.800 ;
        RECT 154.800 151.600 155.600 151.800 ;
        RECT 156.400 151.800 157.800 152.400 ;
        RECT 158.400 151.800 159.400 152.400 ;
        RECT 156.400 151.600 157.200 151.800 ;
        RECT 154.900 150.300 155.500 151.600 ;
        RECT 158.400 150.300 159.000 151.800 ;
        RECT 162.800 151.400 163.600 159.800 ;
        RECT 167.200 156.400 168.000 159.800 ;
        RECT 166.000 155.800 168.000 156.400 ;
        RECT 171.600 155.800 172.400 159.800 ;
        RECT 175.800 155.800 177.000 159.800 ;
        RECT 166.000 155.000 166.800 155.800 ;
        RECT 171.600 155.200 172.200 155.800 ;
        RECT 169.400 154.600 173.000 155.200 ;
        RECT 175.600 155.000 176.400 155.800 ;
        RECT 169.400 154.400 170.200 154.600 ;
        RECT 172.200 154.400 173.000 154.600 ;
        RECT 180.400 154.300 181.200 159.800 ;
        RECT 182.000 154.300 182.800 154.400 ;
        RECT 166.000 153.000 166.800 153.200 ;
        RECT 170.600 153.000 171.400 153.200 ;
        RECT 166.000 152.400 171.400 153.000 ;
        RECT 172.000 153.000 174.200 153.600 ;
        RECT 172.000 151.800 172.600 153.000 ;
        RECT 173.400 152.800 174.200 153.000 ;
        RECT 175.800 153.200 177.200 154.000 ;
        RECT 180.400 153.700 182.800 154.300 ;
        RECT 175.800 152.200 176.400 153.200 ;
        RECT 167.800 151.400 172.600 151.800 ;
        RECT 162.800 151.200 172.600 151.400 ;
        RECT 174.000 151.600 176.400 152.200 ;
        RECT 162.800 151.000 168.600 151.200 ;
        RECT 162.800 150.800 168.400 151.000 ;
        RECT 154.900 149.700 159.000 150.300 ;
        RECT 158.400 148.400 159.000 149.700 ;
        RECT 159.600 148.800 160.400 150.400 ;
        RECT 169.200 150.200 170.000 150.400 ;
        RECT 165.000 149.600 170.000 150.200 ;
        RECT 165.000 149.400 165.800 149.600 ;
        RECT 167.600 149.400 168.400 149.600 ;
        RECT 166.600 148.400 167.400 148.600 ;
        RECT 174.000 148.400 174.600 151.600 ;
        RECT 180.400 151.200 181.200 153.700 ;
        RECT 182.000 153.600 182.800 153.700 ;
        RECT 177.000 150.600 181.200 151.200 ;
        RECT 177.000 150.400 177.800 150.600 ;
        RECT 178.600 149.800 179.400 150.000 ;
        RECT 175.600 149.200 179.400 149.800 ;
        RECT 175.600 149.000 176.400 149.200 ;
        RECT 143.600 147.800 144.600 148.200 ;
        RECT 137.200 147.600 138.200 147.700 ;
        RECT 138.800 147.600 139.600 147.700 ;
        RECT 134.000 146.800 136.600 147.400 ;
        RECT 127.600 146.000 131.600 146.200 ;
        RECT 121.200 145.600 123.000 146.000 ;
        RECT 118.000 143.000 118.800 145.000 ;
        RECT 122.200 143.000 123.000 145.600 ;
        RECT 127.600 142.200 128.400 146.000 ;
        RECT 130.800 142.200 131.600 146.000 ;
        RECT 132.400 142.200 133.200 146.200 ;
        RECT 134.000 142.200 134.800 146.800 ;
        RECT 137.600 146.200 138.200 147.600 ;
        RECT 137.200 145.600 138.200 146.200 ;
        RECT 140.400 147.200 144.600 147.800 ;
        RECT 145.600 147.600 147.600 148.400 ;
        RECT 150.000 148.200 150.800 148.400 ;
        RECT 150.000 147.600 151.600 148.200 ;
        RECT 153.000 147.600 155.600 148.400 ;
        RECT 156.400 147.600 159.000 148.400 ;
        RECT 161.200 148.200 162.000 148.400 ;
        RECT 160.400 147.600 162.000 148.200 ;
        RECT 163.600 147.800 174.600 148.400 ;
        RECT 163.600 147.600 165.200 147.800 ;
        RECT 137.200 142.200 138.000 145.600 ;
        RECT 140.400 145.000 141.000 147.200 ;
        RECT 145.600 147.000 146.200 147.600 ;
        RECT 150.800 147.200 151.600 147.600 ;
        RECT 145.400 146.600 146.200 147.000 ;
        RECT 144.600 146.000 146.200 146.600 ;
        RECT 150.200 146.200 153.800 146.600 ;
        RECT 154.800 146.200 155.400 147.600 ;
        RECT 156.600 146.200 157.200 147.600 ;
        RECT 160.400 147.200 161.200 147.600 ;
        RECT 158.200 146.200 161.800 146.600 ;
        RECT 150.000 146.000 154.000 146.200 ;
        RECT 140.400 143.000 141.200 145.000 ;
        RECT 144.600 143.000 145.400 146.000 ;
        RECT 150.000 142.200 150.800 146.000 ;
        RECT 153.200 142.200 154.000 146.000 ;
        RECT 154.800 142.200 155.600 146.200 ;
        RECT 156.400 142.200 157.200 146.200 ;
        RECT 158.000 146.000 162.000 146.200 ;
        RECT 158.000 142.200 158.800 146.000 ;
        RECT 161.200 142.200 162.000 146.000 ;
        RECT 162.800 142.200 163.600 147.000 ;
        RECT 167.800 145.600 168.400 147.800 ;
        RECT 173.400 147.600 174.200 147.800 ;
        RECT 180.400 147.200 181.200 150.600 ;
        RECT 177.400 146.600 181.200 147.200 ;
        RECT 177.400 146.400 178.200 146.600 ;
        RECT 166.000 144.200 166.800 145.000 ;
        RECT 167.600 144.800 168.400 145.600 ;
        RECT 169.400 145.400 170.200 145.600 ;
        RECT 169.400 144.800 172.200 145.400 ;
        RECT 171.600 144.200 172.200 144.800 ;
        RECT 175.600 144.200 176.400 145.000 ;
        RECT 166.000 143.600 168.000 144.200 ;
        RECT 167.200 142.200 168.000 143.600 ;
        RECT 171.600 142.200 172.400 144.200 ;
        RECT 175.600 143.600 177.000 144.200 ;
        RECT 175.800 142.200 177.000 143.600 ;
        RECT 180.400 142.200 181.200 146.600 ;
        RECT 182.000 144.800 182.800 146.400 ;
        RECT 183.600 142.200 184.400 159.800 ;
        RECT 185.200 155.000 186.000 159.000 ;
        RECT 189.400 158.400 190.200 159.800 ;
        RECT 188.400 157.600 190.200 158.400 ;
        RECT 185.200 151.600 185.800 155.000 ;
        RECT 189.400 152.800 190.200 157.600 ;
        RECT 194.800 155.000 195.600 159.000 ;
        RECT 189.400 152.200 191.000 152.800 ;
        RECT 185.200 151.000 189.000 151.600 ;
        RECT 185.200 148.800 186.000 150.400 ;
        RECT 186.800 148.800 187.600 150.400 ;
        RECT 188.400 149.000 189.000 151.000 ;
        RECT 188.400 148.200 189.800 149.000 ;
        RECT 190.400 148.400 191.000 152.200 ;
        RECT 194.800 151.600 195.400 155.000 ;
        RECT 199.000 152.800 199.800 159.800 ;
        RECT 199.000 152.200 200.600 152.800 ;
        RECT 191.600 149.600 192.400 151.200 ;
        RECT 194.800 151.000 198.600 151.600 ;
        RECT 194.800 148.800 195.600 150.400 ;
        RECT 196.400 148.800 197.200 150.400 ;
        RECT 198.000 149.000 198.600 151.000 ;
        RECT 188.400 147.800 189.400 148.200 ;
        RECT 185.200 147.200 189.400 147.800 ;
        RECT 190.400 147.600 192.400 148.400 ;
        RECT 198.000 148.200 199.400 149.000 ;
        RECT 200.000 148.400 200.600 152.200 ;
        RECT 207.000 152.400 207.800 159.800 ;
        RECT 208.400 153.600 209.200 154.400 ;
        RECT 208.600 152.400 209.200 153.600 ;
        RECT 211.600 153.600 212.400 154.400 ;
        RECT 211.600 152.400 212.200 153.600 ;
        RECT 213.000 152.400 213.800 159.800 ;
        RECT 207.000 151.800 208.000 152.400 ;
        RECT 208.600 151.800 210.000 152.400 ;
        RECT 201.200 149.600 202.000 151.200 ;
        RECT 206.000 148.800 206.800 150.400 ;
        RECT 207.400 150.300 208.000 151.800 ;
        RECT 209.200 151.600 210.000 151.800 ;
        RECT 210.800 151.800 212.200 152.400 ;
        RECT 212.800 151.800 213.800 152.400 ;
        RECT 210.800 151.600 211.600 151.800 ;
        RECT 210.900 150.300 211.500 151.600 ;
        RECT 212.800 150.400 213.400 151.800 ;
        RECT 217.200 151.200 218.000 159.800 ;
        RECT 221.400 155.800 222.600 159.800 ;
        RECT 226.000 155.800 226.800 159.800 ;
        RECT 230.400 156.400 231.200 159.800 ;
        RECT 230.400 155.800 232.400 156.400 ;
        RECT 222.000 155.000 222.800 155.800 ;
        RECT 226.200 155.200 226.800 155.800 ;
        RECT 225.400 154.600 229.000 155.200 ;
        RECT 231.600 155.000 232.400 155.800 ;
        RECT 225.400 154.400 226.200 154.600 ;
        RECT 228.200 154.400 229.000 154.600 ;
        RECT 221.200 153.200 222.600 154.000 ;
        RECT 222.000 152.200 222.600 153.200 ;
        RECT 224.200 153.000 226.400 153.600 ;
        RECT 224.200 152.800 225.000 153.000 ;
        RECT 222.000 151.600 224.400 152.200 ;
        RECT 217.200 150.600 221.400 151.200 ;
        RECT 207.400 149.700 211.500 150.300 ;
        RECT 207.400 148.400 208.000 149.700 ;
        RECT 212.400 149.600 213.400 150.400 ;
        RECT 212.800 148.400 213.400 149.600 ;
        RECT 214.000 148.800 214.800 150.400 ;
        RECT 200.000 148.300 202.000 148.400 ;
        RECT 202.800 148.300 203.600 148.400 ;
        RECT 198.000 147.800 199.000 148.200 ;
        RECT 185.200 145.000 185.800 147.200 ;
        RECT 190.400 147.000 191.000 147.600 ;
        RECT 190.200 146.600 191.000 147.000 ;
        RECT 189.400 146.000 191.000 146.600 ;
        RECT 194.800 147.200 199.000 147.800 ;
        RECT 200.000 147.700 203.600 148.300 ;
        RECT 200.000 147.600 202.000 147.700 ;
        RECT 202.800 147.600 203.600 147.700 ;
        RECT 204.400 148.200 205.200 148.400 ;
        RECT 204.400 147.600 206.000 148.200 ;
        RECT 207.400 147.600 210.000 148.400 ;
        RECT 210.800 147.600 213.400 148.400 ;
        RECT 215.600 148.200 216.400 148.400 ;
        RECT 214.800 147.600 216.400 148.200 ;
        RECT 185.200 143.000 186.000 145.000 ;
        RECT 189.400 143.000 190.200 146.000 ;
        RECT 194.800 145.000 195.400 147.200 ;
        RECT 200.000 147.000 200.600 147.600 ;
        RECT 205.200 147.200 206.000 147.600 ;
        RECT 199.800 146.600 200.600 147.000 ;
        RECT 199.000 146.000 200.600 146.600 ;
        RECT 204.600 146.200 208.200 146.600 ;
        RECT 209.200 146.200 209.800 147.600 ;
        RECT 211.000 146.200 211.600 147.600 ;
        RECT 214.800 147.200 215.600 147.600 ;
        RECT 217.200 147.200 218.000 150.600 ;
        RECT 220.600 150.400 221.400 150.600 ;
        RECT 219.000 149.800 219.800 150.000 ;
        RECT 219.000 149.200 222.800 149.800 ;
        RECT 222.000 149.000 222.800 149.200 ;
        RECT 223.800 148.400 224.400 151.600 ;
        RECT 225.800 151.800 226.400 153.000 ;
        RECT 227.000 153.000 227.800 153.200 ;
        RECT 231.600 153.000 232.400 153.200 ;
        RECT 227.000 152.400 232.400 153.000 ;
        RECT 225.800 151.400 230.600 151.800 ;
        RECT 234.800 151.400 235.600 159.800 ;
        RECT 225.800 151.200 235.600 151.400 ;
        RECT 229.800 151.000 235.600 151.200 ;
        RECT 236.400 155.000 237.200 159.000 ;
        RECT 240.600 158.400 241.400 159.800 ;
        RECT 240.600 157.600 242.000 158.400 ;
        RECT 236.400 151.600 237.000 155.000 ;
        RECT 240.600 152.800 241.400 157.600 ;
        RECT 246.000 155.000 246.800 159.000 ;
        RECT 240.600 152.200 242.200 152.800 ;
        RECT 236.400 151.000 240.200 151.600 ;
        RECT 230.000 150.800 235.600 151.000 ;
        RECT 228.400 150.200 229.200 150.400 ;
        RECT 228.400 149.600 233.400 150.200 ;
        RECT 232.600 149.400 233.400 149.600 ;
        RECT 236.400 148.800 237.200 150.400 ;
        RECT 238.000 148.800 238.800 150.400 ;
        RECT 239.600 149.000 240.200 151.000 ;
        RECT 231.000 148.400 231.800 148.600 ;
        RECT 223.800 147.800 234.800 148.400 ;
        RECT 239.600 148.200 241.000 149.000 ;
        RECT 241.600 148.400 242.200 152.200 ;
        RECT 246.000 151.600 246.600 155.000 ;
        RECT 250.200 152.800 251.000 159.800 ;
        RECT 250.200 152.200 251.800 152.800 ;
        RECT 242.800 149.600 243.600 151.200 ;
        RECT 246.000 151.000 249.800 151.600 ;
        RECT 246.000 148.800 246.800 150.400 ;
        RECT 247.600 148.800 248.400 150.400 ;
        RECT 249.200 149.000 249.800 151.000 ;
        RECT 239.600 147.800 240.600 148.200 ;
        RECT 224.200 147.600 225.000 147.800 ;
        RECT 217.200 146.600 221.000 147.200 ;
        RECT 212.600 146.200 216.200 146.600 ;
        RECT 204.400 146.000 208.400 146.200 ;
        RECT 194.800 143.000 195.600 145.000 ;
        RECT 199.000 143.000 199.800 146.000 ;
        RECT 204.400 142.200 205.200 146.000 ;
        RECT 207.600 142.200 208.400 146.000 ;
        RECT 209.200 142.200 210.000 146.200 ;
        RECT 210.800 142.200 211.600 146.200 ;
        RECT 212.400 146.000 216.400 146.200 ;
        RECT 212.400 142.200 213.200 146.000 ;
        RECT 215.600 142.200 216.400 146.000 ;
        RECT 217.200 142.200 218.000 146.600 ;
        RECT 220.200 146.400 221.000 146.600 ;
        RECT 230.000 145.600 230.600 147.800 ;
        RECT 233.200 147.600 234.800 147.800 ;
        RECT 236.400 147.200 240.600 147.800 ;
        RECT 241.600 147.600 243.600 148.400 ;
        RECT 249.200 148.200 250.600 149.000 ;
        RECT 251.200 148.400 251.800 152.200 ;
        RECT 255.600 152.400 256.400 159.800 ;
        RECT 257.400 152.400 258.200 152.600 ;
        RECT 255.600 151.800 258.200 152.400 ;
        RECT 260.000 151.800 261.600 159.800 ;
        RECT 263.600 152.400 264.400 152.600 ;
        RECT 265.200 152.400 266.000 159.800 ;
        RECT 273.200 156.400 274.000 159.800 ;
        RECT 273.000 155.800 274.000 156.400 ;
        RECT 273.000 155.200 273.600 155.800 ;
        RECT 276.400 155.200 277.200 159.800 ;
        RECT 279.600 157.000 280.400 159.800 ;
        RECT 281.200 157.000 282.000 159.800 ;
        RECT 263.600 151.800 266.000 152.400 ;
        RECT 271.600 154.600 273.600 155.200 ;
        RECT 252.400 150.300 253.200 151.200 ;
        RECT 258.600 150.400 259.400 150.600 ;
        RECT 260.600 150.400 261.200 151.800 ;
        RECT 252.400 149.700 256.300 150.300 ;
        RECT 252.400 149.600 253.200 149.700 ;
        RECT 255.700 148.400 256.300 149.700 ;
        RECT 257.800 149.800 259.400 150.400 ;
        RECT 257.800 149.600 258.600 149.800 ;
        RECT 260.400 149.600 261.200 150.400 ;
        RECT 259.200 148.600 260.000 148.800 ;
        RECT 257.200 148.400 260.000 148.600 ;
        RECT 249.200 147.800 250.200 148.200 ;
        RECT 228.200 145.400 229.000 145.600 ;
        RECT 222.000 144.200 222.800 145.000 ;
        RECT 226.200 144.800 229.000 145.400 ;
        RECT 230.000 144.800 230.800 145.600 ;
        RECT 226.200 144.200 226.800 144.800 ;
        RECT 231.600 144.200 232.400 145.000 ;
        RECT 221.400 143.600 222.800 144.200 ;
        RECT 221.400 142.200 222.600 143.600 ;
        RECT 226.000 142.200 226.800 144.200 ;
        RECT 230.400 143.600 232.400 144.200 ;
        RECT 230.400 142.200 231.200 143.600 ;
        RECT 234.800 142.200 235.600 147.000 ;
        RECT 236.400 145.000 237.000 147.200 ;
        RECT 241.600 147.000 242.200 147.600 ;
        RECT 241.400 146.600 242.200 147.000 ;
        RECT 240.600 146.000 242.200 146.600 ;
        RECT 246.000 147.200 250.200 147.800 ;
        RECT 251.200 147.600 253.200 148.400 ;
        RECT 255.600 148.000 260.000 148.400 ;
        RECT 260.600 148.400 261.200 149.600 ;
        RECT 271.600 149.000 272.400 154.600 ;
        RECT 274.200 154.400 278.400 155.200 ;
        RECT 282.800 155.000 283.600 159.800 ;
        RECT 286.000 155.000 286.800 159.800 ;
        RECT 274.200 154.000 274.800 154.400 ;
        RECT 273.200 153.200 274.800 154.000 ;
        RECT 277.800 153.800 283.600 154.400 ;
        RECT 275.800 153.200 277.200 153.800 ;
        RECT 275.800 153.000 282.000 153.200 ;
        RECT 276.600 152.600 282.000 153.000 ;
        RECT 281.200 152.400 282.000 152.600 ;
        RECT 283.000 153.000 283.600 153.800 ;
        RECT 284.200 153.600 286.800 154.400 ;
        RECT 289.200 153.600 290.000 159.800 ;
        RECT 290.800 157.000 291.600 159.800 ;
        RECT 292.400 157.000 293.200 159.800 ;
        RECT 294.000 157.000 294.800 159.800 ;
        RECT 292.400 154.400 296.600 155.200 ;
        RECT 297.200 154.400 298.000 159.800 ;
        RECT 300.400 155.200 301.200 159.800 ;
        RECT 300.400 154.600 303.000 155.200 ;
        RECT 297.200 153.600 299.800 154.400 ;
        RECT 290.800 153.000 291.600 153.200 ;
        RECT 283.000 152.400 291.600 153.000 ;
        RECT 294.000 153.000 294.800 153.200 ;
        RECT 302.400 153.000 303.000 154.600 ;
        RECT 294.000 152.400 303.000 153.000 ;
        RECT 274.800 151.800 275.600 152.400 ;
        RECT 278.200 151.800 279.000 152.000 ;
        RECT 274.800 151.200 301.800 151.800 ;
        RECT 301.000 151.000 301.800 151.200 ;
        RECT 302.400 150.600 303.000 152.400 ;
        RECT 303.600 154.300 304.400 159.800 ;
        RECT 305.200 154.300 306.000 154.400 ;
        RECT 303.600 153.700 306.000 154.300 ;
        RECT 303.600 152.000 304.400 153.700 ;
        RECT 305.200 153.600 306.000 153.700 ;
        RECT 309.400 152.400 310.200 159.800 ;
        RECT 314.800 156.400 315.600 159.800 ;
        RECT 314.600 155.800 315.600 156.400 ;
        RECT 314.600 155.200 315.200 155.800 ;
        RECT 318.000 155.200 318.800 159.800 ;
        RECT 321.200 157.000 322.000 159.800 ;
        RECT 322.800 157.000 323.600 159.800 ;
        RECT 313.200 154.600 315.200 155.200 ;
        RECT 310.800 153.600 312.400 154.400 ;
        RECT 311.000 152.400 311.600 153.600 ;
        RECT 303.600 151.200 304.600 152.000 ;
        RECT 309.400 151.800 310.400 152.400 ;
        RECT 311.000 151.800 312.400 152.400 ;
        RECT 302.400 150.000 303.200 150.600 ;
        RECT 255.600 147.800 257.800 148.000 ;
        RECT 260.600 147.800 261.600 148.400 ;
        RECT 255.600 147.600 257.200 147.800 ;
        RECT 236.400 143.000 237.200 145.000 ;
        RECT 240.600 143.000 241.400 146.000 ;
        RECT 246.000 145.000 246.600 147.200 ;
        RECT 251.200 147.000 251.800 147.600 ;
        RECT 251.000 146.600 251.800 147.000 ;
        RECT 257.400 146.800 258.200 147.000 ;
        RECT 250.200 146.400 251.800 146.600 ;
        RECT 249.200 146.000 251.800 146.400 ;
        RECT 255.600 146.200 258.200 146.800 ;
        RECT 258.800 146.400 260.400 147.200 ;
        RECT 249.200 145.600 251.000 146.000 ;
        RECT 246.000 143.000 246.800 145.000 ;
        RECT 250.200 143.000 251.000 145.600 ;
        RECT 255.600 142.200 256.400 146.200 ;
        RECT 261.000 145.800 261.600 147.800 ;
        RECT 262.400 147.600 263.200 148.400 ;
        RECT 264.400 147.600 266.000 148.400 ;
        RECT 271.600 148.200 280.400 149.000 ;
        RECT 281.000 148.600 283.000 149.400 ;
        RECT 286.800 148.600 290.000 149.400 ;
        RECT 262.400 147.200 263.000 147.600 ;
        RECT 262.200 146.400 263.000 147.200 ;
        RECT 263.600 146.800 264.400 147.000 ;
        RECT 263.600 146.200 266.000 146.800 ;
        RECT 260.000 142.200 261.600 145.800 ;
        RECT 265.200 142.200 266.000 146.200 ;
        RECT 271.600 142.200 272.400 148.200 ;
        RECT 274.000 146.800 277.000 147.600 ;
        RECT 276.200 146.200 277.000 146.800 ;
        RECT 282.200 146.200 283.000 148.600 ;
        RECT 284.400 146.800 285.200 148.400 ;
        RECT 289.600 147.800 290.400 148.000 ;
        RECT 286.000 147.200 290.400 147.800 ;
        RECT 286.000 147.000 286.800 147.200 ;
        RECT 292.400 146.400 293.200 149.200 ;
        RECT 298.200 148.600 302.000 149.400 ;
        RECT 298.200 147.400 299.000 148.600 ;
        RECT 302.600 148.000 303.200 150.000 ;
        RECT 286.000 146.200 286.800 146.400 ;
        RECT 276.200 145.400 278.800 146.200 ;
        RECT 282.200 145.600 286.800 146.200 ;
        RECT 287.600 145.600 289.200 146.400 ;
        RECT 292.200 145.600 293.200 146.400 ;
        RECT 297.200 146.800 299.000 147.400 ;
        RECT 302.000 147.400 303.200 148.000 ;
        RECT 297.200 146.200 298.000 146.800 ;
        RECT 278.000 142.200 278.800 145.400 ;
        RECT 295.600 145.400 298.000 146.200 ;
        RECT 279.600 142.200 280.400 145.000 ;
        RECT 281.200 142.200 282.000 145.000 ;
        RECT 282.800 142.200 283.600 145.000 ;
        RECT 286.000 142.200 286.800 145.000 ;
        RECT 289.200 142.200 290.000 145.000 ;
        RECT 290.800 142.200 291.600 145.000 ;
        RECT 292.400 142.200 293.200 145.000 ;
        RECT 294.000 142.200 294.800 145.000 ;
        RECT 295.600 142.200 296.400 145.400 ;
        RECT 302.000 142.200 302.800 147.400 ;
        RECT 303.800 146.800 304.600 151.200 ;
        RECT 306.800 150.300 307.600 150.400 ;
        RECT 308.400 150.300 309.200 150.400 ;
        RECT 306.800 149.700 309.200 150.300 ;
        RECT 306.800 149.600 307.600 149.700 ;
        RECT 308.400 148.800 309.200 149.700 ;
        RECT 309.800 148.400 310.400 151.800 ;
        RECT 311.600 151.600 312.400 151.800 ;
        RECT 313.200 149.000 314.000 154.600 ;
        RECT 315.800 154.400 320.000 155.200 ;
        RECT 324.400 155.000 325.200 159.800 ;
        RECT 327.600 155.000 328.400 159.800 ;
        RECT 315.800 154.000 316.400 154.400 ;
        RECT 314.800 153.200 316.400 154.000 ;
        RECT 319.400 153.800 325.200 154.400 ;
        RECT 317.400 153.200 318.800 153.800 ;
        RECT 317.400 153.000 323.600 153.200 ;
        RECT 318.200 152.600 323.600 153.000 ;
        RECT 322.800 152.400 323.600 152.600 ;
        RECT 324.600 153.000 325.200 153.800 ;
        RECT 325.800 153.600 328.400 154.400 ;
        RECT 330.800 153.600 331.600 159.800 ;
        RECT 332.400 157.000 333.200 159.800 ;
        RECT 334.000 157.000 334.800 159.800 ;
        RECT 335.600 157.000 336.400 159.800 ;
        RECT 334.000 154.400 338.200 155.200 ;
        RECT 338.800 154.400 339.600 159.800 ;
        RECT 342.000 155.200 342.800 159.800 ;
        RECT 342.000 154.600 344.600 155.200 ;
        RECT 338.800 153.600 341.400 154.400 ;
        RECT 332.400 153.000 333.200 153.200 ;
        RECT 324.600 152.400 333.200 153.000 ;
        RECT 335.600 153.000 336.400 153.200 ;
        RECT 344.000 153.000 344.600 154.600 ;
        RECT 335.600 152.400 344.600 153.000 ;
        RECT 344.000 150.600 344.600 152.400 ;
        RECT 345.200 152.000 346.000 159.800 ;
        RECT 348.400 154.300 349.200 154.400 ;
        RECT 350.000 154.300 350.800 159.800 ;
        RECT 353.200 155.200 354.000 159.800 ;
        RECT 348.400 153.700 350.800 154.300 ;
        RECT 348.400 153.600 349.200 153.700 ;
        RECT 350.000 152.000 350.800 153.700 ;
        RECT 345.200 151.200 346.200 152.000 ;
        RECT 314.600 150.000 338.000 150.600 ;
        RECT 344.000 150.000 344.800 150.600 ;
        RECT 314.600 149.800 315.400 150.000 ;
        RECT 319.600 149.600 320.400 150.000 ;
        RECT 337.200 149.400 338.000 150.000 ;
        RECT 305.200 148.300 306.000 148.400 ;
        RECT 306.800 148.300 307.600 148.400 ;
        RECT 305.200 148.200 307.600 148.300 ;
        RECT 305.200 147.700 308.400 148.200 ;
        RECT 305.200 147.600 306.000 147.700 ;
        RECT 306.800 147.600 308.400 147.700 ;
        RECT 309.800 147.600 312.400 148.400 ;
        RECT 313.200 148.200 322.000 149.000 ;
        RECT 322.600 148.600 324.600 149.400 ;
        RECT 328.400 148.600 331.600 149.400 ;
        RECT 307.600 147.200 308.400 147.600 ;
        RECT 303.600 146.000 304.600 146.800 ;
        RECT 307.000 146.200 310.600 146.600 ;
        RECT 311.600 146.200 312.200 147.600 ;
        RECT 306.800 146.000 310.800 146.200 ;
        RECT 303.600 142.200 304.400 146.000 ;
        RECT 306.800 142.200 307.600 146.000 ;
        RECT 310.000 142.200 310.800 146.000 ;
        RECT 311.600 142.200 312.400 146.200 ;
        RECT 313.200 142.200 314.000 148.200 ;
        RECT 315.600 146.800 318.600 147.600 ;
        RECT 317.800 146.200 318.600 146.800 ;
        RECT 323.800 146.200 324.600 148.600 ;
        RECT 326.000 146.800 326.800 148.400 ;
        RECT 331.200 147.800 332.000 148.000 ;
        RECT 327.600 147.200 332.000 147.800 ;
        RECT 327.600 147.000 328.400 147.200 ;
        RECT 334.000 146.400 334.800 149.200 ;
        RECT 339.800 148.600 343.600 149.400 ;
        RECT 339.800 147.400 340.600 148.600 ;
        RECT 344.200 148.000 344.800 150.000 ;
        RECT 327.600 146.200 328.400 146.400 ;
        RECT 317.800 145.400 320.400 146.200 ;
        RECT 323.800 145.600 328.400 146.200 ;
        RECT 329.200 145.600 330.800 146.400 ;
        RECT 333.800 145.600 334.800 146.400 ;
        RECT 338.800 146.800 340.600 147.400 ;
        RECT 343.600 147.400 344.800 148.000 ;
        RECT 338.800 146.200 339.600 146.800 ;
        RECT 319.600 142.200 320.400 145.400 ;
        RECT 337.200 145.400 339.600 146.200 ;
        RECT 321.200 142.200 322.000 145.000 ;
        RECT 322.800 142.200 323.600 145.000 ;
        RECT 324.400 142.200 325.200 145.000 ;
        RECT 327.600 142.200 328.400 145.000 ;
        RECT 330.800 142.200 331.600 145.000 ;
        RECT 332.400 142.200 333.200 145.000 ;
        RECT 334.000 142.200 334.800 145.000 ;
        RECT 335.600 142.200 336.400 145.000 ;
        RECT 337.200 142.200 338.000 145.400 ;
        RECT 343.600 142.200 344.400 147.400 ;
        RECT 345.400 146.800 346.200 151.200 ;
        RECT 345.200 146.000 346.200 146.800 ;
        RECT 349.800 151.200 350.800 152.000 ;
        RECT 351.400 154.600 354.000 155.200 ;
        RECT 351.400 153.000 352.000 154.600 ;
        RECT 356.400 154.400 357.200 159.800 ;
        RECT 359.600 157.000 360.400 159.800 ;
        RECT 361.200 157.000 362.000 159.800 ;
        RECT 362.800 157.000 363.600 159.800 ;
        RECT 357.800 154.400 362.000 155.200 ;
        RECT 354.600 153.600 357.200 154.400 ;
        RECT 364.400 153.600 365.200 159.800 ;
        RECT 367.600 155.000 368.400 159.800 ;
        RECT 370.800 155.000 371.600 159.800 ;
        RECT 372.400 157.000 373.200 159.800 ;
        RECT 374.000 157.000 374.800 159.800 ;
        RECT 377.200 155.200 378.000 159.800 ;
        RECT 380.400 156.400 381.200 159.800 ;
        RECT 385.200 156.400 386.000 159.800 ;
        RECT 380.400 155.800 381.400 156.400 ;
        RECT 380.800 155.200 381.400 155.800 ;
        RECT 385.000 155.800 386.000 156.400 ;
        RECT 385.000 155.200 385.600 155.800 ;
        RECT 388.400 155.200 389.200 159.800 ;
        RECT 391.600 157.000 392.400 159.800 ;
        RECT 393.200 157.000 394.000 159.800 ;
        RECT 376.000 154.400 380.200 155.200 ;
        RECT 380.800 154.600 382.800 155.200 ;
        RECT 367.600 153.600 370.200 154.400 ;
        RECT 370.800 153.800 376.600 154.400 ;
        RECT 379.600 154.000 380.200 154.400 ;
        RECT 359.600 153.000 360.400 153.200 ;
        RECT 351.400 152.400 360.400 153.000 ;
        RECT 362.800 153.000 363.600 153.200 ;
        RECT 370.800 153.000 371.400 153.800 ;
        RECT 377.200 153.200 378.600 153.800 ;
        RECT 379.600 153.200 381.200 154.000 ;
        RECT 362.800 152.400 371.400 153.000 ;
        RECT 372.400 153.000 378.600 153.200 ;
        RECT 372.400 152.600 377.800 153.000 ;
        RECT 372.400 152.400 373.200 152.600 ;
        RECT 349.800 146.800 350.600 151.200 ;
        RECT 351.400 150.600 352.000 152.400 ;
        RECT 351.200 150.000 352.000 150.600 ;
        RECT 358.000 150.000 381.400 150.600 ;
        RECT 351.200 148.000 351.800 150.000 ;
        RECT 358.000 149.400 358.800 150.000 ;
        RECT 375.600 149.600 376.400 150.000 ;
        RECT 380.400 149.800 381.400 150.000 ;
        RECT 380.400 149.600 381.200 149.800 ;
        RECT 352.400 148.600 356.200 149.400 ;
        RECT 351.200 147.400 352.400 148.000 ;
        RECT 346.800 146.300 347.600 146.400 ;
        RECT 349.800 146.300 350.800 146.800 ;
        RECT 345.200 142.200 346.000 146.000 ;
        RECT 346.800 145.700 350.800 146.300 ;
        RECT 346.800 145.600 347.600 145.700 ;
        RECT 350.000 142.200 350.800 145.700 ;
        RECT 351.600 142.200 352.400 147.400 ;
        RECT 355.400 147.400 356.200 148.600 ;
        RECT 355.400 146.800 357.200 147.400 ;
        RECT 356.400 146.200 357.200 146.800 ;
        RECT 361.200 146.400 362.000 149.200 ;
        RECT 364.400 148.600 367.600 149.400 ;
        RECT 371.400 148.600 373.400 149.400 ;
        RECT 382.000 149.000 382.800 154.600 ;
        RECT 364.000 147.800 364.800 148.000 ;
        RECT 364.000 147.200 368.400 147.800 ;
        RECT 367.600 147.000 368.400 147.200 ;
        RECT 369.200 146.800 370.000 148.400 ;
        RECT 356.400 145.400 358.800 146.200 ;
        RECT 361.200 145.600 362.200 146.400 ;
        RECT 365.200 145.600 366.800 146.400 ;
        RECT 367.600 146.200 368.400 146.400 ;
        RECT 371.400 146.200 372.200 148.600 ;
        RECT 374.000 148.200 382.800 149.000 ;
        RECT 377.400 146.800 380.400 147.600 ;
        RECT 377.400 146.200 378.200 146.800 ;
        RECT 367.600 145.600 372.200 146.200 ;
        RECT 358.000 142.200 358.800 145.400 ;
        RECT 375.600 145.400 378.200 146.200 ;
        RECT 359.600 142.200 360.400 145.000 ;
        RECT 361.200 142.200 362.000 145.000 ;
        RECT 362.800 142.200 363.600 145.000 ;
        RECT 364.400 142.200 365.200 145.000 ;
        RECT 367.600 142.200 368.400 145.000 ;
        RECT 370.800 142.200 371.600 145.000 ;
        RECT 372.400 142.200 373.200 145.000 ;
        RECT 374.000 142.200 374.800 145.000 ;
        RECT 375.600 142.200 376.400 145.400 ;
        RECT 382.000 142.200 382.800 148.200 ;
        RECT 383.600 154.600 385.600 155.200 ;
        RECT 383.600 149.000 384.400 154.600 ;
        RECT 386.200 154.400 390.400 155.200 ;
        RECT 394.800 155.000 395.600 159.800 ;
        RECT 398.000 155.000 398.800 159.800 ;
        RECT 386.200 154.000 386.800 154.400 ;
        RECT 385.200 153.200 386.800 154.000 ;
        RECT 389.800 153.800 395.600 154.400 ;
        RECT 387.800 153.200 389.200 153.800 ;
        RECT 387.800 153.000 394.000 153.200 ;
        RECT 388.600 152.600 394.000 153.000 ;
        RECT 393.200 152.400 394.000 152.600 ;
        RECT 395.000 153.000 395.600 153.800 ;
        RECT 396.200 153.600 398.800 154.400 ;
        RECT 401.200 153.600 402.000 159.800 ;
        RECT 402.800 157.000 403.600 159.800 ;
        RECT 404.400 157.000 405.200 159.800 ;
        RECT 406.000 157.000 406.800 159.800 ;
        RECT 404.400 154.400 408.600 155.200 ;
        RECT 409.200 154.400 410.000 159.800 ;
        RECT 412.400 155.200 413.200 159.800 ;
        RECT 412.400 154.600 415.000 155.200 ;
        RECT 409.200 153.600 411.800 154.400 ;
        RECT 402.800 153.000 403.600 153.200 ;
        RECT 395.000 152.400 403.600 153.000 ;
        RECT 406.000 153.000 406.800 153.200 ;
        RECT 414.400 153.000 415.000 154.600 ;
        RECT 406.000 152.400 415.000 153.000 ;
        RECT 414.400 150.600 415.000 152.400 ;
        RECT 415.600 152.000 416.400 159.800 ;
        RECT 422.000 158.300 422.800 158.400 ;
        RECT 423.600 158.300 424.400 159.800 ;
        RECT 422.000 157.700 424.400 158.300 ;
        RECT 422.000 157.600 422.800 157.700 ;
        RECT 415.600 151.200 416.600 152.000 ;
        RECT 385.000 150.000 408.400 150.600 ;
        RECT 414.400 150.000 415.200 150.600 ;
        RECT 385.000 149.800 385.800 150.000 ;
        RECT 386.800 149.600 387.600 150.000 ;
        RECT 390.000 149.600 390.800 150.000 ;
        RECT 407.600 149.400 408.400 150.000 ;
        RECT 383.600 148.200 392.400 149.000 ;
        RECT 393.000 148.600 395.000 149.400 ;
        RECT 398.800 148.600 402.000 149.400 ;
        RECT 383.600 142.200 384.400 148.200 ;
        RECT 386.000 146.800 389.000 147.600 ;
        RECT 388.200 146.200 389.000 146.800 ;
        RECT 394.200 146.200 395.000 148.600 ;
        RECT 396.400 146.800 397.200 148.400 ;
        RECT 401.600 147.800 402.400 148.000 ;
        RECT 398.000 147.200 402.400 147.800 ;
        RECT 398.000 147.000 398.800 147.200 ;
        RECT 404.400 146.400 405.200 149.200 ;
        RECT 410.200 148.600 414.000 149.400 ;
        RECT 410.200 147.400 411.000 148.600 ;
        RECT 414.600 148.000 415.200 150.000 ;
        RECT 398.000 146.200 398.800 146.400 ;
        RECT 388.200 145.400 390.800 146.200 ;
        RECT 394.200 145.600 398.800 146.200 ;
        RECT 399.600 145.600 401.200 146.400 ;
        RECT 404.200 145.600 405.200 146.400 ;
        RECT 409.200 146.800 411.000 147.400 ;
        RECT 414.000 147.400 415.200 148.000 ;
        RECT 409.200 146.200 410.000 146.800 ;
        RECT 390.000 142.200 390.800 145.400 ;
        RECT 407.600 145.400 410.000 146.200 ;
        RECT 391.600 142.200 392.400 145.000 ;
        RECT 393.200 142.200 394.000 145.000 ;
        RECT 394.800 142.200 395.600 145.000 ;
        RECT 398.000 142.200 398.800 145.000 ;
        RECT 401.200 142.200 402.000 145.000 ;
        RECT 402.800 142.200 403.600 145.000 ;
        RECT 404.400 142.200 405.200 145.000 ;
        RECT 406.000 142.200 406.800 145.000 ;
        RECT 407.600 142.200 408.400 145.400 ;
        RECT 414.000 142.200 414.800 147.400 ;
        RECT 415.800 146.800 416.600 151.200 ;
        RECT 415.600 146.000 416.600 146.800 ;
        RECT 415.600 142.200 416.400 146.000 ;
        RECT 423.600 142.200 424.400 157.700 ;
        RECT 429.400 152.400 430.200 159.800 ;
        RECT 430.800 153.600 431.600 154.400 ;
        RECT 431.000 152.400 431.600 153.600 ;
        RECT 429.400 151.800 430.400 152.400 ;
        RECT 431.000 151.800 432.400 152.400 ;
        RECT 428.400 148.800 429.200 150.400 ;
        RECT 429.800 148.400 430.400 151.800 ;
        RECT 431.600 151.600 432.400 151.800 ;
        RECT 426.800 148.200 427.600 148.400 ;
        RECT 429.800 148.300 432.400 148.400 ;
        RECT 433.200 148.300 434.000 148.400 ;
        RECT 426.800 147.600 428.400 148.200 ;
        RECT 429.800 147.700 434.000 148.300 ;
        RECT 429.800 147.600 432.400 147.700 ;
        RECT 427.600 147.200 428.400 147.600 ;
        RECT 425.200 144.800 426.000 146.400 ;
        RECT 427.000 146.200 430.600 146.600 ;
        RECT 431.600 146.200 432.200 147.600 ;
        RECT 433.200 146.800 434.000 147.700 ;
        RECT 434.800 146.200 435.600 159.800 ;
        RECT 439.600 156.400 440.400 159.800 ;
        RECT 439.400 155.800 440.400 156.400 ;
        RECT 439.400 155.200 440.000 155.800 ;
        RECT 442.800 155.200 443.600 159.800 ;
        RECT 446.000 157.000 446.800 159.800 ;
        RECT 447.600 157.000 448.400 159.800 ;
        RECT 438.000 154.600 440.000 155.200 ;
        RECT 436.400 151.600 437.200 153.200 ;
        RECT 438.000 149.000 438.800 154.600 ;
        RECT 440.600 154.400 444.800 155.200 ;
        RECT 449.200 155.000 450.000 159.800 ;
        RECT 452.400 155.000 453.200 159.800 ;
        RECT 440.600 154.000 441.200 154.400 ;
        RECT 439.600 153.200 441.200 154.000 ;
        RECT 444.200 153.800 450.000 154.400 ;
        RECT 442.200 153.200 443.600 153.800 ;
        RECT 442.200 153.000 448.400 153.200 ;
        RECT 443.000 152.600 448.400 153.000 ;
        RECT 447.600 152.400 448.400 152.600 ;
        RECT 449.400 153.000 450.000 153.800 ;
        RECT 450.600 153.600 453.200 154.400 ;
        RECT 455.600 153.600 456.400 159.800 ;
        RECT 457.200 157.000 458.000 159.800 ;
        RECT 458.800 157.000 459.600 159.800 ;
        RECT 460.400 157.000 461.200 159.800 ;
        RECT 458.800 154.400 463.000 155.200 ;
        RECT 463.600 154.400 464.400 159.800 ;
        RECT 466.800 155.200 467.600 159.800 ;
        RECT 466.800 154.600 469.400 155.200 ;
        RECT 463.600 153.600 466.200 154.400 ;
        RECT 457.200 153.000 458.000 153.200 ;
        RECT 449.400 152.400 458.000 153.000 ;
        RECT 460.400 153.000 461.200 153.200 ;
        RECT 468.800 153.000 469.400 154.600 ;
        RECT 460.400 152.400 469.400 153.000 ;
        RECT 468.800 150.600 469.400 152.400 ;
        RECT 470.000 152.000 470.800 159.800 ;
        RECT 470.000 151.200 471.000 152.000 ;
        RECT 439.400 150.000 462.800 150.600 ;
        RECT 468.800 150.000 469.600 150.600 ;
        RECT 439.400 149.800 440.200 150.000 ;
        RECT 441.200 149.600 442.000 150.000 ;
        RECT 444.400 149.600 445.200 150.000 ;
        RECT 462.000 149.400 462.800 150.000 ;
        RECT 438.000 148.200 446.800 149.000 ;
        RECT 447.400 148.600 449.400 149.400 ;
        RECT 453.200 148.600 456.400 149.400 ;
        RECT 426.800 146.000 430.800 146.200 ;
        RECT 426.800 142.200 427.600 146.000 ;
        RECT 430.000 142.200 430.800 146.000 ;
        RECT 431.600 142.200 432.400 146.200 ;
        RECT 434.800 145.600 436.600 146.200 ;
        RECT 435.800 144.400 436.600 145.600 ;
        RECT 434.800 143.600 436.600 144.400 ;
        RECT 435.800 142.200 436.600 143.600 ;
        RECT 438.000 142.200 438.800 148.200 ;
        RECT 440.400 146.800 443.400 147.600 ;
        RECT 442.600 146.200 443.400 146.800 ;
        RECT 448.600 146.200 449.400 148.600 ;
        RECT 450.800 146.800 451.600 148.400 ;
        RECT 456.000 147.800 456.800 148.000 ;
        RECT 452.400 147.200 456.800 147.800 ;
        RECT 452.400 147.000 453.200 147.200 ;
        RECT 458.800 146.400 459.600 149.200 ;
        RECT 464.600 148.600 468.400 149.400 ;
        RECT 464.600 147.400 465.400 148.600 ;
        RECT 469.000 148.000 469.600 150.000 ;
        RECT 452.400 146.200 453.200 146.400 ;
        RECT 442.600 145.400 445.200 146.200 ;
        RECT 448.600 145.600 453.200 146.200 ;
        RECT 454.000 145.600 455.600 146.400 ;
        RECT 458.600 145.600 459.600 146.400 ;
        RECT 463.600 146.800 465.400 147.400 ;
        RECT 468.400 147.400 469.600 148.000 ;
        RECT 463.600 146.200 464.400 146.800 ;
        RECT 444.400 142.200 445.200 145.400 ;
        RECT 462.000 145.400 464.400 146.200 ;
        RECT 446.000 142.200 446.800 145.000 ;
        RECT 447.600 142.200 448.400 145.000 ;
        RECT 449.200 142.200 450.000 145.000 ;
        RECT 452.400 142.200 453.200 145.000 ;
        RECT 455.600 142.200 456.400 145.000 ;
        RECT 457.200 142.200 458.000 145.000 ;
        RECT 458.800 142.200 459.600 145.000 ;
        RECT 460.400 142.200 461.200 145.000 ;
        RECT 462.000 142.200 462.800 145.400 ;
        RECT 468.400 142.200 469.200 147.400 ;
        RECT 470.200 146.800 471.000 151.200 ;
        RECT 470.000 146.000 471.000 146.800 ;
        RECT 470.000 142.200 470.800 146.000 ;
        RECT 473.200 142.200 474.000 159.800 ;
        RECT 478.000 156.400 478.800 159.800 ;
        RECT 477.800 155.800 478.800 156.400 ;
        RECT 477.800 155.200 478.400 155.800 ;
        RECT 481.200 155.200 482.000 159.800 ;
        RECT 484.400 157.000 485.200 159.800 ;
        RECT 486.000 157.000 486.800 159.800 ;
        RECT 476.400 154.600 478.400 155.200 ;
        RECT 476.400 149.000 477.200 154.600 ;
        RECT 479.000 154.400 483.200 155.200 ;
        RECT 487.600 155.000 488.400 159.800 ;
        RECT 490.800 155.000 491.600 159.800 ;
        RECT 479.000 154.000 479.600 154.400 ;
        RECT 478.000 153.200 479.600 154.000 ;
        RECT 482.600 153.800 488.400 154.400 ;
        RECT 480.600 153.200 482.000 153.800 ;
        RECT 480.600 153.000 486.800 153.200 ;
        RECT 481.400 152.600 486.800 153.000 ;
        RECT 486.000 152.400 486.800 152.600 ;
        RECT 487.800 153.000 488.400 153.800 ;
        RECT 489.000 153.600 491.600 154.400 ;
        RECT 494.000 153.600 494.800 159.800 ;
        RECT 495.600 157.000 496.400 159.800 ;
        RECT 497.200 157.000 498.000 159.800 ;
        RECT 498.800 157.000 499.600 159.800 ;
        RECT 497.200 154.400 501.400 155.200 ;
        RECT 502.000 154.400 502.800 159.800 ;
        RECT 505.200 155.200 506.000 159.800 ;
        RECT 505.200 154.600 507.800 155.200 ;
        RECT 502.000 153.600 504.600 154.400 ;
        RECT 495.600 153.000 496.400 153.200 ;
        RECT 487.800 152.400 496.400 153.000 ;
        RECT 498.800 153.000 499.600 153.200 ;
        RECT 507.200 153.000 507.800 154.600 ;
        RECT 498.800 152.400 507.800 153.000 ;
        RECT 507.200 150.600 507.800 152.400 ;
        RECT 508.400 152.000 509.200 159.800 ;
        RECT 508.400 151.200 509.400 152.000 ;
        RECT 477.800 150.000 501.200 150.600 ;
        RECT 507.200 150.000 508.000 150.600 ;
        RECT 477.800 149.800 478.600 150.000 ;
        RECT 479.600 149.600 480.400 150.000 ;
        RECT 482.800 149.600 483.600 150.000 ;
        RECT 500.400 149.400 501.200 150.000 ;
        RECT 476.400 148.200 485.200 149.000 ;
        RECT 485.800 148.600 487.800 149.400 ;
        RECT 491.600 148.600 494.800 149.400 ;
        RECT 474.800 144.800 475.600 146.400 ;
        RECT 476.400 142.200 477.200 148.200 ;
        RECT 478.800 146.800 481.800 147.600 ;
        RECT 481.000 146.200 481.800 146.800 ;
        RECT 487.000 146.200 487.800 148.600 ;
        RECT 489.200 146.800 490.000 148.400 ;
        RECT 494.400 147.800 495.200 148.000 ;
        RECT 490.800 147.200 495.200 147.800 ;
        RECT 490.800 147.000 491.600 147.200 ;
        RECT 497.200 146.400 498.000 149.200 ;
        RECT 503.000 148.600 506.800 149.400 ;
        RECT 503.000 147.400 503.800 148.600 ;
        RECT 507.400 148.000 508.000 150.000 ;
        RECT 490.800 146.200 491.600 146.400 ;
        RECT 481.000 145.400 483.600 146.200 ;
        RECT 487.000 145.600 491.600 146.200 ;
        RECT 492.400 145.600 494.000 146.400 ;
        RECT 497.000 145.600 498.000 146.400 ;
        RECT 502.000 146.800 503.800 147.400 ;
        RECT 506.800 147.400 508.000 148.000 ;
        RECT 502.000 146.200 502.800 146.800 ;
        RECT 482.800 142.200 483.600 145.400 ;
        RECT 500.400 145.400 502.800 146.200 ;
        RECT 484.400 142.200 485.200 145.000 ;
        RECT 486.000 142.200 486.800 145.000 ;
        RECT 487.600 142.200 488.400 145.000 ;
        RECT 490.800 142.200 491.600 145.000 ;
        RECT 494.000 142.200 494.800 145.000 ;
        RECT 495.600 142.200 496.400 145.000 ;
        RECT 497.200 142.200 498.000 145.000 ;
        RECT 498.800 142.200 499.600 145.000 ;
        RECT 500.400 142.200 501.200 145.400 ;
        RECT 506.800 142.200 507.600 147.400 ;
        RECT 508.600 146.800 509.400 151.200 ;
        RECT 508.400 146.000 509.400 146.800 ;
        RECT 513.200 150.300 514.000 159.800 ;
        RECT 517.000 158.400 517.800 159.800 ;
        RECT 517.000 157.600 518.800 158.400 ;
        RECT 515.600 153.600 516.400 154.400 ;
        RECT 515.600 152.400 516.200 153.600 ;
        RECT 517.000 152.400 517.800 157.600 ;
        RECT 514.800 151.800 516.200 152.400 ;
        RECT 516.800 151.800 517.800 152.400 ;
        RECT 523.800 152.400 524.600 159.800 ;
        RECT 525.200 153.600 526.000 154.400 ;
        RECT 525.400 152.400 526.000 153.600 ;
        RECT 528.400 153.600 529.200 154.400 ;
        RECT 528.400 152.400 529.000 153.600 ;
        RECT 529.800 152.400 530.600 159.800 ;
        RECT 536.600 152.600 537.400 159.800 ;
        RECT 523.800 151.800 524.800 152.400 ;
        RECT 525.400 151.800 526.800 152.400 ;
        RECT 514.800 151.600 515.600 151.800 ;
        RECT 514.800 150.300 515.600 150.400 ;
        RECT 513.200 149.700 515.600 150.300 ;
        RECT 510.000 146.300 510.800 146.400 ;
        RECT 511.600 146.300 512.400 146.400 ;
        RECT 508.400 142.200 509.200 146.000 ;
        RECT 510.000 145.700 512.400 146.300 ;
        RECT 510.000 145.600 510.800 145.700 ;
        RECT 511.600 144.800 512.400 145.700 ;
        RECT 513.200 142.200 514.000 149.700 ;
        RECT 514.800 149.600 515.600 149.700 ;
        RECT 516.800 148.400 517.400 151.800 ;
        RECT 518.000 148.800 518.800 150.400 ;
        RECT 522.800 148.800 523.600 150.400 ;
        RECT 524.200 148.400 524.800 151.800 ;
        RECT 526.000 151.600 526.800 151.800 ;
        RECT 527.600 151.800 529.000 152.400 ;
        RECT 529.600 151.800 530.600 152.400 ;
        RECT 535.600 151.800 537.400 152.600 ;
        RECT 527.600 151.600 528.400 151.800 ;
        RECT 526.100 150.300 526.700 151.600 ;
        RECT 529.600 150.300 530.200 151.800 ;
        RECT 526.100 149.700 530.200 150.300 ;
        RECT 529.600 148.400 530.200 149.700 ;
        RECT 530.800 148.800 531.600 150.400 ;
        RECT 535.800 148.400 536.400 151.800 ;
        RECT 537.200 150.300 538.000 151.200 ;
        RECT 538.800 150.300 539.600 150.400 ;
        RECT 537.200 149.700 539.600 150.300 ;
        RECT 537.200 149.600 538.000 149.700 ;
        RECT 538.800 149.600 539.600 149.700 ;
        RECT 514.800 147.600 517.400 148.400 ;
        RECT 519.600 148.200 520.400 148.400 ;
        RECT 518.800 147.600 520.400 148.200 ;
        RECT 521.200 148.200 522.000 148.400 ;
        RECT 521.200 147.600 522.800 148.200 ;
        RECT 524.200 147.600 526.800 148.400 ;
        RECT 527.600 147.600 530.200 148.400 ;
        RECT 532.400 148.200 533.200 148.400 ;
        RECT 531.600 147.600 533.200 148.200 ;
        RECT 535.600 147.600 536.400 148.400 ;
        RECT 515.000 146.200 515.600 147.600 ;
        RECT 518.800 147.200 519.600 147.600 ;
        RECT 522.000 147.200 522.800 147.600 ;
        RECT 516.600 146.200 520.200 146.600 ;
        RECT 521.400 146.200 525.000 146.600 ;
        RECT 526.000 146.200 526.600 147.600 ;
        RECT 527.800 146.200 528.400 147.600 ;
        RECT 531.600 147.200 532.400 147.600 ;
        RECT 529.400 146.200 533.000 146.600 ;
        RECT 514.800 142.200 515.600 146.200 ;
        RECT 516.400 146.000 520.400 146.200 ;
        RECT 516.400 142.200 517.200 146.000 ;
        RECT 519.600 142.200 520.400 146.000 ;
        RECT 521.200 146.000 525.200 146.200 ;
        RECT 521.200 142.200 522.000 146.000 ;
        RECT 524.400 142.200 525.200 146.000 ;
        RECT 526.000 142.200 526.800 146.200 ;
        RECT 527.600 142.200 528.400 146.200 ;
        RECT 529.200 146.000 533.200 146.200 ;
        RECT 529.200 142.200 530.000 146.000 ;
        RECT 532.400 142.200 533.200 146.000 ;
        RECT 534.000 144.800 534.800 146.400 ;
        RECT 535.800 144.400 536.400 147.600 ;
        RECT 538.800 144.800 539.600 146.400 ;
        RECT 535.600 142.200 536.400 144.400 ;
        RECT 540.400 142.200 541.200 159.800 ;
        RECT 544.600 152.400 545.400 159.800 ;
        RECT 546.000 153.600 546.800 154.400 ;
        RECT 546.200 152.400 546.800 153.600 ;
        RECT 544.600 151.800 545.600 152.400 ;
        RECT 546.200 151.800 547.600 152.400 ;
        RECT 542.000 150.300 542.800 150.400 ;
        RECT 543.600 150.300 544.400 150.400 ;
        RECT 542.000 149.700 544.400 150.300 ;
        RECT 542.000 149.600 542.800 149.700 ;
        RECT 543.600 148.800 544.400 149.700 ;
        RECT 545.000 148.400 545.600 151.800 ;
        RECT 546.800 151.600 547.600 151.800 ;
        RECT 548.400 150.300 549.200 159.800 ;
        RECT 551.600 151.600 552.400 153.200 ;
        RECT 551.700 150.300 552.300 151.600 ;
        RECT 548.400 149.700 552.300 150.300 ;
        RECT 542.000 148.200 542.800 148.400 ;
        RECT 542.000 147.600 543.600 148.200 ;
        RECT 545.000 147.600 547.600 148.400 ;
        RECT 542.800 147.200 543.600 147.600 ;
        RECT 542.200 146.200 545.800 146.600 ;
        RECT 546.800 146.200 547.400 147.600 ;
        RECT 542.000 146.000 546.000 146.200 ;
        RECT 542.000 142.200 542.800 146.000 ;
        RECT 545.200 142.200 546.000 146.000 ;
        RECT 546.800 142.200 547.600 146.200 ;
        RECT 548.400 142.200 549.200 149.700 ;
        RECT 550.000 146.800 550.800 148.400 ;
        RECT 553.200 146.200 554.000 159.800 ;
        RECT 558.000 152.800 558.800 159.800 ;
        RECT 557.800 151.800 558.800 152.800 ;
        RECT 561.200 152.400 562.000 159.800 ;
        RECT 563.600 153.600 564.400 154.400 ;
        RECT 563.600 152.400 564.200 153.600 ;
        RECT 565.000 152.400 565.800 159.800 ;
        RECT 574.800 153.600 575.600 154.400 ;
        RECT 574.800 152.400 575.400 153.600 ;
        RECT 576.200 152.400 577.000 159.800 ;
        RECT 559.400 151.800 562.000 152.400 ;
        RECT 562.800 151.800 564.200 152.400 ;
        RECT 564.800 151.800 565.800 152.400 ;
        RECT 574.000 151.800 575.400 152.400 ;
        RECT 576.000 151.800 577.000 152.400 ;
        RECT 583.000 152.400 583.800 159.800 ;
        RECT 584.400 153.600 585.200 154.400 ;
        RECT 584.600 152.400 585.200 153.600 ;
        RECT 587.600 153.600 588.400 154.400 ;
        RECT 587.600 152.400 588.200 153.600 ;
        RECT 589.000 152.400 589.800 159.800 ;
        RECT 583.000 151.800 584.000 152.400 ;
        RECT 584.600 151.800 586.000 152.400 ;
        RECT 557.800 148.400 558.400 151.800 ;
        RECT 559.400 149.800 560.000 151.800 ;
        RECT 562.800 151.600 563.600 151.800 ;
        RECT 559.000 149.000 560.000 149.800 ;
        RECT 554.800 148.300 555.600 148.400 ;
        RECT 556.400 148.300 557.200 148.400 ;
        RECT 554.800 147.700 557.200 148.300 ;
        RECT 554.800 146.800 555.600 147.700 ;
        RECT 556.400 147.600 557.200 147.700 ;
        RECT 557.800 147.600 558.800 148.400 ;
        RECT 552.200 145.600 554.000 146.200 ;
        RECT 557.800 146.200 558.400 147.600 ;
        RECT 559.400 147.400 560.000 149.000 ;
        RECT 561.000 149.600 562.000 150.400 ;
        RECT 562.800 150.300 563.600 150.400 ;
        RECT 564.800 150.300 565.400 151.800 ;
        RECT 574.000 151.600 574.800 151.800 ;
        RECT 562.800 149.700 565.400 150.300 ;
        RECT 562.800 149.600 563.600 149.700 ;
        RECT 561.000 148.800 561.800 149.600 ;
        RECT 564.800 148.400 565.400 149.700 ;
        RECT 566.000 150.300 566.800 150.400 ;
        RECT 576.000 150.300 576.600 151.800 ;
        RECT 566.000 149.700 576.600 150.300 ;
        RECT 566.000 148.800 566.800 149.700 ;
        RECT 576.000 148.400 576.600 149.700 ;
        RECT 577.200 148.800 578.000 150.400 ;
        RECT 582.000 148.800 582.800 150.400 ;
        RECT 583.400 150.300 584.000 151.800 ;
        RECT 585.200 151.600 586.000 151.800 ;
        RECT 586.800 151.800 588.200 152.400 ;
        RECT 588.800 151.800 589.800 152.400 ;
        RECT 593.200 155.000 594.000 159.000 ;
        RECT 586.800 151.600 587.600 151.800 ;
        RECT 586.900 150.300 587.500 151.600 ;
        RECT 583.400 149.700 587.500 150.300 ;
        RECT 583.400 148.400 584.000 149.700 ;
        RECT 588.800 148.400 589.400 151.800 ;
        RECT 593.200 151.600 593.800 155.000 ;
        RECT 597.400 152.800 598.200 159.800 ;
        RECT 597.400 152.200 599.000 152.800 ;
        RECT 593.200 151.000 597.000 151.600 ;
        RECT 590.000 148.800 590.800 150.400 ;
        RECT 593.200 148.800 594.000 150.400 ;
        RECT 594.800 148.800 595.600 150.400 ;
        RECT 596.400 149.000 597.000 151.000 ;
        RECT 562.800 147.600 565.400 148.400 ;
        RECT 567.600 148.200 568.400 148.400 ;
        RECT 566.800 147.600 568.400 148.200 ;
        RECT 574.000 147.600 576.600 148.400 ;
        RECT 578.800 148.200 579.600 148.400 ;
        RECT 578.000 147.600 579.600 148.200 ;
        RECT 580.400 148.200 581.200 148.400 ;
        RECT 580.400 147.600 582.000 148.200 ;
        RECT 583.400 147.600 586.000 148.400 ;
        RECT 586.800 147.600 589.400 148.400 ;
        RECT 591.600 148.200 592.400 148.400 ;
        RECT 590.800 147.600 592.400 148.200 ;
        RECT 596.400 148.200 597.800 149.000 ;
        RECT 598.400 148.400 599.000 152.200 ;
        RECT 602.800 152.400 603.600 159.800 ;
        RECT 606.000 152.800 606.800 159.800 ;
        RECT 602.800 151.800 605.400 152.400 ;
        RECT 606.000 151.800 607.000 152.800 ;
        RECT 611.800 152.400 612.600 159.800 ;
        RECT 613.200 153.600 614.000 154.400 ;
        RECT 613.400 152.400 614.000 153.600 ;
        RECT 617.200 152.800 618.000 159.800 ;
        RECT 611.800 151.800 612.800 152.400 ;
        RECT 613.400 151.800 614.800 152.400 ;
        RECT 599.600 149.600 600.400 151.200 ;
        RECT 601.200 150.300 602.000 150.400 ;
        RECT 602.800 150.300 603.800 150.400 ;
        RECT 601.200 149.700 603.800 150.300 ;
        RECT 601.200 149.600 602.000 149.700 ;
        RECT 602.800 149.600 603.800 149.700 ;
        RECT 603.000 148.800 603.800 149.600 ;
        RECT 604.800 149.800 605.400 151.800 ;
        RECT 604.800 149.000 605.800 149.800 ;
        RECT 596.400 147.800 597.400 148.200 ;
        RECT 559.400 146.800 562.000 147.400 ;
        RECT 557.800 145.600 558.800 146.200 ;
        RECT 552.200 144.400 553.000 145.600 ;
        RECT 551.600 143.600 553.000 144.400 ;
        RECT 552.200 142.200 553.000 143.600 ;
        RECT 558.000 142.200 558.800 145.600 ;
        RECT 561.200 142.200 562.000 146.800 ;
        RECT 563.000 146.200 563.600 147.600 ;
        RECT 566.800 147.200 567.600 147.600 ;
        RECT 564.600 146.200 568.200 146.600 ;
        RECT 574.200 146.200 574.800 147.600 ;
        RECT 578.000 147.200 578.800 147.600 ;
        RECT 581.200 147.200 582.000 147.600 ;
        RECT 575.800 146.200 579.400 146.600 ;
        RECT 580.600 146.200 584.200 146.600 ;
        RECT 585.200 146.200 585.800 147.600 ;
        RECT 587.000 146.200 587.600 147.600 ;
        RECT 590.800 147.200 591.600 147.600 ;
        RECT 593.200 147.200 597.400 147.800 ;
        RECT 598.400 147.600 600.400 148.400 ;
        RECT 588.600 146.200 592.200 146.600 ;
        RECT 562.800 142.200 563.600 146.200 ;
        RECT 564.400 146.000 568.400 146.200 ;
        RECT 564.400 142.200 565.200 146.000 ;
        RECT 567.600 142.200 568.400 146.000 ;
        RECT 574.000 142.200 574.800 146.200 ;
        RECT 575.600 146.000 579.600 146.200 ;
        RECT 575.600 142.200 576.400 146.000 ;
        RECT 578.800 142.200 579.600 146.000 ;
        RECT 580.400 146.000 584.400 146.200 ;
        RECT 580.400 142.200 581.200 146.000 ;
        RECT 583.600 142.200 584.400 146.000 ;
        RECT 585.200 142.200 586.000 146.200 ;
        RECT 586.800 142.200 587.600 146.200 ;
        RECT 588.400 146.000 592.400 146.200 ;
        RECT 588.400 142.200 589.200 146.000 ;
        RECT 591.600 142.200 592.400 146.000 ;
        RECT 593.200 145.000 593.800 147.200 ;
        RECT 598.400 147.000 599.000 147.600 ;
        RECT 604.800 147.400 605.400 149.000 ;
        RECT 606.400 148.400 607.000 151.800 ;
        RECT 610.800 148.800 611.600 150.400 ;
        RECT 612.200 148.400 612.800 151.800 ;
        RECT 614.000 151.600 614.800 151.800 ;
        RECT 617.000 151.800 618.000 152.800 ;
        RECT 620.400 152.400 621.200 159.800 ;
        RECT 622.000 155.800 622.800 159.800 ;
        RECT 622.200 155.600 622.800 155.800 ;
        RECT 625.200 155.800 626.000 159.800 ;
        RECT 625.200 155.600 625.800 155.800 ;
        RECT 622.200 155.000 625.800 155.600 ;
        RECT 622.200 154.400 622.800 155.000 ;
        RECT 622.000 153.600 622.800 154.400 ;
        RECT 622.200 152.400 622.800 153.600 ;
        RECT 623.600 152.800 624.400 154.400 ;
        RECT 628.400 152.400 629.200 159.800 ;
        RECT 631.600 152.800 632.400 159.800 ;
        RECT 618.600 151.800 621.200 152.400 ;
        RECT 617.000 148.400 617.600 151.800 ;
        RECT 618.600 149.800 619.200 151.800 ;
        RECT 622.000 151.600 622.800 152.400 ;
        RECT 618.200 149.000 619.200 149.800 ;
        RECT 606.000 147.600 607.000 148.400 ;
        RECT 609.200 148.200 610.000 148.400 ;
        RECT 609.200 147.600 610.800 148.200 ;
        RECT 612.200 147.600 614.800 148.400 ;
        RECT 617.000 147.600 618.000 148.400 ;
        RECT 598.200 146.600 599.000 147.000 ;
        RECT 597.400 146.000 599.000 146.600 ;
        RECT 602.800 146.800 605.400 147.400 ;
        RECT 593.200 143.000 594.000 145.000 ;
        RECT 597.400 144.400 598.200 146.000 ;
        RECT 596.400 143.600 598.200 144.400 ;
        RECT 597.400 143.000 598.200 143.600 ;
        RECT 602.800 142.200 603.600 146.800 ;
        RECT 606.400 146.200 607.000 147.600 ;
        RECT 610.000 147.200 610.800 147.600 ;
        RECT 609.400 146.200 613.000 146.600 ;
        RECT 614.000 146.200 614.600 147.600 ;
        RECT 617.000 146.200 617.600 147.600 ;
        RECT 618.600 147.400 619.200 149.000 ;
        RECT 620.200 149.600 621.200 150.400 ;
        RECT 620.200 148.800 621.000 149.600 ;
        RECT 622.200 148.400 622.800 151.600 ;
        RECT 626.800 150.800 627.600 152.400 ;
        RECT 628.400 151.800 631.000 152.400 ;
        RECT 631.600 151.800 632.600 152.800 ;
        RECT 634.800 152.400 635.600 159.800 ;
        RECT 638.000 152.800 638.800 159.800 ;
        RECT 634.800 151.800 637.400 152.400 ;
        RECT 638.000 151.800 639.000 152.800 ;
        RECT 624.400 149.600 626.000 150.400 ;
        RECT 628.400 149.600 629.400 150.400 ;
        RECT 628.600 148.800 629.400 149.600 ;
        RECT 630.400 149.800 631.000 151.800 ;
        RECT 630.400 149.000 631.400 149.800 ;
        RECT 622.200 148.200 623.800 148.400 ;
        RECT 622.200 147.800 624.000 148.200 ;
        RECT 618.600 146.800 621.200 147.400 ;
        RECT 606.000 145.600 607.000 146.200 ;
        RECT 609.200 146.000 613.200 146.200 ;
        RECT 606.000 142.200 606.800 145.600 ;
        RECT 609.200 142.200 610.000 146.000 ;
        RECT 612.400 142.200 613.200 146.000 ;
        RECT 614.000 142.200 614.800 146.200 ;
        RECT 617.000 145.600 618.000 146.200 ;
        RECT 617.200 142.200 618.000 145.600 ;
        RECT 620.400 142.200 621.200 146.800 ;
        RECT 623.200 142.200 624.000 147.800 ;
        RECT 630.400 147.400 631.000 149.000 ;
        RECT 632.000 148.400 632.600 151.800 ;
        RECT 634.800 149.600 635.800 150.400 ;
        RECT 635.000 148.800 635.800 149.600 ;
        RECT 636.800 149.800 637.400 151.800 ;
        RECT 636.800 149.000 637.800 149.800 ;
        RECT 631.600 147.600 632.600 148.400 ;
        RECT 628.400 146.800 631.000 147.400 ;
        RECT 628.400 142.200 629.200 146.800 ;
        RECT 632.000 146.200 632.600 147.600 ;
        RECT 636.800 147.400 637.400 149.000 ;
        RECT 638.400 148.400 639.000 151.800 ;
        RECT 638.000 147.600 639.000 148.400 ;
        RECT 631.600 145.600 632.600 146.200 ;
        RECT 634.800 146.800 637.400 147.400 ;
        RECT 631.600 142.200 632.400 145.600 ;
        RECT 634.800 142.200 635.600 146.800 ;
        RECT 638.400 146.200 639.000 147.600 ;
        RECT 638.000 145.600 639.000 146.200 ;
        RECT 638.000 142.200 638.800 145.600 ;
        RECT 641.200 142.200 642.000 159.800 ;
        RECT 644.400 155.000 645.200 159.000 ;
        RECT 644.400 151.600 645.000 155.000 ;
        RECT 648.600 152.800 649.400 159.800 ;
        RECT 654.000 155.000 654.800 159.000 ;
        RECT 648.600 152.200 650.200 152.800 ;
        RECT 644.400 151.000 648.200 151.600 ;
        RECT 644.400 148.800 645.200 150.400 ;
        RECT 646.000 148.800 646.800 150.400 ;
        RECT 647.600 149.000 648.200 151.000 ;
        RECT 647.600 148.200 649.000 149.000 ;
        RECT 649.600 148.400 650.200 152.200 ;
        RECT 654.000 151.600 654.600 155.000 ;
        RECT 658.200 152.800 659.000 159.800 ;
        RECT 658.200 152.200 659.800 152.800 ;
        RECT 650.800 149.600 651.600 151.200 ;
        RECT 654.000 151.000 657.800 151.600 ;
        RECT 654.000 148.800 654.800 150.400 ;
        RECT 655.600 148.800 656.400 150.400 ;
        RECT 657.200 149.000 657.800 151.000 ;
        RECT 649.600 148.300 651.600 148.400 ;
        RECT 652.400 148.300 653.200 148.400 ;
        RECT 647.600 147.800 648.600 148.200 ;
        RECT 644.400 147.200 648.600 147.800 ;
        RECT 649.600 147.700 653.200 148.300 ;
        RECT 657.200 148.200 658.600 149.000 ;
        RECT 659.200 148.400 659.800 152.200 ;
        RECT 666.200 152.400 667.000 159.800 ;
        RECT 667.600 153.600 668.400 154.400 ;
        RECT 667.800 152.400 668.400 153.600 ;
        RECT 666.200 151.800 667.200 152.400 ;
        RECT 667.800 151.800 669.200 152.400 ;
        RECT 660.400 149.600 661.200 151.200 ;
        RECT 665.200 150.300 666.000 150.400 ;
        RECT 662.100 149.700 666.000 150.300 ;
        RECT 659.200 148.300 661.200 148.400 ;
        RECT 662.100 148.300 662.700 149.700 ;
        RECT 665.200 148.800 666.000 149.700 ;
        RECT 666.600 150.300 667.200 151.800 ;
        RECT 668.400 151.600 669.200 151.800 ;
        RECT 670.000 151.200 670.800 159.800 ;
        RECT 674.200 155.800 675.400 159.800 ;
        RECT 678.800 155.800 679.600 159.800 ;
        RECT 683.200 156.400 684.000 159.800 ;
        RECT 683.200 155.800 685.200 156.400 ;
        RECT 674.800 155.000 675.600 155.800 ;
        RECT 679.000 155.200 679.600 155.800 ;
        RECT 678.200 154.600 681.800 155.200 ;
        RECT 684.400 155.000 685.200 155.800 ;
        RECT 678.200 154.400 679.000 154.600 ;
        RECT 681.000 154.400 681.800 154.600 ;
        RECT 674.000 153.200 675.400 154.000 ;
        RECT 674.800 152.200 675.400 153.200 ;
        RECT 677.000 153.000 679.200 153.600 ;
        RECT 677.000 152.800 677.800 153.000 ;
        RECT 674.800 151.600 677.200 152.200 ;
        RECT 670.000 150.600 674.200 151.200 ;
        RECT 668.400 150.300 669.200 150.400 ;
        RECT 666.600 149.700 669.200 150.300 ;
        RECT 666.600 148.400 667.200 149.700 ;
        RECT 668.400 149.600 669.200 149.700 ;
        RECT 657.200 147.800 658.200 148.200 ;
        RECT 649.600 147.600 651.600 147.700 ;
        RECT 652.400 147.600 653.200 147.700 ;
        RECT 642.800 144.800 643.600 146.400 ;
        RECT 644.400 145.000 645.000 147.200 ;
        RECT 649.600 147.000 650.200 147.600 ;
        RECT 649.400 146.600 650.200 147.000 ;
        RECT 648.600 146.000 650.200 146.600 ;
        RECT 654.000 147.200 658.200 147.800 ;
        RECT 659.200 147.700 662.700 148.300 ;
        RECT 663.600 148.200 664.400 148.400 ;
        RECT 659.200 147.600 661.200 147.700 ;
        RECT 663.600 147.600 665.200 148.200 ;
        RECT 666.600 147.600 669.200 148.400 ;
        RECT 644.400 143.000 645.200 145.000 ;
        RECT 648.600 143.000 649.400 146.000 ;
        RECT 654.000 145.000 654.600 147.200 ;
        RECT 659.200 147.000 659.800 147.600 ;
        RECT 664.400 147.200 665.200 147.600 ;
        RECT 659.000 146.600 659.800 147.000 ;
        RECT 658.200 146.000 659.800 146.600 ;
        RECT 663.800 146.200 667.400 146.600 ;
        RECT 668.400 146.200 669.000 147.600 ;
        RECT 670.000 147.200 670.800 150.600 ;
        RECT 673.400 150.400 674.200 150.600 ;
        RECT 676.600 150.300 677.200 151.600 ;
        RECT 678.600 151.800 679.200 153.000 ;
        RECT 679.800 153.000 680.600 153.200 ;
        RECT 684.400 153.000 685.200 153.200 ;
        RECT 679.800 152.400 685.200 153.000 ;
        RECT 678.600 151.400 683.400 151.800 ;
        RECT 687.600 151.400 688.400 159.800 ;
        RECT 678.600 151.200 688.400 151.400 ;
        RECT 682.600 151.000 688.400 151.200 ;
        RECT 682.800 150.800 688.400 151.000 ;
        RECT 678.000 150.300 678.800 150.400 ;
        RECT 671.800 149.800 672.600 150.000 ;
        RECT 671.800 149.200 675.600 149.800 ;
        RECT 676.500 149.700 678.800 150.300 ;
        RECT 674.800 149.000 675.600 149.200 ;
        RECT 676.600 148.400 677.200 149.700 ;
        RECT 678.000 149.600 678.800 149.700 ;
        RECT 679.600 150.300 680.400 150.400 ;
        RECT 681.200 150.300 682.000 150.400 ;
        RECT 679.600 150.200 682.000 150.300 ;
        RECT 679.600 149.700 686.200 150.200 ;
        RECT 679.600 149.600 680.400 149.700 ;
        RECT 681.200 149.600 686.200 149.700 ;
        RECT 685.400 149.400 686.200 149.600 ;
        RECT 683.800 148.400 684.600 148.600 ;
        RECT 676.600 147.800 687.600 148.400 ;
        RECT 677.000 147.600 677.800 147.800 ;
        RECT 670.000 146.600 673.800 147.200 ;
        RECT 663.600 146.000 667.600 146.200 ;
        RECT 654.000 143.000 654.800 145.000 ;
        RECT 658.200 143.000 659.000 146.000 ;
        RECT 663.600 142.200 664.400 146.000 ;
        RECT 666.800 142.200 667.600 146.000 ;
        RECT 668.400 142.200 669.200 146.200 ;
        RECT 670.000 142.200 670.800 146.600 ;
        RECT 673.000 146.400 673.800 146.600 ;
        RECT 682.800 146.400 683.400 147.800 ;
        RECT 686.000 147.600 687.600 147.800 ;
        RECT 681.000 145.400 681.800 145.600 ;
        RECT 674.800 144.200 675.600 145.000 ;
        RECT 679.000 144.800 681.800 145.400 ;
        RECT 682.800 144.800 683.600 146.400 ;
        RECT 679.000 144.200 679.600 144.800 ;
        RECT 684.400 144.200 685.200 145.000 ;
        RECT 674.200 143.600 675.600 144.200 ;
        RECT 674.200 142.200 675.400 143.600 ;
        RECT 678.800 142.200 679.600 144.200 ;
        RECT 683.200 143.600 685.200 144.200 ;
        RECT 683.200 142.200 684.000 143.600 ;
        RECT 687.600 142.200 688.400 147.000 ;
        RECT 1.200 135.000 2.000 139.800 ;
        RECT 5.600 138.400 6.400 139.800 ;
        RECT 4.400 137.800 6.400 138.400 ;
        RECT 10.000 137.800 10.800 139.800 ;
        RECT 14.200 138.400 15.400 139.800 ;
        RECT 14.000 137.800 15.400 138.400 ;
        RECT 4.400 137.000 5.200 137.800 ;
        RECT 10.000 137.200 10.600 137.800 ;
        RECT 6.000 136.400 6.800 137.200 ;
        RECT 7.800 136.600 10.600 137.200 ;
        RECT 14.000 137.000 14.800 137.800 ;
        RECT 7.800 136.400 8.600 136.600 ;
        RECT 2.000 134.200 3.600 134.400 ;
        RECT 6.200 134.200 6.800 136.400 ;
        RECT 15.800 135.400 16.600 135.600 ;
        RECT 18.800 135.400 19.600 139.800 ;
        RECT 20.400 135.800 21.200 139.800 ;
        RECT 22.000 136.000 22.800 139.800 ;
        RECT 25.200 136.000 26.000 139.800 ;
        RECT 22.000 135.800 26.000 136.000 ;
        RECT 26.800 135.800 27.600 139.800 ;
        RECT 28.400 136.000 29.200 139.800 ;
        RECT 31.600 136.000 32.400 139.800 ;
        RECT 28.400 135.800 32.400 136.000 ;
        RECT 15.800 134.800 19.600 135.400 ;
        RECT 11.800 134.200 12.600 134.400 ;
        RECT 2.000 133.600 13.000 134.200 ;
        RECT 5.000 133.400 5.800 133.600 ;
        RECT 3.400 132.400 4.200 132.600 ;
        RECT 12.400 132.400 13.000 133.600 ;
        RECT 14.000 132.800 14.800 133.000 ;
        RECT 3.400 131.800 8.400 132.400 ;
        RECT 7.600 131.600 8.400 131.800 ;
        RECT 12.400 131.600 13.200 132.400 ;
        RECT 14.000 132.200 17.800 132.800 ;
        RECT 17.000 132.000 17.800 132.200 ;
        RECT 1.200 131.000 6.800 131.200 ;
        RECT 1.200 130.800 7.000 131.000 ;
        RECT 1.200 130.600 11.000 130.800 ;
        RECT 1.200 122.200 2.000 130.600 ;
        RECT 6.200 130.200 11.000 130.600 ;
        RECT 4.400 129.000 9.800 129.600 ;
        RECT 4.400 128.800 5.200 129.000 ;
        RECT 9.000 128.800 9.800 129.000 ;
        RECT 10.400 129.000 11.000 130.200 ;
        RECT 12.400 130.400 13.000 131.600 ;
        RECT 15.400 131.400 16.200 131.600 ;
        RECT 18.800 131.400 19.600 134.800 ;
        RECT 20.600 134.400 21.200 135.800 ;
        RECT 22.200 135.400 25.800 135.800 ;
        RECT 24.400 134.400 25.200 134.800 ;
        RECT 27.000 134.400 27.600 135.800 ;
        RECT 28.600 135.400 32.200 135.800 ;
        RECT 33.200 135.000 34.000 139.800 ;
        RECT 37.600 138.400 38.400 139.800 ;
        RECT 36.400 137.800 38.400 138.400 ;
        RECT 42.000 137.800 42.800 139.800 ;
        RECT 46.200 138.400 47.400 139.800 ;
        RECT 46.000 137.800 47.400 138.400 ;
        RECT 36.400 137.000 37.200 137.800 ;
        RECT 42.000 137.200 42.600 137.800 ;
        RECT 38.000 135.600 38.800 137.200 ;
        RECT 39.800 136.600 42.600 137.200 ;
        RECT 46.000 137.000 46.800 137.800 ;
        RECT 39.800 136.400 40.600 136.600 ;
        RECT 30.800 134.400 31.600 134.800 ;
        RECT 20.400 133.600 23.000 134.400 ;
        RECT 24.400 133.800 26.000 134.400 ;
        RECT 25.200 133.600 26.000 133.800 ;
        RECT 26.800 133.600 29.400 134.400 ;
        RECT 30.800 133.800 32.400 134.400 ;
        RECT 31.600 133.600 32.400 133.800 ;
        RECT 34.000 134.200 35.600 134.400 ;
        RECT 38.200 134.200 38.800 135.600 ;
        RECT 47.800 135.400 48.600 135.600 ;
        RECT 50.800 135.400 51.600 139.800 ;
        RECT 52.400 136.000 53.200 139.800 ;
        RECT 55.600 136.000 56.400 139.800 ;
        RECT 52.400 135.800 56.400 136.000 ;
        RECT 57.200 135.800 58.000 139.800 ;
        RECT 58.800 135.800 59.600 139.800 ;
        RECT 60.400 136.000 61.200 139.800 ;
        RECT 63.600 136.000 64.400 139.800 ;
        RECT 69.000 136.000 69.800 139.000 ;
        RECT 73.200 137.000 74.000 139.000 ;
        RECT 60.400 135.800 64.400 136.000 ;
        RECT 52.600 135.400 56.200 135.800 ;
        RECT 47.800 134.800 51.600 135.400 ;
        RECT 43.800 134.200 44.600 134.400 ;
        RECT 34.000 133.600 45.000 134.200 ;
        RECT 15.400 130.800 19.600 131.400 ;
        RECT 12.400 129.800 14.800 130.400 ;
        RECT 11.800 129.000 12.600 129.200 ;
        RECT 10.400 128.400 12.600 129.000 ;
        RECT 14.200 128.800 14.800 129.800 ;
        RECT 18.800 130.300 19.600 130.800 ;
        RECT 22.400 130.400 23.000 133.600 ;
        RECT 23.600 132.300 24.400 133.200 ;
        RECT 26.800 132.300 27.600 132.400 ;
        RECT 23.600 131.700 27.600 132.300 ;
        RECT 23.600 131.600 24.400 131.700 ;
        RECT 26.800 131.600 27.600 131.700 ;
        RECT 20.400 130.300 21.200 130.400 ;
        RECT 18.800 130.200 21.200 130.300 ;
        RECT 18.800 129.700 21.800 130.200 ;
        RECT 14.200 128.000 15.600 128.800 ;
        RECT 7.800 127.400 8.600 127.600 ;
        RECT 10.600 127.400 11.400 127.600 ;
        RECT 4.400 126.200 5.200 127.000 ;
        RECT 7.800 126.800 11.400 127.400 ;
        RECT 10.000 126.200 10.600 126.800 ;
        RECT 14.000 126.200 14.800 127.000 ;
        RECT 4.400 125.600 6.400 126.200 ;
        RECT 5.600 122.200 6.400 125.600 ;
        RECT 10.000 122.200 10.800 126.200 ;
        RECT 14.200 122.200 15.400 126.200 ;
        RECT 18.800 122.200 19.600 129.700 ;
        RECT 20.400 129.600 21.800 129.700 ;
        RECT 22.400 129.600 24.400 130.400 ;
        RECT 26.800 130.200 27.600 130.400 ;
        RECT 28.800 130.200 29.400 133.600 ;
        RECT 37.000 133.400 37.800 133.600 ;
        RECT 30.000 131.600 30.800 133.200 ;
        RECT 35.400 132.400 36.200 132.600 ;
        RECT 35.400 131.800 40.400 132.400 ;
        RECT 39.600 131.600 40.400 131.800 ;
        RECT 33.200 131.000 38.800 131.200 ;
        RECT 33.200 130.800 39.000 131.000 ;
        RECT 33.200 130.600 43.000 130.800 ;
        RECT 26.800 129.600 28.200 130.200 ;
        RECT 28.800 129.600 29.800 130.200 ;
        RECT 21.200 128.400 21.800 129.600 ;
        RECT 21.200 127.600 22.000 128.400 ;
        RECT 22.600 122.200 23.400 129.600 ;
        RECT 27.600 128.400 28.200 129.600 ;
        RECT 27.600 127.600 28.400 128.400 ;
        RECT 29.000 122.200 29.800 129.600 ;
        RECT 33.200 122.200 34.000 130.600 ;
        RECT 38.200 130.200 43.000 130.600 ;
        RECT 36.400 129.000 41.800 129.600 ;
        RECT 36.400 128.800 37.200 129.000 ;
        RECT 41.000 128.800 41.800 129.000 ;
        RECT 42.400 129.000 43.000 130.200 ;
        RECT 44.400 130.400 45.000 133.600 ;
        RECT 46.000 132.800 46.800 133.000 ;
        RECT 46.000 132.200 49.800 132.800 ;
        RECT 49.000 132.000 49.800 132.200 ;
        RECT 47.400 131.400 48.200 131.600 ;
        RECT 50.800 131.400 51.600 134.800 ;
        RECT 53.200 134.400 54.000 134.800 ;
        RECT 57.200 134.400 57.800 135.800 ;
        RECT 59.000 134.400 59.600 135.800 ;
        RECT 60.600 135.400 64.200 135.800 ;
        RECT 68.200 135.400 69.800 136.000 ;
        RECT 68.200 135.000 69.000 135.400 ;
        RECT 62.800 134.400 63.600 134.800 ;
        RECT 68.200 134.400 68.800 135.000 ;
        RECT 73.400 134.800 74.000 137.000 ;
        RECT 74.800 136.000 75.600 139.800 ;
        RECT 78.000 136.000 78.800 139.800 ;
        RECT 74.800 135.800 78.800 136.000 ;
        RECT 79.600 135.800 80.400 139.800 ;
        RECT 81.200 135.800 82.000 139.800 ;
        RECT 82.800 136.000 83.600 139.800 ;
        RECT 86.000 136.000 86.800 139.800 ;
        RECT 82.800 135.800 86.800 136.000 ;
        RECT 75.000 135.400 78.600 135.800 ;
        RECT 52.400 133.800 54.000 134.400 ;
        RECT 52.400 133.600 53.200 133.800 ;
        RECT 55.400 133.600 58.000 134.400 ;
        RECT 58.800 133.600 61.400 134.400 ;
        RECT 62.800 133.800 64.400 134.400 ;
        RECT 66.800 134.300 68.800 134.400 ;
        RECT 63.600 133.600 64.400 133.800 ;
        RECT 65.300 133.700 68.800 134.300 ;
        RECT 69.800 134.200 74.000 134.800 ;
        RECT 75.600 134.400 76.400 134.800 ;
        RECT 79.600 134.400 80.200 135.800 ;
        RECT 81.400 134.400 82.000 135.800 ;
        RECT 83.000 135.400 86.600 135.800 ;
        RECT 87.600 135.600 88.400 137.200 ;
        RECT 85.200 134.400 86.000 134.800 ;
        RECT 69.800 133.800 70.800 134.200 ;
        RECT 54.000 131.600 54.800 133.200 ;
        RECT 55.400 132.300 56.000 133.600 ;
        RECT 55.400 131.700 59.500 132.300 ;
        RECT 47.400 130.800 51.600 131.400 ;
        RECT 44.400 129.800 46.800 130.400 ;
        RECT 43.800 129.000 44.600 129.200 ;
        RECT 42.400 128.400 44.600 129.000 ;
        RECT 46.200 128.800 46.800 129.800 ;
        RECT 46.200 128.400 47.600 128.800 ;
        RECT 46.200 128.000 48.400 128.400 ;
        RECT 47.000 127.600 48.400 128.000 ;
        RECT 39.800 127.400 40.600 127.600 ;
        RECT 42.600 127.400 43.400 127.600 ;
        RECT 36.400 126.200 37.200 127.000 ;
        RECT 39.800 126.800 43.400 127.400 ;
        RECT 42.000 126.200 42.600 126.800 ;
        RECT 46.000 126.200 46.800 127.000 ;
        RECT 36.400 125.600 38.400 126.200 ;
        RECT 37.600 122.200 38.400 125.600 ;
        RECT 42.000 122.200 42.800 126.200 ;
        RECT 46.200 122.200 47.400 126.200 ;
        RECT 50.800 122.200 51.600 130.800 ;
        RECT 55.400 130.200 56.000 131.700 ;
        RECT 58.900 130.400 59.500 131.700 ;
        RECT 57.200 130.200 58.000 130.400 ;
        RECT 55.000 129.600 56.000 130.200 ;
        RECT 56.600 129.600 58.000 130.200 ;
        RECT 58.800 130.200 59.600 130.400 ;
        RECT 60.800 130.200 61.400 133.600 ;
        RECT 62.000 132.300 62.800 133.200 ;
        RECT 65.300 132.300 65.900 133.700 ;
        RECT 66.800 133.600 68.800 133.700 ;
        RECT 62.000 131.700 65.900 132.300 ;
        RECT 62.000 131.600 62.800 131.700 ;
        RECT 66.800 130.800 67.600 132.400 ;
        RECT 58.800 129.600 60.200 130.200 ;
        RECT 60.800 129.600 61.800 130.200 ;
        RECT 55.000 122.200 55.800 129.600 ;
        RECT 56.600 128.400 57.200 129.600 ;
        RECT 56.400 127.600 57.200 128.400 ;
        RECT 59.600 128.400 60.200 129.600 ;
        RECT 59.600 127.600 60.400 128.400 ;
        RECT 61.000 122.200 61.800 129.600 ;
        RECT 68.200 129.800 68.800 133.600 ;
        RECT 69.400 133.000 70.800 133.800 ;
        RECT 74.800 133.800 76.400 134.400 ;
        RECT 74.800 133.600 75.600 133.800 ;
        RECT 77.800 133.600 80.400 134.400 ;
        RECT 81.200 133.600 83.800 134.400 ;
        RECT 85.200 133.800 86.800 134.400 ;
        RECT 86.000 133.600 86.800 133.800 ;
        RECT 89.200 134.300 90.000 139.800 ;
        RECT 94.600 136.000 95.400 139.000 ;
        RECT 98.800 137.000 99.600 139.000 ;
        RECT 93.800 135.400 95.400 136.000 ;
        RECT 93.800 135.000 94.600 135.400 ;
        RECT 93.800 134.400 94.400 135.000 ;
        RECT 99.000 134.800 99.600 137.000 ;
        RECT 90.800 134.300 91.600 134.400 ;
        RECT 89.200 133.700 91.600 134.300 ;
        RECT 70.200 131.000 70.800 133.000 ;
        RECT 71.600 131.600 72.400 133.200 ;
        RECT 73.200 131.600 74.000 133.200 ;
        RECT 74.800 132.300 75.600 132.400 ;
        RECT 76.400 132.300 77.200 133.200 ;
        RECT 74.800 131.700 77.200 132.300 ;
        RECT 74.800 131.600 75.600 131.700 ;
        RECT 76.400 131.600 77.200 131.700 ;
        RECT 70.200 130.400 74.000 131.000 ;
        RECT 68.200 129.200 69.800 129.800 ;
        RECT 69.000 122.200 69.800 129.200 ;
        RECT 73.400 127.000 74.000 130.400 ;
        RECT 77.800 130.200 78.400 133.600 ;
        RECT 83.200 132.300 83.800 133.600 ;
        RECT 79.700 131.700 83.800 132.300 ;
        RECT 79.700 130.400 80.300 131.700 ;
        RECT 79.600 130.200 80.400 130.400 ;
        RECT 73.200 123.000 74.000 127.000 ;
        RECT 77.400 129.600 78.400 130.200 ;
        RECT 79.000 129.600 80.400 130.200 ;
        RECT 81.200 130.200 82.000 130.400 ;
        RECT 83.200 130.200 83.800 131.700 ;
        RECT 84.400 131.600 85.200 133.200 ;
        RECT 81.200 129.600 82.600 130.200 ;
        RECT 83.200 129.600 84.200 130.200 ;
        RECT 77.400 124.400 78.200 129.600 ;
        RECT 79.000 128.400 79.600 129.600 ;
        RECT 78.800 127.600 79.600 128.400 ;
        RECT 82.000 128.400 82.600 129.600 ;
        RECT 82.000 127.600 82.800 128.400 ;
        RECT 76.400 123.600 78.200 124.400 ;
        RECT 77.400 122.200 78.200 123.600 ;
        RECT 83.400 122.200 84.200 129.600 ;
        RECT 89.200 122.200 90.000 133.700 ;
        RECT 90.800 133.600 91.600 133.700 ;
        RECT 92.400 133.600 94.400 134.400 ;
        RECT 95.400 134.200 99.600 134.800 ;
        RECT 104.000 134.200 104.800 139.800 ;
        RECT 106.800 135.800 107.600 139.800 ;
        RECT 108.400 136.000 109.200 139.800 ;
        RECT 111.600 136.000 112.400 139.800 ;
        RECT 120.600 136.400 121.400 139.800 ;
        RECT 108.400 135.800 112.400 136.000 ;
        RECT 119.600 135.800 121.400 136.400 ;
        RECT 122.800 135.800 123.600 139.800 ;
        RECT 124.400 136.000 125.200 139.800 ;
        RECT 127.600 136.000 128.400 139.800 ;
        RECT 124.400 135.800 128.400 136.000 ;
        RECT 107.000 134.400 107.600 135.800 ;
        RECT 108.600 135.400 112.200 135.800 ;
        RECT 110.800 134.400 111.600 134.800 ;
        RECT 95.400 133.800 96.400 134.200 ;
        RECT 104.000 133.800 105.800 134.200 ;
        RECT 92.400 130.800 93.200 132.400 ;
        RECT 93.800 129.800 94.400 133.600 ;
        RECT 95.000 133.000 96.400 133.800 ;
        RECT 104.200 133.600 105.800 133.800 ;
        RECT 106.800 133.600 109.400 134.400 ;
        RECT 110.800 133.800 112.400 134.400 ;
        RECT 111.600 133.600 112.400 133.800 ;
        RECT 118.000 133.600 118.800 135.200 ;
        RECT 95.800 131.000 96.400 133.000 ;
        RECT 97.200 131.600 98.000 133.200 ;
        RECT 98.800 131.600 99.600 133.200 ;
        RECT 102.000 131.600 103.600 132.400 ;
        RECT 95.800 130.400 99.600 131.000 ;
        RECT 93.800 129.200 95.400 129.800 ;
        RECT 94.600 124.400 95.400 129.200 ;
        RECT 99.000 127.000 99.600 130.400 ;
        RECT 100.400 129.600 101.200 131.200 ;
        RECT 105.200 130.400 105.800 133.600 ;
        RECT 105.200 130.300 106.000 130.400 ;
        RECT 106.800 130.300 107.600 130.400 ;
        RECT 105.200 130.200 107.600 130.300 ;
        RECT 108.800 130.200 109.400 133.600 ;
        RECT 110.000 131.600 110.800 133.200 ;
        RECT 119.600 132.300 120.400 135.800 ;
        RECT 123.000 134.400 123.600 135.800 ;
        RECT 124.600 135.400 128.200 135.800 ;
        RECT 126.800 134.400 127.600 134.800 ;
        RECT 122.800 133.600 125.400 134.400 ;
        RECT 126.800 134.300 128.400 134.400 ;
        RECT 129.200 134.300 130.000 139.800 ;
        RECT 130.800 135.600 131.600 137.200 ;
        RECT 126.800 133.800 130.000 134.300 ;
        RECT 136.000 134.200 136.800 139.800 ;
        RECT 138.800 135.600 139.600 137.200 ;
        RECT 140.400 134.300 141.200 139.800 ;
        RECT 142.000 136.000 142.800 139.800 ;
        RECT 145.200 136.000 146.000 139.800 ;
        RECT 142.000 135.800 146.000 136.000 ;
        RECT 146.800 135.800 147.600 139.800 ;
        RECT 148.400 135.800 149.200 139.800 ;
        RECT 150.000 136.000 150.800 139.800 ;
        RECT 153.200 136.000 154.000 139.800 ;
        RECT 150.000 135.800 154.000 136.000 ;
        RECT 154.800 136.000 155.600 139.800 ;
        RECT 158.000 136.000 158.800 139.800 ;
        RECT 154.800 135.800 158.800 136.000 ;
        RECT 159.600 135.800 160.400 139.800 ;
        RECT 142.200 135.400 145.800 135.800 ;
        RECT 142.800 134.400 143.600 134.800 ;
        RECT 146.800 134.400 147.400 135.800 ;
        RECT 148.600 134.400 149.200 135.800 ;
        RECT 150.200 135.400 153.800 135.800 ;
        RECT 155.000 135.400 158.600 135.800 ;
        RECT 152.400 134.400 153.200 134.800 ;
        RECT 155.600 134.400 156.400 134.800 ;
        RECT 159.600 134.400 160.200 135.800 ;
        RECT 142.000 134.300 143.600 134.400 ;
        RECT 136.000 133.800 137.800 134.200 ;
        RECT 127.600 133.700 130.000 133.800 ;
        RECT 127.600 133.600 128.400 133.700 ;
        RECT 119.600 131.700 123.500 132.300 ;
        RECT 105.200 129.700 108.200 130.200 ;
        RECT 105.200 129.600 106.000 129.700 ;
        RECT 106.800 129.600 108.200 129.700 ;
        RECT 108.800 129.600 109.800 130.200 ;
        RECT 103.600 127.600 104.400 129.200 ;
        RECT 105.200 127.000 105.800 129.600 ;
        RECT 107.600 128.400 108.200 129.600 ;
        RECT 107.600 127.600 108.400 128.400 ;
        RECT 94.600 123.600 96.400 124.400 ;
        RECT 94.600 122.200 95.400 123.600 ;
        RECT 98.800 123.000 99.600 127.000 ;
        RECT 102.200 126.400 105.800 127.000 ;
        RECT 102.200 126.200 102.800 126.400 ;
        RECT 102.000 122.200 102.800 126.200 ;
        RECT 105.200 126.200 105.800 126.400 ;
        RECT 105.200 122.200 106.000 126.200 ;
        RECT 109.000 122.200 109.800 129.600 ;
        RECT 119.600 122.200 120.400 131.700 ;
        RECT 122.900 130.400 123.500 131.700 ;
        RECT 121.200 128.800 122.000 130.400 ;
        RECT 122.800 130.200 123.600 130.400 ;
        RECT 124.800 130.200 125.400 133.600 ;
        RECT 126.000 131.600 126.800 133.200 ;
        RECT 122.800 129.600 124.200 130.200 ;
        RECT 124.800 129.600 125.800 130.200 ;
        RECT 123.600 128.400 124.200 129.600 ;
        RECT 123.600 127.600 124.400 128.400 ;
        RECT 125.000 124.400 125.800 129.600 ;
        RECT 125.000 123.600 126.800 124.400 ;
        RECT 125.000 122.200 125.800 123.600 ;
        RECT 129.200 122.200 130.000 133.700 ;
        RECT 136.200 133.600 137.800 133.800 ;
        RECT 134.000 131.600 135.600 132.400 ;
        RECT 132.400 129.600 133.200 131.200 ;
        RECT 137.200 130.400 137.800 133.600 ;
        RECT 140.400 133.800 143.600 134.300 ;
        RECT 140.400 133.700 142.800 133.800 ;
        RECT 137.200 129.600 138.000 130.400 ;
        RECT 135.600 127.600 136.400 129.200 ;
        RECT 137.200 127.000 137.800 129.600 ;
        RECT 134.200 126.400 137.800 127.000 ;
        RECT 134.200 126.200 134.800 126.400 ;
        RECT 134.000 122.200 134.800 126.200 ;
        RECT 137.200 126.200 137.800 126.400 ;
        RECT 137.200 122.200 138.000 126.200 ;
        RECT 140.400 122.200 141.200 133.700 ;
        RECT 142.000 133.600 142.800 133.700 ;
        RECT 145.000 133.600 147.600 134.400 ;
        RECT 148.400 133.600 151.000 134.400 ;
        RECT 152.400 133.800 154.000 134.400 ;
        RECT 153.200 133.600 154.000 133.800 ;
        RECT 154.800 133.800 156.400 134.400 ;
        RECT 154.800 133.600 155.600 133.800 ;
        RECT 157.800 133.600 160.400 134.400 ;
        RECT 143.600 131.600 144.400 133.200 ;
        RECT 145.000 132.300 145.600 133.600 ;
        RECT 150.400 132.400 151.000 133.600 ;
        RECT 148.400 132.300 149.200 132.400 ;
        RECT 145.000 131.700 149.200 132.300 ;
        RECT 145.000 130.200 145.600 131.700 ;
        RECT 148.400 131.600 149.200 131.700 ;
        RECT 150.000 131.600 151.000 132.400 ;
        RECT 151.600 131.600 152.400 133.200 ;
        RECT 156.400 131.600 157.200 133.200 ;
        RECT 146.800 130.200 147.600 130.400 ;
        RECT 144.600 129.600 145.600 130.200 ;
        RECT 146.200 129.600 147.600 130.200 ;
        RECT 148.400 130.200 149.200 130.400 ;
        RECT 150.400 130.200 151.000 131.600 ;
        RECT 157.800 130.200 158.400 133.600 ;
        RECT 159.600 130.200 160.400 130.400 ;
        RECT 148.400 129.600 149.800 130.200 ;
        RECT 150.400 129.600 151.400 130.200 ;
        RECT 144.600 122.200 145.400 129.600 ;
        RECT 146.200 128.400 146.800 129.600 ;
        RECT 146.000 127.600 146.800 128.400 ;
        RECT 149.200 128.400 149.800 129.600 ;
        RECT 149.200 127.600 150.000 128.400 ;
        RECT 150.600 122.200 151.400 129.600 ;
        RECT 157.400 129.600 158.400 130.200 ;
        RECT 159.000 129.600 160.400 130.200 ;
        RECT 157.400 122.200 158.200 129.600 ;
        RECT 159.000 128.400 159.600 129.600 ;
        RECT 158.800 127.600 159.600 128.400 ;
        RECT 161.200 122.200 162.000 139.800 ;
        RECT 162.800 135.600 163.600 137.200 ;
        RECT 164.400 135.200 165.200 139.800 ;
        RECT 167.600 136.400 168.400 139.800 ;
        RECT 167.600 135.800 168.600 136.400 ;
        RECT 164.400 134.600 167.000 135.200 ;
        RECT 164.600 132.400 165.400 133.200 ;
        RECT 162.800 132.300 163.600 132.400 ;
        RECT 164.400 132.300 165.400 132.400 ;
        RECT 162.800 131.700 165.400 132.300 ;
        RECT 162.800 131.600 163.600 131.700 ;
        RECT 164.400 131.600 165.400 131.700 ;
        RECT 166.400 133.000 167.000 134.600 ;
        RECT 168.000 134.400 168.600 135.800 ;
        RECT 167.600 133.600 168.600 134.400 ;
        RECT 172.000 134.400 172.800 139.800 ;
        RECT 177.200 135.800 178.000 139.800 ;
        RECT 178.800 136.000 179.600 139.800 ;
        RECT 182.000 136.000 182.800 139.800 ;
        RECT 178.800 135.800 182.800 136.000 ;
        RECT 184.200 136.400 185.000 139.800 ;
        RECT 184.200 135.800 186.000 136.400 ;
        RECT 188.400 135.800 189.200 139.800 ;
        RECT 190.000 136.000 190.800 139.800 ;
        RECT 193.200 136.000 194.000 139.800 ;
        RECT 190.000 135.800 194.000 136.000 ;
        RECT 194.800 136.000 195.600 139.800 ;
        RECT 198.000 136.000 198.800 139.800 ;
        RECT 194.800 135.800 198.800 136.000 ;
        RECT 199.600 135.800 200.400 139.800 ;
        RECT 202.800 136.000 203.600 139.800 ;
        RECT 177.400 134.400 178.000 135.800 ;
        RECT 179.000 135.400 182.600 135.800 ;
        RECT 181.200 134.400 182.000 134.800 ;
        RECT 172.000 134.200 173.200 134.400 ;
        RECT 166.400 132.200 167.400 133.000 ;
        RECT 166.400 130.200 167.000 132.200 ;
        RECT 168.000 130.200 168.600 133.600 ;
        RECT 171.000 133.600 173.200 134.200 ;
        RECT 177.200 133.600 179.800 134.400 ;
        RECT 181.200 134.300 182.800 134.400 ;
        RECT 183.600 134.300 184.400 134.400 ;
        RECT 181.200 133.800 184.400 134.300 ;
        RECT 182.000 133.700 184.400 133.800 ;
        RECT 182.000 133.600 182.800 133.700 ;
        RECT 183.600 133.600 184.400 133.700 ;
        RECT 171.000 130.400 171.600 133.600 ;
        RECT 173.200 131.600 174.800 132.400 ;
        RECT 164.400 129.600 167.000 130.200 ;
        RECT 164.400 122.200 165.200 129.600 ;
        RECT 167.600 129.200 168.600 130.200 ;
        RECT 170.800 129.600 171.600 130.400 ;
        RECT 175.600 129.600 176.400 131.200 ;
        RECT 177.200 130.200 178.000 130.400 ;
        RECT 179.200 130.200 179.800 133.600 ;
        RECT 180.400 131.600 181.200 133.200 ;
        RECT 177.200 129.600 178.600 130.200 ;
        RECT 179.200 129.600 180.200 130.200 ;
        RECT 167.600 122.200 168.400 129.200 ;
        RECT 171.000 127.000 171.600 129.600 ;
        RECT 172.400 127.600 173.200 129.200 ;
        RECT 178.000 128.400 178.600 129.600 ;
        RECT 178.000 127.600 178.800 128.400 ;
        RECT 171.000 126.400 174.600 127.000 ;
        RECT 171.000 126.200 171.600 126.400 ;
        RECT 170.800 122.200 171.600 126.200 ;
        RECT 174.000 126.200 174.600 126.400 ;
        RECT 174.000 122.200 174.800 126.200 ;
        RECT 179.400 122.200 180.200 129.600 ;
        RECT 183.600 128.800 184.400 130.400 ;
        RECT 185.200 130.300 186.000 135.800 ;
        RECT 186.800 133.600 187.600 135.200 ;
        RECT 188.600 134.400 189.200 135.800 ;
        RECT 190.200 135.400 193.800 135.800 ;
        RECT 195.000 135.400 198.600 135.800 ;
        RECT 192.400 134.400 193.200 134.800 ;
        RECT 195.600 134.400 196.400 134.800 ;
        RECT 199.600 134.400 200.200 135.800 ;
        RECT 202.600 135.200 203.600 136.000 ;
        RECT 188.400 133.600 191.000 134.400 ;
        RECT 192.400 133.800 194.000 134.400 ;
        RECT 193.200 133.600 194.000 133.800 ;
        RECT 194.800 133.800 196.400 134.400 ;
        RECT 194.800 133.600 195.600 133.800 ;
        RECT 197.800 133.600 200.400 134.400 ;
        RECT 190.400 130.400 191.000 133.600 ;
        RECT 191.600 131.600 192.400 133.200 ;
        RECT 193.200 132.300 194.000 132.400 ;
        RECT 196.400 132.300 197.200 133.200 ;
        RECT 193.200 131.700 197.200 132.300 ;
        RECT 193.200 131.600 194.000 131.700 ;
        RECT 196.400 131.600 197.200 131.700 ;
        RECT 188.400 130.300 189.200 130.400 ;
        RECT 185.200 130.200 189.200 130.300 ;
        RECT 185.200 129.700 189.800 130.200 ;
        RECT 185.200 122.200 186.000 129.700 ;
        RECT 188.400 129.600 189.800 129.700 ;
        RECT 190.400 129.600 192.400 130.400 ;
        RECT 197.800 130.200 198.400 133.600 ;
        RECT 202.600 130.800 203.400 135.200 ;
        RECT 204.400 134.600 205.200 139.800 ;
        RECT 210.800 136.600 211.600 139.800 ;
        RECT 212.400 137.000 213.200 139.800 ;
        RECT 214.000 137.000 214.800 139.800 ;
        RECT 215.600 137.000 216.400 139.800 ;
        RECT 217.200 137.000 218.000 139.800 ;
        RECT 220.400 137.000 221.200 139.800 ;
        RECT 223.600 137.000 224.400 139.800 ;
        RECT 225.200 137.000 226.000 139.800 ;
        RECT 226.800 137.000 227.600 139.800 ;
        RECT 209.200 135.800 211.600 136.600 ;
        RECT 228.400 136.600 229.200 139.800 ;
        RECT 209.200 135.200 210.000 135.800 ;
        RECT 204.000 134.000 205.200 134.600 ;
        RECT 208.200 134.600 210.000 135.200 ;
        RECT 214.000 135.600 215.000 136.400 ;
        RECT 218.000 135.600 219.600 136.400 ;
        RECT 220.400 135.800 225.000 136.400 ;
        RECT 228.400 135.800 231.000 136.600 ;
        RECT 220.400 135.600 221.200 135.800 ;
        RECT 204.000 132.000 204.600 134.000 ;
        RECT 208.200 133.400 209.000 134.600 ;
        RECT 205.200 132.600 209.000 133.400 ;
        RECT 214.000 132.800 214.800 135.600 ;
        RECT 220.400 134.800 221.200 135.000 ;
        RECT 216.800 134.200 221.200 134.800 ;
        RECT 216.800 134.000 217.600 134.200 ;
        RECT 222.000 133.600 222.800 135.200 ;
        RECT 224.200 133.400 225.000 135.800 ;
        RECT 230.200 135.200 231.000 135.800 ;
        RECT 230.200 134.400 233.200 135.200 ;
        RECT 234.800 133.800 235.600 139.800 ;
        RECT 237.600 134.200 238.400 139.800 ;
        RECT 217.200 132.600 220.400 133.400 ;
        RECT 224.200 132.600 226.200 133.400 ;
        RECT 226.800 133.000 235.600 133.800 ;
        RECT 210.800 132.000 211.600 132.600 ;
        RECT 228.400 132.000 229.200 132.400 ;
        RECT 230.000 132.000 230.800 132.400 ;
        RECT 233.400 132.000 234.200 132.200 ;
        RECT 204.000 131.400 204.800 132.000 ;
        RECT 210.800 131.400 234.200 132.000 ;
        RECT 199.600 130.200 200.400 130.400 ;
        RECT 197.400 129.600 198.400 130.200 ;
        RECT 199.000 129.600 200.400 130.200 ;
        RECT 202.600 130.000 203.600 130.800 ;
        RECT 189.200 128.400 189.800 129.600 ;
        RECT 189.200 127.600 190.000 128.400 ;
        RECT 190.600 122.200 191.400 129.600 ;
        RECT 197.400 126.400 198.200 129.600 ;
        RECT 199.000 128.400 199.600 129.600 ;
        RECT 198.800 127.600 199.600 128.400 ;
        RECT 196.400 125.600 198.200 126.400 ;
        RECT 197.400 122.200 198.200 125.600 ;
        RECT 202.800 122.200 203.600 130.000 ;
        RECT 204.200 129.600 204.800 131.400 ;
        RECT 204.200 129.000 213.200 129.600 ;
        RECT 204.200 127.400 204.800 129.000 ;
        RECT 212.400 128.800 213.200 129.000 ;
        RECT 215.600 129.000 224.200 129.600 ;
        RECT 215.600 128.800 216.400 129.000 ;
        RECT 207.400 127.600 210.000 128.400 ;
        RECT 204.200 126.800 206.800 127.400 ;
        RECT 206.000 122.200 206.800 126.800 ;
        RECT 209.200 122.200 210.000 127.600 ;
        RECT 210.600 126.800 214.800 127.600 ;
        RECT 212.400 122.200 213.200 125.000 ;
        RECT 214.000 122.200 214.800 125.000 ;
        RECT 215.600 122.200 216.400 125.000 ;
        RECT 217.200 122.200 218.000 128.400 ;
        RECT 220.400 127.600 223.000 128.400 ;
        RECT 223.600 128.200 224.200 129.000 ;
        RECT 225.200 129.400 226.000 129.600 ;
        RECT 225.200 129.000 230.600 129.400 ;
        RECT 225.200 128.800 231.400 129.000 ;
        RECT 230.000 128.200 231.400 128.800 ;
        RECT 223.600 127.600 229.400 128.200 ;
        RECT 232.400 128.000 234.000 128.800 ;
        RECT 232.400 127.600 233.000 128.000 ;
        RECT 220.400 122.200 221.200 127.000 ;
        RECT 223.600 122.200 224.400 127.000 ;
        RECT 228.800 126.800 233.000 127.600 ;
        RECT 234.800 127.400 235.600 133.000 ;
        RECT 236.600 133.800 238.400 134.200 ;
        RECT 242.800 135.800 243.600 139.800 ;
        RECT 246.000 137.800 246.800 139.800 ;
        RECT 250.800 137.800 251.600 139.800 ;
        RECT 236.600 133.600 238.200 133.800 ;
        RECT 236.600 130.400 237.200 133.600 ;
        RECT 242.800 132.400 243.400 135.800 ;
        RECT 246.000 135.600 246.600 137.800 ;
        RECT 247.600 136.300 248.400 137.200 ;
        RECT 249.200 136.300 250.000 136.400 ;
        RECT 247.600 135.700 250.000 136.300 ;
        RECT 247.600 135.600 248.400 135.700 ;
        RECT 249.200 135.600 250.000 135.700 ;
        RECT 244.200 135.000 246.600 135.600 ;
        RECT 238.800 131.600 240.400 132.400 ;
        RECT 242.800 131.600 243.600 132.400 ;
        RECT 244.200 132.000 244.800 135.000 ;
        RECT 250.800 134.400 251.400 137.800 ;
        RECT 252.400 135.600 253.200 137.200 ;
        RECT 255.600 135.200 256.400 139.800 ;
        RECT 258.800 135.200 259.600 139.800 ;
        RECT 268.400 136.400 269.200 139.800 ;
        RECT 255.600 134.400 259.600 135.200 ;
        RECT 268.200 135.800 269.200 136.400 ;
        RECT 268.200 134.400 268.800 135.800 ;
        RECT 271.600 135.200 272.400 139.800 ;
        RECT 274.800 136.400 275.600 139.800 ;
        RECT 269.800 134.600 272.400 135.200 ;
        RECT 274.600 135.600 275.600 136.400 ;
        RECT 245.800 133.600 246.800 134.400 ;
        RECT 250.800 133.600 251.600 134.400 ;
        RECT 245.600 132.800 246.400 133.600 ;
        RECT 236.400 129.600 237.200 130.400 ;
        RECT 241.200 129.600 242.000 131.200 ;
        RECT 242.800 130.200 243.400 131.600 ;
        RECT 244.200 131.400 245.000 132.000 ;
        RECT 244.200 131.200 248.400 131.400 ;
        RECT 244.400 130.800 248.400 131.200 ;
        RECT 249.200 130.800 250.000 132.400 ;
        RECT 242.800 129.600 244.200 130.200 ;
        RECT 233.600 126.800 235.600 127.400 ;
        RECT 236.600 127.000 237.200 129.600 ;
        RECT 238.000 127.600 238.800 129.200 ;
        RECT 225.200 122.200 226.000 125.000 ;
        RECT 226.800 122.200 227.600 125.000 ;
        RECT 230.000 122.200 230.800 126.800 ;
        RECT 233.600 126.200 234.200 126.800 ;
        RECT 236.600 126.400 240.200 127.000 ;
        RECT 236.600 126.200 237.200 126.400 ;
        RECT 233.200 125.600 234.200 126.200 ;
        RECT 233.200 122.200 234.000 125.600 ;
        RECT 236.400 122.200 237.200 126.200 ;
        RECT 239.600 126.200 240.200 126.400 ;
        RECT 239.600 122.200 240.400 126.200 ;
        RECT 243.400 124.400 244.200 129.600 ;
        RECT 242.800 123.600 244.200 124.400 ;
        RECT 243.400 122.200 244.200 123.600 ;
        RECT 247.600 122.200 248.400 130.800 ;
        RECT 250.800 130.200 251.400 133.600 ;
        RECT 255.600 131.600 256.400 134.400 ;
        RECT 268.200 133.600 269.200 134.400 ;
        RECT 255.600 130.800 259.600 131.600 ;
        RECT 249.800 129.400 251.600 130.200 ;
        RECT 249.800 124.400 250.600 129.400 ;
        RECT 249.800 123.600 251.600 124.400 ;
        RECT 249.800 122.200 250.600 123.600 ;
        RECT 255.600 122.200 256.400 130.800 ;
        RECT 258.800 122.200 259.600 130.800 ;
        RECT 268.200 130.200 268.800 133.600 ;
        RECT 269.800 133.000 270.400 134.600 ;
        RECT 274.600 134.400 275.200 135.600 ;
        RECT 278.000 135.200 278.800 139.800 ;
        RECT 280.200 138.400 281.000 139.800 ;
        RECT 279.600 137.600 281.000 138.400 ;
        RECT 280.200 136.400 281.000 137.600 ;
        RECT 280.200 135.800 282.000 136.400 ;
        RECT 284.400 135.800 285.200 139.800 ;
        RECT 286.000 136.000 286.800 139.800 ;
        RECT 289.200 136.000 290.000 139.800 ;
        RECT 286.000 135.800 290.000 136.000 ;
        RECT 291.400 136.400 292.200 139.800 ;
        RECT 291.400 135.800 293.200 136.400 ;
        RECT 295.600 136.000 296.400 139.800 ;
        RECT 298.800 136.000 299.600 139.800 ;
        RECT 295.600 135.800 299.600 136.000 ;
        RECT 300.400 135.800 301.200 139.800 ;
        RECT 302.600 138.400 303.400 139.800 ;
        RECT 302.600 137.600 304.400 138.400 ;
        RECT 302.600 136.400 303.400 137.600 ;
        RECT 302.600 135.800 304.400 136.400 ;
        RECT 308.400 136.000 309.200 139.800 ;
        RECT 276.200 134.600 278.800 135.200 ;
        RECT 274.600 133.600 275.600 134.400 ;
        RECT 269.400 132.200 270.400 133.000 ;
        RECT 269.800 130.200 270.400 132.200 ;
        RECT 271.400 132.400 272.200 133.200 ;
        RECT 271.400 131.600 272.400 132.400 ;
        RECT 274.600 130.200 275.200 133.600 ;
        RECT 276.200 133.000 276.800 134.600 ;
        RECT 275.800 132.200 276.800 133.000 ;
        RECT 276.200 130.200 276.800 132.200 ;
        RECT 277.800 132.400 278.600 133.200 ;
        RECT 277.800 132.300 278.800 132.400 ;
        RECT 279.600 132.300 280.400 132.400 ;
        RECT 277.800 131.700 280.400 132.300 ;
        RECT 277.800 131.600 278.800 131.700 ;
        RECT 279.600 131.600 280.400 131.700 ;
        RECT 268.200 129.200 269.200 130.200 ;
        RECT 269.800 129.600 272.400 130.200 ;
        RECT 268.400 122.200 269.200 129.200 ;
        RECT 271.600 122.200 272.400 129.600 ;
        RECT 274.600 129.200 275.600 130.200 ;
        RECT 276.200 129.600 278.800 130.200 ;
        RECT 274.800 122.200 275.600 129.200 ;
        RECT 278.000 122.200 278.800 129.600 ;
        RECT 279.600 128.800 280.400 130.400 ;
        RECT 281.200 122.200 282.000 135.800 ;
        RECT 282.800 134.300 283.600 135.200 ;
        RECT 284.600 134.400 285.200 135.800 ;
        RECT 286.200 135.400 289.800 135.800 ;
        RECT 288.400 134.400 289.200 134.800 ;
        RECT 284.400 134.300 287.000 134.400 ;
        RECT 282.800 133.700 287.000 134.300 ;
        RECT 288.400 133.800 290.000 134.400 ;
        RECT 282.800 133.600 283.600 133.700 ;
        RECT 284.400 133.600 287.000 133.700 ;
        RECT 289.200 133.600 290.000 133.800 ;
        RECT 284.400 130.200 285.200 130.400 ;
        RECT 286.400 130.200 287.000 133.600 ;
        RECT 287.600 131.600 288.400 133.200 ;
        RECT 284.400 129.600 285.800 130.200 ;
        RECT 286.400 129.600 287.400 130.200 ;
        RECT 285.200 128.400 285.800 129.600 ;
        RECT 285.200 127.600 286.000 128.400 ;
        RECT 286.600 122.200 287.400 129.600 ;
        RECT 290.800 128.800 291.600 130.400 ;
        RECT 292.400 128.300 293.200 135.800 ;
        RECT 295.800 135.400 299.400 135.800 ;
        RECT 294.000 133.600 294.800 135.200 ;
        RECT 296.400 134.400 297.200 134.800 ;
        RECT 300.400 134.400 301.000 135.800 ;
        RECT 295.600 133.800 297.200 134.400 ;
        RECT 295.600 133.600 296.400 133.800 ;
        RECT 298.600 133.600 301.200 134.400 ;
        RECT 295.600 132.300 296.400 132.400 ;
        RECT 297.200 132.300 298.000 133.200 ;
        RECT 295.600 131.700 298.000 132.300 ;
        RECT 295.600 131.600 296.400 131.700 ;
        RECT 297.200 131.600 298.000 131.700 ;
        RECT 298.600 130.400 299.200 133.600 ;
        RECT 297.200 129.600 299.200 130.400 ;
        RECT 300.400 130.200 301.200 130.400 ;
        RECT 299.800 129.600 301.200 130.200 ;
        RECT 294.000 128.300 294.800 128.400 ;
        RECT 292.400 127.700 294.800 128.300 ;
        RECT 292.400 122.200 293.200 127.700 ;
        RECT 294.000 127.600 294.800 127.700 ;
        RECT 298.200 122.200 299.000 129.600 ;
        RECT 299.800 128.400 300.400 129.600 ;
        RECT 302.000 128.800 302.800 130.400 ;
        RECT 299.600 127.600 300.400 128.400 ;
        RECT 303.600 122.200 304.400 135.800 ;
        RECT 308.200 135.200 309.200 136.000 ;
        RECT 305.200 133.600 306.000 135.200 ;
        RECT 308.200 130.800 309.000 135.200 ;
        RECT 310.000 134.600 310.800 139.800 ;
        RECT 316.400 136.600 317.200 139.800 ;
        RECT 318.000 137.000 318.800 139.800 ;
        RECT 319.600 137.000 320.400 139.800 ;
        RECT 321.200 137.000 322.000 139.800 ;
        RECT 322.800 137.000 323.600 139.800 ;
        RECT 326.000 137.000 326.800 139.800 ;
        RECT 329.200 137.000 330.000 139.800 ;
        RECT 330.800 137.000 331.600 139.800 ;
        RECT 332.400 137.000 333.200 139.800 ;
        RECT 314.800 135.800 317.200 136.600 ;
        RECT 334.000 136.600 334.800 139.800 ;
        RECT 314.800 135.200 315.600 135.800 ;
        RECT 309.600 134.000 310.800 134.600 ;
        RECT 313.800 134.600 315.600 135.200 ;
        RECT 319.600 135.600 320.600 136.400 ;
        RECT 323.600 135.600 325.200 136.400 ;
        RECT 326.000 135.800 330.600 136.400 ;
        RECT 334.000 135.800 336.600 136.600 ;
        RECT 326.000 135.600 326.800 135.800 ;
        RECT 309.600 132.000 310.200 134.000 ;
        RECT 313.800 133.400 314.600 134.600 ;
        RECT 310.800 132.600 314.600 133.400 ;
        RECT 319.600 132.800 320.400 135.600 ;
        RECT 326.000 134.800 326.800 135.000 ;
        RECT 322.400 134.200 326.800 134.800 ;
        RECT 322.400 134.000 323.200 134.200 ;
        RECT 327.600 133.600 328.400 135.200 ;
        RECT 329.800 133.400 330.600 135.800 ;
        RECT 335.800 135.200 336.600 135.800 ;
        RECT 335.800 134.400 338.800 135.200 ;
        RECT 340.400 133.800 341.200 139.800 ;
        RECT 322.800 132.600 326.000 133.400 ;
        RECT 329.800 132.600 331.800 133.400 ;
        RECT 332.400 133.000 341.200 133.800 ;
        RECT 316.400 132.000 317.200 132.600 ;
        RECT 334.000 132.000 334.800 132.400 ;
        RECT 337.200 132.000 338.000 132.400 ;
        RECT 339.000 132.000 339.800 132.200 ;
        RECT 309.600 131.400 310.400 132.000 ;
        RECT 316.400 131.400 339.800 132.000 ;
        RECT 308.200 130.000 309.200 130.800 ;
        RECT 308.400 122.200 309.200 130.000 ;
        RECT 309.800 129.600 310.400 131.400 ;
        RECT 309.800 129.000 318.800 129.600 ;
        RECT 309.800 127.400 310.400 129.000 ;
        RECT 318.000 128.800 318.800 129.000 ;
        RECT 321.200 129.000 329.800 129.600 ;
        RECT 321.200 128.800 322.000 129.000 ;
        RECT 313.000 127.600 315.600 128.400 ;
        RECT 309.800 126.800 312.400 127.400 ;
        RECT 311.600 122.200 312.400 126.800 ;
        RECT 314.800 122.200 315.600 127.600 ;
        RECT 316.200 126.800 320.400 127.600 ;
        RECT 318.000 122.200 318.800 125.000 ;
        RECT 319.600 122.200 320.400 125.000 ;
        RECT 321.200 122.200 322.000 125.000 ;
        RECT 322.800 122.200 323.600 128.400 ;
        RECT 326.000 127.600 328.600 128.400 ;
        RECT 329.200 128.200 329.800 129.000 ;
        RECT 330.800 129.400 331.600 129.600 ;
        RECT 330.800 129.000 336.200 129.400 ;
        RECT 330.800 128.800 337.000 129.000 ;
        RECT 335.600 128.200 337.000 128.800 ;
        RECT 329.200 127.600 335.000 128.200 ;
        RECT 338.000 128.000 339.600 128.800 ;
        RECT 338.000 127.600 338.600 128.000 ;
        RECT 326.000 122.200 326.800 127.000 ;
        RECT 329.200 122.200 330.000 127.000 ;
        RECT 334.400 126.800 338.600 127.600 ;
        RECT 340.400 127.400 341.200 133.000 ;
        RECT 343.600 137.800 344.400 139.800 ;
        RECT 348.400 137.800 349.200 139.800 ;
        RECT 343.600 134.400 344.200 137.800 ;
        RECT 345.200 135.600 346.000 137.200 ;
        RECT 346.800 135.600 347.600 137.200 ;
        RECT 348.600 134.400 349.200 137.800 ;
        RECT 343.600 133.600 344.400 134.400 ;
        RECT 348.400 133.600 349.200 134.400 ;
        RECT 342.000 130.800 342.800 132.400 ;
        RECT 343.600 130.200 344.200 133.600 ;
        RECT 348.600 130.200 349.200 133.600 ;
        RECT 351.600 133.800 352.400 139.800 ;
        RECT 358.000 136.600 358.800 139.800 ;
        RECT 359.600 137.000 360.400 139.800 ;
        RECT 361.200 137.000 362.000 139.800 ;
        RECT 362.800 137.000 363.600 139.800 ;
        RECT 366.000 137.000 366.800 139.800 ;
        RECT 369.200 137.000 370.000 139.800 ;
        RECT 370.800 137.000 371.600 139.800 ;
        RECT 372.400 137.000 373.200 139.800 ;
        RECT 374.000 137.000 374.800 139.800 ;
        RECT 356.200 135.800 358.800 136.600 ;
        RECT 375.600 136.600 376.400 139.800 ;
        RECT 362.200 135.800 366.800 136.400 ;
        RECT 356.200 135.200 357.000 135.800 ;
        RECT 354.000 134.400 357.000 135.200 ;
        RECT 351.600 133.000 360.400 133.800 ;
        RECT 362.200 133.400 363.000 135.800 ;
        RECT 366.000 135.600 366.800 135.800 ;
        RECT 367.600 135.600 369.200 136.400 ;
        RECT 372.200 135.600 373.200 136.400 ;
        RECT 375.600 135.800 378.000 136.600 ;
        RECT 364.400 133.600 365.200 135.200 ;
        RECT 366.000 134.800 366.800 135.000 ;
        RECT 366.000 134.200 370.400 134.800 ;
        RECT 369.600 134.000 370.400 134.200 ;
        RECT 350.000 130.800 350.800 132.400 ;
        RECT 339.200 126.800 341.200 127.400 ;
        RECT 342.600 129.400 344.400 130.200 ;
        RECT 348.400 129.400 350.200 130.200 ;
        RECT 330.800 122.200 331.600 125.000 ;
        RECT 332.400 122.200 333.200 125.000 ;
        RECT 335.600 122.200 336.400 126.800 ;
        RECT 339.200 126.200 339.800 126.800 ;
        RECT 338.800 125.600 339.800 126.200 ;
        RECT 338.800 122.200 339.600 125.600 ;
        RECT 342.600 124.400 343.400 129.400 ;
        RECT 342.000 123.600 343.400 124.400 ;
        RECT 342.600 122.200 343.400 123.600 ;
        RECT 349.400 124.400 350.200 129.400 ;
        RECT 351.600 127.400 352.400 133.000 ;
        RECT 361.000 132.600 363.000 133.400 ;
        RECT 366.800 132.600 370.000 133.400 ;
        RECT 372.400 132.800 373.200 135.600 ;
        RECT 377.200 135.200 378.000 135.800 ;
        RECT 377.200 134.600 379.000 135.200 ;
        RECT 378.200 133.400 379.000 134.600 ;
        RECT 382.000 134.600 382.800 139.800 ;
        RECT 383.600 136.000 384.400 139.800 ;
        RECT 388.400 136.400 389.200 139.800 ;
        RECT 383.600 135.200 384.600 136.000 ;
        RECT 382.000 134.000 383.200 134.600 ;
        RECT 378.200 132.600 382.000 133.400 ;
        RECT 353.000 132.000 353.800 132.200 ;
        RECT 358.000 132.000 358.800 132.400 ;
        RECT 375.600 132.000 376.400 132.600 ;
        RECT 382.600 132.000 383.200 134.000 ;
        RECT 353.000 131.400 376.400 132.000 ;
        RECT 382.400 131.400 383.200 132.000 ;
        RECT 382.400 129.600 383.000 131.400 ;
        RECT 383.800 130.800 384.600 135.200 ;
        RECT 361.200 129.400 362.000 129.600 ;
        RECT 356.600 129.000 362.000 129.400 ;
        RECT 355.800 128.800 362.000 129.000 ;
        RECT 363.000 129.000 371.600 129.600 ;
        RECT 353.200 128.000 354.800 128.800 ;
        RECT 355.800 128.200 357.200 128.800 ;
        RECT 363.000 128.200 363.600 129.000 ;
        RECT 370.800 128.800 371.600 129.000 ;
        RECT 374.000 129.000 383.000 129.600 ;
        RECT 374.000 128.800 374.800 129.000 ;
        RECT 354.200 127.600 354.800 128.000 ;
        RECT 357.800 127.600 363.600 128.200 ;
        RECT 364.200 127.600 366.800 128.400 ;
        RECT 351.600 126.800 353.600 127.400 ;
        RECT 354.200 126.800 358.400 127.600 ;
        RECT 353.000 126.200 353.600 126.800 ;
        RECT 353.000 125.600 354.000 126.200 ;
        RECT 349.400 123.600 350.800 124.400 ;
        RECT 349.400 122.200 350.200 123.600 ;
        RECT 353.200 122.200 354.000 125.600 ;
        RECT 356.400 122.200 357.200 126.800 ;
        RECT 359.600 122.200 360.400 125.000 ;
        RECT 361.200 122.200 362.000 125.000 ;
        RECT 362.800 122.200 363.600 127.000 ;
        RECT 366.000 122.200 366.800 127.000 ;
        RECT 369.200 122.200 370.000 128.400 ;
        RECT 377.200 127.600 379.800 128.400 ;
        RECT 372.400 126.800 376.600 127.600 ;
        RECT 370.800 122.200 371.600 125.000 ;
        RECT 372.400 122.200 373.200 125.000 ;
        RECT 374.000 122.200 374.800 125.000 ;
        RECT 377.200 122.200 378.000 127.600 ;
        RECT 382.400 127.400 383.000 129.000 ;
        RECT 380.400 126.800 383.000 127.400 ;
        RECT 383.600 130.000 384.600 130.800 ;
        RECT 388.200 135.800 389.200 136.400 ;
        RECT 388.200 134.400 388.800 135.800 ;
        RECT 391.600 135.200 392.400 139.800 ;
        RECT 394.800 136.000 395.600 139.800 ;
        RECT 389.800 134.600 392.400 135.200 ;
        RECT 394.600 135.200 395.600 136.000 ;
        RECT 388.200 133.600 389.200 134.400 ;
        RECT 388.200 130.200 388.800 133.600 ;
        RECT 389.800 133.000 390.400 134.600 ;
        RECT 389.400 132.200 390.400 133.000 ;
        RECT 389.800 130.200 390.400 132.200 ;
        RECT 391.400 132.400 392.200 133.200 ;
        RECT 391.400 131.600 392.400 132.400 ;
        RECT 394.600 130.800 395.400 135.200 ;
        RECT 396.400 134.600 397.200 139.800 ;
        RECT 402.800 136.600 403.600 139.800 ;
        RECT 404.400 137.000 405.200 139.800 ;
        RECT 406.000 137.000 406.800 139.800 ;
        RECT 407.600 137.000 408.400 139.800 ;
        RECT 409.200 137.000 410.000 139.800 ;
        RECT 412.400 137.000 413.200 139.800 ;
        RECT 415.600 137.000 416.400 139.800 ;
        RECT 417.200 137.000 418.000 139.800 ;
        RECT 418.800 137.000 419.600 139.800 ;
        RECT 401.200 135.800 403.600 136.600 ;
        RECT 420.400 136.600 421.200 139.800 ;
        RECT 401.200 135.200 402.000 135.800 ;
        RECT 396.000 134.000 397.200 134.600 ;
        RECT 400.200 134.600 402.000 135.200 ;
        RECT 406.000 135.600 407.000 136.400 ;
        RECT 410.000 135.600 411.600 136.400 ;
        RECT 412.400 135.800 417.000 136.400 ;
        RECT 420.400 135.800 423.000 136.600 ;
        RECT 412.400 135.600 413.200 135.800 ;
        RECT 396.000 132.000 396.600 134.000 ;
        RECT 400.200 133.400 401.000 134.600 ;
        RECT 397.200 132.600 401.000 133.400 ;
        RECT 406.000 132.800 406.800 135.600 ;
        RECT 412.400 134.800 413.200 135.000 ;
        RECT 408.800 134.200 413.200 134.800 ;
        RECT 408.800 134.000 409.600 134.200 ;
        RECT 414.000 133.600 414.800 135.200 ;
        RECT 416.200 133.400 417.000 135.800 ;
        RECT 422.200 135.200 423.000 135.800 ;
        RECT 422.200 134.400 425.200 135.200 ;
        RECT 426.800 133.800 427.600 139.800 ;
        RECT 409.200 132.600 412.400 133.400 ;
        RECT 416.200 132.600 418.200 133.400 ;
        RECT 418.800 133.000 427.600 133.800 ;
        RECT 402.800 132.000 403.600 132.600 ;
        RECT 420.400 132.000 421.200 132.400 ;
        RECT 423.600 132.000 424.400 132.400 ;
        RECT 425.400 132.000 426.200 132.200 ;
        RECT 396.000 131.400 396.800 132.000 ;
        RECT 402.800 131.400 426.200 132.000 ;
        RECT 380.400 122.200 381.200 126.800 ;
        RECT 383.600 122.200 384.400 130.000 ;
        RECT 388.200 129.200 389.200 130.200 ;
        RECT 389.800 129.600 392.400 130.200 ;
        RECT 394.600 130.000 395.600 130.800 ;
        RECT 388.400 122.200 389.200 129.200 ;
        RECT 391.600 122.200 392.400 129.600 ;
        RECT 394.800 122.200 395.600 130.000 ;
        RECT 396.200 129.600 396.800 131.400 ;
        RECT 396.200 129.000 405.200 129.600 ;
        RECT 396.200 127.400 396.800 129.000 ;
        RECT 404.400 128.800 405.200 129.000 ;
        RECT 407.600 129.000 416.200 129.600 ;
        RECT 407.600 128.800 408.400 129.000 ;
        RECT 399.400 127.600 402.000 128.400 ;
        RECT 396.200 126.800 398.800 127.400 ;
        RECT 398.000 122.200 398.800 126.800 ;
        RECT 401.200 122.200 402.000 127.600 ;
        RECT 402.600 126.800 406.800 127.600 ;
        RECT 404.400 122.200 405.200 125.000 ;
        RECT 406.000 122.200 406.800 125.000 ;
        RECT 407.600 122.200 408.400 125.000 ;
        RECT 409.200 122.200 410.000 128.400 ;
        RECT 412.400 127.600 415.000 128.400 ;
        RECT 415.600 128.200 416.200 129.000 ;
        RECT 417.200 129.400 418.000 129.600 ;
        RECT 417.200 129.000 422.600 129.400 ;
        RECT 417.200 128.800 423.400 129.000 ;
        RECT 422.000 128.200 423.400 128.800 ;
        RECT 415.600 127.600 421.400 128.200 ;
        RECT 424.400 128.000 426.000 128.800 ;
        RECT 424.400 127.600 425.000 128.000 ;
        RECT 412.400 122.200 413.200 127.000 ;
        RECT 415.600 122.200 416.400 127.000 ;
        RECT 420.800 126.800 425.000 127.600 ;
        RECT 426.800 127.400 427.600 133.000 ;
        RECT 425.600 126.800 427.600 127.400 ;
        RECT 433.200 132.400 434.000 139.800 ;
        RECT 436.400 135.200 437.200 139.800 ;
        RECT 438.000 135.600 438.800 137.200 ;
        RECT 435.000 134.600 437.200 135.200 ;
        RECT 433.200 130.200 433.800 132.400 ;
        RECT 435.000 131.600 435.600 134.600 ;
        RECT 436.400 131.600 437.200 133.200 ;
        RECT 434.400 130.800 435.600 131.600 ;
        RECT 435.000 130.200 435.600 130.800 ;
        RECT 417.200 122.200 418.000 125.000 ;
        RECT 418.800 122.200 419.600 125.000 ;
        RECT 422.000 122.200 422.800 126.800 ;
        RECT 425.600 126.200 426.200 126.800 ;
        RECT 425.200 125.600 426.200 126.200 ;
        RECT 425.200 122.200 426.000 125.600 ;
        RECT 430.000 124.300 430.800 124.400 ;
        RECT 433.200 124.300 434.000 130.200 ;
        RECT 435.000 129.600 437.200 130.200 ;
        RECT 430.000 123.700 434.000 124.300 ;
        RECT 430.000 123.600 430.800 123.700 ;
        RECT 433.200 122.200 434.000 123.700 ;
        RECT 436.400 122.200 437.200 129.600 ;
        RECT 439.600 122.200 440.400 139.800 ;
        RECT 441.200 133.800 442.000 139.800 ;
        RECT 447.600 136.600 448.400 139.800 ;
        RECT 449.200 137.000 450.000 139.800 ;
        RECT 450.800 137.000 451.600 139.800 ;
        RECT 452.400 137.000 453.200 139.800 ;
        RECT 455.600 137.000 456.400 139.800 ;
        RECT 458.800 137.000 459.600 139.800 ;
        RECT 460.400 137.000 461.200 139.800 ;
        RECT 462.000 137.000 462.800 139.800 ;
        RECT 463.600 137.000 464.400 139.800 ;
        RECT 445.800 135.800 448.400 136.600 ;
        RECT 465.200 136.600 466.000 139.800 ;
        RECT 451.800 135.800 456.400 136.400 ;
        RECT 445.800 135.200 446.600 135.800 ;
        RECT 443.600 134.400 446.600 135.200 ;
        RECT 441.200 133.000 450.000 133.800 ;
        RECT 451.800 133.400 452.600 135.800 ;
        RECT 455.600 135.600 456.400 135.800 ;
        RECT 457.200 135.600 458.800 136.400 ;
        RECT 461.800 135.600 462.800 136.400 ;
        RECT 465.200 135.800 467.600 136.600 ;
        RECT 454.000 133.600 454.800 135.200 ;
        RECT 455.600 134.800 456.400 135.000 ;
        RECT 455.600 134.200 460.000 134.800 ;
        RECT 459.200 134.000 460.000 134.200 ;
        RECT 441.200 127.400 442.000 133.000 ;
        RECT 450.600 132.600 452.600 133.400 ;
        RECT 456.400 132.600 459.600 133.400 ;
        RECT 462.000 132.800 462.800 135.600 ;
        RECT 466.800 135.200 467.600 135.800 ;
        RECT 466.800 134.600 468.600 135.200 ;
        RECT 467.800 133.400 468.600 134.600 ;
        RECT 471.600 134.600 472.400 139.800 ;
        RECT 473.200 136.000 474.000 139.800 ;
        RECT 473.200 135.200 474.200 136.000 ;
        RECT 471.600 134.000 472.800 134.600 ;
        RECT 467.800 132.600 471.600 133.400 ;
        RECT 442.600 132.000 443.400 132.200 ;
        RECT 444.400 132.000 445.200 132.400 ;
        RECT 447.600 132.000 448.400 132.400 ;
        RECT 465.200 132.000 466.000 132.600 ;
        RECT 472.200 132.000 472.800 134.000 ;
        RECT 442.600 131.400 466.000 132.000 ;
        RECT 472.000 131.400 472.800 132.000 ;
        RECT 472.000 129.600 472.600 131.400 ;
        RECT 473.400 130.800 474.200 135.200 ;
        RECT 450.800 129.400 451.600 129.600 ;
        RECT 446.200 129.000 451.600 129.400 ;
        RECT 445.400 128.800 451.600 129.000 ;
        RECT 452.600 129.000 461.200 129.600 ;
        RECT 442.800 128.000 444.400 128.800 ;
        RECT 445.400 128.200 446.800 128.800 ;
        RECT 452.600 128.200 453.200 129.000 ;
        RECT 460.400 128.800 461.200 129.000 ;
        RECT 463.600 129.000 472.600 129.600 ;
        RECT 463.600 128.800 464.400 129.000 ;
        RECT 443.800 127.600 444.400 128.000 ;
        RECT 447.400 127.600 453.200 128.200 ;
        RECT 453.800 127.600 456.400 128.400 ;
        RECT 441.200 126.800 443.200 127.400 ;
        RECT 443.800 126.800 448.000 127.600 ;
        RECT 442.600 126.200 443.200 126.800 ;
        RECT 442.600 125.600 443.600 126.200 ;
        RECT 442.800 122.200 443.600 125.600 ;
        RECT 446.000 122.200 446.800 126.800 ;
        RECT 449.200 122.200 450.000 125.000 ;
        RECT 450.800 122.200 451.600 125.000 ;
        RECT 452.400 122.200 453.200 127.000 ;
        RECT 455.600 122.200 456.400 127.000 ;
        RECT 458.800 122.200 459.600 128.400 ;
        RECT 466.800 127.600 469.400 128.400 ;
        RECT 462.000 126.800 466.200 127.600 ;
        RECT 460.400 122.200 461.200 125.000 ;
        RECT 462.000 122.200 462.800 125.000 ;
        RECT 463.600 122.200 464.400 125.000 ;
        RECT 466.800 122.200 467.600 127.600 ;
        RECT 472.000 127.400 472.600 129.000 ;
        RECT 470.000 126.800 472.600 127.400 ;
        RECT 473.200 130.000 474.200 130.800 ;
        RECT 476.400 133.800 477.200 139.800 ;
        RECT 482.800 136.600 483.600 139.800 ;
        RECT 484.400 137.000 485.200 139.800 ;
        RECT 486.000 137.000 486.800 139.800 ;
        RECT 487.600 137.000 488.400 139.800 ;
        RECT 490.800 137.000 491.600 139.800 ;
        RECT 494.000 137.000 494.800 139.800 ;
        RECT 495.600 137.000 496.400 139.800 ;
        RECT 497.200 137.000 498.000 139.800 ;
        RECT 498.800 137.000 499.600 139.800 ;
        RECT 481.000 135.800 483.600 136.600 ;
        RECT 500.400 136.600 501.200 139.800 ;
        RECT 487.000 135.800 491.600 136.400 ;
        RECT 481.000 135.200 481.800 135.800 ;
        RECT 478.800 134.400 481.800 135.200 ;
        RECT 476.400 133.000 485.200 133.800 ;
        RECT 487.000 133.400 487.800 135.800 ;
        RECT 490.800 135.600 491.600 135.800 ;
        RECT 492.400 135.600 494.000 136.400 ;
        RECT 497.000 135.600 498.000 136.400 ;
        RECT 500.400 135.800 502.800 136.600 ;
        RECT 489.200 133.600 490.000 135.200 ;
        RECT 490.800 134.800 491.600 135.000 ;
        RECT 490.800 134.200 495.200 134.800 ;
        RECT 494.400 134.000 495.200 134.200 ;
        RECT 470.000 122.200 470.800 126.800 ;
        RECT 473.200 122.200 474.000 130.000 ;
        RECT 476.400 127.400 477.200 133.000 ;
        RECT 485.800 132.600 487.800 133.400 ;
        RECT 491.600 132.600 494.800 133.400 ;
        RECT 497.200 132.800 498.000 135.600 ;
        RECT 502.000 135.200 502.800 135.800 ;
        RECT 502.000 134.600 503.800 135.200 ;
        RECT 503.000 133.400 503.800 134.600 ;
        RECT 506.800 134.600 507.600 139.800 ;
        RECT 508.400 136.000 509.200 139.800 ;
        RECT 508.400 135.200 509.400 136.000 ;
        RECT 511.600 135.800 512.400 139.800 ;
        RECT 513.200 136.000 514.000 139.800 ;
        RECT 516.400 136.000 517.200 139.800 ;
        RECT 513.200 135.800 517.200 136.000 ;
        RECT 506.800 134.000 508.000 134.600 ;
        RECT 503.000 132.600 506.800 133.400 ;
        RECT 477.800 132.000 478.600 132.200 ;
        RECT 482.800 132.000 483.600 132.400 ;
        RECT 500.400 132.000 501.200 132.600 ;
        RECT 507.400 132.000 508.000 134.000 ;
        RECT 477.800 131.400 501.200 132.000 ;
        RECT 507.200 131.400 508.000 132.000 ;
        RECT 507.200 129.600 507.800 131.400 ;
        RECT 508.600 130.800 509.400 135.200 ;
        RECT 511.800 134.400 512.400 135.800 ;
        RECT 513.400 135.400 517.000 135.800 ;
        RECT 518.000 135.400 518.800 139.800 ;
        RECT 522.200 138.400 523.400 139.800 ;
        RECT 522.200 137.800 523.600 138.400 ;
        RECT 526.800 137.800 527.600 139.800 ;
        RECT 531.200 138.400 532.000 139.800 ;
        RECT 531.200 137.800 533.200 138.400 ;
        RECT 522.800 137.000 523.600 137.800 ;
        RECT 527.000 137.200 527.600 137.800 ;
        RECT 527.000 136.600 529.800 137.200 ;
        RECT 529.000 136.400 529.800 136.600 ;
        RECT 530.800 136.400 531.600 137.200 ;
        RECT 532.400 137.000 533.200 137.800 ;
        RECT 521.000 135.400 521.800 135.600 ;
        RECT 518.000 134.800 521.800 135.400 ;
        RECT 515.600 134.400 516.400 134.800 ;
        RECT 511.600 133.600 514.200 134.400 ;
        RECT 515.600 133.800 517.200 134.400 ;
        RECT 516.400 133.600 517.200 133.800 ;
        RECT 486.000 129.400 486.800 129.600 ;
        RECT 481.400 129.000 486.800 129.400 ;
        RECT 480.600 128.800 486.800 129.000 ;
        RECT 487.800 129.000 496.400 129.600 ;
        RECT 478.000 128.000 479.600 128.800 ;
        RECT 480.600 128.200 482.000 128.800 ;
        RECT 487.800 128.200 488.400 129.000 ;
        RECT 495.600 128.800 496.400 129.000 ;
        RECT 498.800 129.000 507.800 129.600 ;
        RECT 498.800 128.800 499.600 129.000 ;
        RECT 479.000 127.600 479.600 128.000 ;
        RECT 482.600 127.600 488.400 128.200 ;
        RECT 489.000 127.600 491.600 128.400 ;
        RECT 476.400 126.800 478.400 127.400 ;
        RECT 479.000 126.800 483.200 127.600 ;
        RECT 477.800 126.200 478.400 126.800 ;
        RECT 477.800 125.600 478.800 126.200 ;
        RECT 478.000 122.200 478.800 125.600 ;
        RECT 481.200 122.200 482.000 126.800 ;
        RECT 484.400 122.200 485.200 125.000 ;
        RECT 486.000 122.200 486.800 125.000 ;
        RECT 487.600 122.200 488.400 127.000 ;
        RECT 490.800 122.200 491.600 127.000 ;
        RECT 494.000 122.200 494.800 128.400 ;
        RECT 502.000 127.600 504.600 128.400 ;
        RECT 497.200 126.800 501.400 127.600 ;
        RECT 495.600 122.200 496.400 125.000 ;
        RECT 497.200 122.200 498.000 125.000 ;
        RECT 498.800 122.200 499.600 125.000 ;
        RECT 502.000 122.200 502.800 127.600 ;
        RECT 507.200 127.400 507.800 129.000 ;
        RECT 505.200 126.800 507.800 127.400 ;
        RECT 508.400 130.000 509.400 130.800 ;
        RECT 510.000 130.300 510.800 130.400 ;
        RECT 511.600 130.300 512.400 130.400 ;
        RECT 510.000 130.200 512.400 130.300 ;
        RECT 513.600 130.200 514.200 133.600 ;
        RECT 514.800 131.600 515.600 133.200 ;
        RECT 518.000 131.400 518.800 134.800 ;
        RECT 525.000 134.200 525.800 134.400 ;
        RECT 530.800 134.200 531.400 136.400 ;
        RECT 535.600 135.000 536.400 139.800 ;
        RECT 537.200 135.200 538.000 139.800 ;
        RECT 540.400 136.400 541.200 139.800 ;
        RECT 540.400 135.600 541.400 136.400 ;
        RECT 543.600 136.000 544.400 139.800 ;
        RECT 546.800 136.000 547.600 139.800 ;
        RECT 543.600 135.800 547.600 136.000 ;
        RECT 548.400 135.800 549.200 139.800 ;
        RECT 550.000 135.800 550.800 139.800 ;
        RECT 551.600 136.000 552.400 139.800 ;
        RECT 554.800 136.000 555.600 139.800 ;
        RECT 558.000 137.800 558.800 139.800 ;
        RECT 551.600 135.800 555.600 136.000 ;
        RECT 537.200 134.600 539.800 135.200 ;
        RECT 534.000 134.200 535.600 134.400 ;
        RECT 524.600 133.600 535.600 134.200 ;
        RECT 522.800 132.800 523.600 133.000 ;
        RECT 519.800 132.200 523.600 132.800 ;
        RECT 519.800 132.000 520.600 132.200 ;
        RECT 521.400 131.400 522.200 131.600 ;
        RECT 518.000 130.800 522.200 131.400 ;
        RECT 505.200 122.200 506.000 126.800 ;
        RECT 508.400 122.200 509.200 130.000 ;
        RECT 510.000 129.700 513.000 130.200 ;
        RECT 510.000 129.600 510.800 129.700 ;
        RECT 511.600 129.600 513.000 129.700 ;
        RECT 513.600 129.600 514.600 130.200 ;
        RECT 512.400 128.400 513.000 129.600 ;
        RECT 512.400 127.600 513.200 128.400 ;
        RECT 513.800 122.200 514.600 129.600 ;
        RECT 518.000 122.200 518.800 130.800 ;
        RECT 524.600 130.400 525.200 133.600 ;
        RECT 531.800 133.400 532.600 133.600 ;
        RECT 530.800 132.400 531.600 132.600 ;
        RECT 533.400 132.400 534.200 132.600 ;
        RECT 537.400 132.400 538.200 133.200 ;
        RECT 529.200 131.800 534.200 132.400 ;
        RECT 529.200 131.600 530.000 131.800 ;
        RECT 537.200 131.600 538.200 132.400 ;
        RECT 539.200 133.000 539.800 134.600 ;
        RECT 540.800 134.400 541.400 135.600 ;
        RECT 543.800 135.400 547.400 135.800 ;
        RECT 544.400 134.400 545.200 134.800 ;
        RECT 548.400 134.400 549.000 135.800 ;
        RECT 550.200 134.400 550.800 135.800 ;
        RECT 551.800 135.400 555.400 135.800 ;
        RECT 556.400 135.600 557.200 137.200 ;
        RECT 554.000 134.400 554.800 134.800 ;
        RECT 558.200 134.400 558.800 137.800 ;
        RECT 561.200 135.000 562.000 139.800 ;
        RECT 565.600 138.400 566.400 139.800 ;
        RECT 564.400 137.800 566.400 138.400 ;
        RECT 570.000 137.800 570.800 139.800 ;
        RECT 574.200 138.400 575.400 139.800 ;
        RECT 574.000 137.800 575.400 138.400 ;
        RECT 578.800 138.300 579.600 139.800 ;
        RECT 585.800 138.400 586.600 139.800 ;
        RECT 583.600 138.300 584.400 138.400 ;
        RECT 564.400 137.000 565.200 137.800 ;
        RECT 570.000 137.200 570.600 137.800 ;
        RECT 566.000 136.400 566.800 137.200 ;
        RECT 567.800 136.600 570.600 137.200 ;
        RECT 574.000 137.000 574.800 137.800 ;
        RECT 578.800 137.700 584.400 138.300 ;
        RECT 567.800 136.400 568.600 136.600 ;
        RECT 540.400 133.600 541.400 134.400 ;
        RECT 543.600 133.800 545.200 134.400 ;
        RECT 543.600 133.600 544.400 133.800 ;
        RECT 546.600 133.600 549.200 134.400 ;
        RECT 550.000 133.600 552.600 134.400 ;
        RECT 554.000 133.800 555.600 134.400 ;
        RECT 554.800 133.600 555.600 133.800 ;
        RECT 558.000 133.600 558.800 134.400 ;
        RECT 562.000 134.200 563.600 134.400 ;
        RECT 566.200 134.200 566.800 136.400 ;
        RECT 575.800 135.400 576.600 135.600 ;
        RECT 578.800 135.400 579.600 137.700 ;
        RECT 583.600 137.600 584.400 137.700 ;
        RECT 585.200 137.600 586.600 138.400 ;
        RECT 585.800 136.400 586.600 137.600 ;
        RECT 585.800 135.800 587.600 136.400 ;
        RECT 575.800 134.800 579.600 135.400 ;
        RECT 571.800 134.200 572.600 134.400 ;
        RECT 562.000 133.600 573.000 134.200 ;
        RECT 539.200 132.200 540.200 133.000 ;
        RECT 530.800 131.000 536.400 131.200 ;
        RECT 530.600 130.800 536.400 131.000 ;
        RECT 522.800 129.800 525.200 130.400 ;
        RECT 526.600 130.600 536.400 130.800 ;
        RECT 526.600 130.200 531.400 130.600 ;
        RECT 522.800 128.800 523.400 129.800 ;
        RECT 522.000 128.000 523.400 128.800 ;
        RECT 525.000 129.000 525.800 129.200 ;
        RECT 526.600 129.000 527.200 130.200 ;
        RECT 525.000 128.400 527.200 129.000 ;
        RECT 527.800 129.000 533.200 129.600 ;
        RECT 527.800 128.800 528.600 129.000 ;
        RECT 532.400 128.800 533.200 129.000 ;
        RECT 526.200 127.400 527.000 127.600 ;
        RECT 529.000 127.400 529.800 127.600 ;
        RECT 522.800 126.200 523.600 127.000 ;
        RECT 526.200 126.800 529.800 127.400 ;
        RECT 527.000 126.200 527.600 126.800 ;
        RECT 532.400 126.200 533.200 127.000 ;
        RECT 522.200 122.200 523.400 126.200 ;
        RECT 526.800 122.200 527.600 126.200 ;
        RECT 531.200 125.600 533.200 126.200 ;
        RECT 531.200 122.200 532.000 125.600 ;
        RECT 535.600 122.200 536.400 130.600 ;
        RECT 539.200 130.200 539.800 132.200 ;
        RECT 540.800 130.200 541.400 133.600 ;
        RECT 545.200 131.600 546.000 133.200 ;
        RECT 546.600 132.400 547.200 133.600 ;
        RECT 546.600 131.600 547.600 132.400 ;
        RECT 552.000 132.300 552.600 133.600 ;
        RECT 548.500 131.700 552.600 132.300 ;
        RECT 546.600 130.200 547.200 131.600 ;
        RECT 548.500 130.400 549.100 131.700 ;
        RECT 548.400 130.200 549.200 130.400 ;
        RECT 537.200 129.600 539.800 130.200 ;
        RECT 537.200 122.200 538.000 129.600 ;
        RECT 540.400 129.200 541.400 130.200 ;
        RECT 546.200 129.600 547.200 130.200 ;
        RECT 547.800 129.600 549.200 130.200 ;
        RECT 550.000 130.200 550.800 130.400 ;
        RECT 552.000 130.200 552.600 131.700 ;
        RECT 553.200 131.600 554.000 133.200 ;
        RECT 558.200 130.200 558.800 133.600 ;
        RECT 565.000 133.400 565.800 133.600 ;
        RECT 563.400 132.400 564.200 132.600 ;
        RECT 572.400 132.400 573.000 133.600 ;
        RECT 574.000 132.800 574.800 133.000 ;
        RECT 559.600 130.800 560.400 132.400 ;
        RECT 563.400 131.800 568.400 132.400 ;
        RECT 567.600 131.600 568.400 131.800 ;
        RECT 572.400 131.600 573.200 132.400 ;
        RECT 574.000 132.200 577.800 132.800 ;
        RECT 577.000 132.000 577.800 132.200 ;
        RECT 561.200 131.000 566.800 131.200 ;
        RECT 561.200 130.800 567.000 131.000 ;
        RECT 561.200 130.600 571.000 130.800 ;
        RECT 550.000 129.600 551.400 130.200 ;
        RECT 552.000 129.600 553.000 130.200 ;
        RECT 540.400 122.200 541.200 129.200 ;
        RECT 546.200 122.200 547.000 129.600 ;
        RECT 547.800 128.400 548.400 129.600 ;
        RECT 547.600 127.600 548.400 128.400 ;
        RECT 550.800 128.400 551.400 129.600 ;
        RECT 550.800 127.600 551.600 128.400 ;
        RECT 552.200 122.200 553.000 129.600 ;
        RECT 558.000 129.400 559.800 130.200 ;
        RECT 559.000 124.400 559.800 129.400 ;
        RECT 558.000 123.600 559.800 124.400 ;
        RECT 559.000 122.200 559.800 123.600 ;
        RECT 561.200 122.200 562.000 130.600 ;
        RECT 566.200 130.200 571.000 130.600 ;
        RECT 564.400 129.000 569.800 129.600 ;
        RECT 564.400 128.800 565.200 129.000 ;
        RECT 569.000 128.800 569.800 129.000 ;
        RECT 570.400 129.000 571.000 130.200 ;
        RECT 572.400 130.400 573.000 131.600 ;
        RECT 575.400 131.400 576.200 131.600 ;
        RECT 578.800 131.400 579.600 134.800 ;
        RECT 575.400 130.800 579.600 131.400 ;
        RECT 572.400 129.800 574.800 130.400 ;
        RECT 571.800 129.000 572.600 129.200 ;
        RECT 570.400 128.400 572.600 129.000 ;
        RECT 574.200 128.800 574.800 129.800 ;
        RECT 574.200 128.000 575.600 128.800 ;
        RECT 567.800 127.400 568.600 127.600 ;
        RECT 570.600 127.400 571.400 127.600 ;
        RECT 564.400 126.200 565.200 127.000 ;
        RECT 567.800 126.800 571.400 127.400 ;
        RECT 570.000 126.200 570.600 126.800 ;
        RECT 574.000 126.200 574.800 127.000 ;
        RECT 564.400 125.600 566.400 126.200 ;
        RECT 565.600 122.200 566.400 125.600 ;
        RECT 570.000 122.200 570.800 126.200 ;
        RECT 574.200 122.200 575.400 126.200 ;
        RECT 578.800 122.200 579.600 130.800 ;
        RECT 585.200 128.800 586.000 130.400 ;
        RECT 586.800 122.200 587.600 135.800 ;
        RECT 588.400 133.600 589.200 135.200 ;
        RECT 591.200 134.200 592.000 139.800 ;
        RECT 596.400 135.800 597.200 139.800 ;
        RECT 598.000 136.000 598.800 139.800 ;
        RECT 601.200 136.000 602.000 139.800 ;
        RECT 598.000 135.800 602.000 136.000 ;
        RECT 602.800 137.000 603.600 139.000 ;
        RECT 596.600 134.400 597.200 135.800 ;
        RECT 598.200 135.400 601.800 135.800 ;
        RECT 602.800 134.800 603.400 137.000 ;
        RECT 607.000 136.000 607.800 139.000 ;
        RECT 612.400 136.000 613.200 139.800 ;
        RECT 615.600 136.000 616.400 139.800 ;
        RECT 607.000 135.400 608.600 136.000 ;
        RECT 612.400 135.800 616.400 136.000 ;
        RECT 617.200 135.800 618.000 139.800 ;
        RECT 618.800 136.000 619.600 139.800 ;
        RECT 622.000 136.000 622.800 139.800 ;
        RECT 618.800 135.800 622.800 136.000 ;
        RECT 623.600 135.800 624.400 139.800 ;
        RECT 612.600 135.400 616.200 135.800 ;
        RECT 607.800 135.000 608.600 135.400 ;
        RECT 600.400 134.400 601.200 134.800 ;
        RECT 590.200 133.800 592.000 134.200 ;
        RECT 590.200 133.600 591.800 133.800 ;
        RECT 596.400 133.600 599.000 134.400 ;
        RECT 600.400 133.800 602.000 134.400 ;
        RECT 602.800 134.200 607.000 134.800 ;
        RECT 601.200 133.600 602.000 133.800 ;
        RECT 606.000 133.800 607.000 134.200 ;
        RECT 608.000 134.400 608.600 135.000 ;
        RECT 613.200 134.400 614.000 134.800 ;
        RECT 617.200 134.400 617.800 135.800 ;
        RECT 619.000 135.400 622.600 135.800 ;
        RECT 619.600 134.400 620.400 134.800 ;
        RECT 623.600 134.400 624.200 135.800 ;
        RECT 625.200 135.400 626.000 139.800 ;
        RECT 629.400 138.400 630.600 139.800 ;
        RECT 629.400 137.800 630.800 138.400 ;
        RECT 634.000 137.800 634.800 139.800 ;
        RECT 638.400 138.400 639.200 139.800 ;
        RECT 638.400 137.800 640.400 138.400 ;
        RECT 630.000 137.000 630.800 137.800 ;
        RECT 634.200 137.200 634.800 137.800 ;
        RECT 634.200 136.600 637.000 137.200 ;
        RECT 636.200 136.400 637.000 136.600 ;
        RECT 638.000 136.400 638.800 137.200 ;
        RECT 639.600 137.000 640.400 137.800 ;
        RECT 628.200 135.400 629.000 135.600 ;
        RECT 625.200 134.800 629.000 135.400 ;
        RECT 608.000 134.300 610.000 134.400 ;
        RECT 590.200 130.400 590.800 133.600 ;
        RECT 592.400 131.600 594.000 132.400 ;
        RECT 590.000 129.600 590.800 130.400 ;
        RECT 594.800 129.600 595.600 131.200 ;
        RECT 596.400 130.200 597.200 130.400 ;
        RECT 598.400 130.200 599.000 133.600 ;
        RECT 599.600 131.600 600.400 133.200 ;
        RECT 601.200 132.300 602.000 132.400 ;
        RECT 602.800 132.300 603.600 133.200 ;
        RECT 601.200 131.700 603.600 132.300 ;
        RECT 601.200 131.600 602.000 131.700 ;
        RECT 602.800 131.600 603.600 131.700 ;
        RECT 604.400 131.600 605.200 133.200 ;
        RECT 606.000 133.000 607.400 133.800 ;
        RECT 608.000 133.700 611.500 134.300 ;
        RECT 608.000 133.600 610.000 133.700 ;
        RECT 606.000 131.000 606.600 133.000 ;
        RECT 602.800 130.400 606.600 131.000 ;
        RECT 596.400 129.600 597.800 130.200 ;
        RECT 598.400 129.600 599.400 130.200 ;
        RECT 590.200 127.000 590.800 129.600 ;
        RECT 591.600 128.300 592.400 129.200 ;
        RECT 597.200 128.400 597.800 129.600 ;
        RECT 594.800 128.300 595.600 128.400 ;
        RECT 591.600 127.700 595.600 128.300 ;
        RECT 591.600 127.600 592.400 127.700 ;
        RECT 594.800 127.600 595.600 127.700 ;
        RECT 597.200 127.600 598.000 128.400 ;
        RECT 590.200 126.400 593.800 127.000 ;
        RECT 590.200 126.200 590.800 126.400 ;
        RECT 590.000 122.200 590.800 126.200 ;
        RECT 593.200 126.200 593.800 126.400 ;
        RECT 593.200 122.200 594.000 126.200 ;
        RECT 598.600 122.200 599.400 129.600 ;
        RECT 602.800 127.000 603.400 130.400 ;
        RECT 608.000 129.800 608.600 133.600 ;
        RECT 609.200 130.800 610.000 132.400 ;
        RECT 610.900 132.300 611.500 133.700 ;
        RECT 612.400 133.800 614.000 134.400 ;
        RECT 612.400 133.600 613.200 133.800 ;
        RECT 615.400 133.600 618.000 134.400 ;
        RECT 618.800 133.800 620.400 134.400 ;
        RECT 618.800 133.600 619.600 133.800 ;
        RECT 621.800 133.600 624.400 134.400 ;
        RECT 614.000 132.300 614.800 133.200 ;
        RECT 610.900 131.700 614.800 132.300 ;
        RECT 614.000 131.600 614.800 131.700 ;
        RECT 615.400 130.200 616.000 133.600 ;
        RECT 620.400 131.600 621.200 133.200 ;
        RECT 621.800 130.400 622.400 133.600 ;
        RECT 625.200 131.400 626.000 134.800 ;
        RECT 632.200 134.200 633.000 134.400 ;
        RECT 638.000 134.200 638.600 136.400 ;
        RECT 642.800 135.000 643.600 139.800 ;
        RECT 641.200 134.200 642.800 134.400 ;
        RECT 631.800 133.600 642.800 134.200 ;
        RECT 630.000 132.800 630.800 133.000 ;
        RECT 627.000 132.200 630.800 132.800 ;
        RECT 627.000 132.000 627.800 132.200 ;
        RECT 628.600 131.400 629.400 131.600 ;
        RECT 625.200 130.800 629.400 131.400 ;
        RECT 617.200 130.200 618.000 130.400 ;
        RECT 607.000 129.200 608.600 129.800 ;
        RECT 615.000 129.600 616.000 130.200 ;
        RECT 616.600 129.600 618.000 130.200 ;
        RECT 620.400 129.600 622.400 130.400 ;
        RECT 623.600 130.300 624.400 130.400 ;
        RECT 625.200 130.300 626.000 130.800 ;
        RECT 631.800 130.400 632.400 133.600 ;
        RECT 639.000 133.400 639.800 133.600 ;
        RECT 640.600 132.400 641.400 132.600 ;
        RECT 633.200 132.300 634.000 132.400 ;
        RECT 636.400 132.300 641.400 132.400 ;
        RECT 633.200 131.800 641.400 132.300 ;
        RECT 633.200 131.700 637.200 131.800 ;
        RECT 633.200 131.600 634.000 131.700 ;
        RECT 636.400 131.600 637.200 131.700 ;
        RECT 638.000 131.000 643.600 131.200 ;
        RECT 637.800 130.800 643.600 131.000 ;
        RECT 623.600 130.200 626.000 130.300 ;
        RECT 623.000 129.700 626.000 130.200 ;
        RECT 623.000 129.600 624.400 129.700 ;
        RECT 602.800 123.000 603.600 127.000 ;
        RECT 607.000 122.200 607.800 129.200 ;
        RECT 615.000 122.200 615.800 129.600 ;
        RECT 616.600 128.400 617.200 129.600 ;
        RECT 616.400 127.600 617.200 128.400 ;
        RECT 621.400 122.200 622.200 129.600 ;
        RECT 623.000 128.400 623.600 129.600 ;
        RECT 622.800 127.600 623.600 128.400 ;
        RECT 625.200 122.200 626.000 129.700 ;
        RECT 630.000 129.800 632.400 130.400 ;
        RECT 633.800 130.600 643.600 130.800 ;
        RECT 633.800 130.200 638.600 130.600 ;
        RECT 630.000 128.800 630.600 129.800 ;
        RECT 629.200 128.000 630.600 128.800 ;
        RECT 632.200 129.000 633.000 129.200 ;
        RECT 633.800 129.000 634.400 130.200 ;
        RECT 632.200 128.400 634.400 129.000 ;
        RECT 635.000 129.000 640.400 129.600 ;
        RECT 635.000 128.800 635.800 129.000 ;
        RECT 639.600 128.800 640.400 129.000 ;
        RECT 633.400 127.400 634.200 127.600 ;
        RECT 636.200 127.400 637.000 127.600 ;
        RECT 630.000 126.200 630.800 127.000 ;
        RECT 633.400 126.800 637.000 127.400 ;
        RECT 634.200 126.200 634.800 126.800 ;
        RECT 639.600 126.200 640.400 127.000 ;
        RECT 629.400 122.200 630.600 126.200 ;
        RECT 634.000 122.200 634.800 126.200 ;
        RECT 638.400 125.600 640.400 126.200 ;
        RECT 638.400 122.200 639.200 125.600 ;
        RECT 642.800 122.200 643.600 130.600 ;
        RECT 644.400 122.200 645.200 139.800 ;
        RECT 646.000 135.600 646.800 137.200 ;
        RECT 647.600 137.000 648.400 139.000 ;
        RECT 647.600 134.800 648.200 137.000 ;
        RECT 651.800 136.000 652.600 139.000 ;
        RECT 651.800 135.400 653.400 136.000 ;
        RECT 652.600 135.000 653.400 135.400 ;
        RECT 647.600 134.200 651.800 134.800 ;
        RECT 650.800 133.800 651.800 134.200 ;
        RECT 652.800 134.400 653.400 135.000 ;
        RECT 657.200 135.200 658.000 139.800 ;
        RECT 660.400 136.400 661.200 139.800 ;
        RECT 660.400 135.800 661.400 136.400 ;
        RECT 663.600 136.000 664.400 139.800 ;
        RECT 666.800 136.000 667.600 139.800 ;
        RECT 663.600 135.800 667.600 136.000 ;
        RECT 668.400 135.800 669.200 139.800 ;
        RECT 657.200 134.600 659.800 135.200 ;
        RECT 647.600 131.600 648.400 133.200 ;
        RECT 649.200 131.600 650.000 133.200 ;
        RECT 650.800 133.000 652.200 133.800 ;
        RECT 652.800 133.600 654.800 134.400 ;
        RECT 650.800 131.000 651.400 133.000 ;
        RECT 647.600 130.400 651.400 131.000 ;
        RECT 647.600 127.000 648.200 130.400 ;
        RECT 652.800 129.800 653.400 133.600 ;
        RECT 657.400 132.400 658.200 133.200 ;
        RECT 654.000 130.800 654.800 132.400 ;
        RECT 657.200 131.600 658.200 132.400 ;
        RECT 659.200 133.000 659.800 134.600 ;
        RECT 660.800 134.400 661.400 135.800 ;
        RECT 663.800 135.400 667.400 135.800 ;
        RECT 664.400 134.400 665.200 134.800 ;
        RECT 668.400 134.400 669.000 135.800 ;
        RECT 670.000 135.400 670.800 139.800 ;
        RECT 674.200 138.400 675.400 139.800 ;
        RECT 674.200 137.800 675.600 138.400 ;
        RECT 678.800 137.800 679.600 139.800 ;
        RECT 683.200 138.400 684.000 139.800 ;
        RECT 683.200 137.800 685.200 138.400 ;
        RECT 674.800 137.000 675.600 137.800 ;
        RECT 679.000 137.200 679.600 137.800 ;
        RECT 679.000 136.600 681.800 137.200 ;
        RECT 681.000 136.400 681.800 136.600 ;
        RECT 682.800 135.600 683.600 137.200 ;
        RECT 684.400 137.000 685.200 137.800 ;
        RECT 673.000 135.400 673.800 135.600 ;
        RECT 670.000 134.800 673.800 135.400 ;
        RECT 660.400 134.300 661.400 134.400 ;
        RECT 663.600 134.300 665.200 134.400 ;
        RECT 660.400 133.800 665.200 134.300 ;
        RECT 660.400 133.700 664.400 133.800 ;
        RECT 660.400 133.600 661.400 133.700 ;
        RECT 663.600 133.600 664.400 133.700 ;
        RECT 666.600 133.600 669.200 134.400 ;
        RECT 659.200 132.200 660.200 133.000 ;
        RECT 659.200 130.200 659.800 132.200 ;
        RECT 660.800 130.200 661.400 133.600 ;
        RECT 665.200 131.600 666.000 133.200 ;
        RECT 666.600 132.300 667.200 133.600 ;
        RECT 668.400 132.300 669.200 132.400 ;
        RECT 666.600 131.700 669.200 132.300 ;
        RECT 666.600 130.200 667.200 131.700 ;
        RECT 668.400 131.600 669.200 131.700 ;
        RECT 670.000 131.400 670.800 134.800 ;
        RECT 677.000 134.200 677.800 134.400 ;
        RECT 682.800 134.200 683.400 135.600 ;
        RECT 687.600 135.000 688.400 139.800 ;
        RECT 686.000 134.200 687.600 134.400 ;
        RECT 676.600 133.600 687.600 134.200 ;
        RECT 674.800 132.800 675.600 133.000 ;
        RECT 671.800 132.200 675.600 132.800 ;
        RECT 671.800 132.000 672.600 132.200 ;
        RECT 673.400 131.400 674.200 131.600 ;
        RECT 670.000 130.800 674.200 131.400 ;
        RECT 668.400 130.200 669.200 130.400 ;
        RECT 651.800 129.200 653.400 129.800 ;
        RECT 657.200 129.600 659.800 130.200 ;
        RECT 647.600 123.000 648.400 127.000 ;
        RECT 651.800 124.400 652.600 129.200 ;
        RECT 651.800 123.600 653.200 124.400 ;
        RECT 651.800 122.200 652.600 123.600 ;
        RECT 657.200 122.200 658.000 129.600 ;
        RECT 660.400 129.200 661.400 130.200 ;
        RECT 666.200 129.600 667.200 130.200 ;
        RECT 667.800 129.600 669.200 130.200 ;
        RECT 660.400 122.200 661.200 129.200 ;
        RECT 666.200 122.200 667.000 129.600 ;
        RECT 667.800 128.400 668.400 129.600 ;
        RECT 667.600 127.600 668.400 128.400 ;
        RECT 670.000 122.200 670.800 130.800 ;
        RECT 676.600 130.400 677.200 133.600 ;
        RECT 683.800 133.400 684.600 133.600 ;
        RECT 685.400 132.400 686.200 132.600 ;
        RECT 679.600 132.300 680.400 132.400 ;
        RECT 681.200 132.300 686.200 132.400 ;
        RECT 679.600 131.800 686.200 132.300 ;
        RECT 679.600 131.700 682.000 131.800 ;
        RECT 679.600 131.600 680.400 131.700 ;
        RECT 681.200 131.600 682.000 131.700 ;
        RECT 682.800 131.000 688.400 131.200 ;
        RECT 682.600 130.800 688.400 131.000 ;
        RECT 674.800 129.800 677.200 130.400 ;
        RECT 678.600 130.600 688.400 130.800 ;
        RECT 678.600 130.200 683.400 130.600 ;
        RECT 674.800 128.800 675.400 129.800 ;
        RECT 674.000 128.000 675.400 128.800 ;
        RECT 677.000 129.000 677.800 129.200 ;
        RECT 678.600 129.000 679.200 130.200 ;
        RECT 677.000 128.400 679.200 129.000 ;
        RECT 679.800 129.000 685.200 129.600 ;
        RECT 679.800 128.800 680.600 129.000 ;
        RECT 684.400 128.800 685.200 129.000 ;
        RECT 678.200 127.400 679.000 127.600 ;
        RECT 681.000 127.400 681.800 127.600 ;
        RECT 674.800 126.200 675.600 127.000 ;
        RECT 678.200 126.800 681.800 127.400 ;
        RECT 679.000 126.200 679.600 126.800 ;
        RECT 684.400 126.200 685.200 127.000 ;
        RECT 674.200 122.200 675.400 126.200 ;
        RECT 678.800 122.200 679.600 126.200 ;
        RECT 683.200 125.600 685.200 126.200 ;
        RECT 683.200 122.200 684.000 125.600 ;
        RECT 687.600 122.200 688.400 130.600 ;
        RECT 1.200 111.400 2.000 119.800 ;
        RECT 5.600 116.400 6.400 119.800 ;
        RECT 4.400 115.800 6.400 116.400 ;
        RECT 10.000 115.800 10.800 119.800 ;
        RECT 14.200 115.800 15.400 119.800 ;
        RECT 4.400 115.000 5.200 115.800 ;
        RECT 10.000 115.200 10.600 115.800 ;
        RECT 7.800 114.600 11.400 115.200 ;
        RECT 14.000 115.000 14.800 115.800 ;
        RECT 7.800 114.400 8.600 114.600 ;
        RECT 10.600 114.400 11.400 114.600 ;
        RECT 4.400 113.000 5.200 113.200 ;
        RECT 9.000 113.000 9.800 113.200 ;
        RECT 4.400 112.400 9.800 113.000 ;
        RECT 10.400 113.000 12.600 113.600 ;
        RECT 10.400 111.800 11.000 113.000 ;
        RECT 11.800 112.800 12.600 113.000 ;
        RECT 14.200 113.200 15.600 114.000 ;
        RECT 14.200 112.200 14.800 113.200 ;
        RECT 6.200 111.400 11.000 111.800 ;
        RECT 1.200 111.200 11.000 111.400 ;
        RECT 12.400 111.600 14.800 112.200 ;
        RECT 1.200 111.000 7.000 111.200 ;
        RECT 1.200 110.800 6.800 111.000 ;
        RECT 12.400 110.400 13.000 111.600 ;
        RECT 18.800 111.200 19.600 119.800 ;
        RECT 22.000 112.800 22.800 119.800 ;
        RECT 15.400 110.600 19.600 111.200 ;
        RECT 15.400 110.400 16.200 110.600 ;
        RECT 7.600 110.200 8.400 110.400 ;
        RECT 3.400 109.600 8.400 110.200 ;
        RECT 12.400 109.600 13.200 110.400 ;
        RECT 17.000 109.800 17.800 110.000 ;
        RECT 3.400 109.400 4.200 109.600 ;
        RECT 6.000 109.400 6.800 109.600 ;
        RECT 5.000 108.400 5.800 108.600 ;
        RECT 12.400 108.400 13.000 109.600 ;
        RECT 14.000 109.200 17.800 109.800 ;
        RECT 14.000 109.000 14.800 109.200 ;
        RECT 2.000 107.800 13.000 108.400 ;
        RECT 2.000 107.600 3.600 107.800 ;
        RECT 1.200 102.200 2.000 107.000 ;
        RECT 6.200 105.600 6.800 107.800 ;
        RECT 11.800 107.600 12.600 107.800 ;
        RECT 18.800 107.200 19.600 110.600 ;
        RECT 15.800 106.600 19.600 107.200 ;
        RECT 15.800 106.400 16.600 106.600 ;
        RECT 4.400 104.200 5.200 105.000 ;
        RECT 6.000 104.800 6.800 105.600 ;
        RECT 7.800 105.400 8.600 105.600 ;
        RECT 7.800 104.800 10.600 105.400 ;
        RECT 10.000 104.200 10.600 104.800 ;
        RECT 14.000 104.200 14.800 105.000 ;
        RECT 4.400 103.600 6.400 104.200 ;
        RECT 5.600 102.200 6.400 103.600 ;
        RECT 10.000 102.200 10.800 104.200 ;
        RECT 14.000 103.600 15.400 104.200 ;
        RECT 14.200 102.200 15.400 103.600 ;
        RECT 18.800 102.200 19.600 106.600 ;
        RECT 21.800 111.800 22.800 112.800 ;
        RECT 25.200 112.400 26.000 119.800 ;
        RECT 23.400 111.800 26.000 112.400 ;
        RECT 26.800 115.000 27.600 119.000 ;
        RECT 31.000 118.400 31.800 119.800 ;
        RECT 30.000 117.600 31.800 118.400 ;
        RECT 21.800 108.400 22.400 111.800 ;
        RECT 23.400 109.800 24.000 111.800 ;
        RECT 26.800 111.600 27.400 115.000 ;
        RECT 31.000 112.800 31.800 117.600 ;
        RECT 31.000 112.200 32.600 112.800 ;
        RECT 26.800 111.000 30.600 111.600 ;
        RECT 23.000 109.000 24.000 109.800 ;
        RECT 21.800 107.600 22.800 108.400 ;
        RECT 21.800 106.200 22.400 107.600 ;
        RECT 23.400 107.400 24.000 109.000 ;
        RECT 25.000 109.600 26.000 110.400 ;
        RECT 25.000 108.800 25.800 109.600 ;
        RECT 26.800 108.800 27.600 110.400 ;
        RECT 28.400 108.800 29.200 110.400 ;
        RECT 30.000 109.000 30.600 111.000 ;
        RECT 30.000 108.200 31.400 109.000 ;
        RECT 32.000 108.400 32.600 112.200 ;
        RECT 36.400 112.400 37.200 119.800 ;
        RECT 39.600 112.800 40.400 119.800 ;
        RECT 36.400 111.800 39.000 112.400 ;
        RECT 39.600 111.800 40.600 112.800 ;
        RECT 42.800 112.400 43.600 119.800 ;
        RECT 46.000 112.800 46.800 119.800 ;
        RECT 42.800 111.800 45.400 112.400 ;
        RECT 46.000 111.800 47.000 112.800 ;
        RECT 33.200 110.300 34.000 111.200 ;
        RECT 34.800 110.300 35.600 110.400 ;
        RECT 33.200 109.700 35.600 110.300 ;
        RECT 33.200 109.600 34.000 109.700 ;
        RECT 34.800 109.600 35.600 109.700 ;
        RECT 36.400 109.600 37.400 110.400 ;
        RECT 36.600 108.800 37.400 109.600 ;
        RECT 38.400 109.800 39.000 111.800 ;
        RECT 38.400 109.000 39.400 109.800 ;
        RECT 30.000 107.800 31.000 108.200 ;
        RECT 23.400 106.800 26.000 107.400 ;
        RECT 21.800 105.600 22.800 106.200 ;
        RECT 22.000 102.200 22.800 105.600 ;
        RECT 25.200 102.200 26.000 106.800 ;
        RECT 26.800 107.200 31.000 107.800 ;
        RECT 32.000 107.600 34.000 108.400 ;
        RECT 26.800 105.000 27.400 107.200 ;
        RECT 32.000 107.000 32.600 107.600 ;
        RECT 38.400 107.400 39.000 109.000 ;
        RECT 40.000 108.400 40.600 111.800 ;
        RECT 42.800 109.600 43.800 110.400 ;
        RECT 43.000 108.800 43.800 109.600 ;
        RECT 44.800 109.800 45.400 111.800 ;
        RECT 44.800 109.000 45.800 109.800 ;
        RECT 39.600 108.300 40.600 108.400 ;
        RECT 41.200 108.300 42.000 108.400 ;
        RECT 39.600 107.700 42.000 108.300 ;
        RECT 39.600 107.600 40.600 107.700 ;
        RECT 41.200 107.600 42.000 107.700 ;
        RECT 31.800 106.600 32.600 107.000 ;
        RECT 31.000 106.000 32.600 106.600 ;
        RECT 36.400 106.800 39.000 107.400 ;
        RECT 26.800 103.000 27.600 105.000 ;
        RECT 31.000 103.000 31.800 106.000 ;
        RECT 36.400 102.200 37.200 106.800 ;
        RECT 40.000 106.200 40.600 107.600 ;
        RECT 44.800 107.400 45.400 109.000 ;
        RECT 46.400 108.400 47.000 111.800 ;
        RECT 49.200 111.400 50.000 119.800 ;
        RECT 53.600 116.400 54.400 119.800 ;
        RECT 52.400 115.800 54.400 116.400 ;
        RECT 58.000 115.800 58.800 119.800 ;
        RECT 62.200 115.800 63.400 119.800 ;
        RECT 52.400 115.000 53.200 115.800 ;
        RECT 58.000 115.200 58.600 115.800 ;
        RECT 55.800 114.600 59.400 115.200 ;
        RECT 62.000 115.000 62.800 115.800 ;
        RECT 55.800 114.400 56.600 114.600 ;
        RECT 58.600 114.400 59.400 114.600 ;
        RECT 52.400 113.000 53.200 113.200 ;
        RECT 57.000 113.000 57.800 113.200 ;
        RECT 52.400 112.400 57.800 113.000 ;
        RECT 58.400 113.000 60.600 113.600 ;
        RECT 58.400 111.800 59.000 113.000 ;
        RECT 59.800 112.800 60.600 113.000 ;
        RECT 62.200 113.200 63.600 114.000 ;
        RECT 62.200 112.200 62.800 113.200 ;
        RECT 54.200 111.400 59.000 111.800 ;
        RECT 49.200 111.200 59.000 111.400 ;
        RECT 60.400 111.600 62.800 112.200 ;
        RECT 49.200 111.000 55.000 111.200 ;
        RECT 49.200 110.800 54.800 111.000 ;
        RECT 55.600 110.200 56.400 110.400 ;
        RECT 51.400 109.600 56.400 110.200 ;
        RECT 51.400 109.400 52.200 109.600 ;
        RECT 53.000 108.400 53.800 108.600 ;
        RECT 60.400 108.400 61.000 111.600 ;
        RECT 66.800 111.200 67.600 119.800 ;
        RECT 63.400 110.600 67.600 111.200 ;
        RECT 68.400 115.000 69.200 119.000 ;
        RECT 72.600 118.400 73.400 119.800 ;
        RECT 72.600 117.600 74.000 118.400 ;
        RECT 68.400 111.600 69.000 115.000 ;
        RECT 72.600 112.800 73.400 117.600 ;
        RECT 72.600 112.200 74.200 112.800 ;
        RECT 68.400 111.000 72.200 111.600 ;
        RECT 63.400 110.400 64.200 110.600 ;
        RECT 65.000 109.800 65.800 110.000 ;
        RECT 62.000 109.200 65.800 109.800 ;
        RECT 62.000 109.000 62.800 109.200 ;
        RECT 46.000 107.600 47.000 108.400 ;
        RECT 50.000 107.800 61.000 108.400 ;
        RECT 50.000 107.600 51.600 107.800 ;
        RECT 39.600 105.600 40.600 106.200 ;
        RECT 42.800 106.800 45.400 107.400 ;
        RECT 39.600 102.200 40.400 105.600 ;
        RECT 42.800 102.200 43.600 106.800 ;
        RECT 46.400 106.200 47.000 107.600 ;
        RECT 46.000 105.600 47.000 106.200 ;
        RECT 46.000 102.200 46.800 105.600 ;
        RECT 49.200 102.200 50.000 107.000 ;
        RECT 54.200 105.600 54.800 107.800 ;
        RECT 59.800 107.600 60.600 107.800 ;
        RECT 66.800 107.200 67.600 110.600 ;
        RECT 68.400 108.800 69.200 110.400 ;
        RECT 70.000 108.800 70.800 110.400 ;
        RECT 71.600 109.000 72.200 111.000 ;
        RECT 71.600 108.200 73.000 109.000 ;
        RECT 73.600 108.400 74.200 112.200 ;
        RECT 74.800 110.300 75.600 111.200 ;
        RECT 78.000 110.300 78.800 110.400 ;
        RECT 74.800 109.700 78.800 110.300 ;
        RECT 74.800 109.600 75.600 109.700 ;
        RECT 78.000 109.600 78.800 109.700 ;
        RECT 71.600 107.800 72.600 108.200 ;
        RECT 63.800 106.600 67.600 107.200 ;
        RECT 63.800 106.400 64.600 106.600 ;
        RECT 52.400 104.200 53.200 105.000 ;
        RECT 54.000 104.800 54.800 105.600 ;
        RECT 55.800 105.400 56.600 105.600 ;
        RECT 55.800 104.800 58.600 105.400 ;
        RECT 58.000 104.200 58.600 104.800 ;
        RECT 62.000 104.200 62.800 105.000 ;
        RECT 52.400 103.600 54.400 104.200 ;
        RECT 53.600 102.200 54.400 103.600 ;
        RECT 58.000 102.200 58.800 104.200 ;
        RECT 62.000 103.600 63.400 104.200 ;
        RECT 62.200 102.200 63.400 103.600 ;
        RECT 66.800 102.200 67.600 106.600 ;
        RECT 68.400 107.200 72.600 107.800 ;
        RECT 73.600 107.600 75.600 108.400 ;
        RECT 68.400 105.000 69.000 107.200 ;
        RECT 73.600 107.000 74.200 107.600 ;
        RECT 73.400 106.600 74.200 107.000 ;
        RECT 72.600 106.000 74.200 106.600 ;
        RECT 68.400 103.000 69.200 105.000 ;
        RECT 72.600 103.000 73.400 106.000 ;
        RECT 78.000 104.800 78.800 106.400 ;
        RECT 79.600 102.200 80.400 119.800 ;
        RECT 81.200 111.400 82.000 119.800 ;
        RECT 85.600 116.400 86.400 119.800 ;
        RECT 84.400 115.800 86.400 116.400 ;
        RECT 90.000 115.800 90.800 119.800 ;
        RECT 94.200 115.800 95.400 119.800 ;
        RECT 84.400 115.000 85.200 115.800 ;
        RECT 90.000 115.200 90.600 115.800 ;
        RECT 87.800 114.600 91.400 115.200 ;
        RECT 94.000 115.000 94.800 115.800 ;
        RECT 87.800 114.400 88.600 114.600 ;
        RECT 90.600 114.400 91.400 114.600 ;
        RECT 84.400 113.000 85.200 113.200 ;
        RECT 89.000 113.000 89.800 113.200 ;
        RECT 84.400 112.400 89.800 113.000 ;
        RECT 90.400 113.000 92.600 113.600 ;
        RECT 90.400 111.800 91.000 113.000 ;
        RECT 91.800 112.800 92.600 113.000 ;
        RECT 94.200 113.200 95.600 114.000 ;
        RECT 94.200 112.200 94.800 113.200 ;
        RECT 86.200 111.400 91.000 111.800 ;
        RECT 81.200 111.200 91.000 111.400 ;
        RECT 92.400 111.600 94.800 112.200 ;
        RECT 81.200 111.000 87.000 111.200 ;
        RECT 81.200 110.800 86.800 111.000 ;
        RECT 87.600 110.200 88.400 110.400 ;
        RECT 83.400 109.600 88.400 110.200 ;
        RECT 83.400 109.400 84.200 109.600 ;
        RECT 85.000 108.400 85.800 108.600 ;
        RECT 92.400 108.400 93.000 111.600 ;
        RECT 98.800 111.200 99.600 119.800 ;
        RECT 103.000 112.400 103.800 119.800 ;
        RECT 104.400 113.600 105.200 114.400 ;
        RECT 104.600 112.400 105.200 113.600 ;
        RECT 107.600 113.600 108.400 114.400 ;
        RECT 107.600 112.400 108.200 113.600 ;
        RECT 109.000 112.400 109.800 119.800 ;
        RECT 102.000 111.600 104.000 112.400 ;
        RECT 104.600 111.800 106.000 112.400 ;
        RECT 105.200 111.600 106.000 111.800 ;
        RECT 106.800 111.800 108.200 112.400 ;
        RECT 108.800 111.800 109.800 112.400 ;
        RECT 118.000 112.400 118.800 119.800 ;
        RECT 121.200 112.800 122.000 119.800 ;
        RECT 124.400 114.300 125.200 114.400 ;
        RECT 126.000 114.300 126.800 119.800 ;
        RECT 124.400 113.700 126.800 114.300 ;
        RECT 124.400 113.600 125.200 113.700 ;
        RECT 118.000 111.800 120.600 112.400 ;
        RECT 106.800 111.600 107.600 111.800 ;
        RECT 95.400 110.600 99.600 111.200 ;
        RECT 95.400 110.400 96.200 110.600 ;
        RECT 97.000 109.800 97.800 110.000 ;
        RECT 94.000 109.200 97.800 109.800 ;
        RECT 94.000 109.000 94.800 109.200 ;
        RECT 82.000 107.800 93.000 108.400 ;
        RECT 82.000 107.600 83.600 107.800 ;
        RECT 81.200 102.200 82.000 107.000 ;
        RECT 86.200 105.600 86.800 107.800 ;
        RECT 87.600 107.600 88.400 107.800 ;
        RECT 91.800 107.600 92.600 107.800 ;
        RECT 98.800 107.200 99.600 110.600 ;
        RECT 102.000 108.800 102.800 110.400 ;
        RECT 103.400 108.400 104.000 111.600 ;
        RECT 105.300 110.300 105.900 111.600 ;
        RECT 108.800 110.300 109.400 111.800 ;
        RECT 105.300 109.700 109.400 110.300 ;
        RECT 108.800 108.400 109.400 109.700 ;
        RECT 110.000 110.300 110.800 110.400 ;
        RECT 114.800 110.300 115.600 110.400 ;
        RECT 110.000 109.700 115.600 110.300 ;
        RECT 110.000 108.800 110.800 109.700 ;
        RECT 114.800 109.600 115.600 109.700 ;
        RECT 118.000 109.600 119.000 110.400 ;
        RECT 118.200 108.800 119.000 109.600 ;
        RECT 120.000 109.800 120.600 111.800 ;
        RECT 121.200 111.600 122.200 112.800 ;
        RECT 120.000 109.000 121.000 109.800 ;
        RECT 100.400 108.200 101.200 108.400 ;
        RECT 100.400 107.600 102.000 108.200 ;
        RECT 103.400 107.600 106.000 108.400 ;
        RECT 106.800 107.600 109.400 108.400 ;
        RECT 111.600 108.200 112.400 108.400 ;
        RECT 110.800 107.600 112.400 108.200 ;
        RECT 101.200 107.200 102.000 107.600 ;
        RECT 95.800 106.600 99.600 107.200 ;
        RECT 95.800 106.400 96.600 106.600 ;
        RECT 84.400 104.200 85.200 105.000 ;
        RECT 86.000 104.800 86.800 105.600 ;
        RECT 87.800 105.400 88.600 105.600 ;
        RECT 87.800 104.800 90.600 105.400 ;
        RECT 90.000 104.200 90.600 104.800 ;
        RECT 94.000 104.200 94.800 105.000 ;
        RECT 84.400 103.600 86.400 104.200 ;
        RECT 85.600 102.200 86.400 103.600 ;
        RECT 90.000 102.200 90.800 104.200 ;
        RECT 94.000 103.600 95.400 104.200 ;
        RECT 94.200 102.200 95.400 103.600 ;
        RECT 98.800 102.200 99.600 106.600 ;
        RECT 100.600 106.200 104.200 106.600 ;
        RECT 105.200 106.200 105.800 107.600 ;
        RECT 107.000 106.200 107.600 107.600 ;
        RECT 110.800 107.200 111.600 107.600 ;
        RECT 120.000 107.400 120.600 109.000 ;
        RECT 121.600 108.400 122.200 111.600 ;
        RECT 121.200 108.300 122.200 108.400 ;
        RECT 122.800 108.300 123.600 108.400 ;
        RECT 121.200 107.700 123.600 108.300 ;
        RECT 121.200 107.600 122.200 107.700 ;
        RECT 122.800 107.600 123.600 107.700 ;
        RECT 118.000 106.800 120.600 107.400 ;
        RECT 108.600 106.200 112.200 106.600 ;
        RECT 100.400 106.000 104.400 106.200 ;
        RECT 100.400 102.200 101.200 106.000 ;
        RECT 103.600 102.200 104.400 106.000 ;
        RECT 105.200 102.200 106.000 106.200 ;
        RECT 106.800 102.200 107.600 106.200 ;
        RECT 108.400 106.000 112.400 106.200 ;
        RECT 108.400 102.200 109.200 106.000 ;
        RECT 111.600 102.200 112.400 106.000 ;
        RECT 118.000 102.200 118.800 106.800 ;
        RECT 121.600 106.200 122.200 107.600 ;
        RECT 124.400 106.800 125.200 108.400 ;
        RECT 121.200 105.600 122.200 106.200 ;
        RECT 126.000 106.200 126.800 113.700 ;
        RECT 127.600 111.600 128.400 113.200 ;
        RECT 131.800 112.400 132.600 119.800 ;
        RECT 133.200 113.600 134.000 114.400 ;
        RECT 133.400 112.400 134.000 113.600 ;
        RECT 139.400 112.800 140.200 119.800 ;
        RECT 143.600 115.000 144.400 119.000 ;
        RECT 131.800 111.800 132.800 112.400 ;
        RECT 133.400 111.800 134.800 112.400 ;
        RECT 130.800 108.800 131.600 110.400 ;
        RECT 132.200 108.400 132.800 111.800 ;
        RECT 134.000 111.600 134.800 111.800 ;
        RECT 138.600 112.200 140.200 112.800 ;
        RECT 137.200 109.600 138.000 111.200 ;
        RECT 138.600 110.400 139.200 112.200 ;
        RECT 143.800 111.600 144.400 115.000 ;
        RECT 147.800 112.400 148.600 119.800 ;
        RECT 149.200 113.600 150.000 114.400 ;
        RECT 149.400 112.400 150.000 113.600 ;
        RECT 147.800 111.800 148.800 112.400 ;
        RECT 149.400 111.800 150.800 112.400 ;
        RECT 140.600 111.000 144.400 111.600 ;
        RECT 138.600 109.600 139.600 110.400 ;
        RECT 138.600 108.400 139.200 109.600 ;
        RECT 140.600 109.000 141.200 111.000 ;
        RECT 127.600 108.300 128.400 108.400 ;
        RECT 129.200 108.300 130.000 108.400 ;
        RECT 127.600 108.200 130.000 108.300 ;
        RECT 127.600 107.700 130.800 108.200 ;
        RECT 127.600 107.600 128.400 107.700 ;
        RECT 129.200 107.600 130.800 107.700 ;
        RECT 132.200 107.600 134.800 108.400 ;
        RECT 137.200 107.600 139.200 108.400 ;
        RECT 139.800 108.200 141.200 109.000 ;
        RECT 142.000 108.800 142.800 110.400 ;
        RECT 143.600 108.800 144.400 110.400 ;
        RECT 146.800 108.800 147.600 110.400 ;
        RECT 148.200 110.300 148.800 111.800 ;
        RECT 150.000 111.600 150.800 111.800 ;
        RECT 151.600 111.400 152.400 119.800 ;
        RECT 156.000 116.400 156.800 119.800 ;
        RECT 154.800 115.800 156.800 116.400 ;
        RECT 160.400 115.800 161.200 119.800 ;
        RECT 164.600 115.800 165.800 119.800 ;
        RECT 154.800 115.000 155.600 115.800 ;
        RECT 160.400 115.200 161.000 115.800 ;
        RECT 158.200 114.600 161.800 115.200 ;
        RECT 164.400 115.000 165.200 115.800 ;
        RECT 158.200 114.400 159.000 114.600 ;
        RECT 161.000 114.400 161.800 114.600 ;
        RECT 154.800 113.000 155.600 113.200 ;
        RECT 159.400 113.000 160.200 113.200 ;
        RECT 154.800 112.400 160.200 113.000 ;
        RECT 160.800 113.000 163.000 113.600 ;
        RECT 160.800 111.800 161.400 113.000 ;
        RECT 162.200 112.800 163.000 113.000 ;
        RECT 164.600 113.200 166.000 114.000 ;
        RECT 164.600 112.200 165.200 113.200 ;
        RECT 156.600 111.400 161.400 111.800 ;
        RECT 151.600 111.200 161.400 111.400 ;
        RECT 162.800 111.600 165.200 112.200 ;
        RECT 151.600 111.000 157.400 111.200 ;
        RECT 151.600 110.800 157.200 111.000 ;
        RECT 150.000 110.300 150.800 110.400 ;
        RECT 148.200 109.700 150.800 110.300 ;
        RECT 158.000 110.200 158.800 110.400 ;
        RECT 148.200 108.400 148.800 109.700 ;
        RECT 150.000 109.600 150.800 109.700 ;
        RECT 153.800 109.600 158.800 110.200 ;
        RECT 153.800 109.400 154.600 109.600 ;
        RECT 156.400 109.400 157.200 109.600 ;
        RECT 155.400 108.400 156.200 108.600 ;
        RECT 162.800 108.400 163.400 111.600 ;
        RECT 169.200 111.200 170.000 119.800 ;
        RECT 165.800 110.600 170.000 111.200 ;
        RECT 165.800 110.400 166.600 110.600 ;
        RECT 167.400 109.800 168.200 110.000 ;
        RECT 164.400 109.200 168.200 109.800 ;
        RECT 164.400 109.000 165.200 109.200 ;
        RECT 130.000 107.200 130.800 107.600 ;
        RECT 129.400 106.200 133.000 106.600 ;
        RECT 134.000 106.400 134.600 107.600 ;
        RECT 138.600 107.000 139.200 107.600 ;
        RECT 140.200 107.800 141.200 108.200 ;
        RECT 145.200 108.200 146.000 108.400 ;
        RECT 140.200 107.200 144.400 107.800 ;
        RECT 145.200 107.600 146.800 108.200 ;
        RECT 148.200 107.600 150.800 108.400 ;
        RECT 152.400 107.800 163.400 108.400 ;
        RECT 152.400 107.600 154.000 107.800 ;
        RECT 146.000 107.200 146.800 107.600 ;
        RECT 138.600 106.600 139.400 107.000 ;
        RECT 126.000 105.600 127.800 106.200 ;
        RECT 121.200 102.200 122.000 105.600 ;
        RECT 127.000 102.200 127.800 105.600 ;
        RECT 129.200 106.000 133.200 106.200 ;
        RECT 129.200 102.200 130.000 106.000 ;
        RECT 132.400 102.200 133.200 106.000 ;
        RECT 134.000 102.200 134.800 106.400 ;
        RECT 138.600 106.000 140.200 106.600 ;
        RECT 139.400 103.000 140.200 106.000 ;
        RECT 143.800 105.000 144.400 107.200 ;
        RECT 145.400 106.200 149.000 106.600 ;
        RECT 150.000 106.200 150.600 107.600 ;
        RECT 143.600 103.000 144.400 105.000 ;
        RECT 145.200 106.000 149.200 106.200 ;
        RECT 145.200 102.200 146.000 106.000 ;
        RECT 148.400 102.200 149.200 106.000 ;
        RECT 150.000 102.200 150.800 106.200 ;
        RECT 151.600 102.200 152.400 107.000 ;
        RECT 156.600 105.600 157.200 107.800 ;
        RECT 162.200 107.600 163.000 107.800 ;
        RECT 169.200 107.200 170.000 110.600 ;
        RECT 166.200 106.600 170.000 107.200 ;
        RECT 166.200 106.400 167.000 106.600 ;
        RECT 169.200 106.300 170.000 106.600 ;
        RECT 172.400 108.300 173.200 119.800 ;
        RECT 176.600 112.400 177.400 119.800 ;
        RECT 183.000 116.400 183.800 119.800 ;
        RECT 182.000 115.600 183.800 116.400 ;
        RECT 178.000 113.600 178.800 114.400 ;
        RECT 178.200 112.400 178.800 113.600 ;
        RECT 183.000 112.400 183.800 115.600 ;
        RECT 184.400 113.600 185.200 114.400 ;
        RECT 184.600 112.400 185.200 113.600 ;
        RECT 176.600 111.800 177.600 112.400 ;
        RECT 178.200 111.800 179.600 112.400 ;
        RECT 183.000 111.800 184.000 112.400 ;
        RECT 184.600 111.800 186.000 112.400 ;
        RECT 175.600 108.800 176.400 110.400 ;
        RECT 177.000 110.300 177.600 111.800 ;
        RECT 178.800 111.600 179.600 111.800 ;
        RECT 182.000 110.300 182.800 110.400 ;
        RECT 177.000 109.700 182.800 110.300 ;
        RECT 177.000 108.400 177.600 109.700 ;
        RECT 182.000 108.800 182.800 109.700 ;
        RECT 183.400 108.400 184.000 111.800 ;
        RECT 185.200 111.600 186.000 111.800 ;
        RECT 174.000 108.300 174.800 108.400 ;
        RECT 172.400 108.200 174.800 108.300 ;
        RECT 172.400 107.700 175.600 108.200 ;
        RECT 170.800 106.300 171.600 106.400 ;
        RECT 169.200 105.700 171.600 106.300 ;
        RECT 154.800 104.200 155.600 105.000 ;
        RECT 156.400 104.800 157.200 105.600 ;
        RECT 158.200 105.400 159.000 105.600 ;
        RECT 158.200 104.800 161.000 105.400 ;
        RECT 160.400 104.200 161.000 104.800 ;
        RECT 164.400 104.200 165.200 105.000 ;
        RECT 154.800 103.600 156.800 104.200 ;
        RECT 156.000 102.200 156.800 103.600 ;
        RECT 160.400 102.200 161.200 104.200 ;
        RECT 164.400 103.600 165.800 104.200 ;
        RECT 164.600 102.200 165.800 103.600 ;
        RECT 169.200 102.200 170.000 105.700 ;
        RECT 170.800 104.800 171.600 105.700 ;
        RECT 172.400 102.200 173.200 107.700 ;
        RECT 174.000 107.600 175.600 107.700 ;
        RECT 177.000 107.600 179.600 108.400 ;
        RECT 180.400 108.200 181.200 108.400 ;
        RECT 180.400 107.600 182.000 108.200 ;
        RECT 183.400 107.600 186.000 108.400 ;
        RECT 174.800 107.200 175.600 107.600 ;
        RECT 174.200 106.200 177.800 106.600 ;
        RECT 178.800 106.200 179.400 107.600 ;
        RECT 181.200 107.200 182.000 107.600 ;
        RECT 180.600 106.200 184.200 106.600 ;
        RECT 185.200 106.200 185.800 107.600 ;
        RECT 174.000 106.000 178.000 106.200 ;
        RECT 174.000 102.200 174.800 106.000 ;
        RECT 177.200 102.200 178.000 106.000 ;
        RECT 178.800 102.200 179.600 106.200 ;
        RECT 180.400 106.000 184.400 106.200 ;
        RECT 180.400 102.200 181.200 106.000 ;
        RECT 183.600 102.200 184.400 106.000 ;
        RECT 185.200 102.200 186.000 106.200 ;
        RECT 186.800 102.200 187.600 119.800 ;
        RECT 190.800 113.600 191.600 114.400 ;
        RECT 190.800 112.400 191.400 113.600 ;
        RECT 192.200 112.400 193.000 119.800 ;
        RECT 198.600 118.400 199.400 119.800 ;
        RECT 198.600 117.600 200.400 118.400 ;
        RECT 197.200 113.600 198.000 114.400 ;
        RECT 197.200 112.400 197.800 113.600 ;
        RECT 198.600 112.400 199.400 117.600 ;
        RECT 205.400 112.600 206.200 119.800 ;
        RECT 190.000 111.800 191.400 112.400 ;
        RECT 190.000 111.600 190.800 111.800 ;
        RECT 192.000 111.600 194.000 112.400 ;
        RECT 196.400 111.800 197.800 112.400 ;
        RECT 198.400 111.800 199.400 112.400 ;
        RECT 204.400 111.800 206.200 112.600 ;
        RECT 208.200 112.400 209.000 119.800 ;
        RECT 207.600 111.800 209.000 112.400 ;
        RECT 196.400 111.600 197.200 111.800 ;
        RECT 192.000 108.400 192.600 111.600 ;
        RECT 193.200 108.800 194.000 110.400 ;
        RECT 198.400 108.400 199.000 111.800 ;
        RECT 199.600 108.800 200.400 110.400 ;
        RECT 204.600 108.400 205.200 111.800 ;
        RECT 207.600 111.600 208.400 111.800 ;
        RECT 206.000 110.300 206.800 111.200 ;
        RECT 207.600 110.400 208.200 111.600 ;
        RECT 212.400 111.200 213.200 119.800 ;
        RECT 214.000 111.600 214.800 113.200 ;
        RECT 215.600 112.300 216.400 119.800 ;
        RECT 217.200 112.300 218.000 112.400 ;
        RECT 215.600 111.700 218.000 112.300 ;
        RECT 209.200 110.800 213.200 111.200 ;
        RECT 209.000 110.600 213.200 110.800 ;
        RECT 207.600 110.300 208.400 110.400 ;
        RECT 206.000 109.700 208.400 110.300 ;
        RECT 206.000 109.600 206.800 109.700 ;
        RECT 207.600 109.600 208.400 109.700 ;
        RECT 209.000 110.000 209.800 110.600 ;
        RECT 188.400 106.800 189.200 108.400 ;
        RECT 190.000 107.600 192.600 108.400 ;
        RECT 194.800 108.200 195.600 108.400 ;
        RECT 194.000 107.600 195.600 108.200 ;
        RECT 196.400 107.600 199.000 108.400 ;
        RECT 201.200 108.200 202.000 108.400 ;
        RECT 200.400 107.600 202.000 108.200 ;
        RECT 204.400 107.600 205.200 108.400 ;
        RECT 190.200 106.200 190.800 107.600 ;
        RECT 194.000 107.200 194.800 107.600 ;
        RECT 191.800 106.200 195.400 106.600 ;
        RECT 196.600 106.200 197.200 107.600 ;
        RECT 200.400 107.200 201.200 107.600 ;
        RECT 198.200 106.200 201.800 106.600 ;
        RECT 190.000 102.200 190.800 106.200 ;
        RECT 191.600 106.000 195.600 106.200 ;
        RECT 191.600 102.200 192.400 106.000 ;
        RECT 194.800 102.200 195.600 106.000 ;
        RECT 196.400 102.200 197.200 106.200 ;
        RECT 198.000 106.000 202.000 106.200 ;
        RECT 198.000 102.200 198.800 106.000 ;
        RECT 201.200 102.200 202.000 106.000 ;
        RECT 202.800 104.800 203.600 106.400 ;
        RECT 204.600 104.400 205.200 107.600 ;
        RECT 204.400 102.200 205.200 104.400 ;
        RECT 207.600 106.200 208.200 109.600 ;
        RECT 209.000 107.000 209.600 110.000 ;
        RECT 210.400 108.400 211.200 109.200 ;
        RECT 210.600 107.600 211.600 108.400 ;
        RECT 209.000 106.400 211.400 107.000 ;
        RECT 207.600 102.200 208.400 106.200 ;
        RECT 210.800 104.200 211.400 106.400 ;
        RECT 212.400 104.800 213.200 106.400 ;
        RECT 215.600 106.200 216.400 111.700 ;
        RECT 217.200 111.600 218.000 111.700 ;
        RECT 217.200 110.300 218.000 110.400 ;
        RECT 218.800 110.300 219.600 119.800 ;
        RECT 222.600 118.400 223.400 119.800 ;
        RECT 222.600 117.600 224.400 118.400 ;
        RECT 222.600 112.600 223.400 117.600 ;
        RECT 222.600 111.800 224.400 112.600 ;
        RECT 226.800 112.400 227.600 119.800 ;
        RECT 230.000 112.400 230.800 119.800 ;
        RECT 226.800 111.800 230.800 112.400 ;
        RECT 231.600 111.800 232.400 119.800 ;
        RECT 235.800 112.400 236.600 119.800 ;
        RECT 237.200 113.600 238.000 114.400 ;
        RECT 237.400 112.400 238.000 113.600 ;
        RECT 242.200 112.400 243.000 119.800 ;
        RECT 243.600 113.600 244.400 114.400 ;
        RECT 243.800 112.400 244.400 113.600 ;
        RECT 235.800 111.800 236.800 112.400 ;
        RECT 237.400 111.800 238.800 112.400 ;
        RECT 242.200 111.800 243.200 112.400 ;
        RECT 243.800 111.800 245.200 112.400 ;
        RECT 217.200 109.700 219.600 110.300 ;
        RECT 217.200 109.600 218.000 109.700 ;
        RECT 217.200 106.800 218.000 108.400 ;
        RECT 214.600 105.600 216.400 106.200 ;
        RECT 210.800 102.200 211.600 104.200 ;
        RECT 214.600 102.200 215.400 105.600 ;
        RECT 218.800 102.200 219.600 109.700 ;
        RECT 222.000 109.600 222.800 111.200 ;
        RECT 223.600 108.400 224.200 111.800 ;
        RECT 227.600 110.400 228.400 110.800 ;
        RECT 231.600 110.400 232.200 111.800 ;
        RECT 226.800 109.800 228.400 110.400 ;
        RECT 230.000 110.300 232.400 110.400 ;
        RECT 234.800 110.300 235.600 110.400 ;
        RECT 230.000 109.800 235.600 110.300 ;
        RECT 226.800 109.600 227.600 109.800 ;
        RECT 223.600 107.600 224.400 108.400 ;
        RECT 228.400 107.600 229.200 109.200 ;
        RECT 220.400 104.800 221.200 106.400 ;
        RECT 223.600 104.200 224.200 107.600 ;
        RECT 225.200 104.800 226.000 106.400 ;
        RECT 230.000 106.200 230.600 109.800 ;
        RECT 231.600 109.700 235.600 109.800 ;
        RECT 231.600 109.600 232.400 109.700 ;
        RECT 234.800 108.800 235.600 109.700 ;
        RECT 236.200 110.300 236.800 111.800 ;
        RECT 238.000 111.600 238.800 111.800 ;
        RECT 239.600 110.300 240.400 110.400 ;
        RECT 236.200 109.700 240.400 110.300 ;
        RECT 236.200 108.400 236.800 109.700 ;
        RECT 239.600 109.600 240.400 109.700 ;
        RECT 241.200 108.800 242.000 110.400 ;
        RECT 242.600 108.400 243.200 111.800 ;
        RECT 244.400 111.600 245.200 111.800 ;
        RECT 233.200 108.200 234.000 108.400 ;
        RECT 233.200 107.600 234.800 108.200 ;
        RECT 236.200 107.600 238.800 108.400 ;
        RECT 239.600 108.200 240.400 108.400 ;
        RECT 242.600 108.300 245.200 108.400 ;
        RECT 246.000 108.300 246.800 108.400 ;
        RECT 239.600 107.600 241.200 108.200 ;
        RECT 242.600 107.700 246.800 108.300 ;
        RECT 242.600 107.600 245.200 107.700 ;
        RECT 234.000 107.200 234.800 107.600 ;
        RECT 223.600 102.200 224.400 104.200 ;
        RECT 230.000 102.200 230.800 106.200 ;
        RECT 231.600 105.600 232.400 106.400 ;
        RECT 233.400 106.200 237.000 106.600 ;
        RECT 238.000 106.200 238.600 107.600 ;
        RECT 240.400 107.200 241.200 107.600 ;
        RECT 239.800 106.200 243.400 106.600 ;
        RECT 244.400 106.200 245.000 107.600 ;
        RECT 246.000 106.800 246.800 107.700 ;
        RECT 247.600 106.200 248.400 119.800 ;
        RECT 249.200 111.600 250.000 113.200 ;
        RECT 253.400 112.400 254.200 119.800 ;
        RECT 254.800 114.300 255.600 114.400 ;
        RECT 257.200 114.300 258.000 114.400 ;
        RECT 254.800 113.700 258.000 114.300 ;
        RECT 254.800 113.600 255.600 113.700 ;
        RECT 257.200 113.600 258.000 113.700 ;
        RECT 255.000 112.400 255.600 113.600 ;
        RECT 253.400 111.800 254.400 112.400 ;
        RECT 255.000 111.800 256.400 112.400 ;
        RECT 252.400 108.800 253.200 110.400 ;
        RECT 253.800 108.400 254.400 111.800 ;
        RECT 255.600 111.600 256.400 111.800 ;
        RECT 250.800 108.200 251.600 108.400 ;
        RECT 253.800 108.300 256.400 108.400 ;
        RECT 257.200 108.300 258.000 108.400 ;
        RECT 250.800 107.600 252.400 108.200 ;
        RECT 253.800 107.700 258.000 108.300 ;
        RECT 253.800 107.600 256.400 107.700 ;
        RECT 251.600 107.200 252.400 107.600 ;
        RECT 251.000 106.200 254.600 106.600 ;
        RECT 255.600 106.200 256.200 107.600 ;
        RECT 257.200 106.800 258.000 107.700 ;
        RECT 258.800 108.300 259.600 119.800 ;
        RECT 260.400 111.600 261.200 113.200 ;
        RECT 268.400 112.000 269.200 119.800 ;
        RECT 271.600 115.200 272.400 119.800 ;
        RECT 268.200 111.200 269.200 112.000 ;
        RECT 269.800 114.600 272.400 115.200 ;
        RECT 269.800 113.000 270.400 114.600 ;
        RECT 274.800 114.400 275.600 119.800 ;
        RECT 278.000 117.000 278.800 119.800 ;
        RECT 279.600 117.000 280.400 119.800 ;
        RECT 281.200 117.000 282.000 119.800 ;
        RECT 276.200 114.400 280.400 115.200 ;
        RECT 273.000 113.600 275.600 114.400 ;
        RECT 282.800 113.600 283.600 119.800 ;
        RECT 286.000 115.000 286.800 119.800 ;
        RECT 289.200 115.000 290.000 119.800 ;
        RECT 290.800 117.000 291.600 119.800 ;
        RECT 292.400 117.000 293.200 119.800 ;
        RECT 295.600 115.200 296.400 119.800 ;
        RECT 298.800 116.400 299.600 119.800 ;
        RECT 298.800 115.800 299.800 116.400 ;
        RECT 299.200 115.200 299.800 115.800 ;
        RECT 294.400 114.400 298.600 115.200 ;
        RECT 299.200 114.600 301.200 115.200 ;
        RECT 286.000 113.600 288.600 114.400 ;
        RECT 289.200 113.800 295.000 114.400 ;
        RECT 298.000 114.000 298.600 114.400 ;
        RECT 278.000 113.000 278.800 113.200 ;
        RECT 269.800 112.400 278.800 113.000 ;
        RECT 281.200 113.000 282.000 113.200 ;
        RECT 289.200 113.000 289.800 113.800 ;
        RECT 295.600 113.200 297.000 113.800 ;
        RECT 298.000 113.200 299.600 114.000 ;
        RECT 281.200 112.400 289.800 113.000 ;
        RECT 290.800 113.000 297.000 113.200 ;
        RECT 290.800 112.600 296.200 113.000 ;
        RECT 290.800 112.400 291.600 112.600 ;
        RECT 266.800 108.300 267.600 108.400 ;
        RECT 258.800 107.700 267.600 108.300 ;
        RECT 258.800 106.200 259.600 107.700 ;
        RECT 266.800 107.600 267.600 107.700 ;
        RECT 268.200 106.800 269.000 111.200 ;
        RECT 269.800 110.600 270.400 112.400 ;
        RECT 269.600 110.000 270.400 110.600 ;
        RECT 276.400 110.000 299.800 110.600 ;
        RECT 269.600 108.000 270.200 110.000 ;
        RECT 276.400 109.400 277.200 110.000 ;
        RECT 294.000 109.600 294.800 110.000 ;
        RECT 295.600 109.600 296.400 110.000 ;
        RECT 299.000 109.800 299.800 110.000 ;
        RECT 270.800 108.600 274.600 109.400 ;
        RECT 269.600 107.400 270.800 108.000 ;
        RECT 233.200 106.000 237.200 106.200 ;
        RECT 231.400 104.800 232.200 105.600 ;
        RECT 233.200 102.200 234.000 106.000 ;
        RECT 236.400 102.200 237.200 106.000 ;
        RECT 238.000 102.200 238.800 106.200 ;
        RECT 239.600 106.000 243.600 106.200 ;
        RECT 239.600 102.200 240.400 106.000 ;
        RECT 242.800 102.200 243.600 106.000 ;
        RECT 244.400 102.200 245.200 106.200 ;
        RECT 247.600 105.600 249.400 106.200 ;
        RECT 248.600 104.400 249.400 105.600 ;
        RECT 250.800 106.000 254.800 106.200 ;
        RECT 248.600 103.600 250.000 104.400 ;
        RECT 248.600 102.200 249.400 103.600 ;
        RECT 250.800 102.200 251.600 106.000 ;
        RECT 254.000 102.200 254.800 106.000 ;
        RECT 255.600 102.200 256.400 106.200 ;
        RECT 258.800 105.600 260.600 106.200 ;
        RECT 268.200 106.000 269.200 106.800 ;
        RECT 259.800 102.200 260.600 105.600 ;
        RECT 268.400 102.200 269.200 106.000 ;
        RECT 270.000 102.200 270.800 107.400 ;
        RECT 273.800 107.400 274.600 108.600 ;
        RECT 273.800 106.800 275.600 107.400 ;
        RECT 274.800 106.200 275.600 106.800 ;
        RECT 279.600 106.400 280.400 109.200 ;
        RECT 282.800 108.600 286.000 109.400 ;
        RECT 289.800 108.600 291.800 109.400 ;
        RECT 300.400 109.000 301.200 114.600 ;
        RECT 302.000 112.400 302.800 119.800 ;
        RECT 305.200 112.800 306.000 119.800 ;
        RECT 302.000 111.800 304.600 112.400 ;
        RECT 305.200 111.800 306.200 112.800 ;
        RECT 308.400 112.400 309.200 119.800 ;
        RECT 308.400 111.800 310.600 112.400 ;
        RECT 311.600 111.800 312.400 119.800 ;
        RECT 302.000 109.600 303.000 110.400 ;
        RECT 282.400 107.800 283.200 108.000 ;
        RECT 282.400 107.200 286.800 107.800 ;
        RECT 286.000 107.000 286.800 107.200 ;
        RECT 287.600 106.800 288.400 108.400 ;
        RECT 274.800 105.400 277.200 106.200 ;
        RECT 279.600 105.600 280.600 106.400 ;
        RECT 283.600 105.600 285.200 106.400 ;
        RECT 286.000 106.200 286.800 106.400 ;
        RECT 289.800 106.200 290.600 108.600 ;
        RECT 292.400 108.200 301.200 109.000 ;
        RECT 302.200 108.800 303.000 109.600 ;
        RECT 304.000 109.800 304.600 111.800 ;
        RECT 304.000 109.000 305.000 109.800 ;
        RECT 295.800 106.800 298.800 107.600 ;
        RECT 295.800 106.200 296.600 106.800 ;
        RECT 286.000 105.600 290.600 106.200 ;
        RECT 276.400 102.200 277.200 105.400 ;
        RECT 294.000 105.400 296.600 106.200 ;
        RECT 278.000 102.200 278.800 105.000 ;
        RECT 279.600 102.200 280.400 105.000 ;
        RECT 281.200 102.200 282.000 105.000 ;
        RECT 282.800 102.200 283.600 105.000 ;
        RECT 286.000 102.200 286.800 105.000 ;
        RECT 289.200 102.200 290.000 105.000 ;
        RECT 290.800 102.200 291.600 105.000 ;
        RECT 292.400 102.200 293.200 105.000 ;
        RECT 294.000 102.200 294.800 105.400 ;
        RECT 300.400 102.200 301.200 108.200 ;
        RECT 304.000 107.400 304.600 109.000 ;
        RECT 305.600 108.400 306.200 111.800 ;
        RECT 310.000 111.200 310.600 111.800 ;
        RECT 310.000 110.400 311.200 111.200 ;
        RECT 308.400 108.800 309.200 110.400 ;
        RECT 305.200 108.300 306.200 108.400 ;
        RECT 306.800 108.300 307.600 108.400 ;
        RECT 305.200 107.700 307.600 108.300 ;
        RECT 305.200 107.600 306.200 107.700 ;
        RECT 306.800 107.600 307.600 107.700 ;
        RECT 302.000 106.800 304.600 107.400 ;
        RECT 302.000 102.200 302.800 106.800 ;
        RECT 305.600 106.200 306.200 107.600 ;
        RECT 310.000 107.400 310.600 110.400 ;
        RECT 311.800 109.600 312.400 111.800 ;
        RECT 305.200 105.600 306.200 106.200 ;
        RECT 308.400 106.800 310.600 107.400 ;
        RECT 305.200 102.200 306.000 105.600 ;
        RECT 308.400 102.200 309.200 106.800 ;
        RECT 311.600 102.200 312.400 109.600 ;
        RECT 313.200 102.200 314.000 119.800 ;
        RECT 319.000 112.400 319.800 119.800 ;
        RECT 320.400 114.300 321.200 114.400 ;
        RECT 322.800 114.300 323.600 114.400 ;
        RECT 320.400 113.700 323.600 114.300 ;
        RECT 320.400 113.600 321.200 113.700 ;
        RECT 322.800 113.600 323.600 113.700 ;
        RECT 320.600 112.400 321.200 113.600 ;
        RECT 319.000 111.800 320.000 112.400 ;
        RECT 320.600 111.800 322.000 112.400 ;
        RECT 318.000 108.800 318.800 110.400 ;
        RECT 319.400 108.400 320.000 111.800 ;
        RECT 321.200 111.600 322.000 111.800 ;
        RECT 316.400 108.200 317.200 108.400 ;
        RECT 319.400 108.300 322.000 108.400 ;
        RECT 322.800 108.300 323.600 108.400 ;
        RECT 316.400 107.600 318.000 108.200 ;
        RECT 319.400 107.700 323.600 108.300 ;
        RECT 319.400 107.600 322.000 107.700 ;
        RECT 317.200 107.200 318.000 107.600 ;
        RECT 314.800 104.800 315.600 106.400 ;
        RECT 316.600 106.200 320.200 106.600 ;
        RECT 321.200 106.200 321.800 107.600 ;
        RECT 322.800 106.800 323.600 107.700 ;
        RECT 324.400 108.300 325.200 119.800 ;
        RECT 326.000 111.600 326.800 113.200 ;
        RECT 329.200 112.000 330.000 119.800 ;
        RECT 332.400 115.200 333.200 119.800 ;
        RECT 329.000 111.200 330.000 112.000 ;
        RECT 330.600 114.600 333.200 115.200 ;
        RECT 330.600 113.000 331.200 114.600 ;
        RECT 335.600 114.400 336.400 119.800 ;
        RECT 338.800 117.000 339.600 119.800 ;
        RECT 340.400 117.000 341.200 119.800 ;
        RECT 342.000 117.000 342.800 119.800 ;
        RECT 337.000 114.400 341.200 115.200 ;
        RECT 333.800 113.600 336.400 114.400 ;
        RECT 343.600 113.600 344.400 119.800 ;
        RECT 346.800 115.000 347.600 119.800 ;
        RECT 350.000 115.000 350.800 119.800 ;
        RECT 351.600 117.000 352.400 119.800 ;
        RECT 353.200 117.000 354.000 119.800 ;
        RECT 356.400 115.200 357.200 119.800 ;
        RECT 359.600 116.400 360.400 119.800 ;
        RECT 359.600 115.800 360.600 116.400 ;
        RECT 360.000 115.200 360.600 115.800 ;
        RECT 355.200 114.400 359.400 115.200 ;
        RECT 360.000 114.600 362.000 115.200 ;
        RECT 346.800 113.600 349.400 114.400 ;
        RECT 350.000 113.800 355.800 114.400 ;
        RECT 358.800 114.000 359.400 114.400 ;
        RECT 338.800 113.000 339.600 113.200 ;
        RECT 330.600 112.400 339.600 113.000 ;
        RECT 342.000 113.000 342.800 113.200 ;
        RECT 350.000 113.000 350.600 113.800 ;
        RECT 356.400 113.200 357.800 113.800 ;
        RECT 358.800 113.200 360.400 114.000 ;
        RECT 342.000 112.400 350.600 113.000 ;
        RECT 351.600 113.000 357.800 113.200 ;
        RECT 351.600 112.600 357.000 113.000 ;
        RECT 351.600 112.400 352.400 112.600 ;
        RECT 327.600 108.300 328.400 108.400 ;
        RECT 324.400 107.700 328.400 108.300 ;
        RECT 324.400 106.200 325.200 107.700 ;
        RECT 327.600 107.600 328.400 107.700 ;
        RECT 329.000 106.800 329.800 111.200 ;
        RECT 330.600 110.600 331.200 112.400 ;
        RECT 330.400 110.000 331.200 110.600 ;
        RECT 337.200 110.000 360.600 110.600 ;
        RECT 330.400 108.000 331.000 110.000 ;
        RECT 337.200 109.400 338.000 110.000 ;
        RECT 354.800 109.600 355.600 110.000 ;
        RECT 359.800 109.800 360.600 110.000 ;
        RECT 331.600 108.600 335.400 109.400 ;
        RECT 330.400 107.400 331.600 108.000 ;
        RECT 316.400 106.000 320.400 106.200 ;
        RECT 316.400 102.200 317.200 106.000 ;
        RECT 319.600 102.200 320.400 106.000 ;
        RECT 321.200 102.200 322.000 106.200 ;
        RECT 324.400 105.600 326.200 106.200 ;
        RECT 329.000 106.000 330.000 106.800 ;
        RECT 325.400 102.200 326.200 105.600 ;
        RECT 329.200 102.200 330.000 106.000 ;
        RECT 330.800 102.200 331.600 107.400 ;
        RECT 334.600 107.400 335.400 108.600 ;
        RECT 334.600 106.800 336.400 107.400 ;
        RECT 335.600 106.200 336.400 106.800 ;
        RECT 340.400 106.400 341.200 109.200 ;
        RECT 343.600 108.600 346.800 109.400 ;
        RECT 350.600 108.600 352.600 109.400 ;
        RECT 361.200 109.000 362.000 114.600 ;
        RECT 364.400 112.000 365.200 119.800 ;
        RECT 367.600 115.200 368.400 119.800 ;
        RECT 343.200 107.800 344.000 108.000 ;
        RECT 343.200 107.200 347.600 107.800 ;
        RECT 346.800 107.000 347.600 107.200 ;
        RECT 348.400 106.800 349.200 108.400 ;
        RECT 335.600 105.400 338.000 106.200 ;
        RECT 340.400 105.600 341.400 106.400 ;
        RECT 344.400 105.600 346.000 106.400 ;
        RECT 346.800 106.200 347.600 106.400 ;
        RECT 350.600 106.200 351.400 108.600 ;
        RECT 353.200 108.200 362.000 109.000 ;
        RECT 356.600 106.800 359.600 107.600 ;
        RECT 356.600 106.200 357.400 106.800 ;
        RECT 346.800 105.600 351.400 106.200 ;
        RECT 337.200 102.200 338.000 105.400 ;
        RECT 354.800 105.400 357.400 106.200 ;
        RECT 338.800 102.200 339.600 105.000 ;
        RECT 340.400 102.200 341.200 105.000 ;
        RECT 342.000 102.200 342.800 105.000 ;
        RECT 343.600 102.200 344.400 105.000 ;
        RECT 346.800 102.200 347.600 105.000 ;
        RECT 350.000 102.200 350.800 105.000 ;
        RECT 351.600 102.200 352.400 105.000 ;
        RECT 353.200 102.200 354.000 105.000 ;
        RECT 354.800 102.200 355.600 105.400 ;
        RECT 361.200 102.200 362.000 108.200 ;
        RECT 364.200 111.200 365.200 112.000 ;
        RECT 365.800 114.600 368.400 115.200 ;
        RECT 365.800 113.000 366.400 114.600 ;
        RECT 370.800 114.400 371.600 119.800 ;
        RECT 374.000 117.000 374.800 119.800 ;
        RECT 375.600 117.000 376.400 119.800 ;
        RECT 377.200 117.000 378.000 119.800 ;
        RECT 372.200 114.400 376.400 115.200 ;
        RECT 369.000 113.600 371.600 114.400 ;
        RECT 378.800 113.600 379.600 119.800 ;
        RECT 382.000 115.000 382.800 119.800 ;
        RECT 385.200 115.000 386.000 119.800 ;
        RECT 386.800 117.000 387.600 119.800 ;
        RECT 388.400 117.000 389.200 119.800 ;
        RECT 391.600 115.200 392.400 119.800 ;
        RECT 394.800 116.400 395.600 119.800 ;
        RECT 394.800 115.800 395.800 116.400 ;
        RECT 395.200 115.200 395.800 115.800 ;
        RECT 390.400 114.400 394.600 115.200 ;
        RECT 395.200 114.600 397.200 115.200 ;
        RECT 382.000 113.600 384.600 114.400 ;
        RECT 385.200 113.800 391.000 114.400 ;
        RECT 394.000 114.000 394.600 114.400 ;
        RECT 374.000 113.000 374.800 113.200 ;
        RECT 365.800 112.400 374.800 113.000 ;
        RECT 377.200 113.000 378.000 113.200 ;
        RECT 385.200 113.000 385.800 113.800 ;
        RECT 391.600 113.200 393.000 113.800 ;
        RECT 394.000 113.200 395.600 114.000 ;
        RECT 377.200 112.400 385.800 113.000 ;
        RECT 386.800 113.000 393.000 113.200 ;
        RECT 386.800 112.600 392.200 113.000 ;
        RECT 386.800 112.400 387.600 112.600 ;
        RECT 364.200 106.800 365.000 111.200 ;
        RECT 365.800 110.600 366.400 112.400 ;
        RECT 365.600 110.000 366.400 110.600 ;
        RECT 372.400 110.000 395.800 110.600 ;
        RECT 365.600 108.000 366.200 110.000 ;
        RECT 372.400 109.400 373.200 110.000 ;
        RECT 390.000 109.600 390.800 110.000 ;
        RECT 395.000 109.800 395.800 110.000 ;
        RECT 366.800 108.600 370.600 109.400 ;
        RECT 365.600 107.400 366.800 108.000 ;
        RECT 364.200 106.000 365.200 106.800 ;
        RECT 364.400 102.200 365.200 106.000 ;
        RECT 366.000 102.200 366.800 107.400 ;
        RECT 369.800 107.400 370.600 108.600 ;
        RECT 369.800 106.800 371.600 107.400 ;
        RECT 370.800 106.200 371.600 106.800 ;
        RECT 375.600 106.400 376.400 109.200 ;
        RECT 378.800 108.600 382.000 109.400 ;
        RECT 385.800 108.600 387.800 109.400 ;
        RECT 396.400 109.000 397.200 114.600 ;
        RECT 378.400 107.800 379.200 108.000 ;
        RECT 378.400 107.200 382.800 107.800 ;
        RECT 382.000 107.000 382.800 107.200 ;
        RECT 383.600 106.800 384.400 108.400 ;
        RECT 370.800 105.400 373.200 106.200 ;
        RECT 375.600 105.600 376.600 106.400 ;
        RECT 379.600 105.600 381.200 106.400 ;
        RECT 382.000 106.200 382.800 106.400 ;
        RECT 385.800 106.200 386.600 108.600 ;
        RECT 388.400 108.200 397.200 109.000 ;
        RECT 391.800 106.800 394.800 107.600 ;
        RECT 391.800 106.200 392.600 106.800 ;
        RECT 382.000 105.600 386.600 106.200 ;
        RECT 372.400 102.200 373.200 105.400 ;
        RECT 390.000 105.400 392.600 106.200 ;
        RECT 374.000 102.200 374.800 105.000 ;
        RECT 375.600 102.200 376.400 105.000 ;
        RECT 377.200 102.200 378.000 105.000 ;
        RECT 378.800 102.200 379.600 105.000 ;
        RECT 382.000 102.200 382.800 105.000 ;
        RECT 385.200 102.200 386.000 105.000 ;
        RECT 386.800 102.200 387.600 105.000 ;
        RECT 388.400 102.200 389.200 105.000 ;
        RECT 390.000 102.200 390.800 105.400 ;
        RECT 396.400 102.200 397.200 108.200 ;
        RECT 398.000 102.200 398.800 119.800 ;
        RECT 401.200 113.600 402.800 114.400 ;
        RECT 402.000 112.400 402.600 113.600 ;
        RECT 403.400 112.400 404.200 119.800 ;
        RECT 401.200 111.800 402.600 112.400 ;
        RECT 403.200 111.800 404.200 112.400 ;
        RECT 401.200 111.600 402.000 111.800 ;
        RECT 403.200 108.400 403.800 111.800 ;
        RECT 404.400 108.800 405.200 110.400 ;
        RECT 401.200 107.600 403.800 108.400 ;
        RECT 406.000 108.200 406.800 108.400 ;
        RECT 405.200 107.600 406.800 108.200 ;
        RECT 399.600 104.800 400.400 106.400 ;
        RECT 401.400 106.200 402.000 107.600 ;
        RECT 405.200 107.200 406.000 107.600 ;
        RECT 407.600 106.800 408.400 108.400 ;
        RECT 403.000 106.200 406.600 106.600 ;
        RECT 409.200 106.200 410.000 119.800 ;
        RECT 412.400 113.600 414.000 114.400 ;
        RECT 410.800 111.600 411.600 113.200 ;
        RECT 413.200 112.400 413.800 113.600 ;
        RECT 414.600 112.400 415.400 119.800 ;
        RECT 412.400 111.800 413.800 112.400 ;
        RECT 414.400 111.800 415.400 112.400 ;
        RECT 425.200 112.000 426.000 119.800 ;
        RECT 428.400 115.200 429.200 119.800 ;
        RECT 412.400 111.600 413.200 111.800 ;
        RECT 414.400 108.400 415.000 111.800 ;
        RECT 425.000 111.200 426.000 112.000 ;
        RECT 426.600 114.600 429.200 115.200 ;
        RECT 426.600 113.000 427.200 114.600 ;
        RECT 431.600 114.400 432.400 119.800 ;
        RECT 434.800 117.000 435.600 119.800 ;
        RECT 436.400 117.000 437.200 119.800 ;
        RECT 438.000 117.000 438.800 119.800 ;
        RECT 433.000 114.400 437.200 115.200 ;
        RECT 429.800 113.600 432.400 114.400 ;
        RECT 439.600 113.600 440.400 119.800 ;
        RECT 442.800 115.000 443.600 119.800 ;
        RECT 446.000 115.000 446.800 119.800 ;
        RECT 447.600 117.000 448.400 119.800 ;
        RECT 449.200 117.000 450.000 119.800 ;
        RECT 452.400 115.200 453.200 119.800 ;
        RECT 455.600 116.400 456.400 119.800 ;
        RECT 455.600 115.800 456.600 116.400 ;
        RECT 456.000 115.200 456.600 115.800 ;
        RECT 451.200 114.400 455.400 115.200 ;
        RECT 456.000 114.600 458.000 115.200 ;
        RECT 442.800 113.600 445.400 114.400 ;
        RECT 446.000 113.800 451.800 114.400 ;
        RECT 454.800 114.000 455.400 114.400 ;
        RECT 434.800 113.000 435.600 113.200 ;
        RECT 426.600 112.400 435.600 113.000 ;
        RECT 438.000 113.000 438.800 113.200 ;
        RECT 446.000 113.000 446.600 113.800 ;
        RECT 452.400 113.200 453.800 113.800 ;
        RECT 454.800 113.200 456.400 114.000 ;
        RECT 438.000 112.400 446.600 113.000 ;
        RECT 447.600 113.000 453.800 113.200 ;
        RECT 447.600 112.600 453.000 113.000 ;
        RECT 447.600 112.400 448.400 112.600 ;
        RECT 415.600 108.800 416.400 110.400 ;
        RECT 412.400 107.600 415.000 108.400 ;
        RECT 417.200 108.200 418.000 108.400 ;
        RECT 416.400 107.600 418.000 108.200 ;
        RECT 412.600 106.200 413.200 107.600 ;
        RECT 416.400 107.200 417.200 107.600 ;
        RECT 425.000 106.800 425.800 111.200 ;
        RECT 426.600 110.600 427.200 112.400 ;
        RECT 426.400 110.000 427.200 110.600 ;
        RECT 433.200 110.000 456.600 110.600 ;
        RECT 426.400 108.000 427.000 110.000 ;
        RECT 433.200 109.400 434.000 110.000 ;
        RECT 450.800 109.600 451.600 110.000 ;
        RECT 454.000 109.600 454.800 110.000 ;
        RECT 455.800 109.800 456.600 110.000 ;
        RECT 427.600 108.600 431.400 109.400 ;
        RECT 426.400 107.400 427.600 108.000 ;
        RECT 414.200 106.200 417.800 106.600 ;
        RECT 401.200 102.200 402.000 106.200 ;
        RECT 402.800 106.000 406.800 106.200 ;
        RECT 402.800 102.200 403.600 106.000 ;
        RECT 406.000 102.200 406.800 106.000 ;
        RECT 409.200 105.600 411.000 106.200 ;
        RECT 410.200 102.200 411.000 105.600 ;
        RECT 412.400 102.200 413.200 106.200 ;
        RECT 414.000 106.000 418.000 106.200 ;
        RECT 425.000 106.000 426.000 106.800 ;
        RECT 414.000 102.200 414.800 106.000 ;
        RECT 417.200 102.200 418.000 106.000 ;
        RECT 425.200 102.200 426.000 106.000 ;
        RECT 426.800 102.200 427.600 107.400 ;
        RECT 430.600 107.400 431.400 108.600 ;
        RECT 430.600 106.800 432.400 107.400 ;
        RECT 431.600 106.200 432.400 106.800 ;
        RECT 436.400 106.400 437.200 109.200 ;
        RECT 439.600 108.600 442.800 109.400 ;
        RECT 446.600 108.600 448.600 109.400 ;
        RECT 457.200 109.000 458.000 114.600 ;
        RECT 460.400 112.800 461.200 119.800 ;
        RECT 439.200 107.800 440.000 108.000 ;
        RECT 439.200 107.200 443.600 107.800 ;
        RECT 442.800 107.000 443.600 107.200 ;
        RECT 444.400 106.800 445.200 108.400 ;
        RECT 431.600 105.400 434.000 106.200 ;
        RECT 436.400 105.600 437.400 106.400 ;
        RECT 440.400 105.600 442.000 106.400 ;
        RECT 442.800 106.200 443.600 106.400 ;
        RECT 446.600 106.200 447.400 108.600 ;
        RECT 449.200 108.200 458.000 109.000 ;
        RECT 460.200 111.800 461.200 112.800 ;
        RECT 463.600 112.400 464.400 119.800 ;
        RECT 461.800 111.800 464.400 112.400 ;
        RECT 467.800 112.400 468.600 119.800 ;
        RECT 469.200 114.300 470.000 114.400 ;
        RECT 471.600 114.300 472.400 114.400 ;
        RECT 469.200 113.700 472.400 114.300 ;
        RECT 469.200 113.600 470.000 113.700 ;
        RECT 471.600 113.600 472.400 113.700 ;
        RECT 469.400 112.400 470.000 113.600 ;
        RECT 467.800 111.800 468.800 112.400 ;
        RECT 469.400 111.800 470.800 112.400 ;
        RECT 460.200 108.400 460.800 111.800 ;
        RECT 461.800 109.800 462.400 111.800 ;
        RECT 461.400 109.000 462.400 109.800 ;
        RECT 452.600 106.800 455.600 107.600 ;
        RECT 452.600 106.200 453.400 106.800 ;
        RECT 442.800 105.600 447.400 106.200 ;
        RECT 433.200 102.200 434.000 105.400 ;
        RECT 450.800 105.400 453.400 106.200 ;
        RECT 434.800 102.200 435.600 105.000 ;
        RECT 436.400 102.200 437.200 105.000 ;
        RECT 438.000 102.200 438.800 105.000 ;
        RECT 439.600 102.200 440.400 105.000 ;
        RECT 442.800 102.200 443.600 105.000 ;
        RECT 446.000 102.200 446.800 105.000 ;
        RECT 447.600 102.200 448.400 105.000 ;
        RECT 449.200 102.200 450.000 105.000 ;
        RECT 450.800 102.200 451.600 105.400 ;
        RECT 457.200 102.200 458.000 108.200 ;
        RECT 458.800 108.300 459.600 108.400 ;
        RECT 460.200 108.300 461.200 108.400 ;
        RECT 458.800 107.700 461.200 108.300 ;
        RECT 458.800 107.600 459.600 107.700 ;
        RECT 460.200 107.600 461.200 107.700 ;
        RECT 460.200 106.200 460.800 107.600 ;
        RECT 461.800 107.400 462.400 109.000 ;
        RECT 463.400 109.600 464.400 110.400 ;
        RECT 463.400 108.800 464.200 109.600 ;
        RECT 466.800 108.800 467.600 110.400 ;
        RECT 468.200 108.400 468.800 111.800 ;
        RECT 470.000 111.600 470.800 111.800 ;
        RECT 465.200 108.200 466.000 108.400 ;
        RECT 465.200 107.600 466.800 108.200 ;
        RECT 468.200 107.600 470.800 108.400 ;
        RECT 461.800 106.800 464.400 107.400 ;
        RECT 466.000 107.200 466.800 107.600 ;
        RECT 460.200 105.600 461.200 106.200 ;
        RECT 460.400 102.200 461.200 105.600 ;
        RECT 463.600 102.200 464.400 106.800 ;
        RECT 465.400 106.200 469.000 106.600 ;
        RECT 470.000 106.200 470.600 107.600 ;
        RECT 471.600 106.800 472.400 108.400 ;
        RECT 473.200 106.200 474.000 119.800 ;
        RECT 474.800 111.600 475.600 113.200 ;
        RECT 476.400 106.800 477.200 108.400 ;
        RECT 478.000 108.300 478.800 119.800 ;
        RECT 479.600 111.600 480.400 113.200 ;
        RECT 482.800 112.000 483.600 119.800 ;
        RECT 486.000 115.200 486.800 119.800 ;
        RECT 482.600 111.200 483.600 112.000 ;
        RECT 484.200 114.600 486.800 115.200 ;
        RECT 484.200 113.000 484.800 114.600 ;
        RECT 489.200 114.400 490.000 119.800 ;
        RECT 492.400 117.000 493.200 119.800 ;
        RECT 494.000 117.000 494.800 119.800 ;
        RECT 495.600 117.000 496.400 119.800 ;
        RECT 490.600 114.400 494.800 115.200 ;
        RECT 487.400 113.600 490.000 114.400 ;
        RECT 497.200 113.600 498.000 119.800 ;
        RECT 500.400 115.000 501.200 119.800 ;
        RECT 503.600 115.000 504.400 119.800 ;
        RECT 505.200 117.000 506.000 119.800 ;
        RECT 506.800 117.000 507.600 119.800 ;
        RECT 510.000 115.200 510.800 119.800 ;
        RECT 513.200 116.400 514.000 119.800 ;
        RECT 513.200 115.800 514.200 116.400 ;
        RECT 513.600 115.200 514.200 115.800 ;
        RECT 508.800 114.400 513.000 115.200 ;
        RECT 513.600 114.600 515.600 115.200 ;
        RECT 500.400 113.600 503.000 114.400 ;
        RECT 503.600 113.800 509.400 114.400 ;
        RECT 512.400 114.000 513.000 114.400 ;
        RECT 492.400 113.000 493.200 113.200 ;
        RECT 484.200 112.400 493.200 113.000 ;
        RECT 495.600 113.000 496.400 113.200 ;
        RECT 503.600 113.000 504.200 113.800 ;
        RECT 510.000 113.200 511.400 113.800 ;
        RECT 512.400 113.200 514.000 114.000 ;
        RECT 495.600 112.400 504.200 113.000 ;
        RECT 505.200 113.000 511.400 113.200 ;
        RECT 505.200 112.600 510.600 113.000 ;
        RECT 505.200 112.400 506.000 112.600 ;
        RECT 481.200 108.300 482.000 108.400 ;
        RECT 478.000 107.700 482.000 108.300 ;
        RECT 478.000 106.200 478.800 107.700 ;
        RECT 481.200 107.600 482.000 107.700 ;
        RECT 482.600 106.800 483.400 111.200 ;
        RECT 484.200 110.600 484.800 112.400 ;
        RECT 484.000 110.000 484.800 110.600 ;
        RECT 490.800 110.000 514.200 110.600 ;
        RECT 484.000 108.000 484.600 110.000 ;
        RECT 490.800 109.400 491.600 110.000 ;
        RECT 508.400 109.600 509.200 110.000 ;
        RECT 511.600 109.600 512.400 110.000 ;
        RECT 513.400 109.800 514.200 110.000 ;
        RECT 485.200 108.600 489.000 109.400 ;
        RECT 484.000 107.400 485.200 108.000 ;
        RECT 465.200 106.000 469.200 106.200 ;
        RECT 465.200 102.200 466.000 106.000 ;
        RECT 468.400 102.200 469.200 106.000 ;
        RECT 470.000 102.200 470.800 106.200 ;
        RECT 473.200 105.600 475.000 106.200 ;
        RECT 478.000 105.600 479.800 106.200 ;
        RECT 482.600 106.000 483.600 106.800 ;
        RECT 474.200 104.400 475.000 105.600 ;
        RECT 474.200 103.600 475.600 104.400 ;
        RECT 474.200 102.200 475.000 103.600 ;
        RECT 479.000 102.200 479.800 105.600 ;
        RECT 482.800 102.200 483.600 106.000 ;
        RECT 484.400 102.200 485.200 107.400 ;
        RECT 488.200 107.400 489.000 108.600 ;
        RECT 488.200 106.800 490.000 107.400 ;
        RECT 489.200 106.200 490.000 106.800 ;
        RECT 494.000 106.400 494.800 109.200 ;
        RECT 497.200 108.600 500.400 109.400 ;
        RECT 504.200 108.600 506.200 109.400 ;
        RECT 514.800 109.000 515.600 114.600 ;
        RECT 518.000 112.800 518.800 119.800 ;
        RECT 496.800 107.800 497.600 108.000 ;
        RECT 496.800 107.200 501.200 107.800 ;
        RECT 500.400 107.000 501.200 107.200 ;
        RECT 502.000 106.800 502.800 108.400 ;
        RECT 489.200 105.400 491.600 106.200 ;
        RECT 494.000 105.600 495.000 106.400 ;
        RECT 498.000 105.600 499.600 106.400 ;
        RECT 500.400 106.200 501.200 106.400 ;
        RECT 504.200 106.200 505.000 108.600 ;
        RECT 506.800 108.200 515.600 109.000 ;
        RECT 517.800 111.800 518.800 112.800 ;
        RECT 521.200 112.400 522.000 119.800 ;
        RECT 525.000 114.400 525.800 119.800 ;
        RECT 523.600 113.600 524.400 114.400 ;
        RECT 525.000 113.600 526.800 114.400 ;
        RECT 523.600 112.400 524.200 113.600 ;
        RECT 525.000 112.400 525.800 113.600 ;
        RECT 519.400 111.800 522.000 112.400 ;
        RECT 522.800 111.800 524.200 112.400 ;
        RECT 524.800 111.800 525.800 112.400 ;
        RECT 517.800 108.400 518.400 111.800 ;
        RECT 519.400 109.800 520.000 111.800 ;
        RECT 522.800 111.600 523.600 111.800 ;
        RECT 519.000 109.000 520.000 109.800 ;
        RECT 510.200 106.800 513.200 107.600 ;
        RECT 510.200 106.200 511.000 106.800 ;
        RECT 500.400 105.600 505.000 106.200 ;
        RECT 490.800 102.200 491.600 105.400 ;
        RECT 508.400 105.400 511.000 106.200 ;
        RECT 492.400 102.200 493.200 105.000 ;
        RECT 494.000 102.200 494.800 105.000 ;
        RECT 495.600 102.200 496.400 105.000 ;
        RECT 497.200 102.200 498.000 105.000 ;
        RECT 500.400 102.200 501.200 105.000 ;
        RECT 503.600 102.200 504.400 105.000 ;
        RECT 505.200 102.200 506.000 105.000 ;
        RECT 506.800 102.200 507.600 105.000 ;
        RECT 508.400 102.200 509.200 105.400 ;
        RECT 514.800 102.200 515.600 108.200 ;
        RECT 516.400 108.300 517.200 108.400 ;
        RECT 517.800 108.300 518.800 108.400 ;
        RECT 516.400 107.700 518.800 108.300 ;
        RECT 516.400 107.600 517.200 107.700 ;
        RECT 517.800 107.600 518.800 107.700 ;
        RECT 517.800 106.200 518.400 107.600 ;
        RECT 519.400 107.400 520.000 109.000 ;
        RECT 521.000 109.600 522.000 110.400 ;
        RECT 521.000 108.800 521.800 109.600 ;
        RECT 524.800 108.400 525.400 111.800 ;
        RECT 530.800 111.200 531.600 119.800 ;
        RECT 534.000 111.200 534.800 119.800 ;
        RECT 537.200 111.200 538.000 119.800 ;
        RECT 540.400 111.200 541.200 119.800 ;
        RECT 544.400 113.600 545.200 114.400 ;
        RECT 544.400 112.400 545.000 113.600 ;
        RECT 545.800 112.400 546.600 119.800 ;
        RECT 543.600 111.800 545.000 112.400 ;
        RECT 545.600 111.800 546.600 112.400 ;
        RECT 543.600 111.600 544.400 111.800 ;
        RECT 529.200 110.400 531.600 111.200 ;
        RECT 532.600 110.400 534.800 111.200 ;
        RECT 535.800 110.400 538.000 111.200 ;
        RECT 539.400 110.400 541.200 111.200 ;
        RECT 526.000 108.800 526.800 110.400 ;
        RECT 522.800 107.600 525.400 108.400 ;
        RECT 527.600 108.200 528.400 108.400 ;
        RECT 526.800 107.600 528.400 108.200 ;
        RECT 529.200 107.600 530.000 110.400 ;
        RECT 532.600 109.000 533.400 110.400 ;
        RECT 535.800 109.000 536.600 110.400 ;
        RECT 539.400 109.000 540.200 110.400 ;
        RECT 542.000 110.300 542.800 110.400 ;
        RECT 545.600 110.300 546.200 111.800 ;
        RECT 542.000 109.700 546.200 110.300 ;
        RECT 542.000 109.600 542.800 109.700 ;
        RECT 530.800 108.200 533.400 109.000 ;
        RECT 534.200 108.200 536.600 109.000 ;
        RECT 537.600 108.200 540.200 109.000 ;
        RECT 541.000 108.200 542.800 109.000 ;
        RECT 545.600 108.400 546.200 109.700 ;
        RECT 546.800 108.800 547.600 110.400 ;
        RECT 532.600 107.600 533.400 108.200 ;
        RECT 535.800 107.600 536.600 108.200 ;
        RECT 539.400 107.600 540.200 108.200 ;
        RECT 542.000 107.600 542.800 108.200 ;
        RECT 543.600 107.600 546.200 108.400 ;
        RECT 548.400 108.200 549.200 108.400 ;
        RECT 547.600 107.600 549.200 108.200 ;
        RECT 519.400 106.800 522.000 107.400 ;
        RECT 517.800 105.600 518.800 106.200 ;
        RECT 518.000 102.200 518.800 105.600 ;
        RECT 521.200 102.200 522.000 106.800 ;
        RECT 523.000 106.200 523.600 107.600 ;
        RECT 526.800 107.200 527.600 107.600 ;
        RECT 529.200 106.800 531.600 107.600 ;
        RECT 532.600 106.800 534.800 107.600 ;
        RECT 535.800 106.800 538.000 107.600 ;
        RECT 539.400 106.800 541.200 107.600 ;
        RECT 524.600 106.200 528.200 106.600 ;
        RECT 522.800 102.200 523.600 106.200 ;
        RECT 524.400 106.000 528.400 106.200 ;
        RECT 524.400 102.200 525.200 106.000 ;
        RECT 527.600 102.200 528.400 106.000 ;
        RECT 530.800 102.200 531.600 106.800 ;
        RECT 534.000 102.200 534.800 106.800 ;
        RECT 537.200 102.200 538.000 106.800 ;
        RECT 540.400 102.200 541.200 106.800 ;
        RECT 543.800 106.200 544.400 107.600 ;
        RECT 547.600 107.200 548.400 107.600 ;
        RECT 550.000 106.800 550.800 108.400 ;
        RECT 545.400 106.200 549.000 106.600 ;
        RECT 551.600 106.200 552.400 119.800 ;
        RECT 553.200 111.600 554.000 113.200 ;
        RECT 558.600 112.800 559.400 119.800 ;
        RECT 562.800 115.000 563.600 119.000 ;
        RECT 557.800 112.200 559.400 112.800 ;
        RECT 556.400 109.600 557.200 111.200 ;
        RECT 557.800 108.400 558.400 112.200 ;
        RECT 563.000 111.600 563.600 115.000 ;
        RECT 564.400 112.400 565.200 119.800 ;
        RECT 567.600 112.800 568.400 119.800 ;
        RECT 564.400 111.800 567.000 112.400 ;
        RECT 567.600 111.800 568.600 112.800 ;
        RECT 559.800 111.000 563.600 111.600 ;
        RECT 559.800 109.000 560.400 111.000 ;
        RECT 553.200 108.300 554.000 108.400 ;
        RECT 556.400 108.300 558.400 108.400 ;
        RECT 553.200 107.700 558.400 108.300 ;
        RECT 559.000 108.200 560.400 109.000 ;
        RECT 561.200 108.800 562.000 110.400 ;
        RECT 562.800 108.800 563.600 110.400 ;
        RECT 564.400 109.600 565.400 110.400 ;
        RECT 564.600 108.800 565.400 109.600 ;
        RECT 566.400 109.800 567.000 111.800 ;
        RECT 566.400 109.000 567.400 109.800 ;
        RECT 553.200 107.600 554.000 107.700 ;
        RECT 556.400 107.600 558.400 107.700 ;
        RECT 557.800 107.000 558.400 107.600 ;
        RECT 559.400 107.800 560.400 108.200 ;
        RECT 559.400 107.200 563.600 107.800 ;
        RECT 566.400 107.400 567.000 109.000 ;
        RECT 568.000 108.400 568.600 111.800 ;
        RECT 567.600 107.600 568.600 108.400 ;
        RECT 574.000 108.300 574.800 108.400 ;
        RECT 575.600 108.300 576.400 108.400 ;
        RECT 574.000 107.700 576.400 108.300 ;
        RECT 574.000 107.600 574.800 107.700 ;
        RECT 557.800 106.600 558.600 107.000 ;
        RECT 543.600 102.200 544.400 106.200 ;
        RECT 545.200 106.000 549.200 106.200 ;
        RECT 545.200 102.200 546.000 106.000 ;
        RECT 548.400 102.200 549.200 106.000 ;
        RECT 551.600 105.600 553.400 106.200 ;
        RECT 557.800 106.000 559.400 106.600 ;
        RECT 552.600 102.200 553.400 105.600 ;
        RECT 558.600 103.000 559.400 106.000 ;
        RECT 563.000 105.000 563.600 107.200 ;
        RECT 562.800 103.000 563.600 105.000 ;
        RECT 564.400 106.800 567.000 107.400 ;
        RECT 564.400 102.200 565.200 106.800 ;
        RECT 568.000 106.200 568.600 107.600 ;
        RECT 575.600 106.800 576.400 107.700 ;
        RECT 567.600 105.600 568.600 106.200 ;
        RECT 577.200 106.200 578.000 119.800 ;
        RECT 578.800 112.300 579.600 113.200 ;
        RECT 580.400 112.300 581.200 119.800 ;
        RECT 585.800 118.400 586.600 119.800 ;
        RECT 585.800 117.600 587.600 118.400 ;
        RECT 584.400 113.600 585.200 114.400 ;
        RECT 584.400 112.400 585.000 113.600 ;
        RECT 585.800 112.400 586.600 117.600 ;
        RECT 592.600 112.400 593.400 119.800 ;
        RECT 594.000 113.600 594.800 114.400 ;
        RECT 594.200 112.400 594.800 113.600 ;
        RECT 578.800 111.700 581.200 112.300 ;
        RECT 578.800 111.600 579.600 111.700 ;
        RECT 577.200 105.600 579.000 106.200 ;
        RECT 567.600 102.200 568.400 105.600 ;
        RECT 578.200 104.400 579.000 105.600 ;
        RECT 577.200 103.600 579.000 104.400 ;
        RECT 578.200 102.200 579.000 103.600 ;
        RECT 580.400 102.200 581.200 111.700 ;
        RECT 583.600 111.800 585.000 112.400 ;
        RECT 585.600 111.800 586.600 112.400 ;
        RECT 583.600 111.600 584.400 111.800 ;
        RECT 585.600 108.400 586.200 111.800 ;
        RECT 591.600 111.600 593.600 112.400 ;
        RECT 594.200 111.800 595.600 112.400 ;
        RECT 594.800 111.600 595.600 111.800 ;
        RECT 596.400 111.600 597.200 113.200 ;
        RECT 586.800 108.800 587.600 110.400 ;
        RECT 590.000 110.300 590.800 110.400 ;
        RECT 591.600 110.300 592.400 110.400 ;
        RECT 590.000 109.700 592.400 110.300 ;
        RECT 590.000 109.600 590.800 109.700 ;
        RECT 591.600 108.800 592.400 109.700 ;
        RECT 593.000 108.400 593.600 111.600 ;
        RECT 594.900 110.300 595.500 111.600 ;
        RECT 598.000 110.300 598.800 119.800 ;
        RECT 594.900 109.700 598.800 110.300 ;
        RECT 583.600 107.600 586.200 108.400 ;
        RECT 588.400 108.200 589.200 108.400 ;
        RECT 587.600 107.600 589.200 108.200 ;
        RECT 590.000 108.200 590.800 108.400 ;
        RECT 590.000 107.600 591.600 108.200 ;
        RECT 593.000 107.600 595.600 108.400 ;
        RECT 582.000 104.800 582.800 106.400 ;
        RECT 583.800 106.200 584.400 107.600 ;
        RECT 587.600 107.200 588.400 107.600 ;
        RECT 590.800 107.200 591.600 107.600 ;
        RECT 585.400 106.200 589.000 106.600 ;
        RECT 590.200 106.200 593.800 106.600 ;
        RECT 594.800 106.200 595.400 107.600 ;
        RECT 598.000 106.200 598.800 109.700 ;
        RECT 599.600 106.800 600.400 108.400 ;
        RECT 583.600 102.200 584.400 106.200 ;
        RECT 585.200 106.000 589.200 106.200 ;
        RECT 585.200 102.200 586.000 106.000 ;
        RECT 588.400 102.200 589.200 106.000 ;
        RECT 590.000 106.000 594.000 106.200 ;
        RECT 590.000 102.200 590.800 106.000 ;
        RECT 593.200 102.200 594.000 106.000 ;
        RECT 594.800 102.200 595.600 106.200 ;
        RECT 597.000 105.600 598.800 106.200 ;
        RECT 597.000 102.200 597.800 105.600 ;
        RECT 601.200 102.200 602.000 119.800 ;
        RECT 604.400 111.200 605.200 119.800 ;
        RECT 608.600 115.800 609.800 119.800 ;
        RECT 613.200 115.800 614.000 119.800 ;
        RECT 617.600 116.400 618.400 119.800 ;
        RECT 617.600 115.800 619.600 116.400 ;
        RECT 609.200 115.000 610.000 115.800 ;
        RECT 613.400 115.200 614.000 115.800 ;
        RECT 612.600 114.600 616.200 115.200 ;
        RECT 618.800 115.000 619.600 115.800 ;
        RECT 612.600 114.400 613.400 114.600 ;
        RECT 615.400 114.400 616.200 114.600 ;
        RECT 607.600 114.000 609.000 114.400 ;
        RECT 607.600 113.600 609.800 114.000 ;
        RECT 608.400 113.200 609.800 113.600 ;
        RECT 609.200 112.200 609.800 113.200 ;
        RECT 611.400 113.000 613.600 113.600 ;
        RECT 611.400 112.800 612.200 113.000 ;
        RECT 609.200 111.600 611.600 112.200 ;
        RECT 604.400 110.600 608.600 111.200 ;
        RECT 604.400 107.200 605.200 110.600 ;
        RECT 607.800 110.400 608.600 110.600 ;
        RECT 606.200 109.800 607.000 110.000 ;
        RECT 606.200 109.200 610.000 109.800 ;
        RECT 609.200 109.000 610.000 109.200 ;
        RECT 611.000 108.400 611.600 111.600 ;
        RECT 613.000 111.800 613.600 113.000 ;
        RECT 614.200 113.000 615.000 113.200 ;
        RECT 618.800 113.000 619.600 113.200 ;
        RECT 614.200 112.400 619.600 113.000 ;
        RECT 613.000 111.400 617.800 111.800 ;
        RECT 622.000 111.400 622.800 119.800 ;
        RECT 626.200 114.400 627.000 119.800 ;
        RECT 625.200 113.600 627.000 114.400 ;
        RECT 627.600 113.600 628.400 114.400 ;
        RECT 626.200 112.400 627.000 113.600 ;
        RECT 627.800 112.400 628.400 113.600 ;
        RECT 630.800 113.600 631.600 114.400 ;
        RECT 630.800 112.400 631.400 113.600 ;
        RECT 632.200 112.400 633.000 119.800 ;
        RECT 626.200 111.800 627.200 112.400 ;
        RECT 627.800 111.800 629.200 112.400 ;
        RECT 613.000 111.200 622.800 111.400 ;
        RECT 617.000 111.000 622.800 111.200 ;
        RECT 617.200 110.800 622.800 111.000 ;
        RECT 615.600 110.200 616.400 110.400 ;
        RECT 615.600 109.600 620.600 110.200 ;
        RECT 617.200 109.400 618.000 109.600 ;
        RECT 619.800 109.400 620.600 109.600 ;
        RECT 625.200 108.800 626.000 110.400 ;
        RECT 618.200 108.400 619.000 108.600 ;
        RECT 626.600 108.400 627.200 111.800 ;
        RECT 628.400 111.600 629.200 111.800 ;
        RECT 630.000 111.800 631.400 112.400 ;
        RECT 632.000 111.800 633.000 112.400 ;
        RECT 636.400 115.000 637.200 119.000 ;
        RECT 640.600 118.400 641.400 119.800 ;
        RECT 639.600 117.600 641.400 118.400 ;
        RECT 630.000 111.600 630.800 111.800 ;
        RECT 628.500 110.300 629.100 111.600 ;
        RECT 632.000 110.300 632.600 111.800 ;
        RECT 636.400 111.600 637.000 115.000 ;
        RECT 640.600 112.800 641.400 117.600 ;
        RECT 647.600 112.800 648.400 119.800 ;
        RECT 640.600 112.200 642.200 112.800 ;
        RECT 636.400 111.000 640.200 111.600 ;
        RECT 628.500 109.700 632.600 110.300 ;
        RECT 632.000 108.400 632.600 109.700 ;
        RECT 633.200 110.300 634.000 110.400 ;
        RECT 634.800 110.300 635.600 110.400 ;
        RECT 633.200 109.700 635.600 110.300 ;
        RECT 633.200 108.800 634.000 109.700 ;
        RECT 634.800 109.600 635.600 109.700 ;
        RECT 636.400 108.800 637.200 110.400 ;
        RECT 638.000 108.800 638.800 110.400 ;
        RECT 639.600 109.000 640.200 111.000 ;
        RECT 611.000 107.800 622.000 108.400 ;
        RECT 611.400 107.600 612.200 107.800 ;
        RECT 604.400 106.600 608.200 107.200 ;
        RECT 602.800 106.300 603.600 106.400 ;
        RECT 604.400 106.300 605.200 106.600 ;
        RECT 607.400 106.400 608.200 106.600 ;
        RECT 602.800 105.700 605.200 106.300 ;
        RECT 602.800 104.800 603.600 105.700 ;
        RECT 604.400 102.200 605.200 105.700 ;
        RECT 617.200 105.600 617.800 107.800 ;
        RECT 620.400 107.600 622.000 107.800 ;
        RECT 623.600 108.200 624.400 108.400 ;
        RECT 623.600 107.600 625.200 108.200 ;
        RECT 626.600 107.600 629.200 108.400 ;
        RECT 630.000 107.600 632.600 108.400 ;
        RECT 634.800 108.200 635.600 108.400 ;
        RECT 634.000 107.600 635.600 108.200 ;
        RECT 639.600 108.200 641.000 109.000 ;
        RECT 641.600 108.400 642.200 112.200 ;
        RECT 647.400 111.800 648.400 112.800 ;
        RECT 650.800 112.400 651.600 119.800 ;
        RECT 654.000 112.800 654.800 119.800 ;
        RECT 649.000 111.800 651.600 112.400 ;
        RECT 653.800 111.800 654.800 112.800 ;
        RECT 657.200 112.400 658.000 119.800 ;
        RECT 655.400 111.800 658.000 112.400 ;
        RECT 642.800 109.600 643.600 111.200 ;
        RECT 647.400 108.400 648.000 111.800 ;
        RECT 649.000 109.800 649.600 111.800 ;
        RECT 648.600 109.000 649.600 109.800 ;
        RECT 639.600 107.800 640.600 108.200 ;
        RECT 624.400 107.200 625.200 107.600 ;
        RECT 615.400 105.400 616.200 105.600 ;
        RECT 609.200 104.200 610.000 105.000 ;
        RECT 613.400 104.800 616.200 105.400 ;
        RECT 617.200 104.800 618.000 105.600 ;
        RECT 613.400 104.200 614.000 104.800 ;
        RECT 618.800 104.200 619.600 105.000 ;
        RECT 608.600 103.600 610.000 104.200 ;
        RECT 608.600 102.200 609.800 103.600 ;
        RECT 613.200 102.200 614.000 104.200 ;
        RECT 617.600 103.600 619.600 104.200 ;
        RECT 617.600 102.200 618.400 103.600 ;
        RECT 622.000 102.200 622.800 107.000 ;
        RECT 623.800 106.200 627.400 106.600 ;
        RECT 628.400 106.200 629.000 107.600 ;
        RECT 630.200 106.200 630.800 107.600 ;
        RECT 634.000 107.200 634.800 107.600 ;
        RECT 636.400 107.200 640.600 107.800 ;
        RECT 641.600 107.600 643.600 108.400 ;
        RECT 647.400 107.600 648.400 108.400 ;
        RECT 631.800 106.200 635.400 106.600 ;
        RECT 623.600 106.000 627.600 106.200 ;
        RECT 623.600 102.200 624.400 106.000 ;
        RECT 626.800 102.200 627.600 106.000 ;
        RECT 628.400 102.200 629.200 106.200 ;
        RECT 630.000 102.200 630.800 106.200 ;
        RECT 631.600 106.000 635.600 106.200 ;
        RECT 631.600 102.200 632.400 106.000 ;
        RECT 634.800 102.200 635.600 106.000 ;
        RECT 636.400 105.000 637.000 107.200 ;
        RECT 641.600 107.000 642.200 107.600 ;
        RECT 641.400 106.600 642.200 107.000 ;
        RECT 640.600 106.000 642.200 106.600 ;
        RECT 647.400 106.400 648.000 107.600 ;
        RECT 649.000 107.400 649.600 109.000 ;
        RECT 650.600 110.300 651.600 110.400 ;
        RECT 652.400 110.300 653.200 110.400 ;
        RECT 650.600 109.700 653.200 110.300 ;
        RECT 650.600 109.600 651.600 109.700 ;
        RECT 652.400 109.600 653.200 109.700 ;
        RECT 650.600 108.800 651.400 109.600 ;
        RECT 653.800 108.400 654.400 111.800 ;
        RECT 655.400 109.800 656.000 111.800 ;
        RECT 660.400 111.200 661.200 119.800 ;
        RECT 663.600 111.200 664.400 119.800 ;
        RECT 666.800 111.200 667.600 119.800 ;
        RECT 670.000 111.200 670.800 119.800 ;
        RECT 675.800 112.400 676.600 119.800 ;
        RECT 679.600 115.000 680.400 119.000 ;
        RECT 677.200 113.600 678.000 114.400 ;
        RECT 677.400 112.400 678.000 113.600 ;
        RECT 675.800 111.800 676.800 112.400 ;
        RECT 677.400 111.800 678.800 112.400 ;
        RECT 658.800 110.400 661.200 111.200 ;
        RECT 662.200 110.400 664.400 111.200 ;
        RECT 665.400 110.400 667.600 111.200 ;
        RECT 669.000 110.400 670.800 111.200 ;
        RECT 655.000 109.000 656.000 109.800 ;
        RECT 653.800 107.600 654.800 108.400 ;
        RECT 649.000 106.800 651.600 107.400 ;
        RECT 636.400 103.000 637.200 105.000 ;
        RECT 640.600 103.000 641.400 106.000 ;
        RECT 647.400 105.600 648.400 106.400 ;
        RECT 647.600 102.200 648.400 105.600 ;
        RECT 650.800 102.200 651.600 106.800 ;
        RECT 653.800 106.200 654.400 107.600 ;
        RECT 655.400 107.400 656.000 109.000 ;
        RECT 657.000 109.600 658.000 110.400 ;
        RECT 657.000 108.800 657.800 109.600 ;
        RECT 658.800 107.600 659.600 110.400 ;
        RECT 662.200 109.000 663.000 110.400 ;
        RECT 665.400 109.000 666.200 110.400 ;
        RECT 669.000 109.000 669.800 110.400 ;
        RECT 660.400 108.200 663.000 109.000 ;
        RECT 663.800 108.200 666.200 109.000 ;
        RECT 667.200 108.200 669.800 109.000 ;
        RECT 670.600 108.200 672.400 109.000 ;
        RECT 674.800 108.800 675.600 110.400 ;
        RECT 676.200 108.400 676.800 111.800 ;
        RECT 678.000 111.600 678.800 111.800 ;
        RECT 679.600 111.600 680.200 115.000 ;
        RECT 683.800 112.800 684.600 119.800 ;
        RECT 683.800 112.200 685.400 112.800 ;
        RECT 679.600 111.000 683.400 111.600 ;
        RECT 679.600 108.800 680.400 110.400 ;
        RECT 681.200 108.800 682.000 110.400 ;
        RECT 682.800 109.000 683.400 111.000 ;
        RECT 662.200 107.600 663.000 108.200 ;
        RECT 665.400 107.600 666.200 108.200 ;
        RECT 669.000 107.600 669.800 108.200 ;
        RECT 671.600 107.600 672.400 108.200 ;
        RECT 673.200 108.200 674.000 108.400 ;
        RECT 673.200 107.600 674.800 108.200 ;
        RECT 676.200 107.600 678.800 108.400 ;
        RECT 682.800 108.200 684.200 109.000 ;
        RECT 684.800 108.400 685.400 112.200 ;
        RECT 686.000 109.600 686.800 111.200 ;
        RECT 682.800 107.800 683.800 108.200 ;
        RECT 655.400 106.800 658.000 107.400 ;
        RECT 658.800 106.800 661.200 107.600 ;
        RECT 662.200 106.800 664.400 107.600 ;
        RECT 665.400 106.800 667.600 107.600 ;
        RECT 669.000 106.800 670.800 107.600 ;
        RECT 674.000 107.200 674.800 107.600 ;
        RECT 653.800 105.600 654.800 106.200 ;
        RECT 654.000 102.200 654.800 105.600 ;
        RECT 657.200 102.200 658.000 106.800 ;
        RECT 660.400 102.200 661.200 106.800 ;
        RECT 663.600 102.200 664.400 106.800 ;
        RECT 666.800 102.200 667.600 106.800 ;
        RECT 670.000 102.200 670.800 106.800 ;
        RECT 673.400 106.200 677.000 106.600 ;
        RECT 678.000 106.200 678.600 107.600 ;
        RECT 679.600 107.200 683.800 107.800 ;
        RECT 684.800 107.600 686.800 108.400 ;
        RECT 673.200 106.000 677.200 106.200 ;
        RECT 673.200 102.200 674.000 106.000 ;
        RECT 676.400 102.200 677.200 106.000 ;
        RECT 678.000 102.200 678.800 106.200 ;
        RECT 679.600 105.000 680.200 107.200 ;
        RECT 684.800 107.000 685.400 107.600 ;
        RECT 684.600 106.600 685.400 107.000 ;
        RECT 683.800 106.000 685.400 106.600 ;
        RECT 679.600 103.000 680.400 105.000 ;
        RECT 683.800 104.400 684.600 106.000 ;
        RECT 682.800 103.600 684.600 104.400 ;
        RECT 683.800 103.000 684.600 103.600 ;
        RECT 1.200 95.800 2.000 99.800 ;
        RECT 2.800 96.000 3.600 99.800 ;
        RECT 6.000 96.000 6.800 99.800 ;
        RECT 11.400 96.000 12.200 99.000 ;
        RECT 15.600 97.000 16.400 99.000 ;
        RECT 2.800 95.800 6.800 96.000 ;
        RECT 1.400 94.400 2.000 95.800 ;
        RECT 3.000 95.400 6.600 95.800 ;
        RECT 10.600 95.400 12.200 96.000 ;
        RECT 10.600 95.000 11.400 95.400 ;
        RECT 5.200 94.400 6.000 94.800 ;
        RECT 10.600 94.400 11.200 95.000 ;
        RECT 15.800 94.800 16.400 97.000 ;
        RECT 17.200 95.800 18.000 99.800 ;
        RECT 18.800 96.000 19.600 99.800 ;
        RECT 22.000 96.000 22.800 99.800 ;
        RECT 18.800 95.800 22.800 96.000 ;
        RECT 23.600 95.800 24.400 99.800 ;
        RECT 25.200 96.000 26.000 99.800 ;
        RECT 28.400 96.000 29.200 99.800 ;
        RECT 25.200 95.800 29.200 96.000 ;
        RECT 30.000 96.000 30.800 99.800 ;
        RECT 33.200 96.000 34.000 99.800 ;
        RECT 30.000 95.800 34.000 96.000 ;
        RECT 34.800 95.800 35.600 99.800 ;
        RECT 36.400 96.000 37.200 99.800 ;
        RECT 39.600 96.000 40.400 99.800 ;
        RECT 36.400 95.800 40.400 96.000 ;
        RECT 41.200 95.800 42.000 99.800 ;
        RECT 42.800 96.000 43.600 99.800 ;
        RECT 46.000 96.000 46.800 99.800 ;
        RECT 42.800 95.800 46.800 96.000 ;
        RECT 47.600 95.800 48.400 99.800 ;
        RECT 49.200 95.800 50.000 99.800 ;
        RECT 50.800 96.000 51.600 99.800 ;
        RECT 54.000 96.000 54.800 99.800 ;
        RECT 50.800 95.800 54.800 96.000 ;
        RECT 55.600 97.000 56.400 99.000 ;
        RECT 59.800 98.400 60.600 99.000 ;
        RECT 58.800 97.600 60.600 98.400 ;
        RECT 1.200 93.600 3.800 94.400 ;
        RECT 5.200 93.800 6.800 94.400 ;
        RECT 9.200 94.300 11.200 94.400 ;
        RECT 6.000 93.600 6.800 93.800 ;
        RECT 7.700 93.700 11.200 94.300 ;
        RECT 12.200 94.200 16.400 94.800 ;
        RECT 17.400 94.400 18.000 95.800 ;
        RECT 19.000 95.400 22.600 95.800 ;
        RECT 21.200 94.400 22.000 94.800 ;
        RECT 23.800 94.400 24.400 95.800 ;
        RECT 25.400 95.400 29.000 95.800 ;
        RECT 30.200 95.400 33.800 95.800 ;
        RECT 27.600 94.400 28.400 94.800 ;
        RECT 30.800 94.400 31.600 94.800 ;
        RECT 34.800 94.400 35.400 95.800 ;
        RECT 36.600 95.400 40.200 95.800 ;
        RECT 37.200 94.400 38.000 94.800 ;
        RECT 41.200 94.400 41.800 95.800 ;
        RECT 43.000 95.400 46.600 95.800 ;
        RECT 43.600 94.400 44.400 94.800 ;
        RECT 47.600 94.400 48.200 95.800 ;
        RECT 49.400 94.400 50.000 95.800 ;
        RECT 51.000 95.400 54.600 95.800 ;
        RECT 55.600 94.800 56.200 97.000 ;
        RECT 59.800 96.000 60.600 97.600 ;
        RECT 66.800 96.400 67.600 99.800 ;
        RECT 59.800 95.400 61.400 96.000 ;
        RECT 60.600 95.000 61.400 95.400 ;
        RECT 53.200 94.400 54.000 94.800 ;
        RECT 12.200 93.800 13.200 94.200 ;
        RECT 1.200 90.200 2.000 90.400 ;
        RECT 3.200 90.200 3.800 93.600 ;
        RECT 4.400 92.300 5.200 93.200 ;
        RECT 7.700 92.300 8.300 93.700 ;
        RECT 9.200 93.600 11.200 93.700 ;
        RECT 4.400 91.700 8.300 92.300 ;
        RECT 4.400 91.600 5.200 91.700 ;
        RECT 9.200 90.800 10.000 92.400 ;
        RECT 1.200 89.600 2.600 90.200 ;
        RECT 3.200 89.600 4.200 90.200 ;
        RECT 2.000 88.400 2.600 89.600 ;
        RECT 2.000 87.600 2.800 88.400 ;
        RECT 3.400 82.200 4.200 89.600 ;
        RECT 10.600 89.800 11.200 93.600 ;
        RECT 11.800 93.000 13.200 93.800 ;
        RECT 17.200 93.600 19.800 94.400 ;
        RECT 21.200 93.800 22.800 94.400 ;
        RECT 22.000 93.600 22.800 93.800 ;
        RECT 23.600 93.600 26.200 94.400 ;
        RECT 27.600 94.300 29.200 94.400 ;
        RECT 30.000 94.300 31.600 94.400 ;
        RECT 27.600 93.800 31.600 94.300 ;
        RECT 28.400 93.700 30.800 93.800 ;
        RECT 28.400 93.600 29.200 93.700 ;
        RECT 30.000 93.600 30.800 93.700 ;
        RECT 33.000 93.600 35.600 94.400 ;
        RECT 36.400 93.800 38.000 94.400 ;
        RECT 36.400 93.600 37.200 93.800 ;
        RECT 39.400 93.600 42.000 94.400 ;
        RECT 42.800 93.800 44.400 94.400 ;
        RECT 42.800 93.600 43.600 93.800 ;
        RECT 45.800 93.600 48.400 94.400 ;
        RECT 49.200 93.600 51.800 94.400 ;
        RECT 53.200 93.800 54.800 94.400 ;
        RECT 55.600 94.200 59.800 94.800 ;
        RECT 54.000 93.600 54.800 93.800 ;
        RECT 58.800 93.800 59.800 94.200 ;
        RECT 60.800 94.400 61.400 95.000 ;
        RECT 66.600 95.800 67.600 96.400 ;
        RECT 66.600 94.400 67.200 95.800 ;
        RECT 70.000 95.200 70.800 99.800 ;
        RECT 68.200 94.600 70.800 95.200 ;
        RECT 71.600 95.400 72.400 99.800 ;
        RECT 75.800 98.400 77.000 99.800 ;
        RECT 75.800 97.800 77.200 98.400 ;
        RECT 80.400 97.800 81.200 99.800 ;
        RECT 84.800 98.400 85.600 99.800 ;
        RECT 84.800 97.800 86.800 98.400 ;
        RECT 76.400 97.000 77.200 97.800 ;
        RECT 80.600 97.200 81.200 97.800 ;
        RECT 80.600 96.600 83.400 97.200 ;
        RECT 82.600 96.400 83.400 96.600 ;
        RECT 84.400 96.400 85.200 97.200 ;
        RECT 86.000 97.000 86.800 97.800 ;
        RECT 74.600 95.400 75.400 95.600 ;
        RECT 71.600 94.800 75.400 95.400 ;
        RECT 12.600 91.000 13.200 93.000 ;
        RECT 14.000 91.600 14.800 93.200 ;
        RECT 15.600 91.600 16.400 93.200 ;
        RECT 17.200 92.300 18.000 92.400 ;
        RECT 19.200 92.300 19.800 93.600 ;
        RECT 17.200 91.700 19.800 92.300 ;
        RECT 17.200 91.600 18.000 91.700 ;
        RECT 12.600 90.400 16.400 91.000 ;
        RECT 10.600 89.200 12.200 89.800 ;
        RECT 11.400 82.200 12.200 89.200 ;
        RECT 15.800 87.000 16.400 90.400 ;
        RECT 17.200 90.200 18.000 90.400 ;
        RECT 19.200 90.200 19.800 91.700 ;
        RECT 20.400 91.600 21.200 93.200 ;
        RECT 23.600 90.200 24.400 90.400 ;
        RECT 25.600 90.200 26.200 93.600 ;
        RECT 26.800 91.600 27.600 93.200 ;
        RECT 31.600 91.600 32.400 93.200 ;
        RECT 33.000 90.200 33.600 93.600 ;
        RECT 38.000 91.600 38.800 93.200 ;
        RECT 34.800 90.200 35.600 90.400 ;
        RECT 39.400 90.200 40.000 93.600 ;
        RECT 41.200 92.300 42.000 92.400 ;
        RECT 44.400 92.300 45.200 93.200 ;
        RECT 41.200 91.700 45.200 92.300 ;
        RECT 41.200 91.600 42.000 91.700 ;
        RECT 44.400 91.600 45.200 91.700 ;
        RECT 45.800 92.300 46.400 93.600 ;
        RECT 45.800 91.700 49.900 92.300 ;
        RECT 41.200 90.200 42.000 90.400 ;
        RECT 45.800 90.200 46.400 91.700 ;
        RECT 49.300 90.400 49.900 91.700 ;
        RECT 47.600 90.200 48.400 90.400 ;
        RECT 17.200 89.600 18.600 90.200 ;
        RECT 19.200 89.600 20.200 90.200 ;
        RECT 23.600 89.600 25.000 90.200 ;
        RECT 25.600 89.600 26.600 90.200 ;
        RECT 18.000 88.400 18.600 89.600 ;
        RECT 18.000 87.600 18.800 88.400 ;
        RECT 15.600 83.000 16.400 87.000 ;
        RECT 19.400 82.200 20.200 89.600 ;
        RECT 24.400 88.400 25.000 89.600 ;
        RECT 24.400 87.600 25.200 88.400 ;
        RECT 25.800 86.400 26.600 89.600 ;
        RECT 32.600 89.600 33.600 90.200 ;
        RECT 34.200 89.600 35.600 90.200 ;
        RECT 39.000 89.600 40.000 90.200 ;
        RECT 40.600 89.600 42.000 90.200 ;
        RECT 45.400 89.600 46.400 90.200 ;
        RECT 47.000 89.600 48.400 90.200 ;
        RECT 49.200 90.200 50.000 90.400 ;
        RECT 51.200 90.200 51.800 93.600 ;
        RECT 52.400 91.600 53.200 93.200 ;
        RECT 54.000 92.300 54.800 92.400 ;
        RECT 55.600 92.300 56.400 93.200 ;
        RECT 54.000 91.700 56.400 92.300 ;
        RECT 54.000 91.600 54.800 91.700 ;
        RECT 55.600 91.600 56.400 91.700 ;
        RECT 57.200 91.600 58.000 93.200 ;
        RECT 58.800 93.000 60.200 93.800 ;
        RECT 60.800 93.600 62.800 94.400 ;
        RECT 63.600 94.300 64.400 94.400 ;
        RECT 66.600 94.300 67.600 94.400 ;
        RECT 63.600 93.700 67.600 94.300 ;
        RECT 63.600 93.600 64.400 93.700 ;
        RECT 66.600 93.600 67.600 93.700 ;
        RECT 58.800 91.000 59.400 93.000 ;
        RECT 55.600 90.400 59.400 91.000 ;
        RECT 49.200 89.600 50.600 90.200 ;
        RECT 51.200 89.600 52.200 90.200 ;
        RECT 25.800 85.600 27.600 86.400 ;
        RECT 25.800 82.200 26.600 85.600 ;
        RECT 32.600 82.200 33.400 89.600 ;
        RECT 34.200 88.400 34.800 89.600 ;
        RECT 34.000 87.600 34.800 88.400 ;
        RECT 39.000 84.400 39.800 89.600 ;
        RECT 40.600 88.400 41.200 89.600 ;
        RECT 40.400 87.600 41.200 88.400 ;
        RECT 38.000 83.600 39.800 84.400 ;
        RECT 39.000 82.200 39.800 83.600 ;
        RECT 45.400 82.200 46.200 89.600 ;
        RECT 47.000 88.400 47.600 89.600 ;
        RECT 46.800 87.600 47.600 88.400 ;
        RECT 50.000 88.400 50.600 89.600 ;
        RECT 51.400 88.400 52.200 89.600 ;
        RECT 50.000 87.600 50.800 88.400 ;
        RECT 51.400 87.600 53.200 88.400 ;
        RECT 51.400 82.200 52.200 87.600 ;
        RECT 55.600 87.000 56.200 90.400 ;
        RECT 60.800 89.800 61.400 93.600 ;
        RECT 62.000 92.300 62.800 92.400 ;
        RECT 65.200 92.300 66.000 92.400 ;
        RECT 62.000 91.700 66.000 92.300 ;
        RECT 62.000 90.800 62.800 91.700 ;
        RECT 65.200 91.600 66.000 91.700 ;
        RECT 59.800 89.200 61.400 89.800 ;
        RECT 66.600 90.200 67.200 93.600 ;
        RECT 68.200 93.000 68.800 94.600 ;
        RECT 67.800 92.200 68.800 93.000 ;
        RECT 68.200 90.200 68.800 92.200 ;
        RECT 69.800 92.400 70.600 93.200 ;
        RECT 69.800 91.600 70.800 92.400 ;
        RECT 71.600 91.400 72.400 94.800 ;
        RECT 78.600 94.200 79.400 94.400 ;
        RECT 84.400 94.200 85.000 96.400 ;
        RECT 89.200 95.000 90.000 99.800 ;
        RECT 90.800 95.600 91.600 97.200 ;
        RECT 87.600 94.200 89.200 94.400 ;
        RECT 78.200 93.600 89.200 94.200 ;
        RECT 76.400 92.800 77.200 93.000 ;
        RECT 73.400 92.200 77.200 92.800 ;
        RECT 73.400 92.000 74.200 92.200 ;
        RECT 75.000 91.400 75.800 91.600 ;
        RECT 71.600 90.800 75.800 91.400 ;
        RECT 66.600 89.200 67.600 90.200 ;
        RECT 68.200 89.600 70.800 90.200 ;
        RECT 55.600 83.000 56.400 87.000 ;
        RECT 59.800 82.200 60.600 89.200 ;
        RECT 66.800 82.200 67.600 89.200 ;
        RECT 70.000 82.200 70.800 89.600 ;
        RECT 71.600 82.200 72.400 90.800 ;
        RECT 78.200 90.400 78.800 93.600 ;
        RECT 85.400 93.400 86.200 93.600 ;
        RECT 87.000 92.400 87.800 92.600 ;
        RECT 82.800 91.800 87.800 92.400 ;
        RECT 82.800 91.600 83.600 91.800 ;
        RECT 84.400 91.000 90.000 91.200 ;
        RECT 84.200 90.800 90.000 91.000 ;
        RECT 76.400 89.800 78.800 90.400 ;
        RECT 80.200 90.600 90.000 90.800 ;
        RECT 80.200 90.200 85.000 90.600 ;
        RECT 76.400 88.800 77.000 89.800 ;
        RECT 75.600 88.000 77.000 88.800 ;
        RECT 78.600 89.000 79.400 89.200 ;
        RECT 80.200 89.000 80.800 90.200 ;
        RECT 78.600 88.400 80.800 89.000 ;
        RECT 81.400 89.000 86.800 89.600 ;
        RECT 81.400 88.800 82.200 89.000 ;
        RECT 86.000 88.800 86.800 89.000 ;
        RECT 79.800 87.400 80.600 87.600 ;
        RECT 82.600 87.400 83.400 87.600 ;
        RECT 76.400 86.200 77.200 87.000 ;
        RECT 79.800 86.800 83.400 87.400 ;
        RECT 80.600 86.200 81.200 86.800 ;
        RECT 86.000 86.200 86.800 87.000 ;
        RECT 75.800 82.200 77.000 86.200 ;
        RECT 80.400 82.200 81.200 86.200 ;
        RECT 84.800 85.600 86.800 86.200 ;
        RECT 84.800 82.200 85.600 85.600 ;
        RECT 89.200 82.200 90.000 90.600 ;
        RECT 92.400 82.200 93.200 99.800 ;
        RECT 94.000 95.200 94.800 99.800 ;
        RECT 97.200 96.400 98.000 99.800 ;
        RECT 97.200 95.800 98.200 96.400 ;
        RECT 94.000 94.600 96.600 95.200 ;
        RECT 94.200 92.400 95.000 93.200 ;
        RECT 94.000 91.600 95.000 92.400 ;
        RECT 96.000 93.000 96.600 94.600 ;
        RECT 97.600 94.400 98.200 95.800 ;
        RECT 97.200 93.600 98.200 94.400 ;
        RECT 104.000 94.200 104.800 99.800 ;
        RECT 106.800 95.800 107.600 99.800 ;
        RECT 108.400 96.000 109.200 99.800 ;
        RECT 111.600 96.000 112.400 99.800 ;
        RECT 108.400 95.800 112.400 96.000 ;
        RECT 107.000 94.400 107.600 95.800 ;
        RECT 108.600 95.400 112.200 95.800 ;
        RECT 118.000 95.200 118.800 99.800 ;
        RECT 121.200 96.400 122.000 99.800 ;
        RECT 121.200 95.800 122.200 96.400 ;
        RECT 128.200 96.000 129.000 99.000 ;
        RECT 132.400 97.000 133.200 99.000 ;
        RECT 110.800 94.400 111.600 94.800 ;
        RECT 118.000 94.600 120.600 95.200 ;
        RECT 104.000 93.800 105.800 94.200 ;
        RECT 104.200 93.600 105.800 93.800 ;
        RECT 106.800 93.600 109.400 94.400 ;
        RECT 110.800 93.800 112.400 94.400 ;
        RECT 111.600 93.600 112.400 93.800 ;
        RECT 96.000 92.200 97.000 93.000 ;
        RECT 96.000 90.200 96.600 92.200 ;
        RECT 97.600 90.200 98.200 93.600 ;
        RECT 102.000 91.600 103.600 92.400 ;
        RECT 94.000 89.600 96.600 90.200 ;
        RECT 94.000 82.200 94.800 89.600 ;
        RECT 97.200 89.200 98.200 90.200 ;
        RECT 100.400 89.600 101.200 91.200 ;
        RECT 105.200 90.400 105.800 93.600 ;
        RECT 105.200 90.300 106.000 90.400 ;
        RECT 106.800 90.300 107.600 90.400 ;
        RECT 105.200 90.200 107.600 90.300 ;
        RECT 108.800 90.200 109.400 93.600 ;
        RECT 110.000 91.600 110.800 93.200 ;
        RECT 118.200 92.400 119.000 93.200 ;
        RECT 118.000 91.600 119.000 92.400 ;
        RECT 120.000 93.000 120.600 94.600 ;
        RECT 121.600 94.400 122.200 95.800 ;
        RECT 127.400 95.400 129.000 96.000 ;
        RECT 127.400 95.000 128.200 95.400 ;
        RECT 127.400 94.400 128.000 95.000 ;
        RECT 132.600 94.800 133.200 97.000 ;
        RECT 134.000 96.000 134.800 99.800 ;
        RECT 137.200 96.000 138.000 99.800 ;
        RECT 134.000 95.800 138.000 96.000 ;
        RECT 138.800 95.800 139.600 99.800 ;
        RECT 140.400 95.800 141.200 99.800 ;
        RECT 142.000 96.000 142.800 99.800 ;
        RECT 145.200 96.000 146.000 99.800 ;
        RECT 142.000 95.800 146.000 96.000 ;
        RECT 148.400 97.600 149.200 99.800 ;
        RECT 134.200 95.400 137.800 95.800 ;
        RECT 121.200 93.600 122.200 94.400 ;
        RECT 126.000 93.600 128.000 94.400 ;
        RECT 129.000 94.200 133.200 94.800 ;
        RECT 134.800 94.400 135.600 94.800 ;
        RECT 138.800 94.400 139.400 95.800 ;
        RECT 140.600 94.400 141.200 95.800 ;
        RECT 142.200 95.400 145.800 95.800 ;
        RECT 144.400 94.400 145.200 94.800 ;
        RECT 148.400 94.400 149.000 97.600 ;
        RECT 150.000 95.600 150.800 97.200 ;
        RECT 151.600 95.000 152.400 99.800 ;
        RECT 156.000 98.400 156.800 99.800 ;
        RECT 154.800 97.800 156.800 98.400 ;
        RECT 160.400 97.800 161.200 99.800 ;
        RECT 164.600 98.400 165.800 99.800 ;
        RECT 164.400 97.800 165.800 98.400 ;
        RECT 154.800 97.000 155.600 97.800 ;
        RECT 160.400 97.200 161.000 97.800 ;
        RECT 156.400 96.400 157.200 97.200 ;
        RECT 158.200 96.600 161.000 97.200 ;
        RECT 164.400 97.000 165.200 97.800 ;
        RECT 158.200 96.400 159.000 96.600 ;
        RECT 129.000 93.800 130.000 94.200 ;
        RECT 120.000 92.200 121.000 93.000 ;
        RECT 120.000 90.200 120.600 92.200 ;
        RECT 121.600 90.200 122.200 93.600 ;
        RECT 126.000 90.800 126.800 92.400 ;
        RECT 105.200 89.700 108.200 90.200 ;
        RECT 105.200 89.600 106.000 89.700 ;
        RECT 106.800 89.600 108.200 89.700 ;
        RECT 108.800 89.600 109.800 90.200 ;
        RECT 97.200 82.200 98.000 89.200 ;
        RECT 103.600 87.600 104.400 89.200 ;
        RECT 105.200 87.000 105.800 89.600 ;
        RECT 107.600 88.400 108.200 89.600 ;
        RECT 107.600 87.600 108.400 88.400 ;
        RECT 102.200 86.400 105.800 87.000 ;
        RECT 102.200 86.200 102.800 86.400 ;
        RECT 102.000 82.200 102.800 86.200 ;
        RECT 105.200 86.200 105.800 86.400 ;
        RECT 105.200 82.200 106.000 86.200 ;
        RECT 109.000 84.400 109.800 89.600 ;
        RECT 118.000 89.600 120.600 90.200 ;
        RECT 109.000 83.600 110.800 84.400 ;
        RECT 109.000 82.200 109.800 83.600 ;
        RECT 118.000 82.200 118.800 89.600 ;
        RECT 121.200 89.200 122.200 90.200 ;
        RECT 127.400 89.800 128.000 93.600 ;
        RECT 128.600 93.000 130.000 93.800 ;
        RECT 134.000 93.800 135.600 94.400 ;
        RECT 134.000 93.600 134.800 93.800 ;
        RECT 137.000 93.600 139.600 94.400 ;
        RECT 140.400 93.600 143.000 94.400 ;
        RECT 144.400 93.800 146.000 94.400 ;
        RECT 145.200 93.600 146.000 93.800 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 152.400 94.200 154.000 94.400 ;
        RECT 156.600 94.200 157.200 96.400 ;
        RECT 166.200 95.400 167.000 95.600 ;
        RECT 169.200 95.400 170.000 99.800 ;
        RECT 173.400 98.400 174.200 99.800 ;
        RECT 173.400 97.600 174.800 98.400 ;
        RECT 173.400 96.400 174.200 97.600 ;
        RECT 166.200 94.800 170.000 95.400 ;
        RECT 172.400 95.800 174.200 96.400 ;
        RECT 177.200 96.000 178.000 99.800 ;
        RECT 162.200 94.200 163.000 94.400 ;
        RECT 169.200 94.300 170.000 94.800 ;
        RECT 170.800 94.300 171.600 95.200 ;
        RECT 152.400 93.600 163.400 94.200 ;
        RECT 129.400 91.000 130.000 93.000 ;
        RECT 130.800 91.600 131.600 93.200 ;
        RECT 132.400 91.600 133.200 93.200 ;
        RECT 134.000 92.300 134.800 92.400 ;
        RECT 135.600 92.300 136.400 93.200 ;
        RECT 134.000 91.700 136.400 92.300 ;
        RECT 134.000 91.600 134.800 91.700 ;
        RECT 135.600 91.600 136.400 91.700 ;
        RECT 137.000 92.300 137.600 93.600 ;
        RECT 137.000 91.700 141.100 92.300 ;
        RECT 129.400 90.400 133.200 91.000 ;
        RECT 127.400 89.200 129.000 89.800 ;
        RECT 121.200 82.200 122.000 89.200 ;
        RECT 128.200 84.400 129.000 89.200 ;
        RECT 132.600 87.000 133.200 90.400 ;
        RECT 137.000 90.200 137.600 91.700 ;
        RECT 140.500 90.400 141.100 91.700 ;
        RECT 142.400 90.400 143.000 93.600 ;
        RECT 143.600 91.600 144.400 93.200 ;
        RECT 146.800 92.300 147.600 92.400 ;
        RECT 145.300 91.700 147.600 92.300 ;
        RECT 146.800 90.800 147.600 91.700 ;
        RECT 138.800 90.200 139.600 90.400 ;
        RECT 128.200 83.600 130.000 84.400 ;
        RECT 128.200 82.200 129.000 83.600 ;
        RECT 132.400 83.000 133.200 87.000 ;
        RECT 136.600 89.600 137.600 90.200 ;
        RECT 138.200 89.600 139.600 90.200 ;
        RECT 140.400 90.200 141.200 90.400 ;
        RECT 140.400 89.600 141.800 90.200 ;
        RECT 142.400 89.600 144.400 90.400 ;
        RECT 148.400 90.200 149.000 93.600 ;
        RECT 155.400 93.400 156.200 93.600 ;
        RECT 153.800 92.400 154.600 92.600 ;
        RECT 156.400 92.400 157.200 92.600 ;
        RECT 162.800 92.400 163.400 93.600 ;
        RECT 169.200 93.700 171.600 94.300 ;
        RECT 164.400 92.800 165.200 93.000 ;
        RECT 153.800 91.800 158.800 92.400 ;
        RECT 158.000 91.600 158.800 91.800 ;
        RECT 162.800 91.600 163.600 92.400 ;
        RECT 164.400 92.200 168.200 92.800 ;
        RECT 167.400 92.000 168.200 92.200 ;
        RECT 151.600 91.000 157.200 91.200 ;
        RECT 151.600 90.800 157.400 91.000 ;
        RECT 151.600 90.600 161.400 90.800 ;
        RECT 136.600 82.200 137.400 89.600 ;
        RECT 138.200 88.400 138.800 89.600 ;
        RECT 138.000 87.600 138.800 88.400 ;
        RECT 141.200 88.400 141.800 89.600 ;
        RECT 141.200 87.600 142.000 88.400 ;
        RECT 142.600 82.200 143.400 89.600 ;
        RECT 147.400 89.400 149.200 90.200 ;
        RECT 147.400 88.400 148.200 89.400 ;
        RECT 147.400 87.600 149.200 88.400 ;
        RECT 147.400 82.200 148.200 87.600 ;
        RECT 151.600 82.200 152.400 90.600 ;
        RECT 156.600 90.200 161.400 90.600 ;
        RECT 154.800 89.000 160.200 89.600 ;
        RECT 154.800 88.800 155.600 89.000 ;
        RECT 159.400 88.800 160.200 89.000 ;
        RECT 160.800 89.000 161.400 90.200 ;
        RECT 162.800 90.400 163.400 91.600 ;
        RECT 165.800 91.400 166.600 91.600 ;
        RECT 169.200 91.400 170.000 93.700 ;
        RECT 170.800 93.600 171.600 93.700 ;
        RECT 165.800 90.800 170.000 91.400 ;
        RECT 162.800 89.800 165.200 90.400 ;
        RECT 162.200 89.000 163.000 89.200 ;
        RECT 160.800 88.400 163.000 89.000 ;
        RECT 164.600 88.800 165.200 89.800 ;
        RECT 164.600 88.000 166.000 88.800 ;
        RECT 158.200 87.400 159.000 87.600 ;
        RECT 161.000 87.400 161.800 87.600 ;
        RECT 154.800 86.200 155.600 87.000 ;
        RECT 158.200 86.800 161.800 87.400 ;
        RECT 160.400 86.200 161.000 86.800 ;
        RECT 164.400 86.200 165.200 87.000 ;
        RECT 154.800 85.600 156.800 86.200 ;
        RECT 156.000 82.200 156.800 85.600 ;
        RECT 160.400 82.200 161.200 86.200 ;
        RECT 164.600 82.200 165.800 86.200 ;
        RECT 169.200 82.200 170.000 90.800 ;
        RECT 172.400 82.200 173.200 95.800 ;
        RECT 177.000 95.200 178.000 96.000 ;
        RECT 177.000 90.800 177.800 95.200 ;
        RECT 178.800 94.600 179.600 99.800 ;
        RECT 185.200 96.600 186.000 99.800 ;
        RECT 186.800 97.000 187.600 99.800 ;
        RECT 188.400 97.000 189.200 99.800 ;
        RECT 190.000 97.000 190.800 99.800 ;
        RECT 191.600 97.000 192.400 99.800 ;
        RECT 194.800 97.000 195.600 99.800 ;
        RECT 198.000 97.000 198.800 99.800 ;
        RECT 199.600 97.000 200.400 99.800 ;
        RECT 201.200 97.000 202.000 99.800 ;
        RECT 183.600 95.800 186.000 96.600 ;
        RECT 202.800 96.600 203.600 99.800 ;
        RECT 183.600 95.200 184.400 95.800 ;
        RECT 178.400 94.000 179.600 94.600 ;
        RECT 182.600 94.600 184.400 95.200 ;
        RECT 188.400 95.600 189.400 96.400 ;
        RECT 192.400 95.600 194.000 96.400 ;
        RECT 194.800 95.800 199.400 96.400 ;
        RECT 202.800 95.800 205.400 96.600 ;
        RECT 194.800 95.600 195.600 95.800 ;
        RECT 178.400 92.000 179.000 94.000 ;
        RECT 182.600 93.400 183.400 94.600 ;
        RECT 179.600 92.600 183.400 93.400 ;
        RECT 188.400 92.800 189.200 95.600 ;
        RECT 194.800 94.800 195.600 95.000 ;
        RECT 191.200 94.200 195.600 94.800 ;
        RECT 191.200 94.000 192.000 94.200 ;
        RECT 196.400 93.600 197.200 95.200 ;
        RECT 198.600 93.400 199.400 95.800 ;
        RECT 204.600 95.200 205.400 95.800 ;
        RECT 204.600 94.400 207.600 95.200 ;
        RECT 209.200 93.800 210.000 99.800 ;
        RECT 213.400 98.400 214.200 99.800 ;
        RECT 213.400 97.600 214.800 98.400 ;
        RECT 213.400 96.400 214.200 97.600 ;
        RECT 212.400 95.800 214.200 96.400 ;
        RECT 215.600 96.000 216.400 99.800 ;
        RECT 218.800 96.000 219.600 99.800 ;
        RECT 215.600 95.800 219.600 96.000 ;
        RECT 220.400 96.300 221.200 99.800 ;
        RECT 222.000 96.300 222.800 97.200 ;
        RECT 191.600 92.600 194.800 93.400 ;
        RECT 198.600 92.600 200.600 93.400 ;
        RECT 201.200 93.000 210.000 93.800 ;
        RECT 210.800 93.600 211.600 95.200 ;
        RECT 185.200 92.000 186.000 92.600 ;
        RECT 202.800 92.000 203.600 92.400 ;
        RECT 206.000 92.000 206.800 92.400 ;
        RECT 207.800 92.000 208.600 92.200 ;
        RECT 178.400 91.400 179.200 92.000 ;
        RECT 185.200 91.400 208.600 92.000 ;
        RECT 174.000 88.800 174.800 90.400 ;
        RECT 177.000 90.000 178.000 90.800 ;
        RECT 177.200 82.200 178.000 90.000 ;
        RECT 178.600 89.600 179.200 91.400 ;
        RECT 178.600 89.000 187.600 89.600 ;
        RECT 178.600 87.400 179.200 89.000 ;
        RECT 186.800 88.800 187.600 89.000 ;
        RECT 190.000 89.000 198.600 89.600 ;
        RECT 190.000 88.800 190.800 89.000 ;
        RECT 181.800 87.600 184.400 88.400 ;
        RECT 178.600 86.800 181.200 87.400 ;
        RECT 180.400 82.200 181.200 86.800 ;
        RECT 183.600 82.200 184.400 87.600 ;
        RECT 185.000 86.800 189.200 87.600 ;
        RECT 186.800 82.200 187.600 85.000 ;
        RECT 188.400 82.200 189.200 85.000 ;
        RECT 190.000 82.200 190.800 85.000 ;
        RECT 191.600 82.200 192.400 88.400 ;
        RECT 194.800 87.600 197.400 88.400 ;
        RECT 198.000 88.200 198.600 89.000 ;
        RECT 199.600 89.400 200.400 89.600 ;
        RECT 199.600 89.000 205.000 89.400 ;
        RECT 199.600 88.800 205.800 89.000 ;
        RECT 204.400 88.200 205.800 88.800 ;
        RECT 198.000 87.600 203.800 88.200 ;
        RECT 206.800 88.000 208.400 88.800 ;
        RECT 206.800 87.600 207.400 88.000 ;
        RECT 194.800 82.200 195.600 87.000 ;
        RECT 198.000 82.200 198.800 87.000 ;
        RECT 203.200 86.800 207.400 87.600 ;
        RECT 209.200 87.400 210.000 93.000 ;
        RECT 208.000 86.800 210.000 87.400 ;
        RECT 199.600 82.200 200.400 85.000 ;
        RECT 201.200 82.200 202.000 85.000 ;
        RECT 204.400 82.200 205.200 86.800 ;
        RECT 208.000 86.200 208.600 86.800 ;
        RECT 207.600 85.600 208.600 86.200 ;
        RECT 207.600 82.200 208.400 85.600 ;
        RECT 212.400 82.200 213.200 95.800 ;
        RECT 215.800 95.400 219.400 95.800 ;
        RECT 220.400 95.700 222.800 96.300 ;
        RECT 216.400 94.400 217.200 94.800 ;
        RECT 220.400 94.400 221.000 95.700 ;
        RECT 222.000 95.600 222.800 95.700 ;
        RECT 214.000 94.300 214.800 94.400 ;
        RECT 215.600 94.300 217.200 94.400 ;
        RECT 214.000 93.800 217.200 94.300 ;
        RECT 214.000 93.700 216.400 93.800 ;
        RECT 214.000 93.600 214.800 93.700 ;
        RECT 215.600 93.600 216.400 93.700 ;
        RECT 218.600 93.600 221.200 94.400 ;
        RECT 217.200 92.300 218.000 93.200 ;
        RECT 214.100 91.700 218.000 92.300 ;
        RECT 214.100 90.400 214.700 91.700 ;
        RECT 217.200 91.600 218.000 91.700 ;
        RECT 214.000 88.800 214.800 90.400 ;
        RECT 218.600 90.200 219.200 93.600 ;
        RECT 220.400 90.200 221.200 90.400 ;
        RECT 218.200 89.600 219.200 90.200 ;
        RECT 219.800 89.600 221.200 90.200 ;
        RECT 218.200 82.200 219.000 89.600 ;
        RECT 219.800 88.400 220.400 89.600 ;
        RECT 219.600 87.600 220.400 88.400 ;
        RECT 223.600 82.200 224.400 99.800 ;
        RECT 225.200 95.800 226.000 99.800 ;
        RECT 229.400 98.400 230.200 99.800 ;
        RECT 229.400 97.600 230.800 98.400 ;
        RECT 229.400 96.800 230.200 97.600 ;
        RECT 229.400 95.800 230.800 96.800 ;
        RECT 225.400 95.600 226.000 95.800 ;
        RECT 225.400 95.200 227.200 95.600 ;
        RECT 225.400 95.000 229.600 95.200 ;
        RECT 226.600 94.600 229.600 95.000 ;
        RECT 228.800 94.400 229.600 94.600 ;
        RECT 225.200 92.800 226.000 94.400 ;
        RECT 227.200 93.800 228.000 94.000 ;
        RECT 227.000 93.200 228.000 93.800 ;
        RECT 227.000 92.400 227.600 93.200 ;
        RECT 226.800 91.600 227.600 92.400 ;
        RECT 228.800 91.000 229.400 94.400 ;
        RECT 230.200 92.400 230.800 95.800 ;
        RECT 231.600 95.800 232.400 99.800 ;
        RECT 236.000 96.200 237.600 99.800 ;
        RECT 231.600 95.200 234.000 95.800 ;
        RECT 233.200 95.000 234.000 95.200 ;
        RECT 234.600 94.800 235.400 95.600 ;
        RECT 234.600 94.400 235.200 94.800 ;
        RECT 231.600 93.600 233.200 94.400 ;
        RECT 234.400 93.600 235.200 94.400 ;
        RECT 236.000 94.200 236.600 96.200 ;
        RECT 241.200 95.800 242.000 99.800 ;
        RECT 242.800 95.800 243.600 99.800 ;
        RECT 244.400 96.000 245.200 99.800 ;
        RECT 247.600 96.000 248.400 99.800 ;
        RECT 255.600 96.000 256.400 99.800 ;
        RECT 244.400 95.800 248.400 96.000 ;
        RECT 237.200 94.800 238.800 95.600 ;
        RECT 239.400 95.200 242.000 95.800 ;
        RECT 239.400 95.000 240.200 95.200 ;
        RECT 243.000 94.400 243.600 95.800 ;
        RECT 244.600 95.400 248.200 95.800 ;
        RECT 255.400 95.200 256.400 96.000 ;
        RECT 246.800 94.400 247.600 94.800 ;
        RECT 240.400 94.300 242.000 94.400 ;
        RECT 242.800 94.300 245.400 94.400 ;
        RECT 240.400 94.200 245.400 94.300 ;
        RECT 236.000 93.600 237.000 94.200 ;
        RECT 239.800 94.000 245.400 94.200 ;
        RECT 230.000 91.600 230.800 92.400 ;
        RECT 227.000 90.400 229.400 91.000 ;
        RECT 227.000 86.200 227.600 90.400 ;
        RECT 230.200 90.200 230.800 91.600 ;
        RECT 236.400 92.400 237.000 93.600 ;
        RECT 237.600 93.700 245.400 94.000 ;
        RECT 246.800 94.300 248.400 94.400 ;
        RECT 250.800 94.300 251.600 94.400 ;
        RECT 246.800 93.800 251.600 94.300 ;
        RECT 237.600 93.600 242.000 93.700 ;
        RECT 242.800 93.600 245.400 93.700 ;
        RECT 247.600 93.700 251.600 93.800 ;
        RECT 247.600 93.600 248.400 93.700 ;
        RECT 250.800 93.600 251.600 93.700 ;
        RECT 237.600 93.400 240.400 93.600 ;
        RECT 237.600 93.200 238.400 93.400 ;
        RECT 236.400 91.600 237.200 92.400 ;
        RECT 239.000 92.200 239.800 92.400 ;
        RECT 238.200 91.600 239.800 92.200 ;
        RECT 236.400 90.200 237.000 91.600 ;
        RECT 238.200 91.400 239.000 91.600 ;
        RECT 242.800 90.200 243.600 90.400 ;
        RECT 244.800 90.200 245.400 93.600 ;
        RECT 246.000 92.300 246.800 93.200 ;
        RECT 252.400 92.300 253.200 92.400 ;
        RECT 246.000 91.700 253.200 92.300 ;
        RECT 246.000 91.600 246.800 91.700 ;
        RECT 252.400 91.600 253.200 91.700 ;
        RECT 255.400 90.800 256.200 95.200 ;
        RECT 257.200 94.600 258.000 99.800 ;
        RECT 263.600 96.600 264.400 99.800 ;
        RECT 265.200 97.000 266.000 99.800 ;
        RECT 266.800 97.000 267.600 99.800 ;
        RECT 268.400 97.000 269.200 99.800 ;
        RECT 270.000 97.000 270.800 99.800 ;
        RECT 273.200 97.000 274.000 99.800 ;
        RECT 276.400 97.000 277.200 99.800 ;
        RECT 278.000 97.000 278.800 99.800 ;
        RECT 279.600 97.000 280.400 99.800 ;
        RECT 262.000 95.800 264.400 96.600 ;
        RECT 281.200 96.600 282.000 99.800 ;
        RECT 262.000 95.200 262.800 95.800 ;
        RECT 256.800 94.000 258.000 94.600 ;
        RECT 261.000 94.600 262.800 95.200 ;
        RECT 266.800 95.600 267.800 96.400 ;
        RECT 270.800 95.600 272.400 96.400 ;
        RECT 273.200 95.800 277.800 96.400 ;
        RECT 281.200 95.800 283.800 96.600 ;
        RECT 273.200 95.600 274.000 95.800 ;
        RECT 256.800 92.000 257.400 94.000 ;
        RECT 261.000 93.400 261.800 94.600 ;
        RECT 258.000 92.600 261.800 93.400 ;
        RECT 266.800 92.800 267.600 95.600 ;
        RECT 273.200 94.800 274.000 95.000 ;
        RECT 269.600 94.200 274.000 94.800 ;
        RECT 269.600 94.000 270.400 94.200 ;
        RECT 274.800 93.600 275.600 95.200 ;
        RECT 277.000 93.400 277.800 95.800 ;
        RECT 283.000 95.200 283.800 95.800 ;
        RECT 283.000 94.400 286.000 95.200 ;
        RECT 287.600 93.800 288.400 99.800 ;
        RECT 289.200 95.200 290.000 99.800 ;
        RECT 292.400 96.400 293.200 99.800 ;
        RECT 292.400 95.800 293.400 96.400 ;
        RECT 295.600 96.000 296.400 99.800 ;
        RECT 298.800 96.000 299.600 99.800 ;
        RECT 295.600 95.800 299.600 96.000 ;
        RECT 300.400 95.800 301.200 99.800 ;
        RECT 304.600 96.400 305.400 99.800 ;
        RECT 303.600 95.800 305.400 96.400 ;
        RECT 308.400 96.000 309.200 99.800 ;
        RECT 289.200 94.600 291.800 95.200 ;
        RECT 270.000 92.600 273.200 93.400 ;
        RECT 277.000 92.600 279.000 93.400 ;
        RECT 279.600 93.000 288.400 93.800 ;
        RECT 263.600 92.000 264.400 92.600 ;
        RECT 281.200 92.000 282.000 92.400 ;
        RECT 286.200 92.000 287.000 92.200 ;
        RECT 256.800 91.400 257.600 92.000 ;
        RECT 263.600 91.400 287.000 92.000 ;
        RECT 226.800 82.200 227.600 86.200 ;
        RECT 230.000 82.200 230.800 90.200 ;
        RECT 231.600 89.600 234.000 90.200 ;
        RECT 231.600 82.200 232.400 89.600 ;
        RECT 233.200 89.400 234.000 89.600 ;
        RECT 236.000 84.400 237.600 90.200 ;
        RECT 239.400 89.600 242.000 90.200 ;
        RECT 242.800 89.600 244.200 90.200 ;
        RECT 244.800 89.600 245.800 90.200 ;
        RECT 255.400 90.000 256.400 90.800 ;
        RECT 239.400 89.400 240.200 89.600 ;
        RECT 236.000 83.600 238.800 84.400 ;
        RECT 236.000 82.200 237.600 83.600 ;
        RECT 241.200 82.200 242.000 89.600 ;
        RECT 243.600 88.400 244.200 89.600 ;
        RECT 243.600 87.600 244.400 88.400 ;
        RECT 245.000 82.200 245.800 89.600 ;
        RECT 255.600 82.200 256.400 90.000 ;
        RECT 257.000 89.600 257.600 91.400 ;
        RECT 257.000 89.000 266.000 89.600 ;
        RECT 257.000 87.400 257.600 89.000 ;
        RECT 265.200 88.800 266.000 89.000 ;
        RECT 268.400 89.000 277.000 89.600 ;
        RECT 268.400 88.800 269.200 89.000 ;
        RECT 260.200 87.600 262.800 88.400 ;
        RECT 257.000 86.800 259.600 87.400 ;
        RECT 258.800 82.200 259.600 86.800 ;
        RECT 262.000 82.200 262.800 87.600 ;
        RECT 263.400 86.800 267.600 87.600 ;
        RECT 265.200 82.200 266.000 85.000 ;
        RECT 266.800 82.200 267.600 85.000 ;
        RECT 268.400 82.200 269.200 85.000 ;
        RECT 270.000 82.200 270.800 88.400 ;
        RECT 273.200 87.600 275.800 88.400 ;
        RECT 276.400 88.200 277.000 89.000 ;
        RECT 278.000 89.400 278.800 89.600 ;
        RECT 278.000 89.000 283.400 89.400 ;
        RECT 278.000 88.800 284.200 89.000 ;
        RECT 282.800 88.200 284.200 88.800 ;
        RECT 276.400 87.600 282.200 88.200 ;
        RECT 285.200 88.000 286.800 88.800 ;
        RECT 285.200 87.600 285.800 88.000 ;
        RECT 273.200 82.200 274.000 87.000 ;
        RECT 276.400 82.200 277.200 87.000 ;
        RECT 281.600 86.800 285.800 87.600 ;
        RECT 287.600 87.400 288.400 93.000 ;
        RECT 289.400 92.400 290.200 93.200 ;
        RECT 289.200 91.600 290.200 92.400 ;
        RECT 291.200 93.000 291.800 94.600 ;
        RECT 292.800 94.400 293.400 95.800 ;
        RECT 295.800 95.400 299.400 95.800 ;
        RECT 296.400 94.400 297.200 94.800 ;
        RECT 300.400 94.400 301.000 95.800 ;
        RECT 292.400 93.600 293.400 94.400 ;
        RECT 295.600 93.800 297.200 94.400 ;
        RECT 298.600 94.300 301.200 94.400 ;
        RECT 302.000 94.300 302.800 95.200 ;
        RECT 295.600 93.600 296.400 93.800 ;
        RECT 298.600 93.700 302.800 94.300 ;
        RECT 298.600 93.600 301.200 93.700 ;
        RECT 302.000 93.600 302.800 93.700 ;
        RECT 303.600 94.300 304.400 95.800 ;
        RECT 308.200 95.200 309.200 96.000 ;
        RECT 305.200 94.300 306.000 94.400 ;
        RECT 303.600 93.700 306.000 94.300 ;
        RECT 291.200 92.200 292.200 93.000 ;
        RECT 291.200 90.200 291.800 92.200 ;
        RECT 292.800 90.200 293.400 93.600 ;
        RECT 297.200 91.600 298.000 93.200 ;
        RECT 298.600 90.200 299.200 93.600 ;
        RECT 300.400 90.300 301.200 90.400 ;
        RECT 302.000 90.300 302.800 90.400 ;
        RECT 300.400 90.200 302.800 90.300 ;
        RECT 286.400 86.800 288.400 87.400 ;
        RECT 289.200 89.600 291.800 90.200 ;
        RECT 278.000 82.200 278.800 85.000 ;
        RECT 279.600 82.200 280.400 85.000 ;
        RECT 282.800 82.200 283.600 86.800 ;
        RECT 286.400 86.200 287.000 86.800 ;
        RECT 286.000 85.600 287.000 86.200 ;
        RECT 286.000 82.200 286.800 85.600 ;
        RECT 289.200 82.200 290.000 89.600 ;
        RECT 292.400 89.200 293.400 90.200 ;
        RECT 298.200 89.600 299.200 90.200 ;
        RECT 299.800 89.700 302.800 90.200 ;
        RECT 299.800 89.600 301.200 89.700 ;
        RECT 302.000 89.600 302.800 89.700 ;
        RECT 292.400 82.200 293.200 89.200 ;
        RECT 298.200 82.200 299.000 89.600 ;
        RECT 299.800 88.400 300.400 89.600 ;
        RECT 299.600 87.600 300.400 88.400 ;
        RECT 303.600 82.200 304.400 93.700 ;
        RECT 305.200 93.600 306.000 93.700 ;
        RECT 308.200 90.800 309.000 95.200 ;
        RECT 310.000 94.600 310.800 99.800 ;
        RECT 316.400 96.600 317.200 99.800 ;
        RECT 318.000 97.000 318.800 99.800 ;
        RECT 319.600 97.000 320.400 99.800 ;
        RECT 321.200 97.000 322.000 99.800 ;
        RECT 322.800 97.000 323.600 99.800 ;
        RECT 326.000 97.000 326.800 99.800 ;
        RECT 329.200 97.000 330.000 99.800 ;
        RECT 330.800 97.000 331.600 99.800 ;
        RECT 332.400 97.000 333.200 99.800 ;
        RECT 314.800 95.800 317.200 96.600 ;
        RECT 334.000 96.600 334.800 99.800 ;
        RECT 314.800 95.200 315.600 95.800 ;
        RECT 309.600 94.000 310.800 94.600 ;
        RECT 313.800 94.600 315.600 95.200 ;
        RECT 319.600 95.600 320.600 96.400 ;
        RECT 323.600 95.600 325.200 96.400 ;
        RECT 326.000 95.800 330.600 96.400 ;
        RECT 334.000 95.800 336.600 96.600 ;
        RECT 326.000 95.600 326.800 95.800 ;
        RECT 309.600 92.000 310.200 94.000 ;
        RECT 313.800 93.400 314.600 94.600 ;
        RECT 310.800 92.600 314.600 93.400 ;
        RECT 319.600 92.800 320.400 95.600 ;
        RECT 326.000 94.800 326.800 95.000 ;
        RECT 322.400 94.200 326.800 94.800 ;
        RECT 322.400 94.000 323.200 94.200 ;
        RECT 327.600 93.600 328.400 95.200 ;
        RECT 329.800 93.400 330.600 95.800 ;
        RECT 335.800 95.200 336.600 95.800 ;
        RECT 335.800 94.400 338.800 95.200 ;
        RECT 340.400 93.800 341.200 99.800 ;
        RECT 342.000 95.600 342.800 97.200 ;
        RECT 322.800 92.600 326.000 93.400 ;
        RECT 329.800 92.600 331.800 93.400 ;
        RECT 332.400 93.000 341.200 93.800 ;
        RECT 316.400 92.000 317.200 92.600 ;
        RECT 334.000 92.000 334.800 92.400 ;
        RECT 337.200 92.000 338.000 92.400 ;
        RECT 339.000 92.000 339.800 92.200 ;
        RECT 309.600 91.400 310.400 92.000 ;
        RECT 316.400 91.400 339.800 92.000 ;
        RECT 305.200 88.800 306.000 90.400 ;
        RECT 308.200 90.000 309.200 90.800 ;
        RECT 308.400 82.200 309.200 90.000 ;
        RECT 309.800 89.600 310.400 91.400 ;
        RECT 309.800 89.000 318.800 89.600 ;
        RECT 309.800 87.400 310.400 89.000 ;
        RECT 318.000 88.800 318.800 89.000 ;
        RECT 321.200 89.000 329.800 89.600 ;
        RECT 321.200 88.800 322.000 89.000 ;
        RECT 313.000 87.600 315.600 88.400 ;
        RECT 309.800 86.800 312.400 87.400 ;
        RECT 311.600 82.200 312.400 86.800 ;
        RECT 314.800 82.200 315.600 87.600 ;
        RECT 316.200 86.800 320.400 87.600 ;
        RECT 318.000 82.200 318.800 85.000 ;
        RECT 319.600 82.200 320.400 85.000 ;
        RECT 321.200 82.200 322.000 85.000 ;
        RECT 322.800 82.200 323.600 88.400 ;
        RECT 326.000 87.600 328.600 88.400 ;
        RECT 329.200 88.200 329.800 89.000 ;
        RECT 330.800 89.400 331.600 89.600 ;
        RECT 330.800 89.000 336.200 89.400 ;
        RECT 330.800 88.800 337.000 89.000 ;
        RECT 335.600 88.200 337.000 88.800 ;
        RECT 329.200 87.600 335.000 88.200 ;
        RECT 338.000 88.000 339.600 88.800 ;
        RECT 338.000 87.600 338.600 88.000 ;
        RECT 326.000 82.200 326.800 87.000 ;
        RECT 329.200 82.200 330.000 87.000 ;
        RECT 334.400 86.800 338.600 87.600 ;
        RECT 340.400 87.400 341.200 93.000 ;
        RECT 339.200 86.800 341.200 87.400 ;
        RECT 330.800 82.200 331.600 85.000 ;
        RECT 332.400 82.200 333.200 85.000 ;
        RECT 335.600 82.200 336.400 86.800 ;
        RECT 339.200 86.200 339.800 86.800 ;
        RECT 338.800 85.600 339.800 86.200 ;
        RECT 338.800 82.200 339.600 85.600 ;
        RECT 343.600 82.200 344.400 99.800 ;
        RECT 345.200 93.800 346.000 99.800 ;
        RECT 351.600 96.600 352.400 99.800 ;
        RECT 353.200 97.000 354.000 99.800 ;
        RECT 354.800 97.000 355.600 99.800 ;
        RECT 356.400 97.000 357.200 99.800 ;
        RECT 359.600 97.000 360.400 99.800 ;
        RECT 362.800 97.000 363.600 99.800 ;
        RECT 364.400 97.000 365.200 99.800 ;
        RECT 366.000 97.000 366.800 99.800 ;
        RECT 367.600 97.000 368.400 99.800 ;
        RECT 349.800 95.800 352.400 96.600 ;
        RECT 369.200 96.600 370.000 99.800 ;
        RECT 355.800 95.800 360.400 96.400 ;
        RECT 349.800 95.200 350.600 95.800 ;
        RECT 347.600 94.400 350.600 95.200 ;
        RECT 345.200 93.000 354.000 93.800 ;
        RECT 355.800 93.400 356.600 95.800 ;
        RECT 359.600 95.600 360.400 95.800 ;
        RECT 361.200 95.600 362.800 96.400 ;
        RECT 365.800 95.600 366.800 96.400 ;
        RECT 369.200 95.800 371.600 96.600 ;
        RECT 358.000 93.600 358.800 95.200 ;
        RECT 359.600 94.800 360.400 95.000 ;
        RECT 359.600 94.200 364.000 94.800 ;
        RECT 363.200 94.000 364.000 94.200 ;
        RECT 345.200 87.400 346.000 93.000 ;
        RECT 354.600 92.600 356.600 93.400 ;
        RECT 360.400 92.600 363.600 93.400 ;
        RECT 366.000 92.800 366.800 95.600 ;
        RECT 370.800 95.200 371.600 95.800 ;
        RECT 370.800 94.600 372.600 95.200 ;
        RECT 371.800 93.400 372.600 94.600 ;
        RECT 375.600 94.600 376.400 99.800 ;
        RECT 377.200 96.000 378.000 99.800 ;
        RECT 380.400 96.000 381.200 99.800 ;
        RECT 383.600 96.000 384.400 99.800 ;
        RECT 377.200 95.200 378.200 96.000 ;
        RECT 380.400 95.800 384.400 96.000 ;
        RECT 385.200 95.800 386.000 99.800 ;
        RECT 389.400 96.400 390.200 99.800 ;
        RECT 380.600 95.400 384.200 95.800 ;
        RECT 375.600 94.000 376.800 94.600 ;
        RECT 371.800 92.600 375.600 93.400 ;
        RECT 346.600 92.000 347.400 92.200 ;
        RECT 351.600 92.000 352.400 92.400 ;
        RECT 369.200 92.000 370.000 92.600 ;
        RECT 376.200 92.000 376.800 94.000 ;
        RECT 346.600 91.400 370.000 92.000 ;
        RECT 376.000 91.400 376.800 92.000 ;
        RECT 376.000 89.600 376.600 91.400 ;
        RECT 377.400 90.800 378.200 95.200 ;
        RECT 381.200 94.400 382.000 94.800 ;
        RECT 385.200 94.400 385.800 95.800 ;
        RECT 388.400 95.600 390.800 96.400 ;
        RECT 391.600 96.000 392.400 99.800 ;
        RECT 394.800 96.000 395.600 99.800 ;
        RECT 391.600 95.800 395.600 96.000 ;
        RECT 396.400 95.800 397.200 99.800 ;
        RECT 400.600 96.400 401.400 99.800 ;
        RECT 399.600 95.800 401.400 96.400 ;
        RECT 409.200 96.000 410.000 99.800 ;
        RECT 380.400 93.800 382.000 94.400 ;
        RECT 383.400 94.300 386.000 94.400 ;
        RECT 386.800 94.300 387.600 95.200 ;
        RECT 380.400 93.600 381.200 93.800 ;
        RECT 383.400 93.700 387.600 94.300 ;
        RECT 383.400 93.600 386.000 93.700 ;
        RECT 386.800 93.600 387.600 93.700 ;
        RECT 382.000 91.600 382.800 93.200 ;
        RECT 354.800 89.400 355.600 89.600 ;
        RECT 350.200 89.000 355.600 89.400 ;
        RECT 349.400 88.800 355.600 89.000 ;
        RECT 356.600 89.000 365.200 89.600 ;
        RECT 346.800 88.000 348.400 88.800 ;
        RECT 349.400 88.200 350.800 88.800 ;
        RECT 356.600 88.200 357.200 89.000 ;
        RECT 364.400 88.800 365.200 89.000 ;
        RECT 367.600 89.000 376.600 89.600 ;
        RECT 367.600 88.800 368.400 89.000 ;
        RECT 347.800 87.600 348.400 88.000 ;
        RECT 351.400 87.600 357.200 88.200 ;
        RECT 357.800 87.600 360.400 88.400 ;
        RECT 345.200 86.800 347.200 87.400 ;
        RECT 347.800 86.800 352.000 87.600 ;
        RECT 346.600 86.200 347.200 86.800 ;
        RECT 346.600 85.600 347.600 86.200 ;
        RECT 346.800 82.200 347.600 85.600 ;
        RECT 350.000 82.200 350.800 86.800 ;
        RECT 353.200 82.200 354.000 85.000 ;
        RECT 354.800 82.200 355.600 85.000 ;
        RECT 356.400 82.200 357.200 87.000 ;
        RECT 359.600 82.200 360.400 87.000 ;
        RECT 362.800 82.200 363.600 88.400 ;
        RECT 370.800 87.600 373.400 88.400 ;
        RECT 366.000 86.800 370.200 87.600 ;
        RECT 364.400 82.200 365.200 85.000 ;
        RECT 366.000 82.200 366.800 85.000 ;
        RECT 367.600 82.200 368.400 85.000 ;
        RECT 370.800 82.200 371.600 87.600 ;
        RECT 376.000 87.400 376.600 89.000 ;
        RECT 374.000 86.800 376.600 87.400 ;
        RECT 377.200 90.000 378.200 90.800 ;
        RECT 383.400 90.200 384.000 93.600 ;
        RECT 385.200 90.300 386.000 90.400 ;
        RECT 386.800 90.300 387.600 90.400 ;
        RECT 385.200 90.200 387.600 90.300 ;
        RECT 374.000 82.200 374.800 86.800 ;
        RECT 377.200 82.200 378.000 90.000 ;
        RECT 383.000 89.600 384.000 90.200 ;
        RECT 384.600 89.700 387.600 90.200 ;
        RECT 384.600 89.600 386.000 89.700 ;
        RECT 386.800 89.600 387.600 89.700 ;
        RECT 383.000 82.200 383.800 89.600 ;
        RECT 384.600 88.400 385.200 89.600 ;
        RECT 384.400 87.600 385.200 88.400 ;
        RECT 388.400 82.200 389.200 95.600 ;
        RECT 391.800 95.400 395.400 95.800 ;
        RECT 392.400 94.400 393.200 94.800 ;
        RECT 396.400 94.400 397.000 95.800 ;
        RECT 391.600 93.800 393.200 94.400 ;
        RECT 394.600 94.300 397.200 94.400 ;
        RECT 398.000 94.300 398.800 95.200 ;
        RECT 391.600 93.600 392.400 93.800 ;
        RECT 394.600 93.700 398.800 94.300 ;
        RECT 394.600 93.600 397.200 93.700 ;
        RECT 398.000 93.600 398.800 93.700 ;
        RECT 393.200 91.600 394.000 93.200 ;
        RECT 390.000 88.800 390.800 90.400 ;
        RECT 394.600 90.200 395.200 93.600 ;
        RECT 396.400 90.200 397.200 90.400 ;
        RECT 394.200 89.600 395.200 90.200 ;
        RECT 395.800 89.600 397.200 90.200 ;
        RECT 394.200 82.200 395.000 89.600 ;
        RECT 395.800 88.400 396.400 89.600 ;
        RECT 395.600 88.300 396.400 88.400 ;
        RECT 398.000 88.300 398.800 88.400 ;
        RECT 395.600 87.700 398.800 88.300 ;
        RECT 395.600 87.600 396.400 87.700 ;
        RECT 398.000 87.600 398.800 87.700 ;
        RECT 399.600 82.200 400.400 95.800 ;
        RECT 409.000 95.200 410.000 96.000 ;
        RECT 409.000 90.800 409.800 95.200 ;
        RECT 410.800 94.600 411.600 99.800 ;
        RECT 417.200 96.600 418.000 99.800 ;
        RECT 418.800 97.000 419.600 99.800 ;
        RECT 420.400 97.000 421.200 99.800 ;
        RECT 422.000 97.000 422.800 99.800 ;
        RECT 423.600 97.000 424.400 99.800 ;
        RECT 426.800 97.000 427.600 99.800 ;
        RECT 430.000 97.000 430.800 99.800 ;
        RECT 431.600 97.000 432.400 99.800 ;
        RECT 433.200 97.000 434.000 99.800 ;
        RECT 415.600 95.800 418.000 96.600 ;
        RECT 434.800 96.600 435.600 99.800 ;
        RECT 415.600 95.200 416.400 95.800 ;
        RECT 410.400 94.000 411.600 94.600 ;
        RECT 414.600 94.600 416.400 95.200 ;
        RECT 420.400 95.600 421.400 96.400 ;
        RECT 424.400 95.600 426.000 96.400 ;
        RECT 426.800 95.800 431.400 96.400 ;
        RECT 434.800 95.800 437.400 96.600 ;
        RECT 426.800 95.600 427.600 95.800 ;
        RECT 410.400 92.000 411.000 94.000 ;
        RECT 414.600 93.400 415.400 94.600 ;
        RECT 411.600 92.600 415.400 93.400 ;
        RECT 420.400 92.800 421.200 95.600 ;
        RECT 426.800 94.800 427.600 95.000 ;
        RECT 423.200 94.200 427.600 94.800 ;
        RECT 423.200 94.000 424.000 94.200 ;
        RECT 428.400 93.600 429.200 95.200 ;
        RECT 430.600 93.400 431.400 95.800 ;
        RECT 436.600 95.200 437.400 95.800 ;
        RECT 436.600 94.400 439.600 95.200 ;
        RECT 441.200 93.800 442.000 99.800 ;
        RECT 445.400 98.400 446.200 99.800 ;
        RECT 444.400 97.600 446.200 98.400 ;
        RECT 445.400 96.400 446.200 97.600 ;
        RECT 444.400 95.800 446.200 96.400 ;
        RECT 447.600 95.800 448.400 99.800 ;
        RECT 449.200 96.000 450.000 99.800 ;
        RECT 452.400 96.000 453.200 99.800 ;
        RECT 449.200 95.800 453.200 96.000 ;
        RECT 454.000 95.800 454.800 99.800 ;
        RECT 455.600 96.000 456.400 99.800 ;
        RECT 458.800 96.000 459.600 99.800 ;
        RECT 455.600 95.800 459.600 96.000 ;
        RECT 460.400 96.000 461.200 99.800 ;
        RECT 463.600 96.000 464.400 99.800 ;
        RECT 460.400 95.800 464.400 96.000 ;
        RECT 465.200 95.800 466.000 99.800 ;
        RECT 468.400 96.000 469.200 99.800 ;
        RECT 423.600 92.600 426.800 93.400 ;
        RECT 430.600 92.600 432.600 93.400 ;
        RECT 433.200 93.000 442.000 93.800 ;
        RECT 442.800 93.600 443.600 95.200 ;
        RECT 417.200 92.000 418.000 92.600 ;
        RECT 434.800 92.000 435.600 92.400 ;
        RECT 438.000 92.000 438.800 92.400 ;
        RECT 439.800 92.000 440.600 92.200 ;
        RECT 410.400 91.400 411.200 92.000 ;
        RECT 417.200 91.400 440.600 92.000 ;
        RECT 401.200 88.800 402.000 90.400 ;
        RECT 409.000 90.000 410.000 90.800 ;
        RECT 409.200 82.200 410.000 90.000 ;
        RECT 410.600 89.600 411.200 91.400 ;
        RECT 410.600 89.000 419.600 89.600 ;
        RECT 410.600 87.400 411.200 89.000 ;
        RECT 418.800 88.800 419.600 89.000 ;
        RECT 422.000 89.000 430.600 89.600 ;
        RECT 422.000 88.800 422.800 89.000 ;
        RECT 413.800 87.600 416.400 88.400 ;
        RECT 410.600 86.800 413.200 87.400 ;
        RECT 412.400 82.200 413.200 86.800 ;
        RECT 415.600 82.200 416.400 87.600 ;
        RECT 417.000 86.800 421.200 87.600 ;
        RECT 418.800 82.200 419.600 85.000 ;
        RECT 420.400 82.200 421.200 85.000 ;
        RECT 422.000 82.200 422.800 85.000 ;
        RECT 423.600 82.200 424.400 88.400 ;
        RECT 426.800 87.600 429.400 88.400 ;
        RECT 430.000 88.200 430.600 89.000 ;
        RECT 431.600 89.400 432.400 89.600 ;
        RECT 431.600 89.000 437.000 89.400 ;
        RECT 431.600 88.800 437.800 89.000 ;
        RECT 436.400 88.200 437.800 88.800 ;
        RECT 430.000 87.600 435.800 88.200 ;
        RECT 438.800 88.000 440.400 88.800 ;
        RECT 438.800 87.600 439.400 88.000 ;
        RECT 426.800 82.200 427.600 87.000 ;
        RECT 430.000 82.200 430.800 87.000 ;
        RECT 435.200 86.800 439.400 87.600 ;
        RECT 441.200 87.400 442.000 93.000 ;
        RECT 440.000 86.800 442.000 87.400 ;
        RECT 431.600 82.200 432.400 85.000 ;
        RECT 433.200 82.200 434.000 85.000 ;
        RECT 436.400 82.200 437.200 86.800 ;
        RECT 440.000 86.200 440.600 86.800 ;
        RECT 439.600 85.600 440.600 86.200 ;
        RECT 439.600 82.200 440.400 85.600 ;
        RECT 444.400 82.200 445.200 95.800 ;
        RECT 447.800 94.400 448.400 95.800 ;
        RECT 449.400 95.400 453.000 95.800 ;
        RECT 451.600 94.400 452.400 94.800 ;
        RECT 454.200 94.400 454.800 95.800 ;
        RECT 455.800 95.400 459.400 95.800 ;
        RECT 460.600 95.400 464.200 95.800 ;
        RECT 458.000 94.400 458.800 94.800 ;
        RECT 461.200 94.400 462.000 94.800 ;
        RECT 465.200 94.400 465.800 95.800 ;
        RECT 468.200 95.200 469.200 96.000 ;
        RECT 447.600 93.600 450.200 94.400 ;
        RECT 451.600 93.800 453.200 94.400 ;
        RECT 452.400 93.600 453.200 93.800 ;
        RECT 454.000 93.600 456.600 94.400 ;
        RECT 458.000 93.800 459.600 94.400 ;
        RECT 458.800 93.600 459.600 93.800 ;
        RECT 460.400 93.800 462.000 94.400 ;
        RECT 460.400 93.600 461.200 93.800 ;
        RECT 463.400 93.600 466.000 94.400 ;
        RECT 449.600 92.400 450.200 93.600 ;
        RECT 449.200 91.600 450.200 92.400 ;
        RECT 450.800 91.600 451.600 93.200 ;
        RECT 446.000 88.800 446.800 90.400 ;
        RECT 447.600 90.200 448.400 90.400 ;
        RECT 449.600 90.200 450.200 91.600 ;
        RECT 454.000 90.200 454.800 90.400 ;
        RECT 456.000 90.200 456.600 93.600 ;
        RECT 457.200 91.600 458.000 93.200 ;
        RECT 460.400 92.300 461.200 92.400 ;
        RECT 462.000 92.300 462.800 93.200 ;
        RECT 460.400 91.700 462.800 92.300 ;
        RECT 460.400 91.600 461.200 91.700 ;
        RECT 462.000 91.600 462.800 91.700 ;
        RECT 463.400 90.200 464.000 93.600 ;
        RECT 468.200 90.800 469.000 95.200 ;
        RECT 470.000 94.600 470.800 99.800 ;
        RECT 476.400 96.600 477.200 99.800 ;
        RECT 478.000 97.000 478.800 99.800 ;
        RECT 479.600 97.000 480.400 99.800 ;
        RECT 481.200 97.000 482.000 99.800 ;
        RECT 482.800 97.000 483.600 99.800 ;
        RECT 486.000 97.000 486.800 99.800 ;
        RECT 489.200 97.000 490.000 99.800 ;
        RECT 490.800 97.000 491.600 99.800 ;
        RECT 492.400 97.000 493.200 99.800 ;
        RECT 474.800 95.800 477.200 96.600 ;
        RECT 494.000 96.600 494.800 99.800 ;
        RECT 474.800 95.200 475.600 95.800 ;
        RECT 469.600 94.000 470.800 94.600 ;
        RECT 473.800 94.600 475.600 95.200 ;
        RECT 479.600 95.600 480.600 96.400 ;
        RECT 483.600 95.600 485.200 96.400 ;
        RECT 486.000 95.800 490.600 96.400 ;
        RECT 494.000 95.800 496.600 96.600 ;
        RECT 486.000 95.600 486.800 95.800 ;
        RECT 469.600 92.000 470.200 94.000 ;
        RECT 473.800 93.400 474.600 94.600 ;
        RECT 470.800 92.600 474.600 93.400 ;
        RECT 479.600 92.800 480.400 95.600 ;
        RECT 486.000 94.800 486.800 95.000 ;
        RECT 482.400 94.200 486.800 94.800 ;
        RECT 482.400 94.000 483.200 94.200 ;
        RECT 487.600 93.600 488.400 95.200 ;
        RECT 489.800 93.400 490.600 95.800 ;
        RECT 495.800 95.200 496.600 95.800 ;
        RECT 495.800 94.400 498.800 95.200 ;
        RECT 500.400 93.800 501.200 99.800 ;
        RECT 502.000 96.000 502.800 99.800 ;
        RECT 505.200 96.000 506.000 99.800 ;
        RECT 502.000 95.800 506.000 96.000 ;
        RECT 506.800 95.800 507.600 99.800 ;
        RECT 511.000 98.400 511.800 99.800 ;
        RECT 513.800 98.400 514.600 99.800 ;
        RECT 510.000 97.600 511.800 98.400 ;
        RECT 513.200 97.600 514.600 98.400 ;
        RECT 511.000 96.400 511.800 97.600 ;
        RECT 510.000 95.800 511.800 96.400 ;
        RECT 513.800 96.400 514.600 97.600 ;
        RECT 513.800 95.800 515.600 96.400 ;
        RECT 502.200 95.400 505.800 95.800 ;
        RECT 502.800 94.400 503.600 94.800 ;
        RECT 506.800 94.400 507.400 95.800 ;
        RECT 482.800 92.600 486.000 93.400 ;
        RECT 489.800 92.600 491.800 93.400 ;
        RECT 492.400 93.000 501.200 93.800 ;
        RECT 502.000 93.800 503.600 94.400 ;
        RECT 502.000 93.600 502.800 93.800 ;
        RECT 505.000 93.600 507.600 94.400 ;
        RECT 508.400 93.600 509.200 95.200 ;
        RECT 476.400 92.000 477.200 92.600 ;
        RECT 494.000 92.000 494.800 92.400 ;
        RECT 495.600 92.000 496.400 92.400 ;
        RECT 499.000 92.000 499.800 92.200 ;
        RECT 469.600 91.400 470.400 92.000 ;
        RECT 476.400 91.400 499.800 92.000 ;
        RECT 465.200 90.300 466.000 90.400 ;
        RECT 468.200 90.300 469.200 90.800 ;
        RECT 465.200 90.200 469.200 90.300 ;
        RECT 447.600 89.600 449.000 90.200 ;
        RECT 449.600 89.600 450.600 90.200 ;
        RECT 454.000 89.600 455.400 90.200 ;
        RECT 456.000 89.600 457.000 90.200 ;
        RECT 448.400 88.400 449.000 89.600 ;
        RECT 447.600 87.600 449.200 88.400 ;
        RECT 449.800 82.200 450.600 89.600 ;
        RECT 454.800 88.400 455.400 89.600 ;
        RECT 454.800 87.600 455.600 88.400 ;
        RECT 456.200 84.400 457.000 89.600 ;
        RECT 463.000 89.600 464.000 90.200 ;
        RECT 464.600 89.700 469.200 90.200 ;
        RECT 464.600 89.600 466.000 89.700 ;
        RECT 456.200 83.600 458.000 84.400 ;
        RECT 456.200 82.200 457.000 83.600 ;
        RECT 463.000 82.200 463.800 89.600 ;
        RECT 464.600 88.400 465.200 89.600 ;
        RECT 464.400 87.600 466.000 88.400 ;
        RECT 468.400 82.200 469.200 89.700 ;
        RECT 469.800 89.600 470.400 91.400 ;
        RECT 469.800 89.000 478.800 89.600 ;
        RECT 469.800 87.400 470.400 89.000 ;
        RECT 478.000 88.800 478.800 89.000 ;
        RECT 481.200 89.000 489.800 89.600 ;
        RECT 481.200 88.800 482.000 89.000 ;
        RECT 473.000 87.600 475.600 88.400 ;
        RECT 469.800 86.800 472.400 87.400 ;
        RECT 471.600 82.200 472.400 86.800 ;
        RECT 474.800 82.200 475.600 87.600 ;
        RECT 476.200 86.800 480.400 87.600 ;
        RECT 478.000 82.200 478.800 85.000 ;
        RECT 479.600 82.200 480.400 85.000 ;
        RECT 481.200 82.200 482.000 85.000 ;
        RECT 482.800 82.200 483.600 88.400 ;
        RECT 486.000 87.600 488.600 88.400 ;
        RECT 489.200 88.200 489.800 89.000 ;
        RECT 490.800 89.400 491.600 89.600 ;
        RECT 490.800 89.000 496.200 89.400 ;
        RECT 490.800 88.800 497.000 89.000 ;
        RECT 495.600 88.200 497.000 88.800 ;
        RECT 489.200 87.600 495.000 88.200 ;
        RECT 498.000 88.000 499.600 88.800 ;
        RECT 498.000 87.600 498.600 88.000 ;
        RECT 486.000 82.200 486.800 87.000 ;
        RECT 489.200 82.200 490.000 87.000 ;
        RECT 494.400 86.800 498.600 87.600 ;
        RECT 500.400 87.400 501.200 93.000 ;
        RECT 503.600 91.600 504.400 93.200 ;
        RECT 505.000 90.200 505.600 93.600 ;
        RECT 506.800 90.200 507.600 90.400 ;
        RECT 499.200 86.800 501.200 87.400 ;
        RECT 504.600 89.600 505.600 90.200 ;
        RECT 506.200 89.600 507.600 90.200 ;
        RECT 490.800 82.200 491.600 85.000 ;
        RECT 492.400 82.200 493.200 85.000 ;
        RECT 495.600 82.200 496.400 86.800 ;
        RECT 499.200 86.200 499.800 86.800 ;
        RECT 498.800 85.600 499.800 86.200 ;
        RECT 498.800 82.200 499.600 85.600 ;
        RECT 504.600 82.200 505.400 89.600 ;
        RECT 506.200 88.400 506.800 89.600 ;
        RECT 506.000 87.600 506.800 88.400 ;
        RECT 510.000 82.200 510.800 95.800 ;
        RECT 511.600 87.600 512.400 90.400 ;
        RECT 513.200 87.600 514.000 90.400 ;
        RECT 514.800 82.200 515.600 95.800 ;
        RECT 518.000 95.600 518.800 97.200 ;
        RECT 516.400 94.300 517.200 95.200 ;
        RECT 518.000 94.300 518.800 94.400 ;
        RECT 516.400 93.700 518.800 94.300 ;
        RECT 516.400 93.600 517.200 93.700 ;
        RECT 518.000 93.600 518.800 93.700 ;
        RECT 519.600 92.300 520.400 99.800 ;
        RECT 521.200 96.000 522.000 99.800 ;
        RECT 524.400 96.000 525.200 99.800 ;
        RECT 521.200 95.800 525.200 96.000 ;
        RECT 526.000 95.800 526.800 99.800 ;
        RECT 527.600 95.800 528.400 99.800 ;
        RECT 529.200 96.000 530.000 99.800 ;
        RECT 532.400 96.000 533.200 99.800 ;
        RECT 529.200 95.800 533.200 96.000 ;
        RECT 521.400 95.400 525.000 95.800 ;
        RECT 522.000 94.400 522.800 94.800 ;
        RECT 526.000 94.400 526.600 95.800 ;
        RECT 527.800 94.400 528.400 95.800 ;
        RECT 529.400 95.400 533.000 95.800 ;
        RECT 531.600 94.400 532.400 94.800 ;
        RECT 521.200 93.800 522.800 94.400 ;
        RECT 521.200 93.600 522.000 93.800 ;
        RECT 524.200 93.600 526.800 94.400 ;
        RECT 527.600 93.600 530.200 94.400 ;
        RECT 531.600 94.300 533.200 94.400 ;
        RECT 534.000 94.300 534.800 99.800 ;
        RECT 535.600 95.600 536.400 97.200 ;
        RECT 537.200 95.800 538.000 99.800 ;
        RECT 538.800 96.000 539.600 99.800 ;
        RECT 542.000 96.000 542.800 99.800 ;
        RECT 538.800 95.800 542.800 96.000 ;
        RECT 543.600 95.800 544.400 99.800 ;
        RECT 545.200 96.000 546.000 99.800 ;
        RECT 548.400 96.000 549.200 99.800 ;
        RECT 545.200 95.800 549.200 96.000 ;
        RECT 537.400 94.400 538.000 95.800 ;
        RECT 539.000 95.400 542.600 95.800 ;
        RECT 541.200 94.400 542.000 94.800 ;
        RECT 543.800 94.400 544.400 95.800 ;
        RECT 545.400 95.400 549.000 95.800 ;
        RECT 547.600 94.400 548.400 94.800 ;
        RECT 531.600 93.800 534.800 94.300 ;
        RECT 532.400 93.700 534.800 93.800 ;
        RECT 532.400 93.600 533.200 93.700 ;
        RECT 522.800 92.300 523.600 93.200 ;
        RECT 519.600 91.700 523.600 92.300 ;
        RECT 519.600 82.200 520.400 91.700 ;
        RECT 522.800 91.600 523.600 91.700 ;
        RECT 524.200 90.200 524.800 93.600 ;
        RECT 526.000 90.200 526.800 90.400 ;
        RECT 523.800 89.600 524.800 90.200 ;
        RECT 525.400 89.600 526.800 90.200 ;
        RECT 527.600 90.200 528.400 90.400 ;
        RECT 529.600 90.200 530.200 93.600 ;
        RECT 530.800 91.600 531.600 93.200 ;
        RECT 527.600 89.600 529.000 90.200 ;
        RECT 529.600 89.600 530.600 90.200 ;
        RECT 523.800 86.400 524.600 89.600 ;
        RECT 525.400 88.400 526.000 89.600 ;
        RECT 525.200 87.600 526.000 88.400 ;
        RECT 528.400 88.400 529.000 89.600 ;
        RECT 528.400 87.600 529.200 88.400 ;
        RECT 522.800 85.600 524.600 86.400 ;
        RECT 523.800 82.200 524.600 85.600 ;
        RECT 529.800 82.200 530.600 89.600 ;
        RECT 534.000 82.200 534.800 93.700 ;
        RECT 537.200 93.600 539.800 94.400 ;
        RECT 541.200 93.800 542.800 94.400 ;
        RECT 542.000 93.600 542.800 93.800 ;
        RECT 543.600 93.600 546.200 94.400 ;
        RECT 547.600 94.300 549.200 94.400 ;
        RECT 550.000 94.300 550.800 99.800 ;
        RECT 551.600 95.600 552.400 97.200 ;
        RECT 553.200 95.800 554.000 99.800 ;
        RECT 554.800 96.000 555.600 99.800 ;
        RECT 558.000 96.000 558.800 99.800 ;
        RECT 554.800 95.800 558.800 96.000 ;
        RECT 559.600 95.800 560.400 99.800 ;
        RECT 561.200 96.000 562.000 99.800 ;
        RECT 564.400 96.000 565.200 99.800 ;
        RECT 569.800 96.000 570.600 99.000 ;
        RECT 574.000 97.000 574.800 99.000 ;
        RECT 561.200 95.800 565.200 96.000 ;
        RECT 553.400 94.400 554.000 95.800 ;
        RECT 555.000 95.400 558.600 95.800 ;
        RECT 557.200 94.400 558.000 94.800 ;
        RECT 559.800 94.400 560.400 95.800 ;
        RECT 561.400 95.400 565.000 95.800 ;
        RECT 569.000 95.400 570.600 96.000 ;
        RECT 569.000 95.000 569.800 95.400 ;
        RECT 563.600 94.400 564.400 94.800 ;
        RECT 569.000 94.400 569.600 95.000 ;
        RECT 574.200 94.800 574.800 97.000 ;
        RECT 575.600 96.300 576.400 96.400 ;
        RECT 580.400 96.300 581.200 99.800 ;
        RECT 575.600 95.700 581.200 96.300 ;
        RECT 575.600 95.600 576.400 95.700 ;
        RECT 547.600 93.800 550.800 94.300 ;
        RECT 548.400 93.700 550.800 93.800 ;
        RECT 548.400 93.600 549.200 93.700 ;
        RECT 535.600 92.300 536.400 92.400 ;
        RECT 539.200 92.300 539.800 93.600 ;
        RECT 535.600 91.700 539.800 92.300 ;
        RECT 535.600 91.600 536.400 91.700 ;
        RECT 537.200 90.200 538.000 90.400 ;
        RECT 539.200 90.200 539.800 91.700 ;
        RECT 540.400 92.300 541.200 93.200 ;
        RECT 545.600 92.300 546.200 93.600 ;
        RECT 540.400 91.700 546.200 92.300 ;
        RECT 540.400 91.600 541.200 91.700 ;
        RECT 543.600 90.200 544.400 90.400 ;
        RECT 545.600 90.200 546.200 91.700 ;
        RECT 546.800 91.600 547.600 93.200 ;
        RECT 537.200 89.600 538.600 90.200 ;
        RECT 539.200 89.600 540.200 90.200 ;
        RECT 543.600 89.600 545.000 90.200 ;
        RECT 545.600 89.600 546.600 90.200 ;
        RECT 538.000 88.400 538.600 89.600 ;
        RECT 538.000 87.600 538.800 88.400 ;
        RECT 539.400 82.200 540.200 89.600 ;
        RECT 544.400 88.400 545.000 89.600 ;
        RECT 544.400 87.600 545.200 88.400 ;
        RECT 545.800 82.200 546.600 89.600 ;
        RECT 550.000 82.200 550.800 93.700 ;
        RECT 553.200 93.600 555.800 94.400 ;
        RECT 557.200 93.800 558.800 94.400 ;
        RECT 558.000 93.600 558.800 93.800 ;
        RECT 559.600 93.600 562.200 94.400 ;
        RECT 563.600 93.800 565.200 94.400 ;
        RECT 564.400 93.600 565.200 93.800 ;
        RECT 567.600 93.600 569.600 94.400 ;
        RECT 570.600 94.200 574.800 94.800 ;
        RECT 570.600 93.800 571.600 94.200 ;
        RECT 553.200 90.200 554.000 90.400 ;
        RECT 555.200 90.200 555.800 93.600 ;
        RECT 556.400 92.300 557.200 93.200 ;
        RECT 561.600 92.300 562.200 93.600 ;
        RECT 556.400 91.700 562.200 92.300 ;
        RECT 556.400 91.600 557.200 91.700 ;
        RECT 559.600 90.200 560.400 90.400 ;
        RECT 561.600 90.200 562.200 91.700 ;
        RECT 562.800 91.600 563.600 93.200 ;
        RECT 567.600 90.800 568.400 92.400 ;
        RECT 553.200 89.600 554.600 90.200 ;
        RECT 555.200 89.600 556.200 90.200 ;
        RECT 559.600 89.600 561.000 90.200 ;
        RECT 561.600 89.600 562.600 90.200 ;
        RECT 554.000 88.400 554.600 89.600 ;
        RECT 554.000 87.600 554.800 88.400 ;
        RECT 555.400 84.400 556.200 89.600 ;
        RECT 560.400 88.400 561.000 89.600 ;
        RECT 560.400 87.600 561.200 88.400 ;
        RECT 555.400 83.600 557.200 84.400 ;
        RECT 555.400 82.200 556.200 83.600 ;
        RECT 561.800 82.200 562.600 89.600 ;
        RECT 569.000 89.800 569.600 93.600 ;
        RECT 570.200 93.000 571.600 93.800 ;
        RECT 571.000 91.000 571.600 93.000 ;
        RECT 572.400 91.600 573.200 93.200 ;
        RECT 574.000 91.600 574.800 93.200 ;
        RECT 571.000 90.400 574.800 91.000 ;
        RECT 569.000 89.200 570.600 89.800 ;
        RECT 569.800 84.400 570.600 89.200 ;
        RECT 574.200 87.000 574.800 90.400 ;
        RECT 569.800 83.600 571.600 84.400 ;
        RECT 569.800 82.200 570.600 83.600 ;
        RECT 574.000 83.000 574.800 87.000 ;
        RECT 580.400 82.200 581.200 95.700 ;
        RECT 582.000 96.300 582.800 97.200 ;
        RECT 583.600 96.300 584.400 99.800 ;
        RECT 587.800 98.400 589.000 99.800 ;
        RECT 587.800 97.800 589.200 98.400 ;
        RECT 592.400 97.800 593.200 99.800 ;
        RECT 596.800 98.400 597.600 99.800 ;
        RECT 596.800 97.800 598.800 98.400 ;
        RECT 588.400 97.000 589.200 97.800 ;
        RECT 592.600 97.200 593.200 97.800 ;
        RECT 592.600 96.600 595.400 97.200 ;
        RECT 594.600 96.400 595.400 96.600 ;
        RECT 596.400 96.400 597.200 97.200 ;
        RECT 598.000 97.000 598.800 97.800 ;
        RECT 582.000 95.700 584.400 96.300 ;
        RECT 582.000 95.600 582.800 95.700 ;
        RECT 583.600 95.400 584.400 95.700 ;
        RECT 586.600 95.400 587.400 95.600 ;
        RECT 583.600 94.800 587.400 95.400 ;
        RECT 583.600 91.400 584.400 94.800 ;
        RECT 590.600 94.200 591.400 94.400 ;
        RECT 596.400 94.200 597.000 96.400 ;
        RECT 601.200 95.000 602.000 99.800 ;
        RECT 602.800 97.000 603.600 99.000 ;
        RECT 602.800 94.800 603.400 97.000 ;
        RECT 607.000 96.000 607.800 99.000 ;
        RECT 607.000 95.400 608.600 96.000 ;
        RECT 612.400 95.800 613.200 99.800 ;
        RECT 614.000 96.000 614.800 99.800 ;
        RECT 617.200 96.000 618.000 99.800 ;
        RECT 614.000 95.800 618.000 96.000 ;
        RECT 618.800 96.000 619.600 99.800 ;
        RECT 622.000 96.000 622.800 99.800 ;
        RECT 618.800 95.800 622.800 96.000 ;
        RECT 623.600 95.800 624.400 99.800 ;
        RECT 625.200 95.800 626.000 99.800 ;
        RECT 626.800 96.000 627.600 99.800 ;
        RECT 630.000 96.000 630.800 99.800 ;
        RECT 626.800 95.800 630.800 96.000 ;
        RECT 607.800 95.000 608.600 95.400 ;
        RECT 599.600 94.200 601.200 94.400 ;
        RECT 602.800 94.200 607.000 94.800 ;
        RECT 590.200 93.600 601.200 94.200 ;
        RECT 606.000 93.800 607.000 94.200 ;
        RECT 608.000 94.400 608.600 95.000 ;
        RECT 612.600 94.400 613.200 95.800 ;
        RECT 614.200 95.400 617.800 95.800 ;
        RECT 619.000 95.400 622.600 95.800 ;
        RECT 616.400 94.400 617.200 94.800 ;
        RECT 619.600 94.400 620.400 94.800 ;
        RECT 623.600 94.400 624.200 95.800 ;
        RECT 625.400 94.400 626.000 95.800 ;
        RECT 627.000 95.400 630.600 95.800 ;
        RECT 631.600 95.200 632.400 99.800 ;
        RECT 634.800 96.400 635.600 99.800 ;
        RECT 634.800 95.800 635.800 96.400 ;
        RECT 638.000 96.000 638.800 99.800 ;
        RECT 641.200 96.000 642.000 99.800 ;
        RECT 638.000 95.800 642.000 96.000 ;
        RECT 642.800 95.800 643.600 99.800 ;
        RECT 644.400 96.000 645.200 99.800 ;
        RECT 647.600 96.000 648.400 99.800 ;
        RECT 644.400 95.800 648.400 96.000 ;
        RECT 649.200 95.800 650.000 99.800 ;
        RECT 629.200 94.400 630.000 94.800 ;
        RECT 631.600 94.600 634.200 95.200 ;
        RECT 608.000 94.300 610.000 94.400 ;
        RECT 610.800 94.300 611.600 94.400 ;
        RECT 588.400 92.800 589.200 93.000 ;
        RECT 585.400 92.200 589.200 92.800 ;
        RECT 585.400 92.000 586.200 92.200 ;
        RECT 587.000 91.400 587.800 91.600 ;
        RECT 583.600 90.800 587.800 91.400 ;
        RECT 583.600 82.200 584.400 90.800 ;
        RECT 590.200 90.400 590.800 93.600 ;
        RECT 597.400 93.400 598.200 93.600 ;
        RECT 596.400 92.400 597.200 92.600 ;
        RECT 599.000 92.400 599.800 92.600 ;
        RECT 594.800 91.800 599.800 92.400 ;
        RECT 594.800 91.600 595.600 91.800 ;
        RECT 602.800 91.600 603.600 93.200 ;
        RECT 604.400 91.600 605.200 93.200 ;
        RECT 606.000 93.000 607.400 93.800 ;
        RECT 608.000 93.700 611.600 94.300 ;
        RECT 608.000 93.600 610.000 93.700 ;
        RECT 610.800 93.600 611.600 93.700 ;
        RECT 612.400 93.600 615.000 94.400 ;
        RECT 616.400 93.800 618.000 94.400 ;
        RECT 617.200 93.600 618.000 93.800 ;
        RECT 618.800 93.800 620.400 94.400 ;
        RECT 618.800 93.600 619.600 93.800 ;
        RECT 621.800 93.600 624.400 94.400 ;
        RECT 625.200 93.600 627.800 94.400 ;
        RECT 629.200 93.800 630.800 94.400 ;
        RECT 630.000 93.600 630.800 93.800 ;
        RECT 596.400 91.000 602.000 91.200 ;
        RECT 606.000 91.000 606.600 93.000 ;
        RECT 596.200 90.800 602.000 91.000 ;
        RECT 588.400 89.800 590.800 90.400 ;
        RECT 592.200 90.600 602.000 90.800 ;
        RECT 592.200 90.200 597.000 90.600 ;
        RECT 588.400 88.800 589.000 89.800 ;
        RECT 587.600 88.000 589.000 88.800 ;
        RECT 590.600 89.000 591.400 89.200 ;
        RECT 592.200 89.000 592.800 90.200 ;
        RECT 590.600 88.400 592.800 89.000 ;
        RECT 593.400 89.000 598.800 89.600 ;
        RECT 593.400 88.800 594.200 89.000 ;
        RECT 598.000 88.800 598.800 89.000 ;
        RECT 591.800 87.400 592.600 87.600 ;
        RECT 594.600 87.400 595.400 87.600 ;
        RECT 588.400 86.200 589.200 87.000 ;
        RECT 591.800 86.800 595.400 87.400 ;
        RECT 592.600 86.200 593.200 86.800 ;
        RECT 598.000 86.200 598.800 87.000 ;
        RECT 587.800 82.200 589.000 86.200 ;
        RECT 592.400 82.200 593.200 86.200 ;
        RECT 596.800 85.600 598.800 86.200 ;
        RECT 596.800 82.200 597.600 85.600 ;
        RECT 601.200 82.200 602.000 90.600 ;
        RECT 602.800 90.400 606.600 91.000 ;
        RECT 602.800 87.000 603.400 90.400 ;
        RECT 608.000 89.800 608.600 93.600 ;
        RECT 609.200 90.800 610.000 92.400 ;
        RECT 607.000 89.200 608.600 89.800 ;
        RECT 612.400 90.200 613.200 90.400 ;
        RECT 614.400 90.200 615.000 93.600 ;
        RECT 615.600 91.600 616.400 93.200 ;
        RECT 620.400 91.600 621.200 93.200 ;
        RECT 621.800 90.400 622.400 93.600 ;
        RECT 627.200 92.300 627.800 93.600 ;
        RECT 623.700 91.700 627.800 92.300 ;
        RECT 623.700 90.400 624.300 91.700 ;
        RECT 612.400 89.600 613.800 90.200 ;
        RECT 614.400 89.600 615.400 90.200 ;
        RECT 620.400 89.600 622.400 90.400 ;
        RECT 623.600 90.200 624.400 90.400 ;
        RECT 623.000 89.600 624.400 90.200 ;
        RECT 625.200 90.200 626.000 90.400 ;
        RECT 627.200 90.200 627.800 91.700 ;
        RECT 628.400 92.300 629.200 93.200 ;
        RECT 631.800 92.400 632.600 93.200 ;
        RECT 630.000 92.300 630.800 92.400 ;
        RECT 628.400 91.700 630.800 92.300 ;
        RECT 628.400 91.600 629.200 91.700 ;
        RECT 630.000 91.600 630.800 91.700 ;
        RECT 631.600 91.600 632.600 92.400 ;
        RECT 633.600 93.000 634.200 94.600 ;
        RECT 635.200 94.400 635.800 95.800 ;
        RECT 638.200 95.400 641.800 95.800 ;
        RECT 638.800 94.400 639.600 94.800 ;
        RECT 642.800 94.400 643.400 95.800 ;
        RECT 644.600 95.400 648.200 95.800 ;
        RECT 645.200 94.400 646.000 94.800 ;
        RECT 649.200 94.400 649.800 95.800 ;
        RECT 650.800 95.400 651.600 99.800 ;
        RECT 655.000 98.400 656.200 99.800 ;
        RECT 655.000 97.800 656.400 98.400 ;
        RECT 659.600 97.800 660.400 99.800 ;
        RECT 664.000 98.400 664.800 99.800 ;
        RECT 664.000 97.800 666.000 98.400 ;
        RECT 655.600 97.000 656.400 97.800 ;
        RECT 659.800 97.200 660.400 97.800 ;
        RECT 659.800 96.600 662.600 97.200 ;
        RECT 661.800 96.400 662.600 96.600 ;
        RECT 663.600 96.400 664.400 97.200 ;
        RECT 665.200 97.000 666.000 97.800 ;
        RECT 653.800 95.400 654.600 95.600 ;
        RECT 650.800 94.800 654.600 95.400 ;
        RECT 634.800 93.600 635.800 94.400 ;
        RECT 636.400 94.300 637.200 94.400 ;
        RECT 638.000 94.300 639.600 94.400 ;
        RECT 636.400 93.800 639.600 94.300 ;
        RECT 636.400 93.700 638.800 93.800 ;
        RECT 636.400 93.600 637.200 93.700 ;
        RECT 638.000 93.600 638.800 93.700 ;
        RECT 641.000 93.600 643.600 94.400 ;
        RECT 644.400 93.800 646.000 94.400 ;
        RECT 644.400 93.600 645.200 93.800 ;
        RECT 647.400 93.600 650.000 94.400 ;
        RECT 633.600 92.200 634.600 93.000 ;
        RECT 633.600 90.200 634.200 92.200 ;
        RECT 635.200 90.200 635.800 93.600 ;
        RECT 636.400 92.300 637.200 92.400 ;
        RECT 639.600 92.300 640.400 93.200 ;
        RECT 636.400 91.700 640.400 92.300 ;
        RECT 636.400 91.600 637.200 91.700 ;
        RECT 639.600 91.600 640.400 91.700 ;
        RECT 641.000 92.400 641.600 93.600 ;
        RECT 641.000 91.600 642.000 92.400 ;
        RECT 646.000 91.600 646.800 93.200 ;
        RECT 641.000 90.200 641.600 91.600 ;
        RECT 642.800 90.200 643.600 90.400 ;
        RECT 647.400 90.200 648.000 93.600 ;
        RECT 650.800 91.400 651.600 94.800 ;
        RECT 657.800 94.200 658.600 94.400 ;
        RECT 663.600 94.200 664.200 96.400 ;
        RECT 668.400 95.000 669.200 99.800 ;
        RECT 670.000 95.000 670.800 99.800 ;
        RECT 674.400 98.400 675.200 99.800 ;
        RECT 673.200 97.800 675.200 98.400 ;
        RECT 678.800 97.800 679.600 99.800 ;
        RECT 683.000 98.400 684.200 99.800 ;
        RECT 682.800 97.800 684.200 98.400 ;
        RECT 673.200 97.000 674.000 97.800 ;
        RECT 678.800 97.200 679.400 97.800 ;
        RECT 674.800 96.400 675.600 97.200 ;
        RECT 676.600 96.600 679.400 97.200 ;
        RECT 682.800 97.000 683.600 97.800 ;
        RECT 676.600 96.400 677.400 96.600 ;
        RECT 666.800 94.300 668.400 94.400 ;
        RECT 670.800 94.300 672.400 94.400 ;
        RECT 666.800 94.200 672.400 94.300 ;
        RECT 675.000 94.200 675.600 96.400 ;
        RECT 684.600 95.400 685.400 95.600 ;
        RECT 687.600 95.400 688.400 99.800 ;
        RECT 684.600 94.800 688.400 95.400 ;
        RECT 680.600 94.200 681.400 94.400 ;
        RECT 657.400 93.700 681.800 94.200 ;
        RECT 657.400 93.600 668.400 93.700 ;
        RECT 670.800 93.600 681.800 93.700 ;
        RECT 655.600 92.800 656.400 93.000 ;
        RECT 652.600 92.200 656.400 92.800 ;
        RECT 657.400 92.400 658.000 93.600 ;
        RECT 664.600 93.400 665.400 93.600 ;
        RECT 673.800 93.400 674.600 93.600 ;
        RECT 663.600 92.400 664.400 92.600 ;
        RECT 666.200 92.400 667.000 92.600 ;
        RECT 652.600 92.000 653.400 92.200 ;
        RECT 657.200 91.600 658.000 92.400 ;
        RECT 662.000 91.800 667.000 92.400 ;
        RECT 672.200 92.400 673.000 92.600 ;
        RECT 672.200 92.300 677.200 92.400 ;
        RECT 679.600 92.300 680.400 92.400 ;
        RECT 672.200 91.800 680.400 92.300 ;
        RECT 662.000 91.600 662.800 91.800 ;
        RECT 676.400 91.700 680.400 91.800 ;
        RECT 676.400 91.600 677.200 91.700 ;
        RECT 679.600 91.600 680.400 91.700 ;
        RECT 654.200 91.400 655.000 91.600 ;
        RECT 650.800 90.800 655.000 91.400 ;
        RECT 649.200 90.300 650.000 90.400 ;
        RECT 650.800 90.300 651.600 90.800 ;
        RECT 657.400 90.400 658.000 91.600 ;
        RECT 663.600 91.000 669.200 91.200 ;
        RECT 663.400 90.800 669.200 91.000 ;
        RECT 649.200 90.200 651.600 90.300 ;
        RECT 625.200 89.600 626.600 90.200 ;
        RECT 627.200 89.600 628.200 90.200 ;
        RECT 602.800 83.000 603.600 87.000 ;
        RECT 607.000 82.200 607.800 89.200 ;
        RECT 613.200 88.400 613.800 89.600 ;
        RECT 613.200 87.600 614.000 88.400 ;
        RECT 614.600 82.200 615.400 89.600 ;
        RECT 621.400 82.200 622.200 89.600 ;
        RECT 623.000 88.400 623.600 89.600 ;
        RECT 622.800 87.600 623.600 88.400 ;
        RECT 626.000 88.400 626.600 89.600 ;
        RECT 626.000 87.600 626.800 88.400 ;
        RECT 627.400 82.200 628.200 89.600 ;
        RECT 631.600 89.600 634.200 90.200 ;
        RECT 631.600 82.200 632.400 89.600 ;
        RECT 634.800 89.200 635.800 90.200 ;
        RECT 640.600 89.600 641.600 90.200 ;
        RECT 642.200 89.600 643.600 90.200 ;
        RECT 647.000 89.600 648.000 90.200 ;
        RECT 648.600 89.700 651.600 90.200 ;
        RECT 648.600 89.600 650.000 89.700 ;
        RECT 634.800 82.200 635.600 89.200 ;
        RECT 640.600 82.200 641.400 89.600 ;
        RECT 642.200 88.400 642.800 89.600 ;
        RECT 642.000 87.600 642.800 88.400 ;
        RECT 647.000 84.400 647.800 89.600 ;
        RECT 648.600 88.400 649.200 89.600 ;
        RECT 648.400 87.600 649.200 88.400 ;
        RECT 646.000 83.600 647.800 84.400 ;
        RECT 647.000 82.200 647.800 83.600 ;
        RECT 650.800 82.200 651.600 89.700 ;
        RECT 655.600 89.800 658.000 90.400 ;
        RECT 659.400 90.600 669.200 90.800 ;
        RECT 659.400 90.200 664.200 90.600 ;
        RECT 655.600 88.800 656.200 89.800 ;
        RECT 654.800 88.000 656.200 88.800 ;
        RECT 657.800 89.000 658.600 89.200 ;
        RECT 659.400 89.000 660.000 90.200 ;
        RECT 657.800 88.400 660.000 89.000 ;
        RECT 660.600 89.000 666.000 89.600 ;
        RECT 660.600 88.800 661.400 89.000 ;
        RECT 665.200 88.800 666.000 89.000 ;
        RECT 659.000 87.400 659.800 87.600 ;
        RECT 661.800 87.400 662.600 87.600 ;
        RECT 655.600 86.200 656.400 87.000 ;
        RECT 659.000 86.800 662.600 87.400 ;
        RECT 659.800 86.200 660.400 86.800 ;
        RECT 665.200 86.200 666.000 87.000 ;
        RECT 655.000 82.200 656.200 86.200 ;
        RECT 659.600 82.200 660.400 86.200 ;
        RECT 664.000 85.600 666.000 86.200 ;
        RECT 664.000 82.200 664.800 85.600 ;
        RECT 668.400 82.200 669.200 90.600 ;
        RECT 670.000 91.000 675.600 91.200 ;
        RECT 670.000 90.800 675.800 91.000 ;
        RECT 670.000 90.600 679.800 90.800 ;
        RECT 670.000 82.200 670.800 90.600 ;
        RECT 675.000 90.200 679.800 90.600 ;
        RECT 673.200 89.000 678.600 89.600 ;
        RECT 673.200 88.800 674.000 89.000 ;
        RECT 677.800 88.800 678.600 89.000 ;
        RECT 679.200 89.000 679.800 90.200 ;
        RECT 681.200 90.400 681.800 93.600 ;
        RECT 682.800 92.800 683.600 93.000 ;
        RECT 682.800 92.200 686.600 92.800 ;
        RECT 685.800 92.000 686.600 92.200 ;
        RECT 684.200 91.400 685.000 91.600 ;
        RECT 687.600 91.400 688.400 94.800 ;
        RECT 684.200 90.800 688.400 91.400 ;
        RECT 681.200 89.800 683.600 90.400 ;
        RECT 680.600 89.000 681.400 89.200 ;
        RECT 679.200 88.400 681.400 89.000 ;
        RECT 683.000 88.800 683.600 89.800 ;
        RECT 683.000 88.000 684.400 88.800 ;
        RECT 676.600 87.400 677.400 87.600 ;
        RECT 679.400 87.400 680.200 87.600 ;
        RECT 673.200 86.200 674.000 87.000 ;
        RECT 676.600 86.800 680.200 87.400 ;
        RECT 678.800 86.200 679.400 86.800 ;
        RECT 682.800 86.200 683.600 87.000 ;
        RECT 673.200 85.600 675.200 86.200 ;
        RECT 674.400 82.200 675.200 85.600 ;
        RECT 678.800 82.200 679.600 86.200 ;
        RECT 683.000 82.200 684.200 86.200 ;
        RECT 687.600 82.200 688.400 90.800 ;
        RECT 1.200 71.400 2.000 79.800 ;
        RECT 5.600 76.400 6.400 79.800 ;
        RECT 4.400 75.800 6.400 76.400 ;
        RECT 10.000 75.800 10.800 79.800 ;
        RECT 14.200 75.800 15.400 79.800 ;
        RECT 4.400 75.000 5.200 75.800 ;
        RECT 10.000 75.200 10.600 75.800 ;
        RECT 7.800 74.600 11.400 75.200 ;
        RECT 14.000 75.000 14.800 75.800 ;
        RECT 7.800 74.400 8.600 74.600 ;
        RECT 10.600 74.400 11.400 74.600 ;
        RECT 4.400 73.000 5.200 73.200 ;
        RECT 9.000 73.000 9.800 73.200 ;
        RECT 4.400 72.400 9.800 73.000 ;
        RECT 10.400 73.000 12.600 73.600 ;
        RECT 10.400 71.800 11.000 73.000 ;
        RECT 11.800 72.800 12.600 73.000 ;
        RECT 14.200 73.200 15.600 74.000 ;
        RECT 14.200 72.200 14.800 73.200 ;
        RECT 6.200 71.400 11.000 71.800 ;
        RECT 1.200 71.200 11.000 71.400 ;
        RECT 12.400 71.600 14.800 72.200 ;
        RECT 1.200 71.000 7.000 71.200 ;
        RECT 1.200 70.800 6.800 71.000 ;
        RECT 7.600 70.300 8.400 70.400 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 7.600 70.200 10.000 70.300 ;
        RECT 3.400 69.700 10.000 70.200 ;
        RECT 3.400 69.600 8.400 69.700 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 3.400 69.400 4.200 69.600 ;
        RECT 5.000 68.400 5.800 68.600 ;
        RECT 12.400 68.400 13.000 71.600 ;
        RECT 18.800 71.200 19.600 79.800 ;
        RECT 23.000 72.400 23.800 79.800 ;
        RECT 24.400 73.600 25.200 74.400 ;
        RECT 24.600 72.400 25.200 73.600 ;
        RECT 27.600 73.600 28.400 74.400 ;
        RECT 27.600 72.400 28.200 73.600 ;
        RECT 29.000 72.400 29.800 79.800 ;
        RECT 23.000 71.800 24.000 72.400 ;
        RECT 24.600 71.800 26.000 72.400 ;
        RECT 15.400 70.600 19.600 71.200 ;
        RECT 15.400 70.400 16.200 70.600 ;
        RECT 17.000 69.800 17.800 70.000 ;
        RECT 14.000 69.200 17.800 69.800 ;
        RECT 14.000 69.000 14.800 69.200 ;
        RECT 2.000 67.800 13.000 68.400 ;
        RECT 2.000 67.600 3.600 67.800 ;
        RECT 1.200 62.200 2.000 67.000 ;
        RECT 6.200 66.400 6.800 67.800 ;
        RECT 11.800 67.600 12.600 67.800 ;
        RECT 18.800 67.200 19.600 70.600 ;
        RECT 20.400 70.300 21.200 70.400 ;
        RECT 22.000 70.300 22.800 70.400 ;
        RECT 20.400 69.700 22.800 70.300 ;
        RECT 20.400 69.600 21.200 69.700 ;
        RECT 22.000 68.800 22.800 69.700 ;
        RECT 23.400 70.300 24.000 71.800 ;
        RECT 25.200 71.600 26.000 71.800 ;
        RECT 26.800 71.800 28.200 72.400 ;
        RECT 28.800 71.800 29.800 72.400 ;
        RECT 33.200 75.000 34.000 79.000 ;
        RECT 26.800 71.600 27.600 71.800 ;
        RECT 26.900 70.300 27.500 71.600 ;
        RECT 23.400 69.700 27.500 70.300 ;
        RECT 23.400 68.400 24.000 69.700 ;
        RECT 28.800 68.400 29.400 71.800 ;
        RECT 33.200 71.600 33.800 75.000 ;
        RECT 37.400 72.800 38.200 79.800 ;
        RECT 43.600 73.600 44.400 74.400 ;
        RECT 37.400 72.200 39.000 72.800 ;
        RECT 43.600 72.400 44.200 73.600 ;
        RECT 45.000 72.400 45.800 79.800 ;
        RECT 53.000 72.800 53.800 79.800 ;
        RECT 57.200 75.000 58.000 79.000 ;
        RECT 33.200 71.000 37.000 71.600 ;
        RECT 30.000 68.800 30.800 70.400 ;
        RECT 33.200 68.800 34.000 70.400 ;
        RECT 34.800 68.800 35.600 70.400 ;
        RECT 36.400 69.000 37.000 71.000 ;
        RECT 38.400 70.400 39.000 72.200 ;
        RECT 42.800 71.800 44.200 72.400 ;
        RECT 42.800 71.600 43.600 71.800 ;
        RECT 44.800 71.600 46.800 72.400 ;
        RECT 52.200 72.200 53.800 72.800 ;
        RECT 38.000 69.600 39.000 70.400 ;
        RECT 39.600 70.300 40.400 71.200 ;
        RECT 42.800 70.300 43.600 70.400 ;
        RECT 39.600 69.700 43.600 70.300 ;
        RECT 39.600 69.600 40.400 69.700 ;
        RECT 42.800 69.600 43.600 69.700 ;
        RECT 20.400 68.200 21.200 68.400 ;
        RECT 20.400 67.600 22.000 68.200 ;
        RECT 23.400 67.600 26.000 68.400 ;
        RECT 26.800 67.600 29.400 68.400 ;
        RECT 31.600 68.200 32.400 68.400 ;
        RECT 30.800 67.600 32.400 68.200 ;
        RECT 36.400 68.200 37.800 69.000 ;
        RECT 38.400 68.400 39.000 69.600 ;
        RECT 44.800 68.400 45.400 71.600 ;
        RECT 46.000 70.300 46.800 70.400 ;
        RECT 46.000 69.700 49.900 70.300 ;
        RECT 46.000 68.800 46.800 69.700 ;
        RECT 36.400 67.800 37.400 68.200 ;
        RECT 21.200 67.200 22.000 67.600 ;
        RECT 15.800 66.600 19.600 67.200 ;
        RECT 15.800 66.400 16.600 66.600 ;
        RECT 4.400 64.200 5.200 65.000 ;
        RECT 6.000 64.800 6.800 66.400 ;
        RECT 7.800 65.400 8.600 65.600 ;
        RECT 7.800 64.800 10.600 65.400 ;
        RECT 10.000 64.200 10.600 64.800 ;
        RECT 14.000 64.200 14.800 65.000 ;
        RECT 4.400 63.600 6.400 64.200 ;
        RECT 5.600 62.200 6.400 63.600 ;
        RECT 10.000 62.200 10.800 64.200 ;
        RECT 14.000 63.600 15.400 64.200 ;
        RECT 14.200 62.200 15.400 63.600 ;
        RECT 18.800 62.200 19.600 66.600 ;
        RECT 20.600 66.200 24.200 66.600 ;
        RECT 25.200 66.200 25.800 67.600 ;
        RECT 27.000 66.400 27.600 67.600 ;
        RECT 30.800 67.200 31.600 67.600 ;
        RECT 33.200 67.200 37.400 67.800 ;
        RECT 38.400 67.600 40.400 68.400 ;
        RECT 42.800 67.600 45.400 68.400 ;
        RECT 47.600 68.200 48.400 68.400 ;
        RECT 46.800 67.600 48.400 68.200 ;
        RECT 49.300 68.300 49.900 69.700 ;
        RECT 50.800 69.600 51.600 71.200 ;
        RECT 52.200 68.400 52.800 72.200 ;
        RECT 57.400 71.600 58.000 75.000 ;
        RECT 62.600 72.800 63.400 79.800 ;
        RECT 66.800 75.000 67.600 79.000 ;
        RECT 54.200 71.000 58.000 71.600 ;
        RECT 61.800 72.200 63.400 72.800 ;
        RECT 54.200 69.000 54.800 71.000 ;
        RECT 50.800 68.300 52.800 68.400 ;
        RECT 49.300 67.700 52.800 68.300 ;
        RECT 53.400 68.200 54.800 69.000 ;
        RECT 55.600 68.800 56.400 70.400 ;
        RECT 57.200 70.300 58.000 70.400 ;
        RECT 58.800 70.300 59.600 70.400 ;
        RECT 57.200 69.700 59.600 70.300 ;
        RECT 57.200 68.800 58.000 69.700 ;
        RECT 58.800 69.600 59.600 69.700 ;
        RECT 60.400 69.600 61.200 71.200 ;
        RECT 61.800 68.400 62.400 72.200 ;
        RECT 67.000 71.600 67.600 75.000 ;
        RECT 63.800 71.000 67.600 71.600 ;
        RECT 68.400 71.400 69.200 79.800 ;
        RECT 72.800 76.400 73.600 79.800 ;
        RECT 71.600 75.800 73.600 76.400 ;
        RECT 77.200 75.800 78.000 79.800 ;
        RECT 81.400 75.800 82.600 79.800 ;
        RECT 71.600 75.000 72.400 75.800 ;
        RECT 77.200 75.200 77.800 75.800 ;
        RECT 75.000 74.600 78.600 75.200 ;
        RECT 81.200 75.000 82.000 75.800 ;
        RECT 75.000 74.400 75.800 74.600 ;
        RECT 77.800 74.400 78.600 74.600 ;
        RECT 71.600 73.000 72.400 73.200 ;
        RECT 76.200 73.000 77.000 73.200 ;
        RECT 71.600 72.400 77.000 73.000 ;
        RECT 77.600 73.000 79.800 73.600 ;
        RECT 77.600 71.800 78.200 73.000 ;
        RECT 79.000 72.800 79.800 73.000 ;
        RECT 81.400 73.200 82.800 74.000 ;
        RECT 81.400 72.200 82.000 73.200 ;
        RECT 73.400 71.400 78.200 71.800 ;
        RECT 68.400 71.200 78.200 71.400 ;
        RECT 79.600 71.600 82.000 72.200 ;
        RECT 68.400 71.000 74.200 71.200 ;
        RECT 63.800 69.000 64.400 71.000 ;
        RECT 68.400 70.800 74.000 71.000 ;
        RECT 50.800 67.600 52.800 67.700 ;
        RECT 20.400 66.000 24.400 66.200 ;
        RECT 20.400 62.200 21.200 66.000 ;
        RECT 23.600 62.200 24.400 66.000 ;
        RECT 25.200 62.200 26.000 66.200 ;
        RECT 26.800 62.200 27.600 66.400 ;
        RECT 28.600 66.200 32.200 66.600 ;
        RECT 28.400 66.000 32.400 66.200 ;
        RECT 28.400 62.200 29.200 66.000 ;
        RECT 31.600 62.200 32.400 66.000 ;
        RECT 33.200 65.000 33.800 67.200 ;
        RECT 38.400 67.000 39.000 67.600 ;
        RECT 38.200 66.600 39.000 67.000 ;
        RECT 37.400 66.000 39.000 66.600 ;
        RECT 43.000 66.200 43.600 67.600 ;
        RECT 46.800 67.200 47.600 67.600 ;
        RECT 52.200 67.000 52.800 67.600 ;
        RECT 53.800 67.800 54.800 68.200 ;
        RECT 53.800 67.200 58.000 67.800 ;
        RECT 60.400 67.600 62.400 68.400 ;
        RECT 63.000 68.200 64.400 69.000 ;
        RECT 65.200 68.800 66.000 70.400 ;
        RECT 66.800 68.800 67.600 70.400 ;
        RECT 74.800 70.200 75.600 70.400 ;
        RECT 70.600 69.600 75.600 70.200 ;
        RECT 70.600 69.400 71.400 69.600 ;
        RECT 73.200 69.400 74.000 69.600 ;
        RECT 72.200 68.400 73.000 68.600 ;
        RECT 79.600 68.400 80.200 71.600 ;
        RECT 86.000 71.200 86.800 79.800 ;
        RECT 82.600 70.600 86.800 71.200 ;
        RECT 82.600 70.400 83.400 70.600 ;
        RECT 84.200 69.800 85.000 70.000 ;
        RECT 81.200 69.200 85.000 69.800 ;
        RECT 81.200 69.000 82.000 69.200 ;
        RECT 52.200 66.600 53.000 67.000 ;
        RECT 44.600 66.200 48.200 66.600 ;
        RECT 33.200 63.000 34.000 65.000 ;
        RECT 37.400 63.000 38.200 66.000 ;
        RECT 42.800 62.200 43.600 66.200 ;
        RECT 44.400 66.000 48.400 66.200 ;
        RECT 52.200 66.000 53.800 66.600 ;
        RECT 44.400 62.200 45.200 66.000 ;
        RECT 47.600 62.200 48.400 66.000 ;
        RECT 53.000 63.000 53.800 66.000 ;
        RECT 57.400 65.000 58.000 67.200 ;
        RECT 61.800 67.000 62.400 67.600 ;
        RECT 63.400 67.800 64.400 68.200 ;
        RECT 69.200 67.800 80.200 68.400 ;
        RECT 63.400 67.200 67.600 67.800 ;
        RECT 69.200 67.600 70.800 67.800 ;
        RECT 61.800 66.600 62.600 67.000 ;
        RECT 61.800 66.000 63.400 66.600 ;
        RECT 57.200 63.000 58.000 65.000 ;
        RECT 62.600 64.400 63.400 66.000 ;
        RECT 67.000 65.000 67.600 67.200 ;
        RECT 62.000 63.600 63.400 64.400 ;
        RECT 62.600 63.000 63.400 63.600 ;
        RECT 66.800 63.000 67.600 65.000 ;
        RECT 68.400 62.200 69.200 67.000 ;
        RECT 73.400 65.600 74.000 67.800 ;
        RECT 79.000 67.600 79.800 67.800 ;
        RECT 86.000 67.200 86.800 70.600 ;
        RECT 83.000 66.600 86.800 67.200 ;
        RECT 83.000 66.400 83.800 66.600 ;
        RECT 71.600 64.200 72.400 65.000 ;
        RECT 73.200 64.800 74.000 65.600 ;
        RECT 75.000 65.400 75.800 65.600 ;
        RECT 75.000 64.800 77.800 65.400 ;
        RECT 77.200 64.200 77.800 64.800 ;
        RECT 81.200 64.200 82.000 65.000 ;
        RECT 71.600 63.600 73.600 64.200 ;
        RECT 72.800 62.200 73.600 63.600 ;
        RECT 77.200 62.200 78.000 64.200 ;
        RECT 81.200 63.600 82.600 64.200 ;
        RECT 81.400 62.200 82.600 63.600 ;
        RECT 86.000 62.200 86.800 66.600 ;
        RECT 87.600 64.800 88.400 66.400 ;
        RECT 89.200 62.200 90.000 79.800 ;
        RECT 90.800 66.800 91.600 68.400 ;
        RECT 92.400 66.200 93.200 79.800 ;
        RECT 94.000 71.600 94.800 73.200 ;
        RECT 95.600 71.400 96.400 79.800 ;
        RECT 100.000 76.400 100.800 79.800 ;
        RECT 98.800 75.800 100.800 76.400 ;
        RECT 104.400 75.800 105.200 79.800 ;
        RECT 108.600 75.800 109.800 79.800 ;
        RECT 98.800 75.000 99.600 75.800 ;
        RECT 104.400 75.200 105.000 75.800 ;
        RECT 102.200 74.600 105.800 75.200 ;
        RECT 108.400 75.000 109.200 75.800 ;
        RECT 102.200 74.400 103.000 74.600 ;
        RECT 105.000 74.400 105.800 74.600 ;
        RECT 98.800 73.000 99.600 73.200 ;
        RECT 103.400 73.000 104.200 73.200 ;
        RECT 98.800 72.400 104.200 73.000 ;
        RECT 104.800 73.000 107.000 73.600 ;
        RECT 104.800 71.800 105.400 73.000 ;
        RECT 106.200 72.800 107.000 73.000 ;
        RECT 108.600 73.200 110.000 74.000 ;
        RECT 108.600 72.200 109.200 73.200 ;
        RECT 100.600 71.400 105.400 71.800 ;
        RECT 95.600 71.200 105.400 71.400 ;
        RECT 106.800 71.600 109.200 72.200 ;
        RECT 95.600 71.000 101.400 71.200 ;
        RECT 95.600 70.800 101.200 71.000 ;
        RECT 102.000 70.200 102.800 70.400 ;
        RECT 97.800 69.600 102.800 70.200 ;
        RECT 97.800 69.400 98.600 69.600 ;
        RECT 99.400 68.400 100.200 68.600 ;
        RECT 106.800 68.400 107.400 71.600 ;
        RECT 113.200 71.200 114.000 79.800 ;
        RECT 120.400 73.600 121.200 74.400 ;
        RECT 120.400 72.400 121.000 73.600 ;
        RECT 121.800 72.400 122.600 79.800 ;
        RECT 119.600 71.800 121.000 72.400 ;
        RECT 121.600 71.800 122.600 72.400 ;
        RECT 128.600 72.400 129.400 79.800 ;
        RECT 130.000 73.600 130.800 74.400 ;
        RECT 130.200 72.400 130.800 73.600 ;
        RECT 128.600 71.800 129.600 72.400 ;
        RECT 130.200 71.800 131.600 72.400 ;
        RECT 119.600 71.600 120.400 71.800 ;
        RECT 109.800 70.600 114.000 71.200 ;
        RECT 109.800 70.400 110.600 70.600 ;
        RECT 111.400 69.800 112.200 70.000 ;
        RECT 108.400 69.200 112.200 69.800 ;
        RECT 108.400 69.000 109.200 69.200 ;
        RECT 96.400 67.800 107.400 68.400 ;
        RECT 96.400 67.600 98.000 67.800 ;
        RECT 92.400 65.600 94.200 66.200 ;
        RECT 93.400 64.400 94.200 65.600 ;
        RECT 93.400 63.600 94.800 64.400 ;
        RECT 93.400 62.200 94.200 63.600 ;
        RECT 95.600 62.200 96.400 67.000 ;
        RECT 100.600 65.600 101.200 67.800 ;
        RECT 106.200 67.600 107.000 67.800 ;
        RECT 113.200 67.200 114.000 70.600 ;
        RECT 114.800 70.300 115.600 70.400 ;
        RECT 121.600 70.300 122.200 71.800 ;
        RECT 114.800 69.700 122.200 70.300 ;
        RECT 114.800 69.600 115.600 69.700 ;
        RECT 121.600 68.400 122.200 69.700 ;
        RECT 122.800 68.800 123.600 70.400 ;
        RECT 127.600 68.800 128.400 70.400 ;
        RECT 129.000 68.400 129.600 71.800 ;
        RECT 130.800 71.600 131.600 71.800 ;
        RECT 119.600 67.600 122.200 68.400 ;
        RECT 124.400 68.200 125.200 68.400 ;
        RECT 123.600 67.600 125.200 68.200 ;
        RECT 126.000 68.200 126.800 68.400 ;
        RECT 129.000 68.300 131.600 68.400 ;
        RECT 132.400 68.300 133.200 68.400 ;
        RECT 126.000 67.600 127.600 68.200 ;
        RECT 129.000 67.700 133.200 68.300 ;
        RECT 129.000 67.600 131.600 67.700 ;
        RECT 132.400 67.600 133.200 67.700 ;
        RECT 134.000 68.300 134.800 79.800 ;
        RECT 138.200 72.400 139.000 79.800 ;
        RECT 143.600 75.800 144.400 79.800 ;
        RECT 143.800 75.600 144.400 75.800 ;
        RECT 146.800 75.800 147.600 79.800 ;
        RECT 146.800 75.600 147.400 75.800 ;
        RECT 143.800 75.000 147.400 75.600 ;
        RECT 139.600 73.600 140.400 74.400 ;
        RECT 139.800 72.400 140.400 73.600 ;
        RECT 145.200 72.800 146.000 74.400 ;
        RECT 146.800 72.400 147.400 75.000 ;
        RECT 151.000 72.400 151.800 79.800 ;
        RECT 152.400 73.600 153.200 74.400 ;
        RECT 152.600 72.400 153.200 73.600 ;
        RECT 157.400 72.400 158.200 79.800 ;
        RECT 163.800 78.400 164.600 79.800 ;
        RECT 162.800 77.600 164.600 78.400 ;
        RECT 158.800 73.600 159.600 74.400 ;
        RECT 159.000 72.400 159.600 73.600 ;
        RECT 163.800 72.400 164.600 77.600 ;
        RECT 170.200 74.400 171.000 79.800 ;
        RECT 165.200 73.600 166.000 74.400 ;
        RECT 169.200 73.600 171.000 74.400 ;
        RECT 171.600 73.600 172.400 74.400 ;
        RECT 165.400 72.400 166.000 73.600 ;
        RECT 170.200 72.400 171.000 73.600 ;
        RECT 171.800 72.400 172.400 73.600 ;
        RECT 174.000 72.400 174.800 79.800 ;
        RECT 177.200 72.800 178.000 79.800 ;
        RECT 138.200 71.800 139.200 72.400 ;
        RECT 139.800 71.800 141.200 72.400 ;
        RECT 137.200 68.800 138.000 70.400 ;
        RECT 138.600 70.300 139.200 71.800 ;
        RECT 140.400 71.600 141.200 71.800 ;
        RECT 142.000 70.800 142.800 72.400 ;
        RECT 146.800 71.600 147.600 72.400 ;
        RECT 151.000 71.800 152.000 72.400 ;
        RECT 152.600 71.800 154.000 72.400 ;
        RECT 157.400 71.800 158.400 72.400 ;
        RECT 159.000 71.800 160.400 72.400 ;
        RECT 163.800 71.800 164.800 72.400 ;
        RECT 165.400 71.800 166.800 72.400 ;
        RECT 170.200 71.800 171.200 72.400 ;
        RECT 171.800 71.800 173.200 72.400 ;
        RECT 174.000 71.800 176.600 72.400 ;
        RECT 177.200 71.800 178.200 72.800 ;
        RECT 140.400 70.300 141.200 70.400 ;
        RECT 138.600 69.700 141.200 70.300 ;
        RECT 138.600 68.400 139.200 69.700 ;
        RECT 140.400 69.600 141.200 69.700 ;
        RECT 143.600 69.600 145.200 70.400 ;
        RECT 146.800 68.400 147.400 71.600 ;
        RECT 150.000 68.800 150.800 70.400 ;
        RECT 151.400 68.400 152.000 71.800 ;
        RECT 153.200 71.600 154.000 71.800 ;
        RECT 156.400 68.800 157.200 70.400 ;
        RECT 157.800 68.400 158.400 71.800 ;
        RECT 159.600 71.600 160.400 71.800 ;
        RECT 162.800 68.800 163.600 70.400 ;
        RECT 164.200 68.400 164.800 71.800 ;
        RECT 166.000 71.600 166.800 71.800 ;
        RECT 167.600 70.300 168.400 70.400 ;
        RECT 169.200 70.300 170.000 70.400 ;
        RECT 167.600 69.700 170.000 70.300 ;
        RECT 167.600 69.600 168.400 69.700 ;
        RECT 169.200 68.800 170.000 69.700 ;
        RECT 170.600 68.400 171.200 71.800 ;
        RECT 172.400 71.600 173.200 71.800 ;
        RECT 174.000 69.600 175.000 70.400 ;
        RECT 174.200 68.800 175.000 69.600 ;
        RECT 176.000 69.800 176.600 71.800 ;
        RECT 176.000 69.000 177.000 69.800 ;
        RECT 135.600 68.300 136.400 68.400 ;
        RECT 134.000 68.200 136.400 68.300 ;
        RECT 134.000 67.700 137.200 68.200 ;
        RECT 110.200 66.600 114.000 67.200 ;
        RECT 110.200 66.400 111.000 66.600 ;
        RECT 98.800 64.200 99.600 65.000 ;
        RECT 100.400 64.800 101.200 65.600 ;
        RECT 102.200 65.400 103.000 65.600 ;
        RECT 102.200 64.800 105.000 65.400 ;
        RECT 104.400 64.200 105.000 64.800 ;
        RECT 108.400 64.200 109.200 65.000 ;
        RECT 98.800 63.600 100.800 64.200 ;
        RECT 100.000 62.200 100.800 63.600 ;
        RECT 104.400 62.200 105.200 64.200 ;
        RECT 108.400 63.600 109.800 64.200 ;
        RECT 108.600 62.200 109.800 63.600 ;
        RECT 113.200 62.200 114.000 66.600 ;
        RECT 119.800 66.200 120.400 67.600 ;
        RECT 123.600 67.200 124.400 67.600 ;
        RECT 126.800 67.200 127.600 67.600 ;
        RECT 121.400 66.200 125.000 66.600 ;
        RECT 126.200 66.200 129.800 66.600 ;
        RECT 130.800 66.200 131.400 67.600 ;
        RECT 119.600 62.200 120.400 66.200 ;
        RECT 121.200 66.000 125.200 66.200 ;
        RECT 121.200 62.200 122.000 66.000 ;
        RECT 124.400 62.200 125.200 66.000 ;
        RECT 126.000 66.000 130.000 66.200 ;
        RECT 126.000 62.200 126.800 66.000 ;
        RECT 129.200 62.200 130.000 66.000 ;
        RECT 130.800 62.200 131.600 66.200 ;
        RECT 132.400 64.800 133.200 66.400 ;
        RECT 134.000 62.200 134.800 67.700 ;
        RECT 135.600 67.600 137.200 67.700 ;
        RECT 138.600 67.600 141.200 68.400 ;
        RECT 145.800 68.200 147.400 68.400 ;
        RECT 145.600 67.800 147.400 68.200 ;
        RECT 148.400 68.200 149.200 68.400 ;
        RECT 136.400 67.200 137.200 67.600 ;
        RECT 135.800 66.200 139.400 66.600 ;
        RECT 140.400 66.200 141.000 67.600 ;
        RECT 135.600 66.000 139.600 66.200 ;
        RECT 135.600 62.200 136.400 66.000 ;
        RECT 138.800 62.200 139.600 66.000 ;
        RECT 140.400 62.200 141.200 66.200 ;
        RECT 145.600 62.200 146.400 67.800 ;
        RECT 148.400 67.600 150.000 68.200 ;
        RECT 151.400 67.600 154.000 68.400 ;
        RECT 154.800 68.200 155.600 68.400 ;
        RECT 154.800 67.600 156.400 68.200 ;
        RECT 157.800 67.600 160.400 68.400 ;
        RECT 161.200 68.200 162.000 68.400 ;
        RECT 161.200 67.600 162.800 68.200 ;
        RECT 164.200 67.600 166.800 68.400 ;
        RECT 167.600 68.200 168.400 68.400 ;
        RECT 167.600 67.600 169.200 68.200 ;
        RECT 170.600 67.600 173.200 68.400 ;
        RECT 149.200 67.200 150.000 67.600 ;
        RECT 148.600 66.200 152.200 66.600 ;
        RECT 153.200 66.400 153.800 67.600 ;
        RECT 155.600 67.200 156.400 67.600 ;
        RECT 148.400 66.000 152.400 66.200 ;
        RECT 148.400 62.200 149.200 66.000 ;
        RECT 151.600 62.200 152.400 66.000 ;
        RECT 153.200 62.200 154.000 66.400 ;
        RECT 155.000 66.200 158.600 66.600 ;
        RECT 159.600 66.200 160.200 67.600 ;
        RECT 162.000 67.200 162.800 67.600 ;
        RECT 161.400 66.200 165.000 66.600 ;
        RECT 166.000 66.200 166.600 67.600 ;
        RECT 168.400 67.200 169.200 67.600 ;
        RECT 167.800 66.200 171.400 66.600 ;
        RECT 172.400 66.200 173.000 67.600 ;
        RECT 176.000 67.400 176.600 69.000 ;
        RECT 177.600 68.400 178.200 71.800 ;
        RECT 178.800 70.300 179.600 70.400 ;
        RECT 182.000 70.300 182.800 79.800 ;
        RECT 183.600 71.600 184.400 73.200 ;
        RECT 178.800 69.700 182.800 70.300 ;
        RECT 178.800 69.600 179.600 69.700 ;
        RECT 177.200 67.600 178.200 68.400 ;
        RECT 174.000 66.800 176.600 67.400 ;
        RECT 154.800 66.000 158.800 66.200 ;
        RECT 154.800 62.200 155.600 66.000 ;
        RECT 158.000 62.200 158.800 66.000 ;
        RECT 159.600 62.200 160.400 66.200 ;
        RECT 161.200 66.000 165.200 66.200 ;
        RECT 161.200 62.200 162.000 66.000 ;
        RECT 164.400 62.200 165.200 66.000 ;
        RECT 166.000 62.200 166.800 66.200 ;
        RECT 167.600 66.000 171.600 66.200 ;
        RECT 167.600 62.200 168.400 66.000 ;
        RECT 170.800 62.200 171.600 66.000 ;
        RECT 172.400 62.200 173.200 66.200 ;
        RECT 174.000 62.200 174.800 66.800 ;
        RECT 177.600 66.200 178.200 67.600 ;
        RECT 180.400 66.800 181.200 68.400 ;
        RECT 177.200 65.600 178.200 66.200 ;
        RECT 182.000 66.200 182.800 69.700 ;
        RECT 185.200 66.800 186.000 68.400 ;
        RECT 186.800 66.200 187.600 79.800 ;
        RECT 188.400 72.300 189.200 73.200 ;
        RECT 190.000 72.300 190.800 79.800 ;
        RECT 188.400 71.700 190.800 72.300 ;
        RECT 193.200 72.400 194.000 79.800 ;
        RECT 194.800 72.400 195.600 72.600 ;
        RECT 197.600 72.400 199.200 79.800 ;
        RECT 193.200 71.800 195.600 72.400 ;
        RECT 197.200 71.800 199.200 72.400 ;
        RECT 201.400 72.400 202.200 72.600 ;
        RECT 202.800 72.400 203.600 79.800 ;
        RECT 201.400 71.800 203.600 72.400 ;
        RECT 188.400 71.600 189.200 71.700 ;
        RECT 182.000 65.600 183.800 66.200 ;
        RECT 186.800 65.600 188.600 66.200 ;
        RECT 177.200 62.200 178.000 65.600 ;
        RECT 183.000 64.400 183.800 65.600 ;
        RECT 182.000 63.600 183.800 64.400 ;
        RECT 183.000 62.200 183.800 63.600 ;
        RECT 187.800 62.200 188.600 65.600 ;
        RECT 190.000 62.200 190.800 71.700 ;
        RECT 197.200 70.400 197.800 71.800 ;
        RECT 201.400 71.200 202.000 71.800 ;
        RECT 198.600 70.600 202.000 71.200 ;
        RECT 206.000 71.200 206.800 79.800 ;
        RECT 209.200 71.200 210.000 79.800 ;
        RECT 212.400 71.200 213.200 79.800 ;
        RECT 215.600 71.200 216.400 79.800 ;
        RECT 220.400 72.800 221.200 79.800 ;
        RECT 220.200 71.800 221.200 72.800 ;
        RECT 223.600 72.400 224.400 79.800 ;
        RECT 226.800 72.800 227.600 79.800 ;
        RECT 221.800 71.800 224.400 72.400 ;
        RECT 226.600 71.800 227.600 72.800 ;
        RECT 230.000 72.400 230.800 79.800 ;
        RECT 228.200 71.800 230.800 72.400 ;
        RECT 198.600 70.400 199.400 70.600 ;
        RECT 206.000 70.400 207.800 71.200 ;
        RECT 209.200 70.400 211.400 71.200 ;
        RECT 212.400 70.400 214.600 71.200 ;
        RECT 215.600 70.400 218.000 71.200 ;
        RECT 196.400 69.800 197.800 70.400 ;
        RECT 200.800 69.800 201.600 70.000 ;
        RECT 196.400 69.600 198.200 69.800 ;
        RECT 197.200 69.200 198.200 69.600 ;
        RECT 193.200 67.600 194.800 68.400 ;
        RECT 196.000 67.600 196.800 68.400 ;
        RECT 196.200 67.200 196.800 67.600 ;
        RECT 194.800 66.800 195.600 67.000 ;
        RECT 191.600 64.800 192.400 66.400 ;
        RECT 193.200 66.200 195.600 66.800 ;
        RECT 196.200 66.400 197.000 67.200 ;
        RECT 193.200 62.200 194.000 66.200 ;
        RECT 197.600 65.800 198.200 69.200 ;
        RECT 199.000 69.200 201.600 69.800 ;
        RECT 199.000 68.600 199.600 69.200 ;
        RECT 207.000 69.000 207.800 70.400 ;
        RECT 210.600 69.000 211.400 70.400 ;
        RECT 213.800 69.000 214.600 70.400 ;
        RECT 198.800 67.800 199.600 68.600 ;
        RECT 202.000 68.200 203.600 68.400 ;
        RECT 200.200 67.600 203.600 68.200 ;
        RECT 204.400 68.200 206.200 69.000 ;
        RECT 207.000 68.200 209.600 69.000 ;
        RECT 210.600 68.200 213.000 69.000 ;
        RECT 213.800 68.200 216.400 69.000 ;
        RECT 204.400 67.600 205.200 68.200 ;
        RECT 207.000 67.600 207.800 68.200 ;
        RECT 210.600 67.600 211.400 68.200 ;
        RECT 213.800 67.600 214.600 68.200 ;
        RECT 217.200 67.600 218.000 70.400 ;
        RECT 200.200 67.200 200.800 67.600 ;
        RECT 198.800 66.600 200.800 67.200 ;
        RECT 201.400 66.800 202.200 67.000 ;
        RECT 206.000 66.800 207.800 67.600 ;
        RECT 209.200 66.800 211.400 67.600 ;
        RECT 212.400 66.800 214.600 67.600 ;
        RECT 215.600 66.800 218.000 67.600 ;
        RECT 220.200 68.400 220.800 71.800 ;
        RECT 221.800 69.800 222.400 71.800 ;
        RECT 221.400 69.000 222.400 69.800 ;
        RECT 220.200 67.600 221.200 68.400 ;
        RECT 198.800 66.400 200.400 66.600 ;
        RECT 201.400 66.200 203.600 66.800 ;
        RECT 197.600 64.400 199.200 65.800 ;
        RECT 196.400 63.600 199.200 64.400 ;
        RECT 197.600 62.200 199.200 63.600 ;
        RECT 202.800 62.200 203.600 66.200 ;
        RECT 206.000 62.200 206.800 66.800 ;
        RECT 209.200 62.200 210.000 66.800 ;
        RECT 212.400 62.200 213.200 66.800 ;
        RECT 215.600 62.200 216.400 66.800 ;
        RECT 220.200 66.200 220.800 67.600 ;
        RECT 221.800 67.400 222.400 69.000 ;
        RECT 223.400 69.600 224.400 70.400 ;
        RECT 223.400 68.800 224.200 69.600 ;
        RECT 226.600 68.400 227.200 71.800 ;
        RECT 228.200 69.800 228.800 71.800 ;
        RECT 231.600 71.600 232.400 73.200 ;
        RECT 227.800 69.000 228.800 69.800 ;
        RECT 226.600 67.600 227.600 68.400 ;
        RECT 221.800 66.800 224.400 67.400 ;
        RECT 220.200 65.600 221.200 66.200 ;
        RECT 220.400 62.200 221.200 65.600 ;
        RECT 223.600 62.200 224.400 66.800 ;
        RECT 226.600 66.400 227.200 67.600 ;
        RECT 228.200 67.400 228.800 69.000 ;
        RECT 229.800 69.600 230.800 70.400 ;
        RECT 229.800 68.800 230.600 69.600 ;
        RECT 228.200 66.800 230.800 67.400 ;
        RECT 226.600 65.600 227.600 66.400 ;
        RECT 226.800 62.200 227.600 65.600 ;
        RECT 230.000 62.200 230.800 66.800 ;
        RECT 233.200 66.200 234.000 79.800 ;
        RECT 238.000 76.400 238.800 79.800 ;
        RECT 237.800 75.800 238.800 76.400 ;
        RECT 237.800 75.200 238.400 75.800 ;
        RECT 241.200 75.200 242.000 79.800 ;
        RECT 244.400 77.000 245.200 79.800 ;
        RECT 246.000 77.000 246.800 79.800 ;
        RECT 236.400 74.600 238.400 75.200 ;
        RECT 236.400 69.000 237.200 74.600 ;
        RECT 239.000 74.400 243.200 75.200 ;
        RECT 247.600 75.000 248.400 79.800 ;
        RECT 250.800 75.000 251.600 79.800 ;
        RECT 239.000 74.000 239.600 74.400 ;
        RECT 238.000 73.200 239.600 74.000 ;
        RECT 242.600 73.800 248.400 74.400 ;
        RECT 240.600 73.200 242.000 73.800 ;
        RECT 240.600 73.000 246.800 73.200 ;
        RECT 241.400 72.600 246.800 73.000 ;
        RECT 246.000 72.400 246.800 72.600 ;
        RECT 247.800 73.000 248.400 73.800 ;
        RECT 249.000 73.600 251.600 74.400 ;
        RECT 254.000 73.600 254.800 79.800 ;
        RECT 255.600 77.000 256.400 79.800 ;
        RECT 257.200 77.000 258.000 79.800 ;
        RECT 258.800 77.000 259.600 79.800 ;
        RECT 257.200 74.400 261.400 75.200 ;
        RECT 262.000 74.400 262.800 79.800 ;
        RECT 265.200 75.200 266.000 79.800 ;
        RECT 265.200 74.600 267.800 75.200 ;
        RECT 262.000 73.600 264.600 74.400 ;
        RECT 255.600 73.000 256.400 73.200 ;
        RECT 247.800 72.400 256.400 73.000 ;
        RECT 258.800 73.000 259.600 73.200 ;
        RECT 267.200 73.000 267.800 74.600 ;
        RECT 258.800 72.400 267.800 73.000 ;
        RECT 267.200 70.600 267.800 72.400 ;
        RECT 268.400 72.000 269.200 79.800 ;
        RECT 268.400 71.200 269.400 72.000 ;
        RECT 278.000 71.200 278.800 79.800 ;
        RECT 281.200 71.200 282.000 79.800 ;
        RECT 284.400 71.200 285.200 79.800 ;
        RECT 287.600 71.200 288.400 79.800 ;
        RECT 290.800 71.600 291.600 73.200 ;
        RECT 237.800 70.000 261.200 70.600 ;
        RECT 267.200 70.000 268.000 70.600 ;
        RECT 237.800 69.800 238.600 70.000 ;
        RECT 239.600 69.600 240.400 70.000 ;
        RECT 242.800 69.600 243.600 70.000 ;
        RECT 260.400 69.400 261.200 70.000 ;
        RECT 234.800 66.800 235.600 68.400 ;
        RECT 236.400 68.200 245.200 69.000 ;
        RECT 245.800 68.600 247.800 69.400 ;
        RECT 251.600 68.600 254.800 69.400 ;
        RECT 232.200 65.600 234.000 66.200 ;
        RECT 232.200 64.400 233.000 65.600 ;
        RECT 231.600 63.600 233.000 64.400 ;
        RECT 232.200 62.200 233.000 63.600 ;
        RECT 236.400 62.200 237.200 68.200 ;
        RECT 238.800 66.800 241.800 67.600 ;
        RECT 241.000 66.200 241.800 66.800 ;
        RECT 247.000 66.200 247.800 68.600 ;
        RECT 249.200 66.800 250.000 68.400 ;
        RECT 254.400 67.800 255.200 68.000 ;
        RECT 250.800 67.200 255.200 67.800 ;
        RECT 250.800 67.000 251.600 67.200 ;
        RECT 257.200 66.400 258.000 69.200 ;
        RECT 263.000 68.600 266.800 69.400 ;
        RECT 263.000 67.400 263.800 68.600 ;
        RECT 267.400 68.000 268.000 70.000 ;
        RECT 250.800 66.200 251.600 66.400 ;
        RECT 241.000 65.400 243.600 66.200 ;
        RECT 247.000 65.600 251.600 66.200 ;
        RECT 252.400 65.600 254.000 66.400 ;
        RECT 257.000 65.600 258.000 66.400 ;
        RECT 262.000 66.800 263.800 67.400 ;
        RECT 266.800 67.400 268.000 68.000 ;
        RECT 262.000 66.200 262.800 66.800 ;
        RECT 242.800 62.200 243.600 65.400 ;
        RECT 260.400 65.400 262.800 66.200 ;
        RECT 244.400 62.200 245.200 65.000 ;
        RECT 246.000 62.200 246.800 65.000 ;
        RECT 247.600 62.200 248.400 65.000 ;
        RECT 250.800 62.200 251.600 65.000 ;
        RECT 254.000 62.200 254.800 65.000 ;
        RECT 255.600 62.200 256.400 65.000 ;
        RECT 257.200 62.200 258.000 65.000 ;
        RECT 258.800 62.200 259.600 65.000 ;
        RECT 260.400 62.200 261.200 65.400 ;
        RECT 266.800 62.200 267.600 67.400 ;
        RECT 268.600 66.800 269.400 71.200 ;
        RECT 276.400 70.400 278.800 71.200 ;
        RECT 279.800 70.400 282.000 71.200 ;
        RECT 283.000 70.400 285.200 71.200 ;
        RECT 286.600 70.400 288.400 71.200 ;
        RECT 276.400 67.600 277.200 70.400 ;
        RECT 279.800 69.000 280.600 70.400 ;
        RECT 283.000 69.000 283.800 70.400 ;
        RECT 286.600 69.000 287.400 70.400 ;
        RECT 278.000 68.200 280.600 69.000 ;
        RECT 281.400 68.200 283.800 69.000 ;
        RECT 284.800 68.200 287.400 69.000 ;
        RECT 288.200 68.200 290.000 69.000 ;
        RECT 279.800 67.600 280.600 68.200 ;
        RECT 283.000 67.600 283.800 68.200 ;
        RECT 286.600 67.600 287.400 68.200 ;
        RECT 289.200 67.600 290.000 68.200 ;
        RECT 276.400 66.800 278.800 67.600 ;
        RECT 279.800 66.800 282.000 67.600 ;
        RECT 283.000 66.800 285.200 67.600 ;
        RECT 286.600 66.800 288.400 67.600 ;
        RECT 268.400 66.000 269.400 66.800 ;
        RECT 268.400 62.200 269.200 66.000 ;
        RECT 278.000 62.200 278.800 66.800 ;
        RECT 281.200 62.200 282.000 66.800 ;
        RECT 284.400 62.200 285.200 66.800 ;
        RECT 287.600 62.200 288.400 66.800 ;
        RECT 292.400 66.200 293.200 79.800 ;
        RECT 298.200 72.400 299.000 79.800 ;
        RECT 303.600 76.400 304.400 79.800 ;
        RECT 303.400 75.800 304.400 76.400 ;
        RECT 303.400 75.200 304.000 75.800 ;
        RECT 306.800 75.200 307.600 79.800 ;
        RECT 310.000 77.000 310.800 79.800 ;
        RECT 311.600 77.000 312.400 79.800 ;
        RECT 302.000 74.600 304.000 75.200 ;
        RECT 299.600 73.600 301.200 74.400 ;
        RECT 299.800 72.400 300.400 73.600 ;
        RECT 298.200 71.800 299.200 72.400 ;
        RECT 299.800 71.800 301.200 72.400 ;
        RECT 298.600 70.400 299.200 71.800 ;
        RECT 300.400 71.600 301.200 71.800 ;
        RECT 297.200 68.800 298.000 70.400 ;
        RECT 298.600 69.600 299.600 70.400 ;
        RECT 298.600 68.400 299.200 69.600 ;
        RECT 302.000 69.000 302.800 74.600 ;
        RECT 304.600 74.400 308.800 75.200 ;
        RECT 313.200 75.000 314.000 79.800 ;
        RECT 316.400 75.000 317.200 79.800 ;
        RECT 304.600 74.000 305.200 74.400 ;
        RECT 303.600 73.200 305.200 74.000 ;
        RECT 308.200 73.800 314.000 74.400 ;
        RECT 306.200 73.200 307.600 73.800 ;
        RECT 306.200 73.000 312.400 73.200 ;
        RECT 307.000 72.600 312.400 73.000 ;
        RECT 311.600 72.400 312.400 72.600 ;
        RECT 313.400 73.000 314.000 73.800 ;
        RECT 314.600 73.600 317.200 74.400 ;
        RECT 319.600 73.600 320.400 79.800 ;
        RECT 321.200 77.000 322.000 79.800 ;
        RECT 322.800 77.000 323.600 79.800 ;
        RECT 324.400 77.000 325.200 79.800 ;
        RECT 322.800 74.400 327.000 75.200 ;
        RECT 327.600 74.400 328.400 79.800 ;
        RECT 330.800 75.200 331.600 79.800 ;
        RECT 330.800 74.600 333.400 75.200 ;
        RECT 327.600 73.600 330.200 74.400 ;
        RECT 321.200 73.000 322.000 73.200 ;
        RECT 313.400 72.400 322.000 73.000 ;
        RECT 324.400 73.000 325.200 73.200 ;
        RECT 332.800 73.000 333.400 74.600 ;
        RECT 324.400 72.400 333.400 73.000 ;
        RECT 332.800 70.600 333.400 72.400 ;
        RECT 334.000 72.000 334.800 79.800 ;
        RECT 338.800 76.400 339.600 79.800 ;
        RECT 338.600 75.800 339.600 76.400 ;
        RECT 338.600 75.200 339.200 75.800 ;
        RECT 342.000 75.200 342.800 79.800 ;
        RECT 345.200 77.000 346.000 79.800 ;
        RECT 346.800 77.000 347.600 79.800 ;
        RECT 337.200 74.600 339.200 75.200 ;
        RECT 334.000 71.200 335.000 72.000 ;
        RECT 303.400 70.000 326.800 70.600 ;
        RECT 332.800 70.000 333.600 70.600 ;
        RECT 303.400 69.800 304.200 70.000 ;
        RECT 305.200 69.600 306.000 70.000 ;
        RECT 308.400 69.600 309.200 70.000 ;
        RECT 326.000 69.400 326.800 70.000 ;
        RECT 294.000 66.800 294.800 68.400 ;
        RECT 295.600 68.200 296.400 68.400 ;
        RECT 295.600 67.600 297.200 68.200 ;
        RECT 298.600 67.600 301.200 68.400 ;
        RECT 302.000 68.200 310.800 69.000 ;
        RECT 311.400 68.600 313.400 69.400 ;
        RECT 317.200 68.600 320.400 69.400 ;
        RECT 296.400 67.200 297.200 67.600 ;
        RECT 295.800 66.200 299.400 66.600 ;
        RECT 300.400 66.200 301.000 67.600 ;
        RECT 291.400 65.600 293.200 66.200 ;
        RECT 295.600 66.000 299.600 66.200 ;
        RECT 291.400 62.200 292.200 65.600 ;
        RECT 295.600 62.200 296.400 66.000 ;
        RECT 298.800 62.200 299.600 66.000 ;
        RECT 300.400 62.200 301.200 66.200 ;
        RECT 302.000 62.200 302.800 68.200 ;
        RECT 304.400 66.800 307.400 67.600 ;
        RECT 306.600 66.200 307.400 66.800 ;
        RECT 312.600 66.200 313.400 68.600 ;
        RECT 314.800 66.800 315.600 68.400 ;
        RECT 320.000 67.800 320.800 68.000 ;
        RECT 316.400 67.200 320.800 67.800 ;
        RECT 316.400 67.000 317.200 67.200 ;
        RECT 322.800 66.400 323.600 69.200 ;
        RECT 328.600 68.600 332.400 69.400 ;
        RECT 328.600 67.400 329.400 68.600 ;
        RECT 333.000 68.000 333.600 70.000 ;
        RECT 316.400 66.200 317.200 66.400 ;
        RECT 306.600 65.400 309.200 66.200 ;
        RECT 312.600 65.600 317.200 66.200 ;
        RECT 318.000 65.600 319.600 66.400 ;
        RECT 322.600 65.600 323.600 66.400 ;
        RECT 327.600 66.800 329.400 67.400 ;
        RECT 332.400 67.400 333.600 68.000 ;
        RECT 327.600 66.200 328.400 66.800 ;
        RECT 308.400 62.200 309.200 65.400 ;
        RECT 326.000 65.400 328.400 66.200 ;
        RECT 310.000 62.200 310.800 65.000 ;
        RECT 311.600 62.200 312.400 65.000 ;
        RECT 313.200 62.200 314.000 65.000 ;
        RECT 316.400 62.200 317.200 65.000 ;
        RECT 319.600 62.200 320.400 65.000 ;
        RECT 321.200 62.200 322.000 65.000 ;
        RECT 322.800 62.200 323.600 65.000 ;
        RECT 324.400 62.200 325.200 65.000 ;
        RECT 326.000 62.200 326.800 65.400 ;
        RECT 332.400 62.200 333.200 67.400 ;
        RECT 334.200 66.800 335.000 71.200 ;
        RECT 334.000 66.000 335.000 66.800 ;
        RECT 337.200 69.000 338.000 74.600 ;
        RECT 339.800 74.400 344.000 75.200 ;
        RECT 348.400 75.000 349.200 79.800 ;
        RECT 351.600 75.000 352.400 79.800 ;
        RECT 339.800 74.000 340.400 74.400 ;
        RECT 338.800 73.200 340.400 74.000 ;
        RECT 343.400 73.800 349.200 74.400 ;
        RECT 341.400 73.200 342.800 73.800 ;
        RECT 341.400 73.000 347.600 73.200 ;
        RECT 342.200 72.600 347.600 73.000 ;
        RECT 346.800 72.400 347.600 72.600 ;
        RECT 348.600 73.000 349.200 73.800 ;
        RECT 349.800 73.600 352.400 74.400 ;
        RECT 354.800 73.600 355.600 79.800 ;
        RECT 356.400 77.000 357.200 79.800 ;
        RECT 358.000 77.000 358.800 79.800 ;
        RECT 359.600 77.000 360.400 79.800 ;
        RECT 358.000 74.400 362.200 75.200 ;
        RECT 362.800 74.400 363.600 79.800 ;
        RECT 366.000 75.200 366.800 79.800 ;
        RECT 366.000 74.600 368.600 75.200 ;
        RECT 362.800 73.600 365.400 74.400 ;
        RECT 356.400 73.000 357.200 73.200 ;
        RECT 348.600 72.400 357.200 73.000 ;
        RECT 359.600 73.000 360.400 73.200 ;
        RECT 368.000 73.000 368.600 74.600 ;
        RECT 359.600 72.400 368.600 73.000 ;
        RECT 368.000 70.600 368.600 72.400 ;
        RECT 369.200 72.000 370.000 79.800 ;
        RECT 369.200 71.200 370.200 72.000 ;
        RECT 338.600 70.000 362.000 70.600 ;
        RECT 368.000 70.000 368.800 70.600 ;
        RECT 338.600 69.800 339.400 70.000 ;
        RECT 343.600 69.600 344.400 70.000 ;
        RECT 361.200 69.400 362.000 70.000 ;
        RECT 337.200 68.200 346.000 69.000 ;
        RECT 346.600 68.600 348.600 69.400 ;
        RECT 352.400 68.600 355.600 69.400 ;
        RECT 334.000 62.200 334.800 66.000 ;
        RECT 337.200 62.200 338.000 68.200 ;
        RECT 339.600 66.800 342.600 67.600 ;
        RECT 341.800 66.200 342.600 66.800 ;
        RECT 347.800 66.200 348.600 68.600 ;
        RECT 350.000 66.800 350.800 68.400 ;
        RECT 355.200 67.800 356.000 68.000 ;
        RECT 351.600 67.200 356.000 67.800 ;
        RECT 351.600 67.000 352.400 67.200 ;
        RECT 358.000 66.400 358.800 69.200 ;
        RECT 363.800 68.600 367.600 69.400 ;
        RECT 363.800 67.400 364.600 68.600 ;
        RECT 368.200 68.000 368.800 70.000 ;
        RECT 351.600 66.200 352.400 66.400 ;
        RECT 341.800 65.400 344.400 66.200 ;
        RECT 347.800 65.600 352.400 66.200 ;
        RECT 353.200 65.600 354.800 66.400 ;
        RECT 357.800 65.600 358.800 66.400 ;
        RECT 362.800 66.800 364.600 67.400 ;
        RECT 367.600 67.400 368.800 68.000 ;
        RECT 362.800 66.200 363.600 66.800 ;
        RECT 343.600 62.200 344.400 65.400 ;
        RECT 361.200 65.400 363.600 66.200 ;
        RECT 345.200 62.200 346.000 65.000 ;
        RECT 346.800 62.200 347.600 65.000 ;
        RECT 348.400 62.200 349.200 65.000 ;
        RECT 351.600 62.200 352.400 65.000 ;
        RECT 354.800 62.200 355.600 65.000 ;
        RECT 356.400 62.200 357.200 65.000 ;
        RECT 358.000 62.200 358.800 65.000 ;
        RECT 359.600 62.200 360.400 65.000 ;
        RECT 361.200 62.200 362.000 65.400 ;
        RECT 367.600 62.200 368.400 67.400 ;
        RECT 369.400 66.800 370.200 71.200 ;
        RECT 374.000 71.200 374.800 79.800 ;
        RECT 377.200 71.200 378.000 79.800 ;
        RECT 380.400 71.200 381.200 79.800 ;
        RECT 383.600 71.200 384.400 79.800 ;
        RECT 374.000 70.400 375.800 71.200 ;
        RECT 377.200 70.400 379.400 71.200 ;
        RECT 380.400 70.400 382.600 71.200 ;
        RECT 383.600 70.400 386.000 71.200 ;
        RECT 375.000 69.000 375.800 70.400 ;
        RECT 378.600 69.000 379.400 70.400 ;
        RECT 381.800 69.000 382.600 70.400 ;
        RECT 372.400 68.200 374.200 69.000 ;
        RECT 375.000 68.200 377.600 69.000 ;
        RECT 378.600 68.200 381.000 69.000 ;
        RECT 381.800 68.200 384.400 69.000 ;
        RECT 372.400 67.600 373.200 68.200 ;
        RECT 375.000 67.600 375.800 68.200 ;
        RECT 378.600 67.600 379.400 68.200 ;
        RECT 381.800 67.600 382.600 68.200 ;
        RECT 385.200 67.600 386.000 70.400 ;
        RECT 369.200 66.000 370.200 66.800 ;
        RECT 374.000 66.800 375.800 67.600 ;
        RECT 377.200 66.800 379.400 67.600 ;
        RECT 380.400 66.800 382.600 67.600 ;
        RECT 383.600 66.800 386.000 67.600 ;
        RECT 388.400 70.300 389.200 79.800 ;
        RECT 392.600 72.400 393.400 79.800 ;
        RECT 394.000 73.600 394.800 74.400 ;
        RECT 394.200 72.400 394.800 73.600 ;
        RECT 392.600 71.800 393.600 72.400 ;
        RECT 394.200 71.800 395.600 72.400 ;
        RECT 391.600 70.300 392.400 70.400 ;
        RECT 388.400 69.700 392.400 70.300 ;
        RECT 369.200 62.200 370.000 66.000 ;
        RECT 374.000 62.200 374.800 66.800 ;
        RECT 377.200 62.200 378.000 66.800 ;
        RECT 380.400 62.200 381.200 66.800 ;
        RECT 383.600 62.200 384.400 66.800 ;
        RECT 386.800 64.800 387.600 66.400 ;
        RECT 388.400 62.200 389.200 69.700 ;
        RECT 391.600 68.800 392.400 69.700 ;
        RECT 393.000 68.400 393.600 71.800 ;
        RECT 394.800 71.600 395.600 71.800 ;
        RECT 396.400 71.600 397.200 73.200 ;
        RECT 394.900 70.300 395.500 71.600 ;
        RECT 398.000 70.300 398.800 79.800 ;
        RECT 394.900 69.700 398.800 70.300 ;
        RECT 390.000 68.200 390.800 68.400 ;
        RECT 390.000 67.600 391.600 68.200 ;
        RECT 393.000 67.600 395.600 68.400 ;
        RECT 390.800 67.200 391.600 67.600 ;
        RECT 390.200 66.200 393.800 66.600 ;
        RECT 394.800 66.200 395.400 67.600 ;
        RECT 398.000 66.200 398.800 69.700 ;
        RECT 399.600 68.300 400.400 68.400 ;
        RECT 401.200 68.300 402.000 68.400 ;
        RECT 399.600 67.700 402.000 68.300 ;
        RECT 399.600 66.800 400.400 67.700 ;
        RECT 401.200 66.800 402.000 67.700 ;
        RECT 390.000 66.000 394.000 66.200 ;
        RECT 390.000 62.200 390.800 66.000 ;
        RECT 393.200 62.200 394.000 66.000 ;
        RECT 394.800 62.200 395.600 66.200 ;
        RECT 397.000 65.600 398.800 66.200 ;
        RECT 402.800 66.200 403.600 79.800 ;
        RECT 412.400 74.300 413.200 79.800 ;
        RECT 415.600 75.200 416.400 79.800 ;
        RECT 404.400 73.700 413.200 74.300 ;
        RECT 404.400 71.600 405.200 73.700 ;
        RECT 412.400 72.000 413.200 73.700 ;
        RECT 412.200 71.200 413.200 72.000 ;
        RECT 413.800 74.600 416.400 75.200 ;
        RECT 413.800 73.000 414.400 74.600 ;
        RECT 418.800 74.400 419.600 79.800 ;
        RECT 422.000 77.000 422.800 79.800 ;
        RECT 423.600 77.000 424.400 79.800 ;
        RECT 425.200 77.000 426.000 79.800 ;
        RECT 420.200 74.400 424.400 75.200 ;
        RECT 417.000 73.600 419.600 74.400 ;
        RECT 426.800 73.600 427.600 79.800 ;
        RECT 430.000 75.000 430.800 79.800 ;
        RECT 433.200 75.000 434.000 79.800 ;
        RECT 434.800 77.000 435.600 79.800 ;
        RECT 436.400 77.000 437.200 79.800 ;
        RECT 439.600 75.200 440.400 79.800 ;
        RECT 442.800 76.400 443.600 79.800 ;
        RECT 442.800 75.800 443.800 76.400 ;
        RECT 443.200 75.200 443.800 75.800 ;
        RECT 438.400 74.400 442.600 75.200 ;
        RECT 443.200 74.600 445.200 75.200 ;
        RECT 430.000 73.600 432.600 74.400 ;
        RECT 433.200 73.800 439.000 74.400 ;
        RECT 442.000 74.000 442.600 74.400 ;
        RECT 422.000 73.000 422.800 73.200 ;
        RECT 413.800 72.400 422.800 73.000 ;
        RECT 425.200 73.000 426.000 73.200 ;
        RECT 433.200 73.000 433.800 73.800 ;
        RECT 439.600 73.200 441.000 73.800 ;
        RECT 442.000 73.200 443.600 74.000 ;
        RECT 425.200 72.400 433.800 73.000 ;
        RECT 434.800 73.000 441.000 73.200 ;
        RECT 434.800 72.600 440.200 73.000 ;
        RECT 434.800 72.400 435.600 72.600 ;
        RECT 412.200 66.800 413.000 71.200 ;
        RECT 413.800 70.600 414.400 72.400 ;
        RECT 413.600 70.000 414.400 70.600 ;
        RECT 420.400 70.000 443.800 70.600 ;
        RECT 413.600 68.000 414.200 70.000 ;
        RECT 420.400 69.400 421.200 70.000 ;
        RECT 438.000 69.600 438.800 70.000 ;
        RECT 439.600 69.600 440.400 70.000 ;
        RECT 443.000 69.800 443.800 70.000 ;
        RECT 414.800 68.600 418.600 69.400 ;
        RECT 413.600 67.400 414.800 68.000 ;
        RECT 402.800 65.600 404.600 66.200 ;
        RECT 412.200 66.000 413.200 66.800 ;
        RECT 397.000 62.200 397.800 65.600 ;
        RECT 403.800 64.300 404.600 65.600 ;
        RECT 407.600 64.300 408.400 64.400 ;
        RECT 403.800 63.700 408.400 64.300 ;
        RECT 403.800 62.200 404.600 63.700 ;
        RECT 407.600 63.600 408.400 63.700 ;
        RECT 412.400 62.200 413.200 66.000 ;
        RECT 414.000 62.200 414.800 67.400 ;
        RECT 417.800 67.400 418.600 68.600 ;
        RECT 417.800 66.800 419.600 67.400 ;
        RECT 418.800 66.200 419.600 66.800 ;
        RECT 423.600 66.400 424.400 69.200 ;
        RECT 426.800 68.600 430.000 69.400 ;
        RECT 433.800 68.600 435.800 69.400 ;
        RECT 444.400 69.000 445.200 74.600 ;
        RECT 446.000 71.600 446.800 73.200 ;
        RECT 426.400 67.800 427.200 68.000 ;
        RECT 426.400 67.200 430.800 67.800 ;
        RECT 430.000 67.000 430.800 67.200 ;
        RECT 431.600 66.800 432.400 68.400 ;
        RECT 418.800 65.400 421.200 66.200 ;
        RECT 423.600 65.600 424.600 66.400 ;
        RECT 427.600 65.600 429.200 66.400 ;
        RECT 430.000 66.200 430.800 66.400 ;
        RECT 433.800 66.200 434.600 68.600 ;
        RECT 436.400 68.200 445.200 69.000 ;
        RECT 439.800 66.800 442.800 67.600 ;
        RECT 439.800 66.200 440.600 66.800 ;
        RECT 430.000 65.600 434.600 66.200 ;
        RECT 420.400 62.200 421.200 65.400 ;
        RECT 438.000 65.400 440.600 66.200 ;
        RECT 422.000 62.200 422.800 65.000 ;
        RECT 423.600 62.200 424.400 65.000 ;
        RECT 425.200 62.200 426.000 65.000 ;
        RECT 426.800 62.200 427.600 65.000 ;
        RECT 430.000 62.200 430.800 65.000 ;
        RECT 433.200 62.200 434.000 65.000 ;
        RECT 434.800 62.200 435.600 65.000 ;
        RECT 436.400 62.200 437.200 65.000 ;
        RECT 438.000 62.200 438.800 65.400 ;
        RECT 444.400 62.200 445.200 68.200 ;
        RECT 447.600 66.200 448.400 79.800 ;
        RECT 451.600 73.600 452.400 74.400 ;
        RECT 451.600 72.400 452.200 73.600 ;
        RECT 453.000 72.400 453.800 79.800 ;
        RECT 450.800 71.800 452.200 72.400 ;
        RECT 452.800 71.800 453.800 72.400 ;
        RECT 450.800 71.600 451.600 71.800 ;
        RECT 452.800 68.400 453.400 71.800 ;
        RECT 458.800 71.200 459.600 79.800 ;
        RECT 462.000 71.200 462.800 79.800 ;
        RECT 466.800 76.400 467.600 79.800 ;
        RECT 466.600 75.800 467.600 76.400 ;
        RECT 466.600 75.200 467.200 75.800 ;
        RECT 470.000 75.200 470.800 79.800 ;
        RECT 473.200 77.000 474.000 79.800 ;
        RECT 474.800 77.000 475.600 79.800 ;
        RECT 458.800 70.400 462.800 71.200 ;
        RECT 465.200 74.600 467.200 75.200 ;
        RECT 454.000 68.800 454.800 70.400 ;
        RECT 449.200 66.800 450.000 68.400 ;
        RECT 450.800 67.600 453.400 68.400 ;
        RECT 455.600 68.300 456.400 68.400 ;
        RECT 457.200 68.300 458.000 68.400 ;
        RECT 455.600 68.200 458.000 68.300 ;
        RECT 454.800 67.700 458.000 68.200 ;
        RECT 454.800 67.600 456.400 67.700 ;
        RECT 457.200 67.600 458.000 67.700 ;
        RECT 458.800 67.600 459.600 70.400 ;
        RECT 465.200 69.000 466.000 74.600 ;
        RECT 467.800 74.400 472.000 75.200 ;
        RECT 476.400 75.000 477.200 79.800 ;
        RECT 479.600 75.000 480.400 79.800 ;
        RECT 467.800 74.000 468.400 74.400 ;
        RECT 466.800 73.200 468.400 74.000 ;
        RECT 471.400 73.800 477.200 74.400 ;
        RECT 469.400 73.200 470.800 73.800 ;
        RECT 469.400 73.000 475.600 73.200 ;
        RECT 470.200 72.600 475.600 73.000 ;
        RECT 474.800 72.400 475.600 72.600 ;
        RECT 476.600 73.000 477.200 73.800 ;
        RECT 477.800 73.600 480.400 74.400 ;
        RECT 482.800 73.600 483.600 79.800 ;
        RECT 484.400 77.000 485.200 79.800 ;
        RECT 486.000 77.000 486.800 79.800 ;
        RECT 487.600 77.000 488.400 79.800 ;
        RECT 486.000 74.400 490.200 75.200 ;
        RECT 490.800 74.400 491.600 79.800 ;
        RECT 494.000 75.200 494.800 79.800 ;
        RECT 494.000 74.600 496.600 75.200 ;
        RECT 490.800 73.600 493.400 74.400 ;
        RECT 484.400 73.000 485.200 73.200 ;
        RECT 476.600 72.400 485.200 73.000 ;
        RECT 487.600 73.000 488.400 73.200 ;
        RECT 496.000 73.000 496.600 74.600 ;
        RECT 487.600 72.400 496.600 73.000 ;
        RECT 496.000 70.600 496.600 72.400 ;
        RECT 497.200 72.000 498.000 79.800 ;
        RECT 497.200 71.200 498.200 72.000 ;
        RECT 466.600 70.000 490.000 70.600 ;
        RECT 496.000 70.000 496.800 70.600 ;
        RECT 466.600 69.800 467.400 70.000 ;
        RECT 468.400 69.600 469.200 70.000 ;
        RECT 471.600 69.600 472.400 70.000 ;
        RECT 489.200 69.400 490.000 70.000 ;
        RECT 465.200 68.200 474.000 69.000 ;
        RECT 474.600 68.600 476.600 69.400 ;
        RECT 480.400 68.600 483.600 69.400 ;
        RECT 451.000 66.200 451.600 67.600 ;
        RECT 454.800 67.200 455.600 67.600 ;
        RECT 458.800 66.800 462.800 67.600 ;
        RECT 452.600 66.200 456.200 66.600 ;
        RECT 446.600 65.600 448.400 66.200 ;
        RECT 446.600 64.400 447.400 65.600 ;
        RECT 446.000 63.600 447.400 64.400 ;
        RECT 446.600 62.200 447.400 63.600 ;
        RECT 450.800 62.200 451.600 66.200 ;
        RECT 452.400 66.000 456.400 66.200 ;
        RECT 452.400 62.200 453.200 66.000 ;
        RECT 455.600 62.200 456.400 66.000 ;
        RECT 458.800 62.200 459.600 66.800 ;
        RECT 462.000 62.200 462.800 66.800 ;
        RECT 465.200 62.200 466.000 68.200 ;
        RECT 467.600 66.800 470.600 67.600 ;
        RECT 469.800 66.200 470.600 66.800 ;
        RECT 475.800 66.200 476.600 68.600 ;
        RECT 478.000 66.800 478.800 68.400 ;
        RECT 483.200 67.800 484.000 68.000 ;
        RECT 479.600 67.200 484.000 67.800 ;
        RECT 479.600 67.000 480.400 67.200 ;
        RECT 486.000 66.400 486.800 69.200 ;
        RECT 491.800 68.600 495.600 69.400 ;
        RECT 491.800 67.400 492.600 68.600 ;
        RECT 496.200 68.000 496.800 70.000 ;
        RECT 479.600 66.200 480.400 66.400 ;
        RECT 469.800 65.400 472.400 66.200 ;
        RECT 475.800 65.600 480.400 66.200 ;
        RECT 481.200 65.600 482.800 66.400 ;
        RECT 485.800 65.600 486.800 66.400 ;
        RECT 490.800 66.800 492.600 67.400 ;
        RECT 495.600 67.400 496.800 68.000 ;
        RECT 490.800 66.200 491.600 66.800 ;
        RECT 471.600 62.200 472.400 65.400 ;
        RECT 489.200 65.400 491.600 66.200 ;
        RECT 473.200 62.200 474.000 65.000 ;
        RECT 474.800 62.200 475.600 65.000 ;
        RECT 476.400 62.200 477.200 65.000 ;
        RECT 479.600 62.200 480.400 65.000 ;
        RECT 482.800 62.200 483.600 65.000 ;
        RECT 484.400 62.200 485.200 65.000 ;
        RECT 486.000 62.200 486.800 65.000 ;
        RECT 487.600 62.200 488.400 65.000 ;
        RECT 489.200 62.200 490.000 65.400 ;
        RECT 495.600 62.200 496.400 67.400 ;
        RECT 497.400 66.800 498.200 71.200 ;
        RECT 497.200 66.000 498.200 66.800 ;
        RECT 498.800 66.300 499.600 66.400 ;
        RECT 500.400 66.300 501.200 79.800 ;
        RECT 505.200 68.300 506.000 79.800 ;
        RECT 509.400 72.400 510.200 79.800 ;
        RECT 510.800 73.600 511.600 74.400 ;
        RECT 511.000 72.400 511.600 73.600 ;
        RECT 514.000 73.600 514.800 74.400 ;
        RECT 514.000 72.400 514.600 73.600 ;
        RECT 515.400 72.400 516.200 79.800 ;
        RECT 508.400 71.600 510.400 72.400 ;
        RECT 511.000 71.800 512.400 72.400 ;
        RECT 511.600 71.600 512.400 71.800 ;
        RECT 513.200 71.800 514.600 72.400 ;
        RECT 515.200 71.800 516.200 72.400 ;
        RECT 513.200 71.600 514.000 71.800 ;
        RECT 508.400 68.800 509.200 70.400 ;
        RECT 509.800 68.400 510.400 71.600 ;
        RECT 511.700 70.300 512.300 71.600 ;
        RECT 515.200 70.300 515.800 71.800 ;
        RECT 521.200 71.200 522.000 79.800 ;
        RECT 524.400 71.200 525.200 79.800 ;
        RECT 527.600 71.200 528.400 79.800 ;
        RECT 530.800 71.200 531.600 79.800 ;
        RECT 519.600 70.400 522.000 71.200 ;
        RECT 523.000 70.400 525.200 71.200 ;
        RECT 526.200 70.400 528.400 71.200 ;
        RECT 529.800 70.400 531.600 71.200 ;
        RECT 534.000 71.400 534.800 79.800 ;
        RECT 538.400 76.400 539.200 79.800 ;
        RECT 537.200 75.800 539.200 76.400 ;
        RECT 542.800 75.800 543.600 79.800 ;
        RECT 547.000 75.800 548.200 79.800 ;
        RECT 537.200 75.000 538.000 75.800 ;
        RECT 542.800 75.200 543.400 75.800 ;
        RECT 540.600 74.600 544.200 75.200 ;
        RECT 546.800 75.000 547.600 75.800 ;
        RECT 540.600 74.400 541.400 74.600 ;
        RECT 543.400 74.400 544.200 74.600 ;
        RECT 537.200 73.000 538.000 73.200 ;
        RECT 541.800 73.000 542.600 73.200 ;
        RECT 537.200 72.400 542.600 73.000 ;
        RECT 543.200 73.000 545.400 73.600 ;
        RECT 543.200 71.800 543.800 73.000 ;
        RECT 544.600 72.800 545.400 73.000 ;
        RECT 547.000 73.200 548.400 74.000 ;
        RECT 547.000 72.200 547.600 73.200 ;
        RECT 539.000 71.400 543.800 71.800 ;
        RECT 534.000 71.200 543.800 71.400 ;
        RECT 545.200 71.600 547.600 72.200 ;
        RECT 534.000 71.000 539.800 71.200 ;
        RECT 534.000 70.800 539.600 71.000 ;
        RECT 511.700 69.700 515.800 70.300 ;
        RECT 515.200 68.400 515.800 69.700 ;
        RECT 516.400 68.800 517.200 70.400 ;
        RECT 506.800 68.300 507.600 68.400 ;
        RECT 505.200 68.200 507.600 68.300 ;
        RECT 505.200 67.700 508.400 68.200 ;
        RECT 497.200 62.200 498.000 66.000 ;
        RECT 498.800 65.700 501.200 66.300 ;
        RECT 498.800 65.600 499.600 65.700 ;
        RECT 500.400 62.200 501.200 65.700 ;
        RECT 502.000 64.800 502.800 66.400 ;
        RECT 503.600 64.800 504.400 66.400 ;
        RECT 505.200 62.200 506.000 67.700 ;
        RECT 506.800 67.600 508.400 67.700 ;
        RECT 509.800 67.600 512.400 68.400 ;
        RECT 513.200 67.600 515.800 68.400 ;
        RECT 518.000 68.200 518.800 68.400 ;
        RECT 517.200 67.600 518.800 68.200 ;
        RECT 519.600 67.600 520.400 70.400 ;
        RECT 523.000 69.000 523.800 70.400 ;
        RECT 526.200 69.000 527.000 70.400 ;
        RECT 529.800 69.000 530.600 70.400 ;
        RECT 540.400 70.200 541.200 70.400 ;
        RECT 536.200 69.600 541.200 70.200 ;
        RECT 536.200 69.400 537.000 69.600 ;
        RECT 538.800 69.400 539.600 69.600 ;
        RECT 521.200 68.200 523.800 69.000 ;
        RECT 524.600 68.200 527.000 69.000 ;
        RECT 528.000 68.200 530.600 69.000 ;
        RECT 531.400 68.200 533.200 69.000 ;
        RECT 537.800 68.400 538.600 68.600 ;
        RECT 545.200 68.400 545.800 71.600 ;
        RECT 551.600 71.200 552.400 79.800 ;
        RECT 553.200 75.800 554.000 79.800 ;
        RECT 553.400 75.600 554.000 75.800 ;
        RECT 556.400 75.800 557.200 79.800 ;
        RECT 556.400 75.600 557.000 75.800 ;
        RECT 553.400 75.000 557.000 75.600 ;
        RECT 553.400 72.400 554.000 75.000 ;
        RECT 554.800 72.800 555.600 74.400 ;
        RECT 562.200 72.400 563.000 79.800 ;
        RECT 563.600 73.600 564.400 74.400 ;
        RECT 563.800 72.400 564.400 73.600 ;
        RECT 566.800 73.600 567.600 74.400 ;
        RECT 566.800 72.400 567.400 73.600 ;
        RECT 568.200 72.400 569.000 79.800 ;
        RECT 579.400 76.400 580.200 79.800 ;
        RECT 579.400 75.600 581.200 76.400 ;
        RECT 583.600 75.800 584.400 79.800 ;
        RECT 583.800 75.600 584.400 75.800 ;
        RECT 586.800 75.800 587.600 79.800 ;
        RECT 586.800 75.600 587.400 75.800 ;
        RECT 578.000 73.600 578.800 74.400 ;
        RECT 578.000 72.400 578.600 73.600 ;
        RECT 579.400 72.400 580.200 75.600 ;
        RECT 583.800 75.000 587.400 75.600 ;
        RECT 583.800 74.400 584.400 75.000 ;
        RECT 583.600 73.600 584.400 74.400 ;
        RECT 583.800 72.400 584.400 73.600 ;
        RECT 585.200 72.800 586.000 74.400 ;
        RECT 553.200 71.600 554.000 72.400 ;
        RECT 548.200 70.600 552.400 71.200 ;
        RECT 548.200 70.400 549.000 70.600 ;
        RECT 549.800 69.800 550.600 70.000 ;
        RECT 546.800 69.200 550.600 69.800 ;
        RECT 546.800 69.000 547.600 69.200 ;
        RECT 523.000 67.600 523.800 68.200 ;
        RECT 526.200 67.600 527.000 68.200 ;
        RECT 529.800 67.600 530.600 68.200 ;
        RECT 532.400 67.600 533.200 68.200 ;
        RECT 534.800 67.800 545.800 68.400 ;
        RECT 534.800 67.600 536.400 67.800 ;
        RECT 507.600 67.200 508.400 67.600 ;
        RECT 507.000 66.200 510.600 66.600 ;
        RECT 511.600 66.200 512.200 67.600 ;
        RECT 513.400 66.200 514.000 67.600 ;
        RECT 517.200 67.200 518.000 67.600 ;
        RECT 519.600 66.800 522.000 67.600 ;
        RECT 523.000 66.800 525.200 67.600 ;
        RECT 526.200 66.800 528.400 67.600 ;
        RECT 529.800 66.800 531.600 67.600 ;
        RECT 515.000 66.200 518.600 66.600 ;
        RECT 506.800 66.000 510.800 66.200 ;
        RECT 506.800 62.200 507.600 66.000 ;
        RECT 510.000 62.200 510.800 66.000 ;
        RECT 511.600 62.200 512.400 66.200 ;
        RECT 513.200 62.200 514.000 66.200 ;
        RECT 514.800 66.000 518.800 66.200 ;
        RECT 514.800 62.200 515.600 66.000 ;
        RECT 518.000 62.200 518.800 66.000 ;
        RECT 521.200 62.200 522.000 66.800 ;
        RECT 524.400 62.200 525.200 66.800 ;
        RECT 527.600 62.200 528.400 66.800 ;
        RECT 530.800 62.200 531.600 66.800 ;
        RECT 534.000 62.200 534.800 67.000 ;
        RECT 539.000 65.600 539.600 67.800 ;
        RECT 542.000 67.600 542.800 67.800 ;
        RECT 544.600 67.600 545.400 67.800 ;
        RECT 551.600 67.200 552.400 70.600 ;
        RECT 553.400 68.400 554.000 71.600 ;
        RECT 558.000 70.800 558.800 72.400 ;
        RECT 562.200 71.800 563.200 72.400 ;
        RECT 563.800 71.800 565.200 72.400 ;
        RECT 555.600 69.600 557.200 70.400 ;
        RECT 561.200 68.800 562.000 70.400 ;
        RECT 562.600 70.300 563.200 71.800 ;
        RECT 564.400 71.600 565.200 71.800 ;
        RECT 566.000 71.800 567.400 72.400 ;
        RECT 566.000 71.600 566.800 71.800 ;
        RECT 568.000 71.600 570.000 72.400 ;
        RECT 577.200 71.800 578.600 72.400 ;
        RECT 579.200 71.800 580.200 72.400 ;
        RECT 577.200 71.600 578.000 71.800 ;
        RECT 566.100 70.300 566.700 71.600 ;
        RECT 562.600 69.700 566.700 70.300 ;
        RECT 562.600 68.400 563.200 69.700 ;
        RECT 568.000 68.400 568.600 71.600 ;
        RECT 569.200 70.300 570.000 70.400 ;
        RECT 570.800 70.300 571.600 70.400 ;
        RECT 569.200 69.700 571.600 70.300 ;
        RECT 569.200 68.800 570.000 69.700 ;
        RECT 570.800 69.600 571.600 69.700 ;
        RECT 579.200 68.400 579.800 71.800 ;
        RECT 583.600 71.600 584.400 72.400 ;
        RECT 580.400 68.800 581.200 70.400 ;
        RECT 583.800 68.400 584.400 71.600 ;
        RECT 588.400 70.800 589.200 72.400 ;
        RECT 590.000 71.200 590.800 79.800 ;
        RECT 594.200 75.800 595.400 79.800 ;
        RECT 598.800 75.800 599.600 79.800 ;
        RECT 603.200 76.400 604.000 79.800 ;
        RECT 603.200 75.800 605.200 76.400 ;
        RECT 594.800 75.000 595.600 75.800 ;
        RECT 599.000 75.200 599.600 75.800 ;
        RECT 598.200 74.600 601.800 75.200 ;
        RECT 604.400 75.000 605.200 75.800 ;
        RECT 598.200 74.400 599.000 74.600 ;
        RECT 601.000 74.400 601.800 74.600 ;
        RECT 594.000 73.200 595.400 74.000 ;
        RECT 594.800 72.200 595.400 73.200 ;
        RECT 597.000 73.000 599.200 73.600 ;
        RECT 597.000 72.800 597.800 73.000 ;
        RECT 594.800 71.600 597.200 72.200 ;
        RECT 590.000 70.600 594.200 71.200 ;
        RECT 586.000 69.600 587.600 70.400 ;
        RECT 553.400 68.200 555.000 68.400 ;
        RECT 559.600 68.200 560.400 68.400 ;
        RECT 553.400 67.800 555.200 68.200 ;
        RECT 548.600 66.600 552.400 67.200 ;
        RECT 548.600 66.400 549.400 66.600 ;
        RECT 537.200 64.200 538.000 65.000 ;
        RECT 538.800 64.800 539.600 65.600 ;
        RECT 540.600 65.400 541.400 65.600 ;
        RECT 540.600 64.800 543.400 65.400 ;
        RECT 542.800 64.200 543.400 64.800 ;
        RECT 546.800 64.200 547.600 65.000 ;
        RECT 537.200 63.600 539.200 64.200 ;
        RECT 538.400 62.200 539.200 63.600 ;
        RECT 542.800 62.200 543.600 64.200 ;
        RECT 546.800 63.600 548.200 64.200 ;
        RECT 547.000 62.200 548.200 63.600 ;
        RECT 551.600 62.200 552.400 66.600 ;
        RECT 554.400 62.200 555.200 67.800 ;
        RECT 559.600 67.600 561.200 68.200 ;
        RECT 562.600 67.600 565.200 68.400 ;
        RECT 566.000 67.600 568.600 68.400 ;
        RECT 570.800 68.200 571.600 68.400 ;
        RECT 570.000 67.600 571.600 68.200 ;
        RECT 577.200 67.600 579.800 68.400 ;
        RECT 582.000 68.200 582.800 68.400 ;
        RECT 581.200 67.600 582.800 68.200 ;
        RECT 583.800 68.200 585.400 68.400 ;
        RECT 583.800 67.800 585.600 68.200 ;
        RECT 560.400 67.200 561.200 67.600 ;
        RECT 559.800 66.200 563.400 66.600 ;
        RECT 564.400 66.200 565.000 67.600 ;
        RECT 566.200 66.200 566.800 67.600 ;
        RECT 570.000 67.200 570.800 67.600 ;
        RECT 567.800 66.200 571.400 66.600 ;
        RECT 577.400 66.200 578.000 67.600 ;
        RECT 581.200 67.200 582.000 67.600 ;
        RECT 579.000 66.200 582.600 66.600 ;
        RECT 559.600 66.000 563.600 66.200 ;
        RECT 559.600 62.200 560.400 66.000 ;
        RECT 562.800 62.200 563.600 66.000 ;
        RECT 564.400 62.200 565.200 66.200 ;
        RECT 566.000 62.200 566.800 66.200 ;
        RECT 567.600 66.000 571.600 66.200 ;
        RECT 567.600 62.200 568.400 66.000 ;
        RECT 570.800 62.200 571.600 66.000 ;
        RECT 577.200 62.200 578.000 66.200 ;
        RECT 578.800 66.000 582.800 66.200 ;
        RECT 578.800 62.200 579.600 66.000 ;
        RECT 582.000 62.200 582.800 66.000 ;
        RECT 584.800 62.200 585.600 67.800 ;
        RECT 590.000 67.200 590.800 70.600 ;
        RECT 593.400 70.400 594.200 70.600 ;
        RECT 591.800 69.800 592.600 70.000 ;
        RECT 591.800 69.200 595.600 69.800 ;
        RECT 594.800 69.000 595.600 69.200 ;
        RECT 596.600 68.400 597.200 71.600 ;
        RECT 598.600 71.800 599.200 73.000 ;
        RECT 599.800 73.000 600.600 73.200 ;
        RECT 604.400 73.000 605.200 73.200 ;
        RECT 599.800 72.400 605.200 73.000 ;
        RECT 598.600 71.400 603.400 71.800 ;
        RECT 607.600 71.400 608.400 79.800 ;
        RECT 609.200 75.800 610.000 79.800 ;
        RECT 609.400 75.600 610.000 75.800 ;
        RECT 612.400 75.800 613.200 79.800 ;
        RECT 618.200 78.400 619.000 79.800 ;
        RECT 617.200 77.600 619.000 78.400 ;
        RECT 612.400 75.600 613.000 75.800 ;
        RECT 609.400 75.000 613.000 75.600 ;
        RECT 609.400 72.400 610.000 75.000 ;
        RECT 610.800 72.800 611.600 74.400 ;
        RECT 618.200 72.400 619.000 77.600 ;
        RECT 622.000 75.800 622.800 79.800 ;
        RECT 622.200 75.600 622.800 75.800 ;
        RECT 625.200 75.800 626.000 79.800 ;
        RECT 625.200 75.600 625.800 75.800 ;
        RECT 622.200 75.000 625.800 75.600 ;
        RECT 628.400 75.000 629.200 79.000 ;
        RECT 619.600 73.600 620.400 74.400 ;
        RECT 619.800 72.400 620.400 73.600 ;
        RECT 622.200 72.400 622.800 75.000 ;
        RECT 623.600 72.800 624.400 74.400 ;
        RECT 609.200 71.600 610.000 72.400 ;
        RECT 598.600 71.200 608.400 71.400 ;
        RECT 602.600 71.000 608.400 71.200 ;
        RECT 602.800 70.800 608.400 71.000 ;
        RECT 601.200 70.200 602.000 70.400 ;
        RECT 601.200 69.600 606.200 70.200 ;
        RECT 605.400 69.400 606.200 69.600 ;
        RECT 603.800 68.400 604.600 68.600 ;
        RECT 609.400 68.400 610.000 71.600 ;
        RECT 614.000 70.800 614.800 72.400 ;
        RECT 618.200 71.800 619.200 72.400 ;
        RECT 619.800 72.300 621.200 72.400 ;
        RECT 622.000 72.300 622.800 72.400 ;
        RECT 619.800 71.800 622.800 72.300 ;
        RECT 611.600 69.600 613.200 70.400 ;
        RECT 615.600 70.300 616.400 70.400 ;
        RECT 617.200 70.300 618.000 70.400 ;
        RECT 615.600 69.700 618.000 70.300 ;
        RECT 615.600 69.600 616.400 69.700 ;
        RECT 617.200 68.800 618.000 69.700 ;
        RECT 618.600 68.400 619.200 71.800 ;
        RECT 620.400 71.700 622.800 71.800 ;
        RECT 620.400 71.600 621.200 71.700 ;
        RECT 622.000 71.600 622.800 71.700 ;
        RECT 622.200 68.400 622.800 71.600 ;
        RECT 626.800 70.800 627.600 72.400 ;
        RECT 628.400 71.600 629.000 75.000 ;
        RECT 632.600 72.800 633.400 79.800 ;
        RECT 632.600 72.200 634.200 72.800 ;
        RECT 628.400 71.000 632.200 71.600 ;
        RECT 624.400 69.600 626.000 70.400 ;
        RECT 628.400 68.800 629.200 70.400 ;
        RECT 630.000 68.800 630.800 70.400 ;
        RECT 631.600 69.000 632.200 71.000 ;
        RECT 596.600 67.800 607.600 68.400 ;
        RECT 609.400 68.200 611.000 68.400 ;
        RECT 615.600 68.200 616.400 68.400 ;
        RECT 609.400 67.800 611.200 68.200 ;
        RECT 597.000 67.600 597.800 67.800 ;
        RECT 590.000 66.600 593.800 67.200 ;
        RECT 590.000 62.200 590.800 66.600 ;
        RECT 593.000 66.400 593.800 66.600 ;
        RECT 602.800 65.600 603.400 67.800 ;
        RECT 606.000 67.600 607.600 67.800 ;
        RECT 601.000 65.400 601.800 65.600 ;
        RECT 594.800 64.200 595.600 65.000 ;
        RECT 599.000 64.800 601.800 65.400 ;
        RECT 602.800 64.800 603.600 65.600 ;
        RECT 599.000 64.200 599.600 64.800 ;
        RECT 604.400 64.200 605.200 65.000 ;
        RECT 594.200 63.600 595.600 64.200 ;
        RECT 594.200 62.200 595.400 63.600 ;
        RECT 598.800 62.200 599.600 64.200 ;
        RECT 603.200 63.600 605.200 64.200 ;
        RECT 603.200 62.200 604.000 63.600 ;
        RECT 607.600 62.200 608.400 67.000 ;
        RECT 610.400 62.200 611.200 67.800 ;
        RECT 615.600 67.600 617.200 68.200 ;
        RECT 618.600 67.600 621.200 68.400 ;
        RECT 622.200 68.200 623.800 68.400 ;
        RECT 631.600 68.200 633.000 69.000 ;
        RECT 633.600 68.400 634.200 72.200 ;
        RECT 640.600 72.400 641.400 79.800 ;
        RECT 642.000 73.600 642.800 74.400 ;
        RECT 642.200 72.400 642.800 73.600 ;
        RECT 640.600 71.800 641.600 72.400 ;
        RECT 642.200 71.800 643.600 72.400 ;
        RECT 634.800 70.300 635.600 71.200 ;
        RECT 636.400 70.300 637.200 70.400 ;
        RECT 634.800 69.700 637.200 70.300 ;
        RECT 634.800 69.600 635.600 69.700 ;
        RECT 636.400 69.600 637.200 69.700 ;
        RECT 639.600 68.800 640.400 70.400 ;
        RECT 641.000 70.300 641.600 71.800 ;
        RECT 642.800 71.600 643.600 71.800 ;
        RECT 644.400 71.200 645.200 79.800 ;
        RECT 648.600 75.800 649.800 79.800 ;
        RECT 653.200 75.800 654.000 79.800 ;
        RECT 657.600 76.400 658.400 79.800 ;
        RECT 657.600 75.800 659.600 76.400 ;
        RECT 649.200 75.000 650.000 75.800 ;
        RECT 653.400 75.200 654.000 75.800 ;
        RECT 652.600 74.600 656.200 75.200 ;
        RECT 658.800 75.000 659.600 75.800 ;
        RECT 652.600 74.400 653.400 74.600 ;
        RECT 655.400 74.400 656.200 74.600 ;
        RECT 648.400 73.200 649.800 74.000 ;
        RECT 649.200 72.200 649.800 73.200 ;
        RECT 651.400 73.000 653.600 73.600 ;
        RECT 651.400 72.800 652.200 73.000 ;
        RECT 649.200 71.600 651.600 72.200 ;
        RECT 644.400 70.600 648.600 71.200 ;
        RECT 642.800 70.300 643.600 70.400 ;
        RECT 641.000 69.700 643.600 70.300 ;
        RECT 641.000 68.400 641.600 69.700 ;
        RECT 642.800 69.600 643.600 69.700 ;
        RECT 622.200 67.800 624.000 68.200 ;
        RECT 631.600 67.800 632.600 68.200 ;
        RECT 616.400 67.200 617.200 67.600 ;
        RECT 615.800 66.200 619.400 66.600 ;
        RECT 620.400 66.200 621.000 67.600 ;
        RECT 615.600 66.000 619.600 66.200 ;
        RECT 615.600 62.200 616.400 66.000 ;
        RECT 618.800 62.200 619.600 66.000 ;
        RECT 620.400 62.200 621.200 66.200 ;
        RECT 623.200 62.200 624.000 67.800 ;
        RECT 628.400 67.200 632.600 67.800 ;
        RECT 633.600 67.600 635.600 68.400 ;
        RECT 638.000 68.200 638.800 68.400 ;
        RECT 638.000 67.600 639.600 68.200 ;
        RECT 641.000 67.600 643.600 68.400 ;
        RECT 628.400 65.000 629.000 67.200 ;
        RECT 633.600 67.000 634.200 67.600 ;
        RECT 638.800 67.200 639.600 67.600 ;
        RECT 633.400 66.600 634.200 67.000 ;
        RECT 632.600 66.000 634.200 66.600 ;
        RECT 638.200 66.200 641.800 66.600 ;
        RECT 642.800 66.200 643.400 67.600 ;
        RECT 644.400 67.200 645.200 70.600 ;
        RECT 647.800 70.400 648.600 70.600 ;
        RECT 646.200 69.800 647.000 70.000 ;
        RECT 646.200 69.200 650.000 69.800 ;
        RECT 649.200 69.000 650.000 69.200 ;
        RECT 651.000 68.400 651.600 71.600 ;
        RECT 653.000 71.800 653.600 73.000 ;
        RECT 654.200 73.000 655.000 73.200 ;
        RECT 658.800 73.000 659.600 73.200 ;
        RECT 654.200 72.400 659.600 73.000 ;
        RECT 653.000 71.400 657.800 71.800 ;
        RECT 662.000 71.400 662.800 79.800 ;
        RECT 665.800 78.400 666.600 79.800 ;
        RECT 665.800 77.600 667.600 78.400 ;
        RECT 664.400 73.600 665.200 74.400 ;
        RECT 664.400 72.400 665.000 73.600 ;
        RECT 665.800 72.400 666.600 77.600 ;
        RECT 663.600 71.800 665.000 72.400 ;
        RECT 665.600 71.800 666.600 72.400 ;
        RECT 663.600 71.600 664.400 71.800 ;
        RECT 653.000 71.200 662.800 71.400 ;
        RECT 657.000 71.000 662.800 71.200 ;
        RECT 657.200 70.800 662.800 71.000 ;
        RECT 652.400 70.300 653.200 70.400 ;
        RECT 655.600 70.300 656.400 70.400 ;
        RECT 652.400 70.200 656.400 70.300 ;
        RECT 652.400 69.700 660.600 70.200 ;
        RECT 652.400 69.600 653.200 69.700 ;
        RECT 655.600 69.600 660.600 69.700 ;
        RECT 659.800 69.400 660.600 69.600 ;
        RECT 658.200 68.400 659.000 68.600 ;
        RECT 665.600 68.400 666.200 71.800 ;
        RECT 666.800 68.800 667.600 70.400 ;
        RECT 651.000 67.800 662.000 68.400 ;
        RECT 651.400 67.600 652.200 67.800 ;
        RECT 657.200 67.600 658.000 67.800 ;
        RECT 660.400 67.600 662.000 67.800 ;
        RECT 663.600 67.600 666.200 68.400 ;
        RECT 668.400 68.200 669.200 68.400 ;
        RECT 667.600 67.600 669.200 68.200 ;
        RECT 644.400 66.600 648.200 67.200 ;
        RECT 638.000 66.000 642.000 66.200 ;
        RECT 628.400 63.000 629.200 65.000 ;
        RECT 632.600 63.000 633.400 66.000 ;
        RECT 638.000 62.200 638.800 66.000 ;
        RECT 641.200 62.200 642.000 66.000 ;
        RECT 642.800 62.200 643.600 66.200 ;
        RECT 644.400 62.200 645.200 66.600 ;
        RECT 647.400 66.400 648.200 66.600 ;
        RECT 657.200 65.600 657.800 67.600 ;
        RECT 655.400 65.400 656.200 65.600 ;
        RECT 649.200 64.200 650.000 65.000 ;
        RECT 653.400 64.800 656.200 65.400 ;
        RECT 657.200 64.800 658.000 65.600 ;
        RECT 653.400 64.200 654.000 64.800 ;
        RECT 658.800 64.200 659.600 65.000 ;
        RECT 648.600 63.600 650.000 64.200 ;
        RECT 648.600 62.200 649.800 63.600 ;
        RECT 653.200 62.200 654.000 64.200 ;
        RECT 657.600 63.600 659.600 64.200 ;
        RECT 657.600 62.200 658.400 63.600 ;
        RECT 662.000 62.200 662.800 67.000 ;
        RECT 663.800 66.200 664.400 67.600 ;
        RECT 667.600 67.200 668.400 67.600 ;
        RECT 665.400 66.200 669.000 66.600 ;
        RECT 663.600 62.200 664.400 66.200 ;
        RECT 665.200 66.000 669.200 66.200 ;
        RECT 665.200 62.200 666.000 66.000 ;
        RECT 668.400 62.200 669.200 66.000 ;
        RECT 670.000 62.200 670.800 79.800 ;
        RECT 674.800 71.200 675.600 79.800 ;
        RECT 678.000 71.200 678.800 79.800 ;
        RECT 681.200 71.200 682.000 79.800 ;
        RECT 684.400 71.200 685.200 79.800 ;
        RECT 674.800 70.400 676.600 71.200 ;
        RECT 678.000 70.400 680.200 71.200 ;
        RECT 681.200 70.400 683.400 71.200 ;
        RECT 684.400 70.400 686.800 71.200 ;
        RECT 675.800 69.000 676.600 70.400 ;
        RECT 679.400 69.000 680.200 70.400 ;
        RECT 682.600 69.000 683.400 70.400 ;
        RECT 673.200 68.200 675.000 69.000 ;
        RECT 675.800 68.200 678.400 69.000 ;
        RECT 679.400 68.200 681.800 69.000 ;
        RECT 682.600 68.200 685.200 69.000 ;
        RECT 673.200 67.600 674.000 68.200 ;
        RECT 675.800 67.600 676.600 68.200 ;
        RECT 679.400 67.600 680.200 68.200 ;
        RECT 682.600 67.600 683.400 68.200 ;
        RECT 686.000 67.600 686.800 70.400 ;
        RECT 674.800 66.800 676.600 67.600 ;
        RECT 678.000 66.800 680.200 67.600 ;
        RECT 681.200 66.800 683.400 67.600 ;
        RECT 684.400 66.800 686.800 67.600 ;
        RECT 671.600 64.800 672.400 66.400 ;
        RECT 674.800 62.200 675.600 66.800 ;
        RECT 678.000 62.200 678.800 66.800 ;
        RECT 681.200 62.200 682.000 66.800 ;
        RECT 684.400 62.200 685.200 66.800 ;
        RECT 1.200 55.000 2.000 59.800 ;
        RECT 5.600 58.400 6.400 59.800 ;
        RECT 4.400 57.800 6.400 58.400 ;
        RECT 10.000 57.800 10.800 59.800 ;
        RECT 14.200 58.400 15.400 59.800 ;
        RECT 14.000 57.800 15.400 58.400 ;
        RECT 4.400 57.000 5.200 57.800 ;
        RECT 10.000 57.200 10.600 57.800 ;
        RECT 6.000 55.600 6.800 57.200 ;
        RECT 7.800 56.600 10.600 57.200 ;
        RECT 14.000 57.000 14.800 57.800 ;
        RECT 7.800 56.400 8.600 56.600 ;
        RECT 2.000 54.200 3.600 54.400 ;
        RECT 6.200 54.200 6.800 55.600 ;
        RECT 15.800 55.400 16.600 55.600 ;
        RECT 18.800 55.400 19.600 59.800 ;
        RECT 20.400 56.000 21.200 59.800 ;
        RECT 23.600 56.000 24.400 59.800 ;
        RECT 20.400 55.800 24.400 56.000 ;
        RECT 25.200 55.800 26.000 59.800 ;
        RECT 26.800 55.800 27.600 59.800 ;
        RECT 28.400 56.000 29.200 59.800 ;
        RECT 31.600 56.000 32.400 59.800 ;
        RECT 28.400 55.800 32.400 56.000 ;
        RECT 33.800 58.400 34.600 59.800 ;
        RECT 40.600 58.400 41.400 59.800 ;
        RECT 33.800 57.600 35.600 58.400 ;
        RECT 39.600 57.600 41.400 58.400 ;
        RECT 33.800 56.400 34.600 57.600 ;
        RECT 40.600 56.400 41.400 57.600 ;
        RECT 33.800 55.800 35.600 56.400 ;
        RECT 20.600 55.400 24.200 55.800 ;
        RECT 15.800 54.800 19.600 55.400 ;
        RECT 11.800 54.200 12.600 54.400 ;
        RECT 2.000 53.600 13.000 54.200 ;
        RECT 5.000 53.400 5.800 53.600 ;
        RECT 3.400 52.400 4.200 52.600 ;
        RECT 12.400 52.400 13.000 53.600 ;
        RECT 14.000 52.800 14.800 53.000 ;
        RECT 3.400 52.300 8.400 52.400 ;
        RECT 9.200 52.300 10.000 52.400 ;
        RECT 3.400 51.800 10.000 52.300 ;
        RECT 7.600 51.700 10.000 51.800 ;
        RECT 7.600 51.600 8.400 51.700 ;
        RECT 9.200 51.600 10.000 51.700 ;
        RECT 12.400 51.600 13.200 52.400 ;
        RECT 14.000 52.200 17.800 52.800 ;
        RECT 17.000 52.000 17.800 52.200 ;
        RECT 1.200 51.000 6.800 51.200 ;
        RECT 1.200 50.800 7.000 51.000 ;
        RECT 1.200 50.600 11.000 50.800 ;
        RECT 1.200 42.200 2.000 50.600 ;
        RECT 6.200 50.200 11.000 50.600 ;
        RECT 4.400 49.000 9.800 49.600 ;
        RECT 4.400 48.800 5.200 49.000 ;
        RECT 9.000 48.800 9.800 49.000 ;
        RECT 10.400 49.000 11.000 50.200 ;
        RECT 12.400 50.400 13.000 51.600 ;
        RECT 15.400 51.400 16.200 51.600 ;
        RECT 18.800 51.400 19.600 54.800 ;
        RECT 21.200 54.400 22.000 54.800 ;
        RECT 25.200 54.400 25.800 55.800 ;
        RECT 27.000 54.400 27.600 55.800 ;
        RECT 28.600 55.400 32.200 55.800 ;
        RECT 30.800 54.400 31.600 54.800 ;
        RECT 20.400 53.800 22.000 54.400 ;
        RECT 20.400 53.600 21.200 53.800 ;
        RECT 23.400 53.600 26.000 54.400 ;
        RECT 26.800 53.600 29.400 54.400 ;
        RECT 30.800 53.800 32.400 54.400 ;
        RECT 31.600 53.600 32.400 53.800 ;
        RECT 22.000 51.600 22.800 53.200 ;
        RECT 23.400 52.300 24.000 53.600 ;
        RECT 23.400 51.700 27.500 52.300 ;
        RECT 15.400 50.800 19.600 51.400 ;
        RECT 12.400 49.800 14.800 50.400 ;
        RECT 11.800 49.000 12.600 49.200 ;
        RECT 10.400 48.400 12.600 49.000 ;
        RECT 14.200 48.800 14.800 49.800 ;
        RECT 14.200 48.000 15.600 48.800 ;
        RECT 7.800 47.400 8.600 47.600 ;
        RECT 10.600 47.400 11.400 47.600 ;
        RECT 4.400 46.200 5.200 47.000 ;
        RECT 7.800 46.800 11.400 47.400 ;
        RECT 10.000 46.200 10.600 46.800 ;
        RECT 14.000 46.200 14.800 47.000 ;
        RECT 4.400 45.600 6.400 46.200 ;
        RECT 5.600 42.200 6.400 45.600 ;
        RECT 10.000 42.200 10.800 46.200 ;
        RECT 14.200 42.200 15.400 46.200 ;
        RECT 18.800 42.200 19.600 50.800 ;
        RECT 23.400 50.200 24.000 51.700 ;
        RECT 26.900 50.400 27.500 51.700 ;
        RECT 25.200 50.200 26.000 50.400 ;
        RECT 23.000 49.600 24.000 50.200 ;
        RECT 24.600 49.600 26.000 50.200 ;
        RECT 26.800 50.200 27.600 50.400 ;
        RECT 28.800 50.200 29.400 53.600 ;
        RECT 30.000 51.600 30.800 53.200 ;
        RECT 26.800 49.600 28.200 50.200 ;
        RECT 28.800 49.600 29.800 50.200 ;
        RECT 23.000 42.200 23.800 49.600 ;
        RECT 24.600 48.400 25.200 49.600 ;
        RECT 24.400 47.600 25.200 48.400 ;
        RECT 27.600 48.400 28.200 49.600 ;
        RECT 27.600 47.600 28.400 48.400 ;
        RECT 29.000 42.200 29.800 49.600 ;
        RECT 33.200 47.600 34.000 50.400 ;
        RECT 34.800 42.200 35.600 55.800 ;
        RECT 39.600 55.800 41.400 56.400 ;
        RECT 46.600 56.000 47.400 59.000 ;
        RECT 50.800 57.000 51.600 59.000 ;
        RECT 36.400 54.300 37.200 55.200 ;
        RECT 38.000 54.300 38.800 55.200 ;
        RECT 36.400 53.700 38.800 54.300 ;
        RECT 36.400 53.600 37.200 53.700 ;
        RECT 38.000 53.600 38.800 53.700 ;
        RECT 39.600 42.200 40.400 55.800 ;
        RECT 45.800 55.400 47.400 56.000 ;
        RECT 45.800 55.000 46.600 55.400 ;
        RECT 45.800 54.400 46.400 55.000 ;
        RECT 51.000 54.800 51.600 57.000 ;
        RECT 52.400 56.000 53.200 59.800 ;
        RECT 55.600 56.000 56.400 59.800 ;
        RECT 52.400 55.800 56.400 56.000 ;
        RECT 57.200 55.800 58.000 59.800 ;
        RECT 58.800 55.800 59.600 59.800 ;
        RECT 60.400 56.000 61.200 59.800 ;
        RECT 63.600 56.000 64.400 59.800 ;
        RECT 60.400 55.800 64.400 56.000 ;
        RECT 52.600 55.400 56.200 55.800 ;
        RECT 41.200 54.300 42.000 54.400 ;
        RECT 44.400 54.300 46.400 54.400 ;
        RECT 41.200 53.700 46.400 54.300 ;
        RECT 47.400 54.200 51.600 54.800 ;
        RECT 53.200 54.400 54.000 54.800 ;
        RECT 57.200 54.400 57.800 55.800 ;
        RECT 59.000 54.400 59.600 55.800 ;
        RECT 60.600 55.400 64.200 55.800 ;
        RECT 65.200 55.000 66.000 59.800 ;
        RECT 69.600 58.400 70.400 59.800 ;
        RECT 68.400 57.800 70.400 58.400 ;
        RECT 74.000 57.800 74.800 59.800 ;
        RECT 78.200 58.400 79.400 59.800 ;
        RECT 78.000 57.800 79.400 58.400 ;
        RECT 68.400 57.000 69.200 57.800 ;
        RECT 74.000 57.200 74.600 57.800 ;
        RECT 70.000 55.600 70.800 57.200 ;
        RECT 71.800 56.600 74.600 57.200 ;
        RECT 78.000 57.000 78.800 57.800 ;
        RECT 71.800 56.400 72.600 56.600 ;
        RECT 62.800 54.400 63.600 54.800 ;
        RECT 47.400 53.800 48.400 54.200 ;
        RECT 41.200 53.600 42.000 53.700 ;
        RECT 44.400 53.600 46.400 53.700 ;
        RECT 44.400 50.800 45.200 52.400 ;
        RECT 41.200 47.600 42.000 50.400 ;
        RECT 45.800 49.800 46.400 53.600 ;
        RECT 47.000 53.000 48.400 53.800 ;
        RECT 52.400 53.800 54.000 54.400 ;
        RECT 52.400 53.600 53.200 53.800 ;
        RECT 55.400 53.600 58.000 54.400 ;
        RECT 58.800 53.600 61.400 54.400 ;
        RECT 62.800 53.800 64.400 54.400 ;
        RECT 63.600 53.600 64.400 53.800 ;
        RECT 66.000 54.200 67.600 54.400 ;
        RECT 70.200 54.200 70.800 55.600 ;
        RECT 79.800 55.400 80.600 55.600 ;
        RECT 82.800 55.400 83.600 59.800 ;
        RECT 87.000 58.400 87.800 59.800 ;
        RECT 86.000 57.600 87.800 58.400 ;
        RECT 87.000 56.400 87.800 57.600 ;
        RECT 79.800 54.800 83.600 55.400 ;
        RECT 86.000 55.800 87.800 56.400 ;
        RECT 89.800 56.400 90.600 59.800 ;
        RECT 94.000 57.000 94.800 59.000 ;
        RECT 89.800 55.800 91.600 56.400 ;
        RECT 75.800 54.200 76.600 54.400 ;
        RECT 66.000 53.600 77.000 54.200 ;
        RECT 47.800 51.000 48.400 53.000 ;
        RECT 49.200 51.600 50.000 53.200 ;
        RECT 50.800 51.600 51.600 53.200 ;
        RECT 54.000 51.600 54.800 53.200 ;
        RECT 55.400 52.300 56.000 53.600 ;
        RECT 60.800 52.400 61.400 53.600 ;
        RECT 69.000 53.400 69.800 53.600 ;
        RECT 55.400 51.700 59.500 52.300 ;
        RECT 47.800 50.400 51.600 51.000 ;
        RECT 45.800 49.200 47.400 49.800 ;
        RECT 46.600 42.200 47.400 49.200 ;
        RECT 51.000 47.000 51.600 50.400 ;
        RECT 55.400 50.200 56.000 51.700 ;
        RECT 58.900 50.400 59.500 51.700 ;
        RECT 60.400 51.600 61.400 52.400 ;
        RECT 62.000 51.600 62.800 53.200 ;
        RECT 67.400 52.400 68.200 52.600 ;
        RECT 70.000 52.400 70.800 52.600 ;
        RECT 67.400 51.800 72.400 52.400 ;
        RECT 71.600 51.600 72.400 51.800 ;
        RECT 57.200 50.200 58.000 50.400 ;
        RECT 50.800 43.000 51.600 47.000 ;
        RECT 55.000 49.600 56.000 50.200 ;
        RECT 56.600 49.600 58.000 50.200 ;
        RECT 58.800 50.200 59.600 50.400 ;
        RECT 60.800 50.200 61.400 51.600 ;
        RECT 65.200 51.000 70.800 51.200 ;
        RECT 65.200 50.800 71.000 51.000 ;
        RECT 65.200 50.600 75.000 50.800 ;
        RECT 58.800 49.600 60.200 50.200 ;
        RECT 60.800 49.600 61.800 50.200 ;
        RECT 55.000 42.200 55.800 49.600 ;
        RECT 56.600 48.400 57.200 49.600 ;
        RECT 56.400 47.600 57.200 48.400 ;
        RECT 59.600 48.400 60.200 49.600 ;
        RECT 59.600 47.600 60.400 48.400 ;
        RECT 61.000 42.200 61.800 49.600 ;
        RECT 65.200 42.200 66.000 50.600 ;
        RECT 70.200 50.200 75.000 50.600 ;
        RECT 68.400 49.000 73.800 49.600 ;
        RECT 68.400 48.800 69.200 49.000 ;
        RECT 73.000 48.800 73.800 49.000 ;
        RECT 74.400 49.000 75.000 50.200 ;
        RECT 76.400 50.400 77.000 53.600 ;
        RECT 78.000 52.800 78.800 53.000 ;
        RECT 78.000 52.200 81.800 52.800 ;
        RECT 81.000 52.000 81.800 52.200 ;
        RECT 79.400 51.400 80.200 51.600 ;
        RECT 82.800 51.400 83.600 54.800 ;
        RECT 84.400 53.600 85.200 55.200 ;
        RECT 79.400 50.800 83.600 51.400 ;
        RECT 76.400 49.800 78.800 50.400 ;
        RECT 75.800 49.000 76.600 49.200 ;
        RECT 74.400 48.400 76.600 49.000 ;
        RECT 78.200 48.800 78.800 49.800 ;
        RECT 78.200 48.000 79.600 48.800 ;
        RECT 71.800 47.400 72.600 47.600 ;
        RECT 74.600 47.400 75.400 47.600 ;
        RECT 68.400 46.200 69.200 47.000 ;
        RECT 71.800 46.800 75.400 47.400 ;
        RECT 74.000 46.200 74.600 46.800 ;
        RECT 78.000 46.200 78.800 47.000 ;
        RECT 68.400 45.600 70.400 46.200 ;
        RECT 69.600 42.200 70.400 45.600 ;
        RECT 74.000 42.200 74.800 46.200 ;
        RECT 78.200 42.200 79.400 46.200 ;
        RECT 82.800 42.200 83.600 50.800 ;
        RECT 86.000 42.200 86.800 55.800 ;
        RECT 87.600 48.800 88.400 50.400 ;
        RECT 89.200 48.800 90.000 50.400 ;
        RECT 90.800 42.200 91.600 55.800 ;
        RECT 92.400 53.600 93.200 55.200 ;
        RECT 94.000 54.800 94.600 57.000 ;
        RECT 98.200 56.000 99.000 59.000 ;
        RECT 107.400 58.400 108.200 59.000 ;
        RECT 106.800 57.600 108.200 58.400 ;
        RECT 107.400 56.000 108.200 57.600 ;
        RECT 111.600 57.000 112.400 59.000 ;
        RECT 98.200 55.400 99.800 56.000 ;
        RECT 99.000 55.000 99.800 55.400 ;
        RECT 94.000 54.200 98.200 54.800 ;
        RECT 97.200 53.800 98.200 54.200 ;
        RECT 99.200 54.400 99.800 55.000 ;
        RECT 106.600 55.400 108.200 56.000 ;
        RECT 106.600 55.000 107.400 55.400 ;
        RECT 106.600 54.400 107.200 55.000 ;
        RECT 111.800 54.800 112.400 57.000 ;
        RECT 118.000 56.000 118.800 59.800 ;
        RECT 121.200 56.000 122.000 59.800 ;
        RECT 118.000 55.800 122.000 56.000 ;
        RECT 122.800 55.800 123.600 59.800 ;
        RECT 124.400 56.000 125.200 59.800 ;
        RECT 127.600 56.000 128.400 59.800 ;
        RECT 124.400 55.800 128.400 56.000 ;
        RECT 129.200 55.800 130.000 59.800 ;
        RECT 130.800 56.000 131.600 59.800 ;
        RECT 134.000 56.000 134.800 59.800 ;
        RECT 130.800 55.800 134.800 56.000 ;
        RECT 135.600 55.800 136.400 59.800 ;
        RECT 137.200 57.000 138.000 59.000 ;
        RECT 118.200 55.400 121.800 55.800 ;
        RECT 94.000 51.600 94.800 53.200 ;
        RECT 95.600 51.600 96.400 53.200 ;
        RECT 97.200 53.000 98.600 53.800 ;
        RECT 99.200 53.600 101.200 54.400 ;
        RECT 105.200 53.600 107.200 54.400 ;
        RECT 108.200 54.200 112.400 54.800 ;
        RECT 118.800 54.400 119.600 54.800 ;
        RECT 122.800 54.400 123.400 55.800 ;
        RECT 124.600 55.400 128.200 55.800 ;
        RECT 125.200 54.400 126.000 54.800 ;
        RECT 129.200 54.400 129.800 55.800 ;
        RECT 131.000 55.400 134.600 55.800 ;
        RECT 131.600 54.400 132.400 54.800 ;
        RECT 135.600 54.400 136.200 55.800 ;
        RECT 137.200 54.800 137.800 57.000 ;
        RECT 141.400 56.400 142.200 59.000 ;
        RECT 140.400 56.000 142.200 56.400 ;
        RECT 140.400 55.600 143.000 56.000 ;
        RECT 146.800 55.600 147.600 57.200 ;
        RECT 141.400 55.400 143.000 55.600 ;
        RECT 142.200 55.000 143.000 55.400 ;
        RECT 108.200 53.800 109.200 54.200 ;
        RECT 97.200 51.000 97.800 53.000 ;
        RECT 94.000 50.400 97.800 51.000 ;
        RECT 94.000 47.000 94.600 50.400 ;
        RECT 99.200 49.800 99.800 53.600 ;
        RECT 100.400 50.800 101.200 52.400 ;
        RECT 105.200 50.800 106.000 52.400 ;
        RECT 98.200 49.200 99.800 49.800 ;
        RECT 106.600 49.800 107.200 53.600 ;
        RECT 107.800 53.000 109.200 53.800 ;
        RECT 118.000 53.800 119.600 54.400 ;
        RECT 118.000 53.600 118.800 53.800 ;
        RECT 121.000 53.600 123.600 54.400 ;
        RECT 124.400 53.800 126.000 54.400 ;
        RECT 124.400 53.600 125.200 53.800 ;
        RECT 127.400 53.600 130.000 54.400 ;
        RECT 130.800 53.800 132.400 54.400 ;
        RECT 130.800 53.600 131.600 53.800 ;
        RECT 133.800 53.600 136.400 54.400 ;
        RECT 137.200 54.200 141.400 54.800 ;
        RECT 140.400 53.800 141.400 54.200 ;
        RECT 142.400 54.400 143.000 55.000 ;
        RECT 108.600 51.000 109.200 53.000 ;
        RECT 110.000 51.600 110.800 53.200 ;
        RECT 111.600 52.300 112.400 53.200 ;
        RECT 118.000 52.300 118.800 52.400 ;
        RECT 111.600 51.700 118.800 52.300 ;
        RECT 111.600 51.600 112.400 51.700 ;
        RECT 118.000 51.600 118.800 51.700 ;
        RECT 119.600 51.600 120.400 53.200 ;
        RECT 108.600 50.400 112.400 51.000 ;
        RECT 106.600 49.200 108.200 49.800 ;
        RECT 94.000 43.000 94.800 47.000 ;
        RECT 98.200 44.400 99.000 49.200 ;
        RECT 98.200 43.600 99.600 44.400 ;
        RECT 98.200 42.200 99.000 43.600 ;
        RECT 107.400 42.200 108.200 49.200 ;
        RECT 111.800 47.000 112.400 50.400 ;
        RECT 121.000 50.200 121.600 53.600 ;
        RECT 126.000 51.600 126.800 53.200 ;
        RECT 127.400 52.400 128.000 53.600 ;
        RECT 127.400 51.600 128.400 52.400 ;
        RECT 132.400 51.600 133.200 53.200 ;
        RECT 122.800 50.200 123.600 50.400 ;
        RECT 127.400 50.200 128.000 51.600 ;
        RECT 129.200 50.200 130.000 50.400 ;
        RECT 133.800 50.200 134.400 53.600 ;
        RECT 137.200 51.600 138.000 53.200 ;
        RECT 138.800 51.600 139.600 53.200 ;
        RECT 140.400 53.000 141.800 53.800 ;
        RECT 142.400 53.600 144.400 54.400 ;
        RECT 140.400 51.000 141.000 53.000 ;
        RECT 137.200 50.400 141.000 51.000 ;
        RECT 135.600 50.200 136.400 50.400 ;
        RECT 111.600 43.000 112.400 47.000 ;
        RECT 120.600 49.600 121.600 50.200 ;
        RECT 122.200 49.600 123.600 50.200 ;
        RECT 127.000 49.600 128.000 50.200 ;
        RECT 128.600 49.600 130.000 50.200 ;
        RECT 133.400 49.600 134.400 50.200 ;
        RECT 135.000 49.600 136.400 50.200 ;
        RECT 120.600 42.200 121.400 49.600 ;
        RECT 122.200 48.400 122.800 49.600 ;
        RECT 122.000 47.600 122.800 48.400 ;
        RECT 127.000 42.200 127.800 49.600 ;
        RECT 128.600 48.400 129.200 49.600 ;
        RECT 133.400 48.400 134.200 49.600 ;
        RECT 135.000 48.400 135.600 49.600 ;
        RECT 128.400 47.600 129.200 48.400 ;
        RECT 132.400 47.600 134.200 48.400 ;
        RECT 134.800 47.600 135.600 48.400 ;
        RECT 133.400 42.200 134.200 47.600 ;
        RECT 137.200 47.000 137.800 50.400 ;
        RECT 142.400 49.800 143.000 53.600 ;
        RECT 143.600 50.800 144.400 52.400 ;
        RECT 141.400 49.200 143.000 49.800 ;
        RECT 137.200 43.000 138.000 47.000 ;
        RECT 141.400 42.200 142.200 49.200 ;
        RECT 148.400 42.200 149.200 59.800 ;
        RECT 153.800 56.000 154.600 59.000 ;
        RECT 158.000 57.000 158.800 59.000 ;
        RECT 153.000 55.400 154.600 56.000 ;
        RECT 153.000 55.000 153.800 55.400 ;
        RECT 153.000 54.400 153.600 55.000 ;
        RECT 158.200 54.800 158.800 57.000 ;
        RECT 159.600 55.600 160.400 57.200 ;
        RECT 151.600 53.600 153.600 54.400 ;
        RECT 154.600 54.200 158.800 54.800 ;
        RECT 161.200 54.300 162.000 59.800 ;
        RECT 162.800 56.000 163.600 59.800 ;
        RECT 166.000 56.000 166.800 59.800 ;
        RECT 162.800 55.800 166.800 56.000 ;
        RECT 167.600 55.800 168.400 59.800 ;
        RECT 163.000 55.400 166.600 55.800 ;
        RECT 163.600 54.400 164.400 54.800 ;
        RECT 167.600 54.400 168.200 55.800 ;
        RECT 162.800 54.300 164.400 54.400 ;
        RECT 154.600 53.800 155.600 54.200 ;
        RECT 151.600 50.800 152.400 52.400 ;
        RECT 153.000 49.800 153.600 53.600 ;
        RECT 154.200 53.000 155.600 53.800 ;
        RECT 161.200 53.800 164.400 54.300 ;
        RECT 161.200 53.700 163.600 53.800 ;
        RECT 155.000 51.000 155.600 53.000 ;
        RECT 156.400 51.600 157.200 53.200 ;
        RECT 158.000 51.600 158.800 53.200 ;
        RECT 155.000 50.400 158.800 51.000 ;
        RECT 153.000 49.200 154.600 49.800 ;
        RECT 153.800 44.400 154.600 49.200 ;
        RECT 158.200 47.000 158.800 50.400 ;
        RECT 153.200 43.600 154.600 44.400 ;
        RECT 153.800 42.200 154.600 43.600 ;
        RECT 158.000 43.000 158.800 47.000 ;
        RECT 161.200 42.200 162.000 53.700 ;
        RECT 162.800 53.600 163.600 53.700 ;
        RECT 165.800 53.600 168.400 54.400 ;
        RECT 172.800 54.200 173.600 59.800 ;
        RECT 175.600 56.300 176.400 56.400 ;
        RECT 177.200 56.300 178.000 59.800 ;
        RECT 175.600 55.700 178.000 56.300 ;
        RECT 175.600 55.600 176.400 55.700 ;
        RECT 177.000 55.200 178.000 55.700 ;
        RECT 172.800 53.800 174.600 54.200 ;
        RECT 173.000 53.600 174.600 53.800 ;
        RECT 164.400 51.600 165.200 53.200 ;
        RECT 165.800 50.200 166.400 53.600 ;
        RECT 170.800 51.600 172.400 52.400 ;
        RECT 167.600 50.200 168.400 50.400 ;
        RECT 165.400 49.600 166.400 50.200 ;
        RECT 167.000 49.600 168.400 50.200 ;
        RECT 169.200 49.600 170.000 51.200 ;
        RECT 174.000 50.400 174.600 53.600 ;
        RECT 177.000 50.800 177.800 55.200 ;
        RECT 178.800 54.600 179.600 59.800 ;
        RECT 185.200 56.600 186.000 59.800 ;
        RECT 186.800 57.000 187.600 59.800 ;
        RECT 188.400 57.000 189.200 59.800 ;
        RECT 190.000 57.000 190.800 59.800 ;
        RECT 191.600 57.000 192.400 59.800 ;
        RECT 194.800 57.000 195.600 59.800 ;
        RECT 198.000 57.000 198.800 59.800 ;
        RECT 199.600 57.000 200.400 59.800 ;
        RECT 201.200 57.000 202.000 59.800 ;
        RECT 183.600 55.800 186.000 56.600 ;
        RECT 202.800 56.600 203.600 59.800 ;
        RECT 183.600 55.200 184.400 55.800 ;
        RECT 178.400 54.000 179.600 54.600 ;
        RECT 182.600 54.600 184.400 55.200 ;
        RECT 188.400 55.600 189.400 56.400 ;
        RECT 192.400 55.600 194.000 56.400 ;
        RECT 194.800 55.800 199.400 56.400 ;
        RECT 202.800 55.800 205.400 56.600 ;
        RECT 194.800 55.600 195.600 55.800 ;
        RECT 178.400 52.000 179.000 54.000 ;
        RECT 182.600 53.400 183.400 54.600 ;
        RECT 179.600 52.600 183.400 53.400 ;
        RECT 188.400 52.800 189.200 55.600 ;
        RECT 194.800 54.800 195.600 55.000 ;
        RECT 191.200 54.200 195.600 54.800 ;
        RECT 191.200 54.000 192.000 54.200 ;
        RECT 196.400 53.600 197.200 55.200 ;
        RECT 198.600 53.400 199.400 55.800 ;
        RECT 204.600 55.200 205.400 55.800 ;
        RECT 204.600 54.400 207.600 55.200 ;
        RECT 209.200 53.800 210.000 59.800 ;
        RECT 212.400 56.400 213.200 59.800 ;
        RECT 191.600 52.600 194.800 53.400 ;
        RECT 198.600 52.600 200.600 53.400 ;
        RECT 201.200 53.000 210.000 53.800 ;
        RECT 185.200 52.000 186.000 52.600 ;
        RECT 202.800 52.000 203.600 52.400 ;
        RECT 206.000 52.000 206.800 52.400 ;
        RECT 207.800 52.000 208.600 52.200 ;
        RECT 178.400 51.400 179.200 52.000 ;
        RECT 185.200 51.400 208.600 52.000 ;
        RECT 174.000 49.600 174.800 50.400 ;
        RECT 177.000 50.000 178.000 50.800 ;
        RECT 165.400 42.200 166.200 49.600 ;
        RECT 167.000 48.400 167.600 49.600 ;
        RECT 166.800 47.600 167.600 48.400 ;
        RECT 172.400 47.600 173.200 49.200 ;
        RECT 174.000 47.000 174.600 49.600 ;
        RECT 171.000 46.400 174.600 47.000 ;
        RECT 170.800 42.200 171.600 46.400 ;
        RECT 174.000 46.200 174.600 46.400 ;
        RECT 174.000 42.200 174.800 46.200 ;
        RECT 177.200 42.200 178.000 50.000 ;
        RECT 178.600 49.600 179.200 51.400 ;
        RECT 178.600 49.000 187.600 49.600 ;
        RECT 178.600 47.400 179.200 49.000 ;
        RECT 186.800 48.800 187.600 49.000 ;
        RECT 190.000 49.000 198.600 49.600 ;
        RECT 190.000 48.800 190.800 49.000 ;
        RECT 181.800 47.600 184.400 48.400 ;
        RECT 178.600 46.800 181.200 47.400 ;
        RECT 180.400 42.200 181.200 46.800 ;
        RECT 183.600 42.200 184.400 47.600 ;
        RECT 185.000 46.800 189.200 47.600 ;
        RECT 186.800 42.200 187.600 45.000 ;
        RECT 188.400 42.200 189.200 45.000 ;
        RECT 190.000 42.200 190.800 45.000 ;
        RECT 191.600 42.200 192.400 48.400 ;
        RECT 194.800 47.600 197.400 48.400 ;
        RECT 198.000 48.200 198.600 49.000 ;
        RECT 199.600 49.400 200.400 49.600 ;
        RECT 199.600 49.000 205.000 49.400 ;
        RECT 199.600 48.800 205.800 49.000 ;
        RECT 204.400 48.200 205.800 48.800 ;
        RECT 198.000 47.600 203.800 48.200 ;
        RECT 206.800 48.000 208.400 48.800 ;
        RECT 206.800 47.600 207.400 48.000 ;
        RECT 194.800 42.200 195.600 47.000 ;
        RECT 198.000 42.200 198.800 47.000 ;
        RECT 203.200 46.800 207.400 47.600 ;
        RECT 209.200 47.400 210.000 53.000 ;
        RECT 212.200 55.800 213.200 56.400 ;
        RECT 212.200 54.400 212.800 55.800 ;
        RECT 215.600 55.200 216.400 59.800 ;
        RECT 213.800 54.600 216.400 55.200 ;
        RECT 212.200 53.600 213.200 54.400 ;
        RECT 212.200 50.200 212.800 53.600 ;
        RECT 213.800 53.000 214.400 54.600 ;
        RECT 213.400 52.200 214.400 53.000 ;
        RECT 213.800 50.200 214.400 52.200 ;
        RECT 217.200 53.800 218.000 59.800 ;
        RECT 223.600 56.600 224.400 59.800 ;
        RECT 225.200 57.000 226.000 59.800 ;
        RECT 226.800 57.000 227.600 59.800 ;
        RECT 228.400 57.000 229.200 59.800 ;
        RECT 231.600 57.000 232.400 59.800 ;
        RECT 234.800 57.000 235.600 59.800 ;
        RECT 236.400 57.000 237.200 59.800 ;
        RECT 238.000 57.000 238.800 59.800 ;
        RECT 239.600 57.000 240.400 59.800 ;
        RECT 221.800 55.800 224.400 56.600 ;
        RECT 241.200 56.600 242.000 59.800 ;
        RECT 227.800 55.800 232.400 56.400 ;
        RECT 221.800 55.200 222.600 55.800 ;
        RECT 219.600 54.400 222.600 55.200 ;
        RECT 217.200 53.000 226.000 53.800 ;
        RECT 227.800 53.400 228.600 55.800 ;
        RECT 231.600 55.600 232.400 55.800 ;
        RECT 233.200 55.600 234.800 56.400 ;
        RECT 237.800 55.600 238.800 56.400 ;
        RECT 241.200 55.800 243.600 56.600 ;
        RECT 230.000 53.600 230.800 55.200 ;
        RECT 231.600 54.800 232.400 55.000 ;
        RECT 231.600 54.200 236.000 54.800 ;
        RECT 235.200 54.000 236.000 54.200 ;
        RECT 212.200 49.200 213.200 50.200 ;
        RECT 213.800 49.600 216.400 50.200 ;
        RECT 208.000 46.800 210.000 47.400 ;
        RECT 199.600 42.200 200.400 45.000 ;
        RECT 201.200 42.200 202.000 45.000 ;
        RECT 204.400 42.200 205.200 46.800 ;
        RECT 208.000 46.200 208.600 46.800 ;
        RECT 207.600 45.600 208.600 46.200 ;
        RECT 207.600 42.200 208.400 45.600 ;
        RECT 212.400 42.200 213.200 49.200 ;
        RECT 215.600 42.200 216.400 49.600 ;
        RECT 217.200 47.400 218.000 53.000 ;
        RECT 226.600 52.600 228.600 53.400 ;
        RECT 232.400 52.600 235.600 53.400 ;
        RECT 238.000 52.800 238.800 55.600 ;
        RECT 242.800 55.200 243.600 55.800 ;
        RECT 242.800 54.600 244.600 55.200 ;
        RECT 243.800 53.400 244.600 54.600 ;
        RECT 247.600 54.600 248.400 59.800 ;
        RECT 249.200 56.000 250.000 59.800 ;
        RECT 249.200 55.200 250.200 56.000 ;
        RECT 252.400 55.800 253.200 59.800 ;
        RECT 254.000 56.000 254.800 59.800 ;
        RECT 257.200 56.000 258.000 59.800 ;
        RECT 254.000 55.800 258.000 56.000 ;
        RECT 247.600 54.000 248.800 54.600 ;
        RECT 243.800 52.600 247.600 53.400 ;
        RECT 218.800 52.200 219.600 52.400 ;
        RECT 218.600 52.000 219.600 52.200 ;
        RECT 220.400 52.000 221.200 52.400 ;
        RECT 223.600 52.000 224.400 52.400 ;
        RECT 241.200 52.000 242.000 52.600 ;
        RECT 248.200 52.000 248.800 54.000 ;
        RECT 218.600 51.400 242.000 52.000 ;
        RECT 248.000 51.400 248.800 52.000 ;
        RECT 248.000 49.600 248.600 51.400 ;
        RECT 249.400 50.800 250.200 55.200 ;
        RECT 252.600 54.400 253.200 55.800 ;
        RECT 254.200 55.400 257.800 55.800 ;
        RECT 256.400 54.400 257.200 54.800 ;
        RECT 252.400 53.600 255.000 54.400 ;
        RECT 256.400 53.800 258.000 54.400 ;
        RECT 257.200 53.600 258.000 53.800 ;
        RECT 263.600 53.800 264.400 59.800 ;
        RECT 270.000 56.600 270.800 59.800 ;
        RECT 271.600 57.000 272.400 59.800 ;
        RECT 273.200 57.000 274.000 59.800 ;
        RECT 274.800 57.000 275.600 59.800 ;
        RECT 278.000 57.000 278.800 59.800 ;
        RECT 281.200 57.000 282.000 59.800 ;
        RECT 282.800 57.000 283.600 59.800 ;
        RECT 284.400 57.000 285.200 59.800 ;
        RECT 286.000 57.000 286.800 59.800 ;
        RECT 268.200 55.800 270.800 56.600 ;
        RECT 287.600 56.600 288.400 59.800 ;
        RECT 274.200 55.800 278.800 56.400 ;
        RECT 268.200 55.200 269.000 55.800 ;
        RECT 266.000 54.400 269.000 55.200 ;
        RECT 226.800 49.400 227.600 49.600 ;
        RECT 222.200 49.000 227.600 49.400 ;
        RECT 221.400 48.800 227.600 49.000 ;
        RECT 228.600 49.000 237.200 49.600 ;
        RECT 218.800 48.000 220.400 48.800 ;
        RECT 221.400 48.200 222.800 48.800 ;
        RECT 228.600 48.200 229.200 49.000 ;
        RECT 236.400 48.800 237.200 49.000 ;
        RECT 239.600 49.000 248.600 49.600 ;
        RECT 239.600 48.800 240.400 49.000 ;
        RECT 219.800 47.600 220.400 48.000 ;
        RECT 223.400 47.600 229.200 48.200 ;
        RECT 229.800 47.600 232.400 48.400 ;
        RECT 217.200 46.800 219.200 47.400 ;
        RECT 219.800 46.800 224.000 47.600 ;
        RECT 218.600 46.200 219.200 46.800 ;
        RECT 218.600 45.600 219.600 46.200 ;
        RECT 218.800 42.200 219.600 45.600 ;
        RECT 222.000 42.200 222.800 46.800 ;
        RECT 225.200 42.200 226.000 45.000 ;
        RECT 226.800 42.200 227.600 45.000 ;
        RECT 228.400 42.200 229.200 47.000 ;
        RECT 231.600 42.200 232.400 47.000 ;
        RECT 234.800 42.200 235.600 48.400 ;
        RECT 242.800 47.600 245.400 48.400 ;
        RECT 238.000 46.800 242.200 47.600 ;
        RECT 236.400 42.200 237.200 45.000 ;
        RECT 238.000 42.200 238.800 45.000 ;
        RECT 239.600 42.200 240.400 45.000 ;
        RECT 242.800 42.200 243.600 47.600 ;
        RECT 248.000 47.400 248.600 49.000 ;
        RECT 246.000 46.800 248.600 47.400 ;
        RECT 249.200 50.300 250.200 50.800 ;
        RECT 252.400 50.300 253.200 50.400 ;
        RECT 249.200 50.200 253.200 50.300 ;
        RECT 254.400 50.200 255.000 53.600 ;
        RECT 255.600 51.600 256.400 53.200 ;
        RECT 263.600 53.000 272.400 53.800 ;
        RECT 274.200 53.400 275.000 55.800 ;
        RECT 278.000 55.600 278.800 55.800 ;
        RECT 279.600 55.600 281.200 56.400 ;
        RECT 284.200 55.600 285.200 56.400 ;
        RECT 287.600 55.800 290.000 56.600 ;
        RECT 276.400 53.600 277.200 55.200 ;
        RECT 278.000 54.800 278.800 55.000 ;
        RECT 278.000 54.200 282.400 54.800 ;
        RECT 281.600 54.000 282.400 54.200 ;
        RECT 249.200 49.700 253.800 50.200 ;
        RECT 246.000 42.200 246.800 46.800 ;
        RECT 249.200 42.200 250.000 49.700 ;
        RECT 252.400 49.600 253.800 49.700 ;
        RECT 254.400 49.600 255.400 50.200 ;
        RECT 253.200 48.400 253.800 49.600 ;
        RECT 252.400 47.600 254.000 48.400 ;
        RECT 254.600 42.200 255.400 49.600 ;
        RECT 263.600 47.400 264.400 53.000 ;
        RECT 273.000 52.600 275.000 53.400 ;
        RECT 278.800 52.600 282.000 53.400 ;
        RECT 284.400 52.800 285.200 55.600 ;
        RECT 289.200 55.200 290.000 55.800 ;
        RECT 289.200 54.600 291.000 55.200 ;
        RECT 290.200 53.400 291.000 54.600 ;
        RECT 294.000 54.600 294.800 59.800 ;
        RECT 295.600 56.000 296.400 59.800 ;
        RECT 299.400 56.400 300.200 59.800 ;
        RECT 295.600 55.200 296.600 56.000 ;
        RECT 299.400 55.800 301.200 56.400 ;
        RECT 303.600 55.800 304.400 59.800 ;
        RECT 305.200 56.000 306.000 59.800 ;
        RECT 308.400 56.000 309.200 59.800 ;
        RECT 312.600 56.400 313.400 59.800 ;
        RECT 305.200 55.800 309.200 56.000 ;
        RECT 311.600 55.800 313.400 56.400 ;
        RECT 316.400 56.000 317.200 59.800 ;
        RECT 294.000 54.000 295.200 54.600 ;
        RECT 290.200 52.600 294.000 53.400 ;
        RECT 265.000 52.000 265.800 52.200 ;
        RECT 266.800 52.000 267.600 52.400 ;
        RECT 270.000 52.000 270.800 52.400 ;
        RECT 287.600 52.000 288.400 52.600 ;
        RECT 294.600 52.000 295.200 54.000 ;
        RECT 265.000 51.400 288.400 52.000 ;
        RECT 294.400 51.400 295.200 52.000 ;
        RECT 294.400 49.600 295.000 51.400 ;
        RECT 295.800 50.800 296.600 55.200 ;
        RECT 297.200 54.300 298.000 54.400 ;
        RECT 300.400 54.300 301.200 55.800 ;
        RECT 297.200 53.700 301.200 54.300 ;
        RECT 297.200 53.600 298.000 53.700 ;
        RECT 273.200 49.400 274.000 49.600 ;
        RECT 268.600 49.000 274.000 49.400 ;
        RECT 267.800 48.800 274.000 49.000 ;
        RECT 275.000 49.000 283.600 49.600 ;
        RECT 265.200 48.000 266.800 48.800 ;
        RECT 267.800 48.200 269.200 48.800 ;
        RECT 275.000 48.200 275.600 49.000 ;
        RECT 282.800 48.800 283.600 49.000 ;
        RECT 286.000 49.000 295.000 49.600 ;
        RECT 286.000 48.800 286.800 49.000 ;
        RECT 266.200 47.600 266.800 48.000 ;
        RECT 269.800 47.600 275.600 48.200 ;
        RECT 276.200 47.600 278.800 48.400 ;
        RECT 263.600 46.800 265.600 47.400 ;
        RECT 266.200 46.800 270.400 47.600 ;
        RECT 265.000 46.200 265.600 46.800 ;
        RECT 265.000 45.600 266.000 46.200 ;
        RECT 265.200 42.200 266.000 45.600 ;
        RECT 268.400 42.200 269.200 46.800 ;
        RECT 271.600 42.200 272.400 45.000 ;
        RECT 273.200 42.200 274.000 45.000 ;
        RECT 274.800 42.200 275.600 47.000 ;
        RECT 278.000 42.200 278.800 47.000 ;
        RECT 281.200 42.200 282.000 48.400 ;
        RECT 289.200 47.600 291.800 48.400 ;
        RECT 284.400 46.800 288.600 47.600 ;
        RECT 282.800 42.200 283.600 45.000 ;
        RECT 284.400 42.200 285.200 45.000 ;
        RECT 286.000 42.200 286.800 45.000 ;
        RECT 289.200 42.200 290.000 47.600 ;
        RECT 294.400 47.400 295.000 49.000 ;
        RECT 292.400 46.800 295.000 47.400 ;
        RECT 295.600 50.000 296.600 50.800 ;
        RECT 292.400 42.200 293.200 46.800 ;
        RECT 295.600 42.200 296.400 50.000 ;
        RECT 298.800 48.800 299.600 50.400 ;
        RECT 300.400 42.200 301.200 53.700 ;
        RECT 302.000 54.300 302.800 55.200 ;
        RECT 303.800 54.400 304.400 55.800 ;
        RECT 305.400 55.400 309.000 55.800 ;
        RECT 307.600 54.400 308.400 54.800 ;
        RECT 303.600 54.300 306.200 54.400 ;
        RECT 302.000 53.700 306.200 54.300 ;
        RECT 307.600 53.800 309.200 54.400 ;
        RECT 302.000 53.600 302.800 53.700 ;
        RECT 303.600 53.600 306.200 53.700 ;
        RECT 308.400 53.600 309.200 53.800 ;
        RECT 310.000 53.600 310.800 55.200 ;
        RECT 302.000 50.300 302.800 50.400 ;
        RECT 303.600 50.300 304.400 50.400 ;
        RECT 302.000 50.200 304.400 50.300 ;
        RECT 305.600 50.200 306.200 53.600 ;
        RECT 306.800 51.600 307.600 53.200 ;
        RECT 302.000 49.700 305.000 50.200 ;
        RECT 302.000 49.600 302.800 49.700 ;
        RECT 303.600 49.600 305.000 49.700 ;
        RECT 305.600 49.600 306.600 50.200 ;
        RECT 304.400 48.400 305.000 49.600 ;
        RECT 304.400 47.600 305.200 48.400 ;
        RECT 305.800 42.200 306.600 49.600 ;
        RECT 311.600 42.200 312.400 55.800 ;
        RECT 316.200 55.200 317.200 56.000 ;
        RECT 316.200 50.800 317.000 55.200 ;
        RECT 318.000 54.600 318.800 59.800 ;
        RECT 324.400 56.600 325.200 59.800 ;
        RECT 326.000 57.000 326.800 59.800 ;
        RECT 327.600 57.000 328.400 59.800 ;
        RECT 329.200 57.000 330.000 59.800 ;
        RECT 330.800 57.000 331.600 59.800 ;
        RECT 334.000 57.000 334.800 59.800 ;
        RECT 337.200 57.000 338.000 59.800 ;
        RECT 338.800 57.000 339.600 59.800 ;
        RECT 340.400 57.000 341.200 59.800 ;
        RECT 322.800 55.800 325.200 56.600 ;
        RECT 342.000 56.600 342.800 59.800 ;
        RECT 322.800 55.200 323.600 55.800 ;
        RECT 317.600 54.000 318.800 54.600 ;
        RECT 321.800 54.600 323.600 55.200 ;
        RECT 327.600 55.600 328.600 56.400 ;
        RECT 331.600 55.600 333.200 56.400 ;
        RECT 334.000 55.800 338.600 56.400 ;
        RECT 342.000 55.800 344.600 56.600 ;
        RECT 334.000 55.600 334.800 55.800 ;
        RECT 317.600 52.000 318.200 54.000 ;
        RECT 321.800 53.400 322.600 54.600 ;
        RECT 318.800 52.600 322.600 53.400 ;
        RECT 327.600 52.800 328.400 55.600 ;
        RECT 334.000 54.800 334.800 55.000 ;
        RECT 330.400 54.200 334.800 54.800 ;
        RECT 330.400 54.000 331.200 54.200 ;
        RECT 335.600 53.600 336.400 55.200 ;
        RECT 337.800 53.400 338.600 55.800 ;
        RECT 343.800 55.200 344.600 55.800 ;
        RECT 343.800 54.400 346.800 55.200 ;
        RECT 348.400 53.800 349.200 59.800 ;
        RECT 330.800 52.600 334.000 53.400 ;
        RECT 337.800 52.600 339.800 53.400 ;
        RECT 340.400 53.000 349.200 53.800 ;
        RECT 324.400 52.000 325.200 52.600 ;
        RECT 342.000 52.000 342.800 52.400 ;
        RECT 343.600 52.000 344.400 52.400 ;
        RECT 347.000 52.000 347.800 52.200 ;
        RECT 317.600 51.400 318.400 52.000 ;
        RECT 324.400 51.400 347.800 52.000 ;
        RECT 313.200 50.300 314.000 50.400 ;
        RECT 316.200 50.300 317.200 50.800 ;
        RECT 313.200 49.700 317.200 50.300 ;
        RECT 313.200 47.600 314.000 49.700 ;
        RECT 316.400 42.200 317.200 49.700 ;
        RECT 317.800 49.600 318.400 51.400 ;
        RECT 317.800 49.000 326.800 49.600 ;
        RECT 317.800 47.400 318.400 49.000 ;
        RECT 326.000 48.800 326.800 49.000 ;
        RECT 329.200 49.000 337.800 49.600 ;
        RECT 329.200 48.800 330.000 49.000 ;
        RECT 321.000 47.600 323.600 48.400 ;
        RECT 317.800 46.800 320.400 47.400 ;
        RECT 319.600 42.200 320.400 46.800 ;
        RECT 322.800 42.200 323.600 47.600 ;
        RECT 324.200 46.800 328.400 47.600 ;
        RECT 326.000 42.200 326.800 45.000 ;
        RECT 327.600 42.200 328.400 45.000 ;
        RECT 329.200 42.200 330.000 45.000 ;
        RECT 330.800 42.200 331.600 48.400 ;
        RECT 334.000 47.600 336.600 48.400 ;
        RECT 337.200 48.200 337.800 49.000 ;
        RECT 338.800 49.400 339.600 49.600 ;
        RECT 338.800 49.000 344.200 49.400 ;
        RECT 338.800 48.800 345.000 49.000 ;
        RECT 343.600 48.200 345.000 48.800 ;
        RECT 337.200 47.600 343.000 48.200 ;
        RECT 346.000 48.000 347.600 48.800 ;
        RECT 346.000 47.600 346.600 48.000 ;
        RECT 334.000 42.200 334.800 47.000 ;
        RECT 337.200 42.200 338.000 47.000 ;
        RECT 342.400 46.800 346.600 47.600 ;
        RECT 348.400 47.400 349.200 53.000 ;
        RECT 347.200 46.800 349.200 47.400 ;
        RECT 351.600 55.200 352.400 59.800 ;
        RECT 354.800 55.200 355.600 59.800 ;
        RECT 359.600 56.000 360.400 59.800 ;
        RECT 351.600 54.400 355.600 55.200 ;
        RECT 359.400 55.200 360.400 56.000 ;
        RECT 351.600 51.600 352.400 54.400 ;
        RECT 358.000 52.300 358.800 52.400 ;
        RECT 354.800 51.700 358.800 52.300 ;
        RECT 354.800 51.600 355.600 51.700 ;
        RECT 358.000 51.600 358.800 51.700 ;
        RECT 351.600 50.800 355.600 51.600 ;
        RECT 338.800 42.200 339.600 45.000 ;
        RECT 340.400 42.200 341.200 45.000 ;
        RECT 343.600 42.200 344.400 46.800 ;
        RECT 347.200 46.200 347.800 46.800 ;
        RECT 346.800 45.600 347.800 46.200 ;
        RECT 346.800 42.200 347.600 45.600 ;
        RECT 351.600 42.200 352.400 50.800 ;
        RECT 354.800 42.200 355.600 50.800 ;
        RECT 359.400 50.800 360.200 55.200 ;
        RECT 361.200 54.600 362.000 59.800 ;
        RECT 367.600 56.600 368.400 59.800 ;
        RECT 369.200 57.000 370.000 59.800 ;
        RECT 370.800 57.000 371.600 59.800 ;
        RECT 372.400 57.000 373.200 59.800 ;
        RECT 374.000 57.000 374.800 59.800 ;
        RECT 377.200 57.000 378.000 59.800 ;
        RECT 380.400 57.000 381.200 59.800 ;
        RECT 382.000 57.000 382.800 59.800 ;
        RECT 383.600 57.000 384.400 59.800 ;
        RECT 366.000 55.800 368.400 56.600 ;
        RECT 385.200 56.600 386.000 59.800 ;
        RECT 366.000 55.200 366.800 55.800 ;
        RECT 360.800 54.000 362.000 54.600 ;
        RECT 365.000 54.600 366.800 55.200 ;
        RECT 370.800 55.600 371.800 56.400 ;
        RECT 374.800 55.600 376.400 56.400 ;
        RECT 377.200 55.800 381.800 56.400 ;
        RECT 385.200 55.800 387.800 56.600 ;
        RECT 377.200 55.600 378.000 55.800 ;
        RECT 360.800 52.000 361.400 54.000 ;
        RECT 365.000 53.400 365.800 54.600 ;
        RECT 362.000 52.600 365.800 53.400 ;
        RECT 370.800 52.800 371.600 55.600 ;
        RECT 377.200 54.800 378.000 55.000 ;
        RECT 373.600 54.200 378.000 54.800 ;
        RECT 373.600 54.000 374.400 54.200 ;
        RECT 378.800 53.600 379.600 55.200 ;
        RECT 381.000 53.400 381.800 55.800 ;
        RECT 387.000 55.200 387.800 55.800 ;
        RECT 387.000 54.400 390.000 55.200 ;
        RECT 391.600 53.800 392.400 59.800 ;
        RECT 395.800 56.400 396.600 59.800 ;
        RECT 394.800 55.800 396.600 56.400 ;
        RECT 399.600 56.000 400.400 59.800 ;
        RECT 374.000 52.600 377.200 53.400 ;
        RECT 381.000 52.600 383.000 53.400 ;
        RECT 383.600 53.000 392.400 53.800 ;
        RECT 393.200 53.600 394.000 55.200 ;
        RECT 367.600 52.000 368.400 52.600 ;
        RECT 378.800 52.000 379.600 52.400 ;
        RECT 385.200 52.000 386.000 52.400 ;
        RECT 390.200 52.000 391.000 52.200 ;
        RECT 360.800 51.400 361.600 52.000 ;
        RECT 367.600 51.400 391.000 52.000 ;
        RECT 359.400 50.000 360.400 50.800 ;
        RECT 359.600 42.200 360.400 50.000 ;
        RECT 361.000 49.600 361.600 51.400 ;
        RECT 361.000 49.000 370.000 49.600 ;
        RECT 361.000 47.400 361.600 49.000 ;
        RECT 369.200 48.800 370.000 49.000 ;
        RECT 372.400 49.000 381.000 49.600 ;
        RECT 372.400 48.800 373.200 49.000 ;
        RECT 364.200 47.600 366.800 48.400 ;
        RECT 361.000 46.800 363.600 47.400 ;
        RECT 362.800 42.200 363.600 46.800 ;
        RECT 366.000 42.200 366.800 47.600 ;
        RECT 367.400 46.800 371.600 47.600 ;
        RECT 369.200 42.200 370.000 45.000 ;
        RECT 370.800 42.200 371.600 45.000 ;
        RECT 372.400 42.200 373.200 45.000 ;
        RECT 374.000 42.200 374.800 48.400 ;
        RECT 377.200 47.600 379.800 48.400 ;
        RECT 380.400 48.200 381.000 49.000 ;
        RECT 382.000 49.400 382.800 49.600 ;
        RECT 382.000 49.000 387.400 49.400 ;
        RECT 382.000 48.800 388.200 49.000 ;
        RECT 386.800 48.200 388.200 48.800 ;
        RECT 380.400 47.600 386.200 48.200 ;
        RECT 389.200 48.000 390.800 48.800 ;
        RECT 389.200 47.600 389.800 48.000 ;
        RECT 377.200 42.200 378.000 47.000 ;
        RECT 380.400 42.200 381.200 47.000 ;
        RECT 385.600 46.800 389.800 47.600 ;
        RECT 391.600 47.400 392.400 53.000 ;
        RECT 390.400 46.800 392.400 47.400 ;
        RECT 382.000 42.200 382.800 45.000 ;
        RECT 383.600 42.200 384.400 45.000 ;
        RECT 386.800 42.200 387.600 46.800 ;
        RECT 390.400 46.200 391.000 46.800 ;
        RECT 390.000 45.600 391.000 46.200 ;
        RECT 390.000 42.200 390.800 45.600 ;
        RECT 394.800 42.200 395.600 55.800 ;
        RECT 399.400 55.200 400.400 56.000 ;
        RECT 399.400 50.800 400.200 55.200 ;
        RECT 401.200 54.600 402.000 59.800 ;
        RECT 407.600 56.600 408.400 59.800 ;
        RECT 409.200 57.000 410.000 59.800 ;
        RECT 410.800 57.000 411.600 59.800 ;
        RECT 412.400 57.000 413.200 59.800 ;
        RECT 414.000 57.000 414.800 59.800 ;
        RECT 417.200 57.000 418.000 59.800 ;
        RECT 420.400 57.000 421.200 59.800 ;
        RECT 422.000 57.000 422.800 59.800 ;
        RECT 423.600 57.000 424.400 59.800 ;
        RECT 406.000 55.800 408.400 56.600 ;
        RECT 425.200 56.600 426.000 59.800 ;
        RECT 406.000 55.200 406.800 55.800 ;
        RECT 400.800 54.000 402.000 54.600 ;
        RECT 405.000 54.600 406.800 55.200 ;
        RECT 410.800 55.600 411.800 56.400 ;
        RECT 414.800 55.600 416.400 56.400 ;
        RECT 417.200 55.800 421.800 56.400 ;
        RECT 425.200 55.800 427.800 56.600 ;
        RECT 417.200 55.600 418.000 55.800 ;
        RECT 400.800 52.000 401.400 54.000 ;
        RECT 405.000 53.400 405.800 54.600 ;
        RECT 402.000 52.600 405.800 53.400 ;
        RECT 410.800 52.800 411.600 55.600 ;
        RECT 417.200 54.800 418.000 55.000 ;
        RECT 413.600 54.200 418.000 54.800 ;
        RECT 413.600 54.000 414.400 54.200 ;
        RECT 418.800 53.600 419.600 55.200 ;
        RECT 421.000 53.400 421.800 55.800 ;
        RECT 427.000 55.200 427.800 55.800 ;
        RECT 427.000 54.400 430.000 55.200 ;
        RECT 431.600 53.800 432.400 59.800 ;
        RECT 438.600 56.400 439.400 59.800 ;
        RECT 444.400 57.800 445.200 59.800 ;
        RECT 438.600 55.800 440.400 56.400 ;
        RECT 414.000 52.600 417.200 53.400 ;
        RECT 421.000 52.600 423.000 53.400 ;
        RECT 423.600 53.000 432.400 53.800 ;
        RECT 407.600 52.000 408.400 52.600 ;
        RECT 425.200 52.000 426.000 52.400 ;
        RECT 428.400 52.000 429.200 52.400 ;
        RECT 430.200 52.000 431.000 52.200 ;
        RECT 400.800 51.400 401.600 52.000 ;
        RECT 407.600 51.400 431.000 52.000 ;
        RECT 396.400 50.300 397.200 50.400 ;
        RECT 399.400 50.300 400.400 50.800 ;
        RECT 396.400 49.700 400.400 50.300 ;
        RECT 396.400 48.800 397.200 49.700 ;
        RECT 399.600 42.200 400.400 49.700 ;
        RECT 401.000 49.600 401.600 51.400 ;
        RECT 401.000 49.000 410.000 49.600 ;
        RECT 401.000 47.400 401.600 49.000 ;
        RECT 409.200 48.800 410.000 49.000 ;
        RECT 412.400 49.000 421.000 49.600 ;
        RECT 412.400 48.800 413.200 49.000 ;
        RECT 404.200 47.600 406.800 48.400 ;
        RECT 401.000 46.800 403.600 47.400 ;
        RECT 402.800 42.200 403.600 46.800 ;
        RECT 406.000 42.200 406.800 47.600 ;
        RECT 407.400 46.800 411.600 47.600 ;
        RECT 409.200 42.200 410.000 45.000 ;
        RECT 410.800 42.200 411.600 45.000 ;
        RECT 412.400 42.200 413.200 45.000 ;
        RECT 414.000 42.200 414.800 48.400 ;
        RECT 417.200 47.600 419.800 48.400 ;
        RECT 420.400 48.200 421.000 49.000 ;
        RECT 422.000 49.400 422.800 49.600 ;
        RECT 422.000 49.000 427.400 49.400 ;
        RECT 422.000 48.800 428.200 49.000 ;
        RECT 426.800 48.200 428.200 48.800 ;
        RECT 420.400 47.600 426.200 48.200 ;
        RECT 429.200 48.000 430.800 48.800 ;
        RECT 429.200 47.600 429.800 48.000 ;
        RECT 417.200 42.200 418.000 47.000 ;
        RECT 420.400 42.200 421.200 47.000 ;
        RECT 425.600 46.800 429.800 47.600 ;
        RECT 431.600 47.400 432.400 53.000 ;
        RECT 434.800 52.300 435.600 52.400 ;
        RECT 439.600 52.300 440.400 55.800 ;
        RECT 442.800 55.600 443.600 57.200 ;
        RECT 444.600 55.600 445.200 57.800 ;
        RECT 447.600 55.800 448.400 59.800 ;
        RECT 451.800 58.400 452.600 59.800 ;
        RECT 456.600 58.400 457.400 59.800 ;
        RECT 451.800 57.600 453.200 58.400 ;
        RECT 455.600 57.600 457.400 58.400 ;
        RECT 451.800 56.400 452.600 57.600 ;
        RECT 456.600 56.400 457.400 57.600 ;
        RECT 441.200 53.600 442.000 55.200 ;
        RECT 444.600 55.000 447.000 55.600 ;
        RECT 444.400 53.600 445.400 54.400 ;
        RECT 444.800 52.800 445.600 53.600 ;
        RECT 434.800 51.700 440.400 52.300 ;
        RECT 446.400 52.000 447.000 55.000 ;
        RECT 447.800 52.400 448.400 55.800 ;
        RECT 450.800 55.800 452.600 56.400 ;
        RECT 455.600 55.800 457.400 56.400 ;
        RECT 449.200 53.600 450.000 55.200 ;
        RECT 434.800 51.600 435.600 51.700 ;
        RECT 433.200 48.300 434.000 48.400 ;
        RECT 438.000 48.300 438.800 50.400 ;
        RECT 433.200 47.700 438.800 48.300 ;
        RECT 433.200 47.600 434.000 47.700 ;
        RECT 430.400 46.800 432.400 47.400 ;
        RECT 422.000 42.200 422.800 45.000 ;
        RECT 423.600 42.200 424.400 45.000 ;
        RECT 426.800 42.200 427.600 46.800 ;
        RECT 430.400 46.200 431.000 46.800 ;
        RECT 430.000 45.600 431.000 46.200 ;
        RECT 430.000 42.200 430.800 45.600 ;
        RECT 439.600 42.200 440.400 51.700 ;
        RECT 446.200 51.400 447.000 52.000 ;
        RECT 447.600 51.600 448.400 52.400 ;
        RECT 442.800 51.200 447.000 51.400 ;
        RECT 442.800 50.800 446.800 51.200 ;
        RECT 442.800 42.200 443.600 50.800 ;
        RECT 447.800 50.200 448.400 51.600 ;
        RECT 447.000 49.600 448.400 50.200 ;
        RECT 447.000 44.400 447.800 49.600 ;
        RECT 447.000 43.600 448.400 44.400 ;
        RECT 447.000 42.200 447.800 43.600 ;
        RECT 450.800 42.200 451.600 55.800 ;
        RECT 454.000 53.600 454.800 55.200 ;
        RECT 452.400 48.300 453.200 50.400 ;
        RECT 454.000 48.300 454.800 48.400 ;
        RECT 452.400 47.700 454.800 48.300 ;
        RECT 454.000 47.600 454.800 47.700 ;
        RECT 455.600 42.200 456.400 55.800 ;
        RECT 458.800 53.800 459.600 59.800 ;
        RECT 465.200 56.600 466.000 59.800 ;
        RECT 466.800 57.000 467.600 59.800 ;
        RECT 468.400 57.000 469.200 59.800 ;
        RECT 470.000 57.000 470.800 59.800 ;
        RECT 473.200 57.000 474.000 59.800 ;
        RECT 476.400 57.000 477.200 59.800 ;
        RECT 478.000 57.000 478.800 59.800 ;
        RECT 479.600 57.000 480.400 59.800 ;
        RECT 481.200 57.000 482.000 59.800 ;
        RECT 463.400 55.800 466.000 56.600 ;
        RECT 482.800 56.600 483.600 59.800 ;
        RECT 469.400 55.800 474.000 56.400 ;
        RECT 463.400 55.200 464.200 55.800 ;
        RECT 461.200 54.400 464.200 55.200 ;
        RECT 458.800 53.000 467.600 53.800 ;
        RECT 469.400 53.400 470.200 55.800 ;
        RECT 473.200 55.600 474.000 55.800 ;
        RECT 474.800 55.600 476.400 56.400 ;
        RECT 479.400 55.600 480.400 56.400 ;
        RECT 482.800 55.800 485.200 56.600 ;
        RECT 471.600 53.600 472.400 55.200 ;
        RECT 473.200 54.800 474.000 55.000 ;
        RECT 473.200 54.200 477.600 54.800 ;
        RECT 476.800 54.000 477.600 54.200 ;
        RECT 457.200 47.600 458.000 50.400 ;
        RECT 458.800 47.400 459.600 53.000 ;
        RECT 468.200 52.600 470.200 53.400 ;
        RECT 474.000 52.600 477.200 53.400 ;
        RECT 479.600 52.800 480.400 55.600 ;
        RECT 484.400 55.200 485.200 55.800 ;
        RECT 484.400 54.600 486.200 55.200 ;
        RECT 485.400 53.400 486.200 54.600 ;
        RECT 489.200 54.600 490.000 59.800 ;
        RECT 490.800 56.000 491.600 59.800 ;
        RECT 490.800 55.200 491.800 56.000 ;
        RECT 494.000 55.800 494.800 59.800 ;
        RECT 495.600 56.000 496.400 59.800 ;
        RECT 498.800 56.000 499.600 59.800 ;
        RECT 495.600 55.800 499.600 56.000 ;
        RECT 500.400 55.800 501.200 59.800 ;
        RECT 502.000 56.000 502.800 59.800 ;
        RECT 505.200 56.000 506.000 59.800 ;
        RECT 507.400 58.400 508.200 59.800 ;
        RECT 506.800 57.600 508.200 58.400 ;
        RECT 502.000 55.800 506.000 56.000 ;
        RECT 507.400 56.400 508.200 57.600 ;
        RECT 507.400 55.800 509.200 56.400 ;
        RECT 511.600 55.800 512.400 59.800 ;
        RECT 513.200 56.000 514.000 59.800 ;
        RECT 516.400 56.000 517.200 59.800 ;
        RECT 519.600 56.400 520.400 59.800 ;
        RECT 513.200 55.800 517.200 56.000 ;
        RECT 489.200 54.000 490.400 54.600 ;
        RECT 485.400 52.600 489.200 53.400 ;
        RECT 460.200 52.000 461.000 52.200 ;
        RECT 462.000 52.000 462.800 52.400 ;
        RECT 465.200 52.000 466.000 52.400 ;
        RECT 482.800 52.000 483.600 52.600 ;
        RECT 489.800 52.000 490.400 54.000 ;
        RECT 460.200 51.400 483.600 52.000 ;
        RECT 489.600 51.400 490.400 52.000 ;
        RECT 489.600 49.600 490.200 51.400 ;
        RECT 491.000 50.800 491.800 55.200 ;
        RECT 494.200 54.400 494.800 55.800 ;
        RECT 495.800 55.400 499.400 55.800 ;
        RECT 498.000 54.400 498.800 54.800 ;
        RECT 500.600 54.400 501.200 55.800 ;
        RECT 502.200 55.400 505.800 55.800 ;
        RECT 504.400 54.400 505.200 54.800 ;
        RECT 492.400 54.300 493.200 54.400 ;
        RECT 494.000 54.300 496.600 54.400 ;
        RECT 492.400 53.700 496.600 54.300 ;
        RECT 498.000 53.800 499.600 54.400 ;
        RECT 492.400 53.600 493.200 53.700 ;
        RECT 494.000 53.600 496.600 53.700 ;
        RECT 498.800 53.600 499.600 53.800 ;
        RECT 500.400 53.600 503.000 54.400 ;
        RECT 504.400 53.800 506.000 54.400 ;
        RECT 505.200 53.600 506.000 53.800 ;
        RECT 468.400 49.400 469.200 49.600 ;
        RECT 463.800 49.000 469.200 49.400 ;
        RECT 463.000 48.800 469.200 49.000 ;
        RECT 470.200 49.000 478.800 49.600 ;
        RECT 460.400 48.000 462.000 48.800 ;
        RECT 463.000 48.200 464.400 48.800 ;
        RECT 470.200 48.200 470.800 49.000 ;
        RECT 478.000 48.800 478.800 49.000 ;
        RECT 481.200 49.000 490.200 49.600 ;
        RECT 481.200 48.800 482.000 49.000 ;
        RECT 461.400 47.600 462.000 48.000 ;
        RECT 465.000 47.600 470.800 48.200 ;
        RECT 471.400 47.600 474.000 48.400 ;
        RECT 458.800 46.800 460.800 47.400 ;
        RECT 461.400 46.800 465.600 47.600 ;
        RECT 460.200 46.200 460.800 46.800 ;
        RECT 460.200 45.600 461.200 46.200 ;
        RECT 460.400 42.200 461.200 45.600 ;
        RECT 463.600 42.200 464.400 46.800 ;
        RECT 466.800 42.200 467.600 45.000 ;
        RECT 468.400 42.200 469.200 45.000 ;
        RECT 470.000 42.200 470.800 47.000 ;
        RECT 473.200 42.200 474.000 47.000 ;
        RECT 476.400 42.200 477.200 48.400 ;
        RECT 484.400 47.600 487.000 48.400 ;
        RECT 479.600 46.800 483.800 47.600 ;
        RECT 478.000 42.200 478.800 45.000 ;
        RECT 479.600 42.200 480.400 45.000 ;
        RECT 481.200 42.200 482.000 45.000 ;
        RECT 484.400 42.200 485.200 47.600 ;
        RECT 489.600 47.400 490.200 49.000 ;
        RECT 487.600 46.800 490.200 47.400 ;
        RECT 490.800 50.000 491.800 50.800 ;
        RECT 494.000 50.200 494.800 50.400 ;
        RECT 496.000 50.200 496.600 53.600 ;
        RECT 497.200 52.300 498.000 53.200 ;
        RECT 498.800 52.300 499.600 52.400 ;
        RECT 497.200 51.700 499.600 52.300 ;
        RECT 497.200 51.600 498.000 51.700 ;
        RECT 498.800 51.600 499.600 51.700 ;
        RECT 500.400 50.200 501.200 50.400 ;
        RECT 502.400 50.200 503.000 53.600 ;
        RECT 503.600 51.600 504.400 53.200 ;
        RECT 487.600 42.200 488.400 46.800 ;
        RECT 490.800 42.200 491.600 50.000 ;
        RECT 494.000 49.600 495.400 50.200 ;
        RECT 496.000 49.600 497.000 50.200 ;
        RECT 500.400 49.600 501.800 50.200 ;
        RECT 502.400 49.600 503.400 50.200 ;
        RECT 494.800 48.400 495.400 49.600 ;
        RECT 494.800 47.600 495.600 48.400 ;
        RECT 496.200 42.200 497.000 49.600 ;
        RECT 501.200 48.400 501.800 49.600 ;
        RECT 501.200 47.600 502.000 48.400 ;
        RECT 502.600 42.200 503.400 49.600 ;
        RECT 506.800 47.600 507.600 50.400 ;
        RECT 508.400 42.200 509.200 55.800 ;
        RECT 510.000 53.600 510.800 55.200 ;
        RECT 511.800 54.400 512.400 55.800 ;
        RECT 513.400 55.400 517.000 55.800 ;
        RECT 519.400 55.600 520.400 56.400 ;
        RECT 515.600 54.400 516.400 54.800 ;
        RECT 519.400 54.400 520.000 55.600 ;
        RECT 522.800 55.200 523.600 59.800 ;
        RECT 527.000 58.400 527.800 59.800 ;
        RECT 526.000 57.600 527.800 58.400 ;
        RECT 527.000 56.400 527.800 57.600 ;
        RECT 526.000 55.800 527.800 56.400 ;
        RECT 529.200 56.000 530.000 59.800 ;
        RECT 532.400 56.000 533.200 59.800 ;
        RECT 529.200 55.800 533.200 56.000 ;
        RECT 534.000 55.800 534.800 59.800 ;
        RECT 535.600 55.800 536.400 59.800 ;
        RECT 537.200 56.000 538.000 59.800 ;
        RECT 540.400 56.000 541.200 59.800 ;
        RECT 545.800 56.000 546.600 59.000 ;
        RECT 550.000 57.000 550.800 59.000 ;
        RECT 537.200 55.800 541.200 56.000 ;
        RECT 521.000 54.600 523.600 55.200 ;
        RECT 511.600 53.600 514.200 54.400 ;
        RECT 515.600 54.300 517.200 54.400 ;
        RECT 519.400 54.300 520.400 54.400 ;
        RECT 515.600 53.800 520.400 54.300 ;
        RECT 516.400 53.700 520.400 53.800 ;
        RECT 516.400 53.600 517.200 53.700 ;
        RECT 519.400 53.600 520.400 53.700 ;
        RECT 511.600 50.200 512.400 50.400 ;
        RECT 513.600 50.200 514.200 53.600 ;
        RECT 514.800 51.600 515.600 53.200 ;
        RECT 519.400 50.200 520.000 53.600 ;
        RECT 521.000 53.000 521.600 54.600 ;
        RECT 524.400 53.600 525.200 55.200 ;
        RECT 520.600 52.200 521.600 53.000 ;
        RECT 521.000 50.200 521.600 52.200 ;
        RECT 522.600 52.400 523.400 53.200 ;
        RECT 522.600 51.600 523.600 52.400 ;
        RECT 511.600 49.600 513.000 50.200 ;
        RECT 513.600 49.600 514.600 50.200 ;
        RECT 512.400 48.400 513.000 49.600 ;
        RECT 512.400 47.600 513.200 48.400 ;
        RECT 513.800 44.400 514.600 49.600 ;
        RECT 519.400 49.200 520.400 50.200 ;
        RECT 521.000 49.600 523.600 50.200 ;
        RECT 513.800 43.600 515.600 44.400 ;
        RECT 513.800 42.200 514.600 43.600 ;
        RECT 519.600 42.200 520.400 49.200 ;
        RECT 522.800 42.200 523.600 49.600 ;
        RECT 526.000 42.200 526.800 55.800 ;
        RECT 529.400 55.400 533.000 55.800 ;
        RECT 530.000 54.400 530.800 54.800 ;
        RECT 534.000 54.400 534.600 55.800 ;
        RECT 535.800 54.400 536.400 55.800 ;
        RECT 537.400 55.400 541.000 55.800 ;
        RECT 545.000 55.400 546.600 56.000 ;
        RECT 545.000 55.000 545.800 55.400 ;
        RECT 539.600 54.400 540.400 54.800 ;
        RECT 545.000 54.400 545.600 55.000 ;
        RECT 550.200 54.800 550.800 57.000 ;
        RECT 551.600 56.000 552.400 59.800 ;
        RECT 554.800 56.000 555.600 59.800 ;
        RECT 551.600 55.800 555.600 56.000 ;
        RECT 556.400 55.800 557.200 59.800 ;
        RECT 560.600 58.400 561.400 59.800 ;
        RECT 560.600 57.600 562.000 58.400 ;
        RECT 560.600 56.400 561.400 57.600 ;
        RECT 559.600 55.800 561.400 56.400 ;
        RECT 562.800 55.800 563.600 59.800 ;
        RECT 564.400 56.000 565.200 59.800 ;
        RECT 567.600 56.000 568.400 59.800 ;
        RECT 564.400 55.800 568.400 56.000 ;
        RECT 574.000 55.800 574.800 59.800 ;
        RECT 578.400 58.400 580.000 59.800 ;
        RECT 578.400 57.600 581.200 58.400 ;
        RECT 578.400 56.200 580.000 57.600 ;
        RECT 551.800 55.400 555.400 55.800 ;
        RECT 529.200 53.800 530.800 54.400 ;
        RECT 529.200 53.600 530.000 53.800 ;
        RECT 532.200 53.600 534.800 54.400 ;
        RECT 535.600 53.600 538.200 54.400 ;
        RECT 539.600 53.800 541.200 54.400 ;
        RECT 540.400 53.600 541.200 53.800 ;
        RECT 543.600 53.600 545.600 54.400 ;
        RECT 546.600 54.200 550.800 54.800 ;
        RECT 552.400 54.400 553.200 54.800 ;
        RECT 556.400 54.400 557.000 55.800 ;
        RECT 546.600 53.800 547.600 54.200 ;
        RECT 530.800 51.600 531.600 53.200 ;
        RECT 532.200 52.300 532.800 53.600 ;
        RECT 532.200 51.700 536.300 52.300 ;
        RECT 527.600 47.600 528.400 50.400 ;
        RECT 532.200 50.200 532.800 51.700 ;
        RECT 535.700 50.400 536.300 51.700 ;
        RECT 534.000 50.200 534.800 50.400 ;
        RECT 531.800 49.600 532.800 50.200 ;
        RECT 533.400 49.600 534.800 50.200 ;
        RECT 535.600 50.200 536.400 50.400 ;
        RECT 537.600 50.200 538.200 53.600 ;
        RECT 538.800 51.600 539.600 53.200 ;
        RECT 540.400 52.300 541.200 52.400 ;
        RECT 542.000 52.300 542.800 52.400 ;
        RECT 543.600 52.300 544.400 52.400 ;
        RECT 540.400 51.700 544.400 52.300 ;
        RECT 540.400 51.600 541.200 51.700 ;
        RECT 542.000 51.600 542.800 51.700 ;
        RECT 543.600 50.800 544.400 51.700 ;
        RECT 535.600 49.600 537.000 50.200 ;
        RECT 537.600 49.600 538.600 50.200 ;
        RECT 531.800 42.200 532.600 49.600 ;
        RECT 533.400 48.400 534.000 49.600 ;
        RECT 533.200 47.600 534.000 48.400 ;
        RECT 536.400 48.400 537.000 49.600 ;
        RECT 536.400 47.600 537.200 48.400 ;
        RECT 537.800 42.200 538.600 49.600 ;
        RECT 545.000 49.800 545.600 53.600 ;
        RECT 546.200 53.000 547.600 53.800 ;
        RECT 551.600 53.800 553.200 54.400 ;
        RECT 551.600 53.600 552.400 53.800 ;
        RECT 554.600 53.600 557.200 54.400 ;
        RECT 558.000 53.600 558.800 55.200 ;
        RECT 547.000 51.000 547.600 53.000 ;
        RECT 548.400 51.600 549.200 53.200 ;
        RECT 550.000 51.600 550.800 53.200 ;
        RECT 553.200 51.600 554.000 53.200 ;
        RECT 554.600 52.400 555.200 53.600 ;
        RECT 554.600 51.600 555.600 52.400 ;
        RECT 547.000 50.400 550.800 51.000 ;
        RECT 545.000 49.200 546.600 49.800 ;
        RECT 545.800 42.200 546.600 49.200 ;
        RECT 550.200 47.000 550.800 50.400 ;
        RECT 554.600 50.200 555.200 51.600 ;
        RECT 556.400 50.200 557.200 50.400 ;
        RECT 550.000 43.000 550.800 47.000 ;
        RECT 554.200 49.600 555.200 50.200 ;
        RECT 555.800 49.600 557.200 50.200 ;
        RECT 554.200 42.200 555.000 49.600 ;
        RECT 555.800 48.400 556.400 49.600 ;
        RECT 555.600 47.600 556.400 48.400 ;
        RECT 559.600 42.200 560.400 55.800 ;
        RECT 563.000 54.400 563.600 55.800 ;
        RECT 564.600 55.400 568.200 55.800 ;
        RECT 574.000 55.200 576.400 55.800 ;
        RECT 575.600 55.000 576.400 55.200 ;
        RECT 577.000 54.800 577.800 55.600 ;
        RECT 566.800 54.400 567.600 54.800 ;
        RECT 577.000 54.400 577.600 54.800 ;
        RECT 562.800 53.600 565.400 54.400 ;
        RECT 566.800 53.800 568.400 54.400 ;
        RECT 567.600 53.600 568.400 53.800 ;
        RECT 569.200 54.300 570.000 54.400 ;
        RECT 574.000 54.300 575.600 54.400 ;
        RECT 569.200 53.700 575.600 54.300 ;
        RECT 569.200 53.600 570.000 53.700 ;
        RECT 574.000 53.600 575.600 53.700 ;
        RECT 576.800 53.600 577.600 54.400 ;
        RECT 578.400 54.200 579.000 56.200 ;
        RECT 583.600 55.800 584.400 59.800 ;
        RECT 585.800 58.400 586.600 59.800 ;
        RECT 585.200 57.600 586.600 58.400 ;
        RECT 585.800 56.400 586.600 57.600 ;
        RECT 585.800 55.800 587.600 56.400 ;
        RECT 593.800 56.000 594.600 59.000 ;
        RECT 598.000 57.000 598.800 59.000 ;
        RECT 579.600 54.800 581.200 55.600 ;
        RECT 581.800 55.200 584.400 55.800 ;
        RECT 581.800 55.000 582.600 55.200 ;
        RECT 582.800 54.200 584.400 54.400 ;
        RECT 578.400 53.600 579.400 54.200 ;
        RECT 582.200 54.000 584.400 54.200 ;
        RECT 561.200 48.800 562.000 50.400 ;
        RECT 562.800 50.200 563.600 50.400 ;
        RECT 564.800 50.200 565.400 53.600 ;
        RECT 566.000 51.600 566.800 53.200 ;
        RECT 578.800 52.400 579.400 53.600 ;
        RECT 580.000 53.600 584.400 54.000 ;
        RECT 580.000 53.400 582.800 53.600 ;
        RECT 580.000 53.200 580.800 53.400 ;
        RECT 578.800 51.600 579.600 52.400 ;
        RECT 581.400 52.200 582.200 52.400 ;
        RECT 580.600 51.600 582.200 52.200 ;
        RECT 578.800 50.200 579.400 51.600 ;
        RECT 580.600 51.400 581.400 51.600 ;
        RECT 562.800 49.600 564.200 50.200 ;
        RECT 564.800 49.600 565.800 50.200 ;
        RECT 563.600 48.400 564.200 49.600 ;
        RECT 563.600 47.600 564.400 48.400 ;
        RECT 565.000 44.400 565.800 49.600 ;
        RECT 574.000 49.600 576.400 50.200 ;
        RECT 565.000 43.600 566.800 44.400 ;
        RECT 565.000 42.200 565.800 43.600 ;
        RECT 574.000 42.200 574.800 49.600 ;
        RECT 575.600 49.400 576.400 49.600 ;
        RECT 578.400 42.200 580.000 50.200 ;
        RECT 581.800 49.600 584.400 50.200 ;
        RECT 581.800 49.400 582.600 49.600 ;
        RECT 583.600 42.200 584.400 49.600 ;
        RECT 585.200 48.800 586.000 50.400 ;
        RECT 586.800 42.200 587.600 55.800 ;
        RECT 593.000 55.400 594.600 56.000 ;
        RECT 588.400 53.600 589.200 55.200 ;
        RECT 593.000 55.000 593.800 55.400 ;
        RECT 593.000 54.400 593.600 55.000 ;
        RECT 598.200 54.800 598.800 57.000 ;
        RECT 591.600 53.600 593.600 54.400 ;
        RECT 594.600 54.200 598.800 54.800 ;
        RECT 599.600 55.400 600.400 59.800 ;
        RECT 603.800 58.400 605.000 59.800 ;
        RECT 603.800 57.800 605.200 58.400 ;
        RECT 608.400 57.800 609.200 59.800 ;
        RECT 612.800 58.400 613.600 59.800 ;
        RECT 612.800 57.800 614.800 58.400 ;
        RECT 604.400 57.000 605.200 57.800 ;
        RECT 608.600 57.200 609.200 57.800 ;
        RECT 608.600 56.600 611.400 57.200 ;
        RECT 610.600 56.400 611.400 56.600 ;
        RECT 612.400 55.600 613.200 57.200 ;
        RECT 614.000 57.000 614.800 57.800 ;
        RECT 602.600 55.400 603.400 55.600 ;
        RECT 599.600 54.800 603.400 55.400 ;
        RECT 594.600 53.800 595.600 54.200 ;
        RECT 591.600 50.800 592.400 52.400 ;
        RECT 593.000 49.800 593.600 53.600 ;
        RECT 594.200 53.000 595.600 53.800 ;
        RECT 595.000 51.000 595.600 53.000 ;
        RECT 596.400 51.600 597.200 53.200 ;
        RECT 598.000 51.600 598.800 53.200 ;
        RECT 599.600 51.400 600.400 54.800 ;
        RECT 606.600 54.200 607.400 54.400 ;
        RECT 612.400 54.200 613.000 55.600 ;
        RECT 617.200 55.000 618.000 59.800 ;
        RECT 618.800 57.000 619.600 59.000 ;
        RECT 618.800 54.800 619.400 57.000 ;
        RECT 623.000 56.000 623.800 59.000 ;
        RECT 630.000 56.400 630.800 59.800 ;
        RECT 623.000 55.400 624.600 56.000 ;
        RECT 623.800 55.000 624.600 55.400 ;
        RECT 615.600 54.200 617.200 54.400 ;
        RECT 618.800 54.200 623.000 54.800 ;
        RECT 606.200 53.600 617.200 54.200 ;
        RECT 622.000 53.800 623.000 54.200 ;
        RECT 624.000 54.400 624.600 55.000 ;
        RECT 629.800 55.800 630.800 56.400 ;
        RECT 629.800 54.400 630.400 55.800 ;
        RECT 633.200 55.200 634.000 59.800 ;
        RECT 631.400 54.600 634.000 55.200 ;
        RECT 634.800 57.000 635.600 59.000 ;
        RECT 634.800 54.800 635.400 57.000 ;
        RECT 639.000 56.000 639.800 59.000 ;
        RECT 639.000 55.400 640.600 56.000 ;
        RECT 644.400 55.800 645.200 59.800 ;
        RECT 646.000 56.000 646.800 59.800 ;
        RECT 649.200 56.000 650.000 59.800 ;
        RECT 646.000 55.800 650.000 56.000 ;
        RECT 650.800 55.800 651.600 59.800 ;
        RECT 652.400 56.000 653.200 59.800 ;
        RECT 655.600 56.000 656.400 59.800 ;
        RECT 661.000 56.000 661.800 59.000 ;
        RECT 665.200 57.000 666.000 59.000 ;
        RECT 652.400 55.800 656.400 56.000 ;
        RECT 639.800 55.000 640.600 55.400 ;
        RECT 624.000 54.300 626.000 54.400 ;
        RECT 626.800 54.300 627.600 54.400 ;
        RECT 604.400 52.800 605.200 53.000 ;
        RECT 601.400 52.200 605.200 52.800 ;
        RECT 601.400 52.000 602.200 52.200 ;
        RECT 603.000 51.400 603.800 51.600 ;
        RECT 595.000 50.400 598.800 51.000 ;
        RECT 593.000 49.200 594.600 49.800 ;
        RECT 593.800 44.400 594.600 49.200 ;
        RECT 598.200 47.000 598.800 50.400 ;
        RECT 593.200 43.600 594.600 44.400 ;
        RECT 593.800 42.200 594.600 43.600 ;
        RECT 598.000 43.000 598.800 47.000 ;
        RECT 599.600 50.800 603.800 51.400 ;
        RECT 599.600 42.200 600.400 50.800 ;
        RECT 606.200 50.400 606.800 53.600 ;
        RECT 613.400 53.400 614.200 53.600 ;
        RECT 612.400 52.400 613.200 52.600 ;
        RECT 615.000 52.400 615.800 52.600 ;
        RECT 610.800 51.800 615.800 52.400 ;
        RECT 610.800 51.600 611.600 51.800 ;
        RECT 618.800 51.600 619.600 53.200 ;
        RECT 620.400 51.600 621.200 53.200 ;
        RECT 622.000 53.000 623.400 53.800 ;
        RECT 624.000 53.700 627.600 54.300 ;
        RECT 624.000 53.600 626.000 53.700 ;
        RECT 626.800 53.600 627.600 53.700 ;
        RECT 629.800 53.600 630.800 54.400 ;
        RECT 612.400 51.000 618.000 51.200 ;
        RECT 622.000 51.000 622.600 53.000 ;
        RECT 612.200 50.800 618.000 51.000 ;
        RECT 604.400 49.800 606.800 50.400 ;
        RECT 608.200 50.600 618.000 50.800 ;
        RECT 608.200 50.200 613.000 50.600 ;
        RECT 604.400 48.800 605.000 49.800 ;
        RECT 603.600 48.000 605.000 48.800 ;
        RECT 606.600 49.000 607.400 49.200 ;
        RECT 608.200 49.000 608.800 50.200 ;
        RECT 606.600 48.400 608.800 49.000 ;
        RECT 609.400 49.000 614.800 49.600 ;
        RECT 609.400 48.800 610.200 49.000 ;
        RECT 614.000 48.800 614.800 49.000 ;
        RECT 607.800 47.400 608.600 47.600 ;
        RECT 610.600 47.400 611.400 47.600 ;
        RECT 604.400 46.200 605.200 47.000 ;
        RECT 607.800 46.800 611.400 47.400 ;
        RECT 608.600 46.200 609.200 46.800 ;
        RECT 614.000 46.200 614.800 47.000 ;
        RECT 603.800 42.200 605.000 46.200 ;
        RECT 608.400 42.200 609.200 46.200 ;
        RECT 612.800 45.600 614.800 46.200 ;
        RECT 612.800 42.200 613.600 45.600 ;
        RECT 617.200 42.200 618.000 50.600 ;
        RECT 618.800 50.400 622.600 51.000 ;
        RECT 618.800 47.000 619.400 50.400 ;
        RECT 624.000 49.800 624.600 53.600 ;
        RECT 625.200 50.800 626.000 52.400 ;
        RECT 623.000 49.200 624.600 49.800 ;
        RECT 629.800 50.200 630.400 53.600 ;
        RECT 631.400 53.000 632.000 54.600 ;
        RECT 634.800 54.200 639.000 54.800 ;
        RECT 638.000 53.800 639.000 54.200 ;
        RECT 640.000 54.400 640.600 55.000 ;
        RECT 644.600 54.400 645.200 55.800 ;
        RECT 646.200 55.400 649.800 55.800 ;
        RECT 648.400 54.400 649.200 54.800 ;
        RECT 651.000 54.400 651.600 55.800 ;
        RECT 652.600 55.400 656.200 55.800 ;
        RECT 660.200 55.400 661.800 56.000 ;
        RECT 660.200 55.000 661.000 55.400 ;
        RECT 654.800 54.400 655.600 54.800 ;
        RECT 660.200 54.400 660.800 55.000 ;
        RECT 665.400 54.800 666.000 57.000 ;
        RECT 631.000 52.200 632.000 53.000 ;
        RECT 631.400 50.200 632.000 52.200 ;
        RECT 633.000 52.400 633.800 53.200 ;
        RECT 633.000 51.600 634.000 52.400 ;
        RECT 634.800 51.600 635.600 53.200 ;
        RECT 636.400 51.600 637.200 53.200 ;
        RECT 638.000 53.000 639.400 53.800 ;
        RECT 640.000 53.600 642.000 54.400 ;
        RECT 644.400 53.600 647.000 54.400 ;
        RECT 648.400 53.800 650.000 54.400 ;
        RECT 649.200 53.600 650.000 53.800 ;
        RECT 650.800 53.600 653.400 54.400 ;
        RECT 654.800 53.800 656.400 54.400 ;
        RECT 655.600 53.600 656.400 53.800 ;
        RECT 658.800 53.600 660.800 54.400 ;
        RECT 661.800 54.200 666.000 54.800 ;
        RECT 666.800 57.000 667.600 59.000 ;
        RECT 666.800 54.800 667.400 57.000 ;
        RECT 671.000 56.000 671.800 59.000 ;
        RECT 676.400 56.000 677.200 59.800 ;
        RECT 679.600 56.000 680.400 59.800 ;
        RECT 671.000 55.400 672.600 56.000 ;
        RECT 676.400 55.800 680.400 56.000 ;
        RECT 681.200 55.800 682.000 59.800 ;
        RECT 682.800 55.800 683.600 59.800 ;
        RECT 684.400 56.000 685.200 59.800 ;
        RECT 687.600 56.000 688.400 59.800 ;
        RECT 684.400 55.800 688.400 56.000 ;
        RECT 676.600 55.400 680.200 55.800 ;
        RECT 671.800 55.000 672.600 55.400 ;
        RECT 666.800 54.200 671.000 54.800 ;
        RECT 661.800 53.800 662.800 54.200 ;
        RECT 638.000 51.000 638.600 53.000 ;
        RECT 634.800 50.400 638.600 51.000 ;
        RECT 629.800 49.200 630.800 50.200 ;
        RECT 631.400 49.600 634.000 50.200 ;
        RECT 618.800 43.000 619.600 47.000 ;
        RECT 623.000 42.200 623.800 49.200 ;
        RECT 630.000 42.200 630.800 49.200 ;
        RECT 633.200 42.200 634.000 49.600 ;
        RECT 634.800 47.000 635.400 50.400 ;
        RECT 640.000 49.800 640.600 53.600 ;
        RECT 641.200 50.800 642.000 52.400 ;
        RECT 639.000 49.200 640.600 49.800 ;
        RECT 644.400 50.200 645.200 50.400 ;
        RECT 646.400 50.200 647.000 53.600 ;
        RECT 647.600 52.300 648.400 53.200 ;
        RECT 650.800 52.300 651.600 52.400 ;
        RECT 647.600 51.700 651.600 52.300 ;
        RECT 647.600 51.600 648.400 51.700 ;
        RECT 650.800 51.600 651.600 51.700 ;
        RECT 650.800 50.200 651.600 50.400 ;
        RECT 652.800 50.200 653.400 53.600 ;
        RECT 654.000 51.600 654.800 53.200 ;
        RECT 658.800 50.800 659.600 52.400 ;
        RECT 644.400 49.600 645.800 50.200 ;
        RECT 646.400 49.600 647.400 50.200 ;
        RECT 650.800 49.600 652.200 50.200 ;
        RECT 652.800 49.600 653.800 50.200 ;
        RECT 634.800 43.000 635.600 47.000 ;
        RECT 639.000 44.400 639.800 49.200 ;
        RECT 645.200 48.400 645.800 49.600 ;
        RECT 646.600 48.400 647.400 49.600 ;
        RECT 651.600 48.400 652.200 49.600 ;
        RECT 645.200 47.600 646.000 48.400 ;
        RECT 646.600 47.600 648.400 48.400 ;
        RECT 651.600 47.600 652.400 48.400 ;
        RECT 639.000 43.600 640.400 44.400 ;
        RECT 639.000 42.200 639.800 43.600 ;
        RECT 646.600 42.200 647.400 47.600 ;
        RECT 653.000 42.200 653.800 49.600 ;
        RECT 660.200 49.800 660.800 53.600 ;
        RECT 661.400 53.000 662.800 53.800 ;
        RECT 670.000 53.800 671.000 54.200 ;
        RECT 672.000 54.400 672.600 55.000 ;
        RECT 677.200 54.400 678.000 54.800 ;
        RECT 681.200 54.400 681.800 55.800 ;
        RECT 683.000 54.400 683.600 55.800 ;
        RECT 684.600 55.400 688.200 55.800 ;
        RECT 686.800 54.400 687.600 54.800 ;
        RECT 662.200 51.000 662.800 53.000 ;
        RECT 663.600 51.600 664.400 53.200 ;
        RECT 665.200 51.600 666.000 53.200 ;
        RECT 666.800 51.600 667.600 53.200 ;
        RECT 668.400 51.600 669.200 53.200 ;
        RECT 670.000 53.000 671.400 53.800 ;
        RECT 672.000 53.600 674.000 54.400 ;
        RECT 674.800 54.300 675.600 54.400 ;
        RECT 676.400 54.300 678.000 54.400 ;
        RECT 674.800 53.800 678.000 54.300 ;
        RECT 674.800 53.700 677.200 53.800 ;
        RECT 674.800 53.600 675.600 53.700 ;
        RECT 676.400 53.600 677.200 53.700 ;
        RECT 679.400 53.600 682.000 54.400 ;
        RECT 682.800 53.600 685.400 54.400 ;
        RECT 686.800 53.800 688.400 54.400 ;
        RECT 687.600 53.600 688.400 53.800 ;
        RECT 670.000 51.000 670.600 53.000 ;
        RECT 662.200 50.400 666.000 51.000 ;
        RECT 660.200 49.200 661.800 49.800 ;
        RECT 661.000 44.400 661.800 49.200 ;
        RECT 665.400 47.000 666.000 50.400 ;
        RECT 661.000 43.600 662.800 44.400 ;
        RECT 661.000 42.200 661.800 43.600 ;
        RECT 665.200 43.000 666.000 47.000 ;
        RECT 666.800 50.400 670.600 51.000 ;
        RECT 666.800 47.000 667.400 50.400 ;
        RECT 672.000 49.800 672.600 53.600 ;
        RECT 673.200 52.300 674.000 52.400 ;
        RECT 676.400 52.300 677.200 52.400 ;
        RECT 673.200 51.700 677.200 52.300 ;
        RECT 673.200 50.800 674.000 51.700 ;
        RECT 676.400 51.600 677.200 51.700 ;
        RECT 678.000 51.600 678.800 53.200 ;
        RECT 679.400 52.300 680.000 53.600 ;
        RECT 679.400 51.700 683.500 52.300 ;
        RECT 679.400 50.200 680.000 51.700 ;
        RECT 682.900 50.400 683.500 51.700 ;
        RECT 681.200 50.200 682.000 50.400 ;
        RECT 671.000 49.200 672.600 49.800 ;
        RECT 679.000 49.600 680.000 50.200 ;
        RECT 680.600 49.600 682.000 50.200 ;
        RECT 682.800 50.200 683.600 50.400 ;
        RECT 684.800 50.200 685.400 53.600 ;
        RECT 686.000 51.600 686.800 53.200 ;
        RECT 682.800 49.600 684.200 50.200 ;
        RECT 684.800 49.600 685.800 50.200 ;
        RECT 666.800 43.000 667.600 47.000 ;
        RECT 671.000 42.200 671.800 49.200 ;
        RECT 679.000 42.200 679.800 49.600 ;
        RECT 680.600 48.400 681.200 49.600 ;
        RECT 680.400 47.600 681.200 48.400 ;
        RECT 683.600 48.400 684.200 49.600 ;
        RECT 683.600 47.600 684.400 48.400 ;
        RECT 685.000 42.200 685.800 49.600 ;
        RECT 2.800 36.400 3.600 39.800 ;
        RECT 2.600 35.800 3.600 36.400 ;
        RECT 2.600 35.200 3.200 35.800 ;
        RECT 6.000 35.200 6.800 39.800 ;
        RECT 9.200 37.000 10.000 39.800 ;
        RECT 10.800 37.000 11.600 39.800 ;
        RECT 1.200 34.600 3.200 35.200 ;
        RECT 1.200 29.000 2.000 34.600 ;
        RECT 3.800 34.400 8.000 35.200 ;
        RECT 12.400 35.000 13.200 39.800 ;
        RECT 15.600 35.000 16.400 39.800 ;
        RECT 3.800 34.000 4.400 34.400 ;
        RECT 2.800 33.200 4.400 34.000 ;
        RECT 7.400 33.800 13.200 34.400 ;
        RECT 5.400 33.200 6.800 33.800 ;
        RECT 5.400 33.000 11.600 33.200 ;
        RECT 6.200 32.600 11.600 33.000 ;
        RECT 10.800 32.400 11.600 32.600 ;
        RECT 12.600 33.000 13.200 33.800 ;
        RECT 13.800 33.600 16.400 34.400 ;
        RECT 18.800 33.600 19.600 39.800 ;
        RECT 20.400 37.000 21.200 39.800 ;
        RECT 22.000 37.000 22.800 39.800 ;
        RECT 23.600 37.000 24.400 39.800 ;
        RECT 22.000 34.400 26.200 35.200 ;
        RECT 26.800 34.400 27.600 39.800 ;
        RECT 30.000 35.200 30.800 39.800 ;
        RECT 30.000 34.600 32.600 35.200 ;
        RECT 26.800 33.600 29.400 34.400 ;
        RECT 20.400 33.000 21.200 33.200 ;
        RECT 12.600 32.400 21.200 33.000 ;
        RECT 23.600 33.000 24.400 33.200 ;
        RECT 32.000 33.000 32.600 34.600 ;
        RECT 23.600 32.400 32.600 33.000 ;
        RECT 32.000 30.600 32.600 32.400 ;
        RECT 33.200 32.000 34.000 39.800 ;
        RECT 33.200 31.200 34.200 32.000 ;
        RECT 2.600 30.000 26.000 30.600 ;
        RECT 32.000 30.000 32.800 30.600 ;
        RECT 2.600 29.800 3.400 30.000 ;
        RECT 7.600 29.600 8.400 30.000 ;
        RECT 25.200 29.400 26.000 30.000 ;
        RECT 1.200 28.200 10.000 29.000 ;
        RECT 10.600 28.600 12.600 29.400 ;
        RECT 16.400 28.600 19.600 29.400 ;
        RECT 1.200 22.200 2.000 28.200 ;
        RECT 3.600 26.800 6.600 27.600 ;
        RECT 5.800 26.200 6.600 26.800 ;
        RECT 11.800 26.200 12.600 28.600 ;
        RECT 14.000 26.800 14.800 28.400 ;
        RECT 19.200 27.800 20.000 28.000 ;
        RECT 15.600 27.200 20.000 27.800 ;
        RECT 15.600 27.000 16.400 27.200 ;
        RECT 22.000 26.400 22.800 29.200 ;
        RECT 27.800 28.600 31.600 29.400 ;
        RECT 27.800 27.400 28.600 28.600 ;
        RECT 32.200 28.000 32.800 30.000 ;
        RECT 15.600 26.200 16.400 26.400 ;
        RECT 5.800 25.400 8.400 26.200 ;
        RECT 11.800 25.600 16.400 26.200 ;
        RECT 17.200 25.600 18.800 26.400 ;
        RECT 21.800 25.600 22.800 26.400 ;
        RECT 26.800 26.800 28.600 27.400 ;
        RECT 31.600 27.400 32.800 28.000 ;
        RECT 26.800 26.200 27.600 26.800 ;
        RECT 7.600 22.200 8.400 25.400 ;
        RECT 25.200 25.400 27.600 26.200 ;
        RECT 9.200 22.200 10.000 25.000 ;
        RECT 10.800 22.200 11.600 25.000 ;
        RECT 12.400 22.200 13.200 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 18.800 22.200 19.600 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 22.000 22.200 22.800 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.400 ;
        RECT 31.600 22.200 32.400 27.400 ;
        RECT 33.400 26.800 34.200 31.200 ;
        RECT 33.200 26.000 34.200 26.800 ;
        RECT 38.000 28.300 38.800 39.800 ;
        RECT 42.200 32.400 43.000 39.800 ;
        RECT 43.600 33.600 44.400 34.400 ;
        RECT 43.800 32.400 44.400 33.600 ;
        RECT 46.800 33.600 47.600 34.400 ;
        RECT 46.800 32.400 47.400 33.600 ;
        RECT 48.200 32.400 49.000 39.800 ;
        RECT 42.200 31.800 43.200 32.400 ;
        RECT 43.800 31.800 45.200 32.400 ;
        RECT 41.200 28.800 42.000 30.400 ;
        RECT 42.600 28.400 43.200 31.800 ;
        RECT 44.400 31.600 45.200 31.800 ;
        RECT 46.000 31.800 47.400 32.400 ;
        RECT 48.000 31.800 49.000 32.400 ;
        RECT 55.000 32.400 55.800 39.800 ;
        RECT 56.400 33.600 57.200 34.400 ;
        RECT 56.600 32.400 57.200 33.600 ;
        RECT 61.400 32.400 62.200 39.800 ;
        RECT 62.800 33.600 63.600 34.400 ;
        RECT 63.000 32.400 63.600 33.600 ;
        RECT 55.000 31.800 56.000 32.400 ;
        RECT 56.600 31.800 58.000 32.400 ;
        RECT 61.400 31.800 62.400 32.400 ;
        RECT 63.000 31.800 64.400 32.400 ;
        RECT 46.000 31.600 46.800 31.800 ;
        RECT 44.500 30.300 45.100 31.600 ;
        RECT 48.000 30.300 48.600 31.800 ;
        RECT 44.500 29.700 48.600 30.300 ;
        RECT 48.000 28.400 48.600 29.700 ;
        RECT 49.200 30.300 50.000 30.400 ;
        RECT 50.800 30.300 51.600 30.400 ;
        RECT 54.000 30.300 54.800 30.400 ;
        RECT 49.200 29.700 54.800 30.300 ;
        RECT 49.200 28.800 50.000 29.700 ;
        RECT 50.800 29.600 51.600 29.700 ;
        RECT 54.000 28.800 54.800 29.700 ;
        RECT 55.400 30.300 56.000 31.800 ;
        RECT 57.200 31.600 58.000 31.800 ;
        RECT 58.800 30.300 59.600 30.400 ;
        RECT 55.400 29.700 59.600 30.300 ;
        RECT 55.400 28.400 56.000 29.700 ;
        RECT 58.800 29.600 59.600 29.700 ;
        RECT 60.400 28.800 61.200 30.400 ;
        RECT 61.800 28.400 62.400 31.800 ;
        RECT 63.600 31.600 64.400 31.800 ;
        RECT 66.800 31.200 67.600 39.800 ;
        RECT 70.000 31.200 70.800 39.800 ;
        RECT 73.200 31.200 74.000 39.800 ;
        RECT 76.400 31.200 77.200 39.800 ;
        RECT 65.200 30.400 67.600 31.200 ;
        RECT 68.600 30.400 70.800 31.200 ;
        RECT 71.800 30.400 74.000 31.200 ;
        RECT 75.400 30.400 77.200 31.200 ;
        RECT 81.200 31.200 82.000 39.800 ;
        RECT 84.400 31.200 85.200 39.800 ;
        RECT 87.600 31.200 88.400 39.800 ;
        RECT 90.800 31.200 91.600 39.800 ;
        RECT 94.800 33.600 95.600 34.400 ;
        RECT 94.800 32.400 95.400 33.600 ;
        RECT 96.200 32.400 97.000 39.800 ;
        RECT 102.600 36.400 103.400 39.800 ;
        RECT 102.600 35.600 104.400 36.400 ;
        RECT 101.200 33.600 102.000 34.400 ;
        RECT 101.200 32.400 101.800 33.600 ;
        RECT 102.600 32.400 103.400 35.600 ;
        RECT 107.600 33.600 108.400 34.400 ;
        RECT 107.600 32.400 108.200 33.600 ;
        RECT 109.000 32.400 109.800 39.800 ;
        RECT 94.000 31.800 95.400 32.400 ;
        RECT 96.000 31.800 97.000 32.400 ;
        RECT 100.400 31.800 101.800 32.400 ;
        RECT 102.400 31.800 103.400 32.400 ;
        RECT 106.800 31.800 108.200 32.400 ;
        RECT 94.000 31.600 94.800 31.800 ;
        RECT 81.200 30.400 83.000 31.200 ;
        RECT 84.400 30.400 86.600 31.200 ;
        RECT 87.600 30.400 89.800 31.200 ;
        RECT 90.800 30.400 93.200 31.200 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 38.000 28.200 40.400 28.300 ;
        RECT 38.000 27.700 41.200 28.200 ;
        RECT 33.200 22.200 34.000 26.000 ;
        RECT 38.000 22.200 38.800 27.700 ;
        RECT 39.600 27.600 41.200 27.700 ;
        RECT 42.600 27.600 45.200 28.400 ;
        RECT 46.000 27.600 48.600 28.400 ;
        RECT 50.800 28.300 51.600 28.400 ;
        RECT 52.400 28.300 53.200 28.400 ;
        RECT 50.800 28.200 53.200 28.300 ;
        RECT 50.000 27.700 54.000 28.200 ;
        RECT 50.000 27.600 51.600 27.700 ;
        RECT 52.400 27.600 54.000 27.700 ;
        RECT 55.400 27.600 58.000 28.400 ;
        RECT 58.800 28.200 59.600 28.400 ;
        RECT 58.800 27.600 60.400 28.200 ;
        RECT 61.800 27.600 64.400 28.400 ;
        RECT 65.200 27.600 66.000 30.400 ;
        RECT 68.600 29.000 69.400 30.400 ;
        RECT 71.800 29.000 72.600 30.400 ;
        RECT 75.400 29.000 76.200 30.400 ;
        RECT 82.200 29.000 83.000 30.400 ;
        RECT 85.800 29.000 86.600 30.400 ;
        RECT 89.000 29.000 89.800 30.400 ;
        RECT 66.800 28.200 69.400 29.000 ;
        RECT 70.200 28.200 72.600 29.000 ;
        RECT 73.600 28.200 76.200 29.000 ;
        RECT 77.000 28.300 78.800 29.000 ;
        RECT 79.600 28.300 81.400 29.000 ;
        RECT 77.000 28.200 81.400 28.300 ;
        RECT 82.200 28.200 84.800 29.000 ;
        RECT 85.800 28.200 88.200 29.000 ;
        RECT 89.000 28.200 91.600 29.000 ;
        RECT 68.600 27.600 69.400 28.200 ;
        RECT 71.800 27.600 72.600 28.200 ;
        RECT 75.400 27.600 76.200 28.200 ;
        RECT 78.000 27.700 80.400 28.200 ;
        RECT 78.000 27.600 78.800 27.700 ;
        RECT 79.600 27.600 80.400 27.700 ;
        RECT 82.200 27.600 83.000 28.200 ;
        RECT 85.800 27.600 86.600 28.200 ;
        RECT 89.000 27.600 89.800 28.200 ;
        RECT 92.400 27.600 93.200 30.400 ;
        RECT 96.000 28.400 96.600 31.800 ;
        RECT 100.400 31.600 101.200 31.800 ;
        RECT 97.200 28.800 98.000 30.400 ;
        RECT 102.400 28.400 103.000 31.800 ;
        RECT 106.800 31.600 107.600 31.800 ;
        RECT 108.800 31.600 110.800 32.400 ;
        RECT 103.600 28.800 104.400 30.400 ;
        RECT 108.800 28.400 109.400 31.600 ;
        RECT 118.000 31.400 118.800 39.800 ;
        RECT 122.400 36.400 123.200 39.800 ;
        RECT 121.200 35.800 123.200 36.400 ;
        RECT 126.800 35.800 127.600 39.800 ;
        RECT 131.000 35.800 132.200 39.800 ;
        RECT 121.200 35.000 122.000 35.800 ;
        RECT 126.800 35.200 127.400 35.800 ;
        RECT 124.600 34.600 128.200 35.200 ;
        RECT 130.800 35.000 131.600 35.800 ;
        RECT 124.600 34.400 125.400 34.600 ;
        RECT 127.400 34.400 128.200 34.600 ;
        RECT 121.200 33.000 122.000 33.200 ;
        RECT 125.800 33.000 126.600 33.200 ;
        RECT 121.200 32.400 126.600 33.000 ;
        RECT 127.200 33.000 129.400 33.600 ;
        RECT 127.200 31.800 127.800 33.000 ;
        RECT 128.600 32.800 129.400 33.000 ;
        RECT 131.000 33.200 132.400 34.000 ;
        RECT 131.000 32.200 131.600 33.200 ;
        RECT 123.000 31.400 127.800 31.800 ;
        RECT 118.000 31.200 127.800 31.400 ;
        RECT 129.200 31.600 131.600 32.200 ;
        RECT 118.000 31.000 123.800 31.200 ;
        RECT 118.000 30.800 123.600 31.000 ;
        RECT 110.000 28.800 110.800 30.400 ;
        RECT 124.400 30.200 125.200 30.400 ;
        RECT 120.200 29.600 125.200 30.200 ;
        RECT 120.200 29.400 121.000 29.600 ;
        RECT 122.800 29.400 123.600 29.600 ;
        RECT 121.800 28.400 122.600 28.600 ;
        RECT 129.200 28.400 129.800 31.600 ;
        RECT 135.600 31.200 136.400 39.800 ;
        RECT 139.800 32.400 140.600 39.800 ;
        RECT 141.200 33.600 142.000 34.400 ;
        RECT 141.400 32.400 142.000 33.600 ;
        RECT 139.800 31.800 140.800 32.400 ;
        RECT 141.400 31.800 142.800 32.400 ;
        RECT 132.200 30.600 136.400 31.200 ;
        RECT 132.200 30.400 133.000 30.600 ;
        RECT 133.800 29.800 134.600 30.000 ;
        RECT 130.800 29.200 134.600 29.800 ;
        RECT 130.800 29.000 131.600 29.200 ;
        RECT 94.000 27.600 96.600 28.400 ;
        RECT 98.800 28.200 99.600 28.400 ;
        RECT 98.000 27.600 99.600 28.200 ;
        RECT 100.400 27.600 103.000 28.400 ;
        RECT 105.200 28.200 106.000 28.400 ;
        RECT 104.400 27.600 106.000 28.200 ;
        RECT 106.800 27.600 109.400 28.400 ;
        RECT 111.600 28.200 112.400 28.400 ;
        RECT 110.800 27.600 112.400 28.200 ;
        RECT 118.800 27.800 129.800 28.400 ;
        RECT 118.800 27.600 120.400 27.800 ;
        RECT 40.400 27.200 41.200 27.600 ;
        RECT 39.800 26.200 43.400 26.600 ;
        RECT 44.400 26.200 45.000 27.600 ;
        RECT 46.200 26.200 46.800 27.600 ;
        RECT 50.000 27.200 50.800 27.600 ;
        RECT 53.200 27.200 54.000 27.600 ;
        RECT 47.800 26.200 51.400 26.600 ;
        RECT 52.600 26.200 56.200 26.600 ;
        RECT 57.200 26.200 57.800 27.600 ;
        RECT 59.600 27.200 60.400 27.600 ;
        RECT 59.000 26.200 62.600 26.600 ;
        RECT 63.600 26.200 64.200 27.600 ;
        RECT 65.200 26.800 67.600 27.600 ;
        RECT 68.600 26.800 70.800 27.600 ;
        RECT 71.800 26.800 74.000 27.600 ;
        RECT 75.400 26.800 77.200 27.600 ;
        RECT 39.600 26.000 43.600 26.200 ;
        RECT 39.600 22.200 40.400 26.000 ;
        RECT 42.800 22.200 43.600 26.000 ;
        RECT 44.400 22.200 45.200 26.200 ;
        RECT 46.000 22.200 46.800 26.200 ;
        RECT 47.600 26.000 51.600 26.200 ;
        RECT 47.600 22.200 48.400 26.000 ;
        RECT 50.800 22.200 51.600 26.000 ;
        RECT 52.400 26.000 56.400 26.200 ;
        RECT 52.400 22.200 53.200 26.000 ;
        RECT 55.600 22.200 56.400 26.000 ;
        RECT 57.200 22.200 58.000 26.200 ;
        RECT 58.800 26.000 62.800 26.200 ;
        RECT 58.800 22.200 59.600 26.000 ;
        RECT 62.000 22.200 62.800 26.000 ;
        RECT 63.600 22.200 64.400 26.200 ;
        RECT 66.800 22.200 67.600 26.800 ;
        RECT 70.000 22.200 70.800 26.800 ;
        RECT 73.200 22.200 74.000 26.800 ;
        RECT 76.400 22.200 77.200 26.800 ;
        RECT 81.200 26.800 83.000 27.600 ;
        RECT 84.400 26.800 86.600 27.600 ;
        RECT 87.600 26.800 89.800 27.600 ;
        RECT 90.800 26.800 93.200 27.600 ;
        RECT 81.200 22.200 82.000 26.800 ;
        RECT 84.400 22.200 85.200 26.800 ;
        RECT 87.600 22.200 88.400 26.800 ;
        RECT 90.800 22.200 91.600 26.800 ;
        RECT 94.200 26.200 94.800 27.600 ;
        RECT 98.000 27.200 98.800 27.600 ;
        RECT 95.800 26.200 99.400 26.600 ;
        RECT 100.600 26.200 101.200 27.600 ;
        RECT 104.400 27.200 105.200 27.600 ;
        RECT 102.200 26.200 105.800 26.600 ;
        RECT 107.000 26.200 107.600 27.600 ;
        RECT 110.800 27.200 111.600 27.600 ;
        RECT 108.600 26.200 112.200 26.600 ;
        RECT 94.000 22.200 94.800 26.200 ;
        RECT 95.600 26.000 99.600 26.200 ;
        RECT 95.600 22.200 96.400 26.000 ;
        RECT 98.800 22.200 99.600 26.000 ;
        RECT 100.400 22.200 101.200 26.200 ;
        RECT 102.000 26.000 106.000 26.200 ;
        RECT 102.000 22.200 102.800 26.000 ;
        RECT 105.200 22.200 106.000 26.000 ;
        RECT 106.800 22.200 107.600 26.200 ;
        RECT 108.400 26.000 112.400 26.200 ;
        RECT 108.400 22.200 109.200 26.000 ;
        RECT 111.600 22.200 112.400 26.000 ;
        RECT 118.000 22.200 118.800 27.000 ;
        RECT 123.000 25.600 123.600 27.800 ;
        RECT 124.400 27.600 125.200 27.800 ;
        RECT 128.600 27.600 129.400 27.800 ;
        RECT 135.600 27.200 136.400 30.600 ;
        RECT 137.200 30.300 138.000 30.400 ;
        RECT 138.800 30.300 139.600 30.400 ;
        RECT 137.200 29.700 139.600 30.300 ;
        RECT 137.200 29.600 138.000 29.700 ;
        RECT 138.800 28.800 139.600 29.700 ;
        RECT 140.200 30.300 140.800 31.800 ;
        RECT 142.000 31.600 142.800 31.800 ;
        RECT 143.600 31.600 144.400 33.200 ;
        RECT 143.600 30.300 144.400 30.400 ;
        RECT 140.200 29.700 144.400 30.300 ;
        RECT 140.200 28.400 140.800 29.700 ;
        RECT 143.600 29.600 144.400 29.700 ;
        RECT 137.200 28.200 138.000 28.400 ;
        RECT 137.200 27.600 138.800 28.200 ;
        RECT 140.200 27.600 142.800 28.400 ;
        RECT 138.000 27.200 138.800 27.600 ;
        RECT 132.600 26.600 136.400 27.200 ;
        RECT 132.600 26.400 133.400 26.600 ;
        RECT 121.200 24.200 122.000 25.000 ;
        RECT 122.800 24.800 123.600 25.600 ;
        RECT 124.600 25.400 125.400 25.600 ;
        RECT 124.600 24.800 127.400 25.400 ;
        RECT 126.800 24.200 127.400 24.800 ;
        RECT 130.800 24.200 131.600 25.000 ;
        RECT 121.200 23.600 123.200 24.200 ;
        RECT 122.400 22.200 123.200 23.600 ;
        RECT 126.800 22.200 127.600 24.200 ;
        RECT 130.800 23.600 132.200 24.200 ;
        RECT 131.000 22.200 132.200 23.600 ;
        RECT 135.600 22.200 136.400 26.600 ;
        RECT 137.400 26.200 141.000 26.600 ;
        RECT 142.000 26.200 142.600 27.600 ;
        RECT 145.200 26.200 146.000 39.800 ;
        RECT 149.200 33.600 150.000 34.400 ;
        RECT 149.200 32.400 149.800 33.600 ;
        RECT 150.600 32.400 151.400 39.800 ;
        RECT 148.400 31.800 149.800 32.400 ;
        RECT 150.400 31.800 151.400 32.400 ;
        RECT 148.400 31.600 149.200 31.800 ;
        RECT 150.400 30.400 151.000 31.800 ;
        RECT 154.800 31.400 155.600 39.800 ;
        RECT 159.200 36.400 160.000 39.800 ;
        RECT 158.000 35.800 160.000 36.400 ;
        RECT 163.600 35.800 164.400 39.800 ;
        RECT 167.800 35.800 169.000 39.800 ;
        RECT 158.000 35.000 158.800 35.800 ;
        RECT 163.600 35.200 164.200 35.800 ;
        RECT 161.400 34.600 165.000 35.200 ;
        RECT 167.600 35.000 168.400 35.800 ;
        RECT 161.400 34.400 162.200 34.600 ;
        RECT 164.200 34.400 165.000 34.600 ;
        RECT 158.000 33.000 158.800 33.200 ;
        RECT 162.600 33.000 163.400 33.200 ;
        RECT 158.000 32.400 163.400 33.000 ;
        RECT 164.000 33.000 166.200 33.600 ;
        RECT 164.000 31.800 164.600 33.000 ;
        RECT 165.400 32.800 166.200 33.000 ;
        RECT 167.800 33.200 169.200 34.000 ;
        RECT 167.800 32.200 168.400 33.200 ;
        RECT 159.800 31.400 164.600 31.800 ;
        RECT 154.800 31.200 164.600 31.400 ;
        RECT 166.000 31.600 168.400 32.200 ;
        RECT 154.800 31.000 160.600 31.200 ;
        RECT 154.800 30.800 160.400 31.000 ;
        RECT 166.000 30.400 166.600 31.600 ;
        RECT 172.400 31.200 173.200 39.800 ;
        RECT 176.600 38.400 177.400 39.800 ;
        RECT 175.600 37.600 177.400 38.400 ;
        RECT 176.600 32.600 177.400 37.600 ;
        RECT 175.600 31.800 177.400 32.600 ;
        RECT 169.000 30.600 173.200 31.200 ;
        RECT 169.000 30.400 169.800 30.600 ;
        RECT 150.000 29.600 151.000 30.400 ;
        RECT 150.400 28.400 151.000 29.600 ;
        RECT 151.600 30.300 152.400 30.400 ;
        RECT 153.200 30.300 154.000 30.400 ;
        RECT 151.600 29.700 154.000 30.300 ;
        RECT 161.200 30.200 162.000 30.400 ;
        RECT 151.600 28.800 152.400 29.700 ;
        RECT 153.200 29.600 154.000 29.700 ;
        RECT 157.000 29.600 162.000 30.200 ;
        RECT 166.000 29.600 166.800 30.400 ;
        RECT 170.600 29.800 171.400 30.000 ;
        RECT 157.000 29.400 157.800 29.600 ;
        RECT 159.600 29.400 160.400 29.600 ;
        RECT 158.600 28.400 159.400 28.600 ;
        RECT 166.000 28.400 166.600 29.600 ;
        RECT 167.600 29.200 171.400 29.800 ;
        RECT 167.600 29.000 168.400 29.200 ;
        RECT 146.800 26.800 147.600 28.400 ;
        RECT 148.400 27.600 151.000 28.400 ;
        RECT 153.200 28.200 154.000 28.400 ;
        RECT 152.400 27.600 154.000 28.200 ;
        RECT 155.600 27.800 166.600 28.400 ;
        RECT 155.600 27.600 157.200 27.800 ;
        RECT 148.600 26.200 149.200 27.600 ;
        RECT 152.400 27.200 153.200 27.600 ;
        RECT 150.200 26.200 153.800 26.600 ;
        RECT 137.200 26.000 141.200 26.200 ;
        RECT 137.200 22.200 138.000 26.000 ;
        RECT 140.400 22.200 141.200 26.000 ;
        RECT 142.000 22.200 142.800 26.200 ;
        RECT 144.200 25.600 146.000 26.200 ;
        RECT 144.200 22.200 145.000 25.600 ;
        RECT 148.400 22.200 149.200 26.200 ;
        RECT 150.000 26.000 154.000 26.200 ;
        RECT 150.000 22.200 150.800 26.000 ;
        RECT 153.200 22.200 154.000 26.000 ;
        RECT 154.800 22.200 155.600 27.000 ;
        RECT 159.800 25.600 160.400 27.800 ;
        RECT 165.400 27.600 166.200 27.800 ;
        RECT 172.400 27.200 173.200 30.600 ;
        RECT 175.800 28.400 176.400 31.800 ;
        RECT 177.200 30.300 178.000 31.200 ;
        RECT 178.800 30.300 179.600 39.800 ;
        RECT 184.600 38.400 185.400 39.800 ;
        RECT 183.600 37.600 185.400 38.400 ;
        RECT 184.600 32.600 185.400 37.600 ;
        RECT 183.600 31.800 185.400 32.600 ;
        RECT 186.800 32.400 187.600 39.800 ;
        RECT 188.200 32.400 189.000 32.600 ;
        RECT 186.800 31.800 189.000 32.400 ;
        RECT 191.200 32.400 192.800 39.800 ;
        RECT 194.800 32.400 195.600 32.600 ;
        RECT 196.400 32.400 197.200 39.800 ;
        RECT 191.200 31.800 193.200 32.400 ;
        RECT 194.800 31.800 197.200 32.400 ;
        RECT 199.600 32.000 200.400 39.800 ;
        RECT 202.800 35.200 203.600 39.800 ;
        RECT 177.200 29.700 179.600 30.300 ;
        RECT 177.200 29.600 178.000 29.700 ;
        RECT 175.600 27.600 176.400 28.400 ;
        RECT 169.400 26.600 173.200 27.200 ;
        RECT 169.400 26.400 170.200 26.600 ;
        RECT 158.000 24.200 158.800 25.000 ;
        RECT 159.600 24.800 160.400 25.600 ;
        RECT 161.400 25.400 162.200 25.600 ;
        RECT 161.400 24.800 164.200 25.400 ;
        RECT 163.600 24.200 164.200 24.800 ;
        RECT 167.600 24.200 168.400 25.000 ;
        RECT 158.000 23.600 160.000 24.200 ;
        RECT 159.200 22.200 160.000 23.600 ;
        RECT 163.600 22.200 164.400 24.200 ;
        RECT 167.600 23.600 169.000 24.200 ;
        RECT 167.800 22.200 169.000 23.600 ;
        RECT 172.400 22.200 173.200 26.600 ;
        RECT 174.000 24.800 174.800 26.400 ;
        RECT 175.800 24.200 176.400 27.600 ;
        RECT 175.600 22.200 176.400 24.200 ;
        RECT 178.800 22.200 179.600 29.700 ;
        RECT 183.800 28.400 184.400 31.800 ;
        RECT 188.400 31.200 189.000 31.800 ;
        RECT 185.200 29.600 186.000 31.200 ;
        RECT 188.400 30.600 191.800 31.200 ;
        RECT 191.000 30.400 191.800 30.600 ;
        RECT 192.600 30.400 193.200 31.800 ;
        RECT 199.400 31.200 200.400 32.000 ;
        RECT 201.000 34.600 203.600 35.200 ;
        RECT 201.000 33.000 201.600 34.600 ;
        RECT 206.000 34.400 206.800 39.800 ;
        RECT 209.200 37.000 210.000 39.800 ;
        RECT 210.800 37.000 211.600 39.800 ;
        RECT 212.400 37.000 213.200 39.800 ;
        RECT 207.400 34.400 211.600 35.200 ;
        RECT 204.200 33.600 206.800 34.400 ;
        RECT 214.000 33.600 214.800 39.800 ;
        RECT 217.200 35.000 218.000 39.800 ;
        RECT 220.400 35.000 221.200 39.800 ;
        RECT 222.000 37.000 222.800 39.800 ;
        RECT 223.600 37.000 224.400 39.800 ;
        RECT 226.800 35.200 227.600 39.800 ;
        RECT 230.000 36.400 230.800 39.800 ;
        RECT 234.800 36.400 235.600 39.800 ;
        RECT 230.000 35.800 231.000 36.400 ;
        RECT 230.400 35.200 231.000 35.800 ;
        RECT 234.600 35.800 235.600 36.400 ;
        RECT 234.600 35.200 235.200 35.800 ;
        RECT 238.000 35.200 238.800 39.800 ;
        RECT 241.200 37.000 242.000 39.800 ;
        RECT 242.800 37.000 243.600 39.800 ;
        RECT 225.600 34.400 229.800 35.200 ;
        RECT 230.400 34.600 232.400 35.200 ;
        RECT 217.200 33.600 219.800 34.400 ;
        RECT 220.400 33.800 226.200 34.400 ;
        RECT 229.200 34.000 229.800 34.400 ;
        RECT 209.200 33.000 210.000 33.200 ;
        RECT 201.000 32.400 210.000 33.000 ;
        RECT 212.400 33.000 213.200 33.200 ;
        RECT 220.400 33.000 221.000 33.800 ;
        RECT 226.800 33.200 228.200 33.800 ;
        RECT 229.200 33.200 230.800 34.000 ;
        RECT 212.400 32.400 221.000 33.000 ;
        RECT 222.000 33.000 228.200 33.200 ;
        RECT 222.000 32.600 227.400 33.000 ;
        RECT 222.000 32.400 222.800 32.600 ;
        RECT 192.600 30.300 194.000 30.400 ;
        RECT 198.000 30.300 198.800 30.400 ;
        RECT 188.800 29.800 189.600 30.000 ;
        RECT 192.600 29.800 198.800 30.300 ;
        RECT 188.800 29.200 191.400 29.800 ;
        RECT 190.800 28.600 191.400 29.200 ;
        RECT 192.200 29.700 198.800 29.800 ;
        RECT 192.200 29.600 194.000 29.700 ;
        RECT 198.000 29.600 198.800 29.700 ;
        RECT 192.200 29.200 193.200 29.600 ;
        RECT 183.600 27.600 184.400 28.400 ;
        RECT 186.800 28.200 188.400 28.400 ;
        RECT 186.800 27.600 190.200 28.200 ;
        RECT 190.800 27.800 191.600 28.600 ;
        RECT 180.400 24.800 181.200 26.400 ;
        RECT 182.000 24.800 182.800 26.400 ;
        RECT 183.800 24.200 184.400 27.600 ;
        RECT 189.600 27.200 190.200 27.600 ;
        RECT 188.200 26.800 189.000 27.000 ;
        RECT 183.600 22.200 184.400 24.200 ;
        RECT 186.800 26.200 189.000 26.800 ;
        RECT 189.600 26.600 191.600 27.200 ;
        RECT 190.000 26.400 191.600 26.600 ;
        RECT 186.800 22.200 187.600 26.200 ;
        RECT 192.200 25.800 192.800 29.200 ;
        RECT 193.600 27.600 194.400 28.400 ;
        RECT 195.600 28.300 197.200 28.400 ;
        RECT 199.400 28.300 200.200 31.200 ;
        RECT 201.000 30.600 201.600 32.400 ;
        RECT 195.600 27.700 200.200 28.300 ;
        RECT 195.600 27.600 197.200 27.700 ;
        RECT 193.600 27.200 194.200 27.600 ;
        RECT 193.400 26.400 194.200 27.200 ;
        RECT 194.800 26.800 195.600 27.000 ;
        RECT 199.400 26.800 200.200 27.700 ;
        RECT 200.800 30.000 201.600 30.600 ;
        RECT 207.600 30.000 231.000 30.600 ;
        RECT 200.800 28.000 201.400 30.000 ;
        RECT 207.600 29.400 208.400 30.000 ;
        RECT 218.800 29.600 219.600 30.000 ;
        RECT 225.200 29.600 226.000 30.000 ;
        RECT 230.200 29.800 231.000 30.000 ;
        RECT 202.000 28.600 205.800 29.400 ;
        RECT 200.800 27.400 202.000 28.000 ;
        RECT 194.800 26.200 197.200 26.800 ;
        RECT 191.200 22.200 192.800 25.800 ;
        RECT 196.400 22.200 197.200 26.200 ;
        RECT 199.400 26.000 200.400 26.800 ;
        RECT 199.600 22.200 200.400 26.000 ;
        RECT 201.200 22.200 202.000 27.400 ;
        RECT 205.000 27.400 205.800 28.600 ;
        RECT 205.000 26.800 206.800 27.400 ;
        RECT 206.000 26.200 206.800 26.800 ;
        RECT 210.800 26.400 211.600 29.200 ;
        RECT 214.000 28.600 217.200 29.400 ;
        RECT 221.000 28.600 223.000 29.400 ;
        RECT 231.600 29.000 232.400 34.600 ;
        RECT 213.600 27.800 214.400 28.000 ;
        RECT 213.600 27.200 218.000 27.800 ;
        RECT 217.200 27.000 218.000 27.200 ;
        RECT 218.800 26.800 219.600 28.400 ;
        RECT 206.000 25.400 208.400 26.200 ;
        RECT 210.800 25.600 211.800 26.400 ;
        RECT 214.800 25.600 216.400 26.400 ;
        RECT 217.200 26.200 218.000 26.400 ;
        RECT 221.000 26.200 221.800 28.600 ;
        RECT 223.600 28.200 232.400 29.000 ;
        RECT 227.000 26.800 230.000 27.600 ;
        RECT 227.000 26.200 227.800 26.800 ;
        RECT 217.200 25.600 221.800 26.200 ;
        RECT 207.600 22.200 208.400 25.400 ;
        RECT 225.200 25.400 227.800 26.200 ;
        RECT 209.200 22.200 210.000 25.000 ;
        RECT 210.800 22.200 211.600 25.000 ;
        RECT 212.400 22.200 213.200 25.000 ;
        RECT 214.000 22.200 214.800 25.000 ;
        RECT 217.200 22.200 218.000 25.000 ;
        RECT 220.400 22.200 221.200 25.000 ;
        RECT 222.000 22.200 222.800 25.000 ;
        RECT 223.600 22.200 224.400 25.000 ;
        RECT 225.200 22.200 226.000 25.400 ;
        RECT 231.600 22.200 232.400 28.200 ;
        RECT 233.200 34.600 235.200 35.200 ;
        RECT 233.200 29.000 234.000 34.600 ;
        RECT 235.800 34.400 240.000 35.200 ;
        RECT 244.400 35.000 245.200 39.800 ;
        RECT 247.600 35.000 248.400 39.800 ;
        RECT 235.800 34.000 236.400 34.400 ;
        RECT 234.800 33.200 236.400 34.000 ;
        RECT 239.400 33.800 245.200 34.400 ;
        RECT 237.400 33.200 238.800 33.800 ;
        RECT 237.400 33.000 243.600 33.200 ;
        RECT 238.200 32.600 243.600 33.000 ;
        RECT 242.800 32.400 243.600 32.600 ;
        RECT 244.600 33.000 245.200 33.800 ;
        RECT 245.800 33.600 248.400 34.400 ;
        RECT 250.800 33.600 251.600 39.800 ;
        RECT 252.400 37.000 253.200 39.800 ;
        RECT 254.000 37.000 254.800 39.800 ;
        RECT 255.600 37.000 256.400 39.800 ;
        RECT 254.000 34.400 258.200 35.200 ;
        RECT 258.800 34.400 259.600 39.800 ;
        RECT 262.000 35.200 262.800 39.800 ;
        RECT 262.000 34.600 264.600 35.200 ;
        RECT 258.800 33.600 261.400 34.400 ;
        RECT 252.400 33.000 253.200 33.200 ;
        RECT 244.600 32.400 253.200 33.000 ;
        RECT 255.600 33.000 256.400 33.200 ;
        RECT 264.000 33.000 264.600 34.600 ;
        RECT 255.600 32.400 264.600 33.000 ;
        RECT 264.000 30.600 264.600 32.400 ;
        RECT 265.200 32.000 266.000 39.800 ;
        RECT 275.800 32.400 276.600 39.800 ;
        RECT 277.200 33.600 278.000 34.400 ;
        RECT 277.400 32.400 278.000 33.600 ;
        RECT 265.200 31.200 266.200 32.000 ;
        RECT 275.800 31.800 276.800 32.400 ;
        RECT 277.400 31.800 278.800 32.400 ;
        RECT 234.600 30.000 258.000 30.600 ;
        RECT 264.000 30.000 264.800 30.600 ;
        RECT 234.600 29.800 235.600 30.000 ;
        RECT 234.800 29.600 235.600 29.800 ;
        RECT 239.600 29.600 240.400 30.000 ;
        RECT 257.200 29.400 258.000 30.000 ;
        RECT 233.200 28.200 242.000 29.000 ;
        RECT 242.600 28.600 244.600 29.400 ;
        RECT 248.400 28.600 251.600 29.400 ;
        RECT 233.200 22.200 234.000 28.200 ;
        RECT 235.600 26.800 238.600 27.600 ;
        RECT 237.800 26.200 238.600 26.800 ;
        RECT 243.800 26.200 244.600 28.600 ;
        RECT 246.000 26.800 246.800 28.400 ;
        RECT 251.200 27.800 252.000 28.000 ;
        RECT 247.600 27.200 252.000 27.800 ;
        RECT 247.600 27.000 248.400 27.200 ;
        RECT 254.000 26.400 254.800 29.200 ;
        RECT 259.800 28.600 263.600 29.400 ;
        RECT 259.800 27.400 260.600 28.600 ;
        RECT 264.200 28.000 264.800 30.000 ;
        RECT 247.600 26.200 248.400 26.400 ;
        RECT 237.800 25.400 240.400 26.200 ;
        RECT 243.800 25.600 248.400 26.200 ;
        RECT 249.200 25.600 250.800 26.400 ;
        RECT 253.800 25.600 254.800 26.400 ;
        RECT 258.800 26.800 260.600 27.400 ;
        RECT 263.600 27.400 264.800 28.000 ;
        RECT 258.800 26.200 259.600 26.800 ;
        RECT 239.600 22.200 240.400 25.400 ;
        RECT 257.200 25.400 259.600 26.200 ;
        RECT 241.200 22.200 242.000 25.000 ;
        RECT 242.800 22.200 243.600 25.000 ;
        RECT 244.400 22.200 245.200 25.000 ;
        RECT 247.600 22.200 248.400 25.000 ;
        RECT 250.800 22.200 251.600 25.000 ;
        RECT 252.400 22.200 253.200 25.000 ;
        RECT 254.000 22.200 254.800 25.000 ;
        RECT 255.600 22.200 256.400 25.000 ;
        RECT 257.200 22.200 258.000 25.400 ;
        RECT 263.600 22.200 264.400 27.400 ;
        RECT 265.400 26.800 266.200 31.200 ;
        RECT 276.200 30.400 276.800 31.800 ;
        RECT 278.000 31.600 278.800 31.800 ;
        RECT 279.600 31.600 280.400 33.200 ;
        RECT 271.600 30.300 272.400 30.400 ;
        RECT 274.800 30.300 275.600 30.400 ;
        RECT 271.600 29.700 275.600 30.300 ;
        RECT 271.600 29.600 272.400 29.700 ;
        RECT 274.800 28.800 275.600 29.700 ;
        RECT 276.200 29.600 277.200 30.400 ;
        RECT 278.100 30.300 278.700 31.600 ;
        RECT 281.200 30.300 282.000 39.800 ;
        RECT 278.100 29.700 282.000 30.300 ;
        RECT 276.200 28.400 276.800 29.600 ;
        RECT 273.200 28.200 274.000 28.400 ;
        RECT 273.200 27.600 274.800 28.200 ;
        RECT 276.200 27.600 278.800 28.400 ;
        RECT 274.000 27.200 274.800 27.600 ;
        RECT 265.200 26.000 266.200 26.800 ;
        RECT 273.400 26.200 277.000 26.600 ;
        RECT 278.000 26.200 278.600 27.600 ;
        RECT 281.200 26.200 282.000 29.700 ;
        RECT 282.800 28.300 283.600 28.400 ;
        RECT 284.400 28.300 285.200 28.400 ;
        RECT 282.800 27.700 285.200 28.300 ;
        RECT 282.800 26.800 283.600 27.700 ;
        RECT 284.400 26.800 285.200 27.700 ;
        RECT 273.200 26.000 277.200 26.200 ;
        RECT 265.200 22.200 266.000 26.000 ;
        RECT 273.200 22.200 274.000 26.000 ;
        RECT 276.400 22.200 277.200 26.000 ;
        RECT 278.000 22.200 278.800 26.200 ;
        RECT 280.200 25.600 282.000 26.200 ;
        RECT 286.000 26.200 286.800 39.800 ;
        RECT 287.600 31.600 288.400 33.200 ;
        RECT 290.800 31.200 291.600 39.800 ;
        RECT 294.000 31.200 294.800 39.800 ;
        RECT 297.200 31.200 298.000 39.800 ;
        RECT 300.400 31.200 301.200 39.800 ;
        RECT 306.200 32.400 307.000 39.800 ;
        RECT 307.600 33.600 308.400 34.400 ;
        RECT 307.800 32.400 308.400 33.600 ;
        RECT 306.200 31.800 307.200 32.400 ;
        RECT 307.800 31.800 309.200 32.400 ;
        RECT 289.200 30.400 291.600 31.200 ;
        RECT 292.600 30.400 294.800 31.200 ;
        RECT 295.800 30.400 298.000 31.200 ;
        RECT 299.400 30.400 301.200 31.200 ;
        RECT 289.200 27.600 290.000 30.400 ;
        RECT 292.600 29.000 293.400 30.400 ;
        RECT 295.800 29.000 296.600 30.400 ;
        RECT 299.400 29.000 300.200 30.400 ;
        RECT 290.800 28.200 293.400 29.000 ;
        RECT 294.200 28.200 296.600 29.000 ;
        RECT 297.600 28.200 300.200 29.000 ;
        RECT 301.000 28.200 302.800 29.000 ;
        RECT 305.200 28.800 306.000 30.400 ;
        RECT 306.600 28.400 307.200 31.800 ;
        RECT 308.400 31.600 309.200 31.800 ;
        RECT 308.400 30.300 309.200 30.400 ;
        RECT 310.000 30.300 310.800 39.800 ;
        RECT 314.800 32.000 315.600 39.800 ;
        RECT 318.000 35.200 318.800 39.800 ;
        RECT 308.400 29.700 310.800 30.300 ;
        RECT 308.400 29.600 309.200 29.700 ;
        RECT 292.600 27.600 293.400 28.200 ;
        RECT 295.800 27.600 296.600 28.200 ;
        RECT 299.400 27.600 300.200 28.200 ;
        RECT 302.000 27.600 302.800 28.200 ;
        RECT 303.600 28.200 304.400 28.400 ;
        RECT 303.600 27.600 305.200 28.200 ;
        RECT 306.600 27.600 309.200 28.400 ;
        RECT 289.200 26.800 291.600 27.600 ;
        RECT 292.600 26.800 294.800 27.600 ;
        RECT 295.800 26.800 298.000 27.600 ;
        RECT 299.400 26.800 301.200 27.600 ;
        RECT 304.400 27.200 305.200 27.600 ;
        RECT 286.000 25.600 287.800 26.200 ;
        RECT 280.200 22.200 281.000 25.600 ;
        RECT 287.000 24.400 287.800 25.600 ;
        RECT 286.000 23.600 287.800 24.400 ;
        RECT 287.000 22.200 287.800 23.600 ;
        RECT 290.800 22.200 291.600 26.800 ;
        RECT 294.000 22.200 294.800 26.800 ;
        RECT 297.200 22.200 298.000 26.800 ;
        RECT 300.400 22.200 301.200 26.800 ;
        RECT 303.800 26.200 307.400 26.600 ;
        RECT 308.400 26.400 309.000 27.600 ;
        RECT 303.600 26.000 307.600 26.200 ;
        RECT 303.600 22.200 304.400 26.000 ;
        RECT 306.800 22.200 307.600 26.000 ;
        RECT 308.400 22.200 309.200 26.400 ;
        RECT 310.000 22.200 310.800 29.700 ;
        RECT 314.600 31.200 315.600 32.000 ;
        RECT 316.200 34.600 318.800 35.200 ;
        RECT 316.200 33.000 316.800 34.600 ;
        RECT 321.200 34.400 322.000 39.800 ;
        RECT 324.400 37.000 325.200 39.800 ;
        RECT 326.000 37.000 326.800 39.800 ;
        RECT 327.600 37.000 328.400 39.800 ;
        RECT 322.600 34.400 326.800 35.200 ;
        RECT 319.400 33.600 322.000 34.400 ;
        RECT 329.200 33.600 330.000 39.800 ;
        RECT 332.400 35.000 333.200 39.800 ;
        RECT 335.600 35.000 336.400 39.800 ;
        RECT 337.200 37.000 338.000 39.800 ;
        RECT 338.800 37.000 339.600 39.800 ;
        RECT 342.000 35.200 342.800 39.800 ;
        RECT 345.200 36.400 346.000 39.800 ;
        RECT 345.200 35.800 346.200 36.400 ;
        RECT 345.600 35.200 346.200 35.800 ;
        RECT 340.800 34.400 345.000 35.200 ;
        RECT 345.600 34.600 347.600 35.200 ;
        RECT 332.400 33.600 335.000 34.400 ;
        RECT 335.600 33.800 341.400 34.400 ;
        RECT 344.400 34.000 345.000 34.400 ;
        RECT 324.400 33.000 325.200 33.200 ;
        RECT 316.200 32.400 325.200 33.000 ;
        RECT 327.600 33.000 328.400 33.200 ;
        RECT 335.600 33.000 336.200 33.800 ;
        RECT 342.000 33.200 343.400 33.800 ;
        RECT 344.400 33.200 346.000 34.000 ;
        RECT 327.600 32.400 336.200 33.000 ;
        RECT 337.200 33.000 343.400 33.200 ;
        RECT 337.200 32.600 342.600 33.000 ;
        RECT 337.200 32.400 338.000 32.600 ;
        RECT 314.600 26.800 315.400 31.200 ;
        RECT 316.200 30.600 316.800 32.400 ;
        RECT 316.000 30.000 316.800 30.600 ;
        RECT 322.800 30.000 346.200 30.600 ;
        RECT 316.000 28.000 316.600 30.000 ;
        RECT 322.800 29.400 323.600 30.000 ;
        RECT 340.400 29.600 341.200 30.000 ;
        RECT 343.600 29.600 344.400 30.000 ;
        RECT 345.400 29.800 346.200 30.000 ;
        RECT 317.200 28.600 321.000 29.400 ;
        RECT 316.000 27.400 317.200 28.000 ;
        RECT 311.600 26.300 312.400 26.400 ;
        RECT 314.600 26.300 315.600 26.800 ;
        RECT 311.600 25.700 315.600 26.300 ;
        RECT 311.600 24.800 312.400 25.700 ;
        RECT 314.800 22.200 315.600 25.700 ;
        RECT 316.400 22.200 317.200 27.400 ;
        RECT 320.200 27.400 321.000 28.600 ;
        RECT 320.200 26.800 322.000 27.400 ;
        RECT 321.200 26.200 322.000 26.800 ;
        RECT 326.000 26.400 326.800 29.200 ;
        RECT 329.200 28.600 332.400 29.400 ;
        RECT 336.200 28.600 338.200 29.400 ;
        RECT 346.800 29.000 347.600 34.600 ;
        RECT 350.000 31.200 350.800 39.800 ;
        RECT 353.200 31.200 354.000 39.800 ;
        RECT 356.400 31.200 357.200 39.800 ;
        RECT 359.600 31.200 360.400 39.800 ;
        RECT 350.000 30.400 351.800 31.200 ;
        RECT 353.200 30.400 355.400 31.200 ;
        RECT 356.400 30.400 358.600 31.200 ;
        RECT 359.600 30.400 362.000 31.200 ;
        RECT 351.000 29.000 351.800 30.400 ;
        RECT 354.600 29.000 355.400 30.400 ;
        RECT 357.800 29.000 358.600 30.400 ;
        RECT 328.800 27.800 329.600 28.000 ;
        RECT 328.800 27.200 333.200 27.800 ;
        RECT 332.400 27.000 333.200 27.200 ;
        RECT 334.000 26.800 334.800 28.400 ;
        RECT 321.200 25.400 323.600 26.200 ;
        RECT 326.000 25.600 327.000 26.400 ;
        RECT 330.000 25.600 331.600 26.400 ;
        RECT 332.400 26.200 333.200 26.400 ;
        RECT 336.200 26.200 337.000 28.600 ;
        RECT 338.800 28.200 347.600 29.000 ;
        RECT 342.200 26.800 345.200 27.600 ;
        RECT 342.200 26.200 343.000 26.800 ;
        RECT 332.400 25.600 337.000 26.200 ;
        RECT 322.800 22.200 323.600 25.400 ;
        RECT 340.400 25.400 343.000 26.200 ;
        RECT 324.400 22.200 325.200 25.000 ;
        RECT 326.000 22.200 326.800 25.000 ;
        RECT 327.600 22.200 328.400 25.000 ;
        RECT 329.200 22.200 330.000 25.000 ;
        RECT 332.400 22.200 333.200 25.000 ;
        RECT 335.600 22.200 336.400 25.000 ;
        RECT 337.200 22.200 338.000 25.000 ;
        RECT 338.800 22.200 339.600 25.000 ;
        RECT 340.400 22.200 341.200 25.400 ;
        RECT 346.800 22.200 347.600 28.200 ;
        RECT 348.400 28.200 350.200 29.000 ;
        RECT 351.000 28.200 353.600 29.000 ;
        RECT 354.600 28.200 357.000 29.000 ;
        RECT 357.800 28.200 360.400 29.000 ;
        RECT 348.400 27.600 349.200 28.200 ;
        RECT 351.000 27.600 351.800 28.200 ;
        RECT 354.600 27.600 355.400 28.200 ;
        RECT 357.800 27.600 358.600 28.200 ;
        RECT 361.200 27.600 362.000 30.400 ;
        RECT 350.000 26.800 351.800 27.600 ;
        RECT 353.200 26.800 355.400 27.600 ;
        RECT 356.400 26.800 358.600 27.600 ;
        RECT 359.600 26.800 362.000 27.600 ;
        RECT 364.400 30.300 365.200 39.800 ;
        RECT 368.600 32.400 369.400 39.800 ;
        RECT 374.000 36.400 374.800 39.800 ;
        RECT 373.800 35.800 374.800 36.400 ;
        RECT 373.800 35.200 374.400 35.800 ;
        RECT 377.200 35.200 378.000 39.800 ;
        RECT 380.400 37.000 381.200 39.800 ;
        RECT 382.000 37.000 382.800 39.800 ;
        RECT 372.400 34.600 374.400 35.200 ;
        RECT 370.000 33.600 370.800 34.400 ;
        RECT 370.200 32.400 370.800 33.600 ;
        RECT 368.600 31.800 369.600 32.400 ;
        RECT 370.200 31.800 371.600 32.400 ;
        RECT 367.600 30.300 368.400 30.400 ;
        RECT 364.400 29.700 368.400 30.300 ;
        RECT 350.000 22.200 350.800 26.800 ;
        RECT 353.200 22.200 354.000 26.800 ;
        RECT 356.400 22.200 357.200 26.800 ;
        RECT 359.600 22.200 360.400 26.800 ;
        RECT 362.800 24.800 363.600 26.400 ;
        RECT 364.400 22.200 365.200 29.700 ;
        RECT 367.600 28.800 368.400 29.700 ;
        RECT 369.000 28.400 369.600 31.800 ;
        RECT 370.800 31.600 371.600 31.800 ;
        RECT 372.400 29.000 373.200 34.600 ;
        RECT 375.000 34.400 379.200 35.200 ;
        RECT 383.600 35.000 384.400 39.800 ;
        RECT 386.800 35.000 387.600 39.800 ;
        RECT 375.000 34.000 375.600 34.400 ;
        RECT 374.000 33.200 375.600 34.000 ;
        RECT 378.600 33.800 384.400 34.400 ;
        RECT 376.600 33.200 378.000 33.800 ;
        RECT 376.600 33.000 382.800 33.200 ;
        RECT 377.400 32.600 382.800 33.000 ;
        RECT 382.000 32.400 382.800 32.600 ;
        RECT 383.800 33.000 384.400 33.800 ;
        RECT 385.000 33.600 387.600 34.400 ;
        RECT 390.000 33.600 390.800 39.800 ;
        RECT 391.600 37.000 392.400 39.800 ;
        RECT 393.200 37.000 394.000 39.800 ;
        RECT 394.800 37.000 395.600 39.800 ;
        RECT 393.200 34.400 397.400 35.200 ;
        RECT 398.000 34.400 398.800 39.800 ;
        RECT 401.200 35.200 402.000 39.800 ;
        RECT 401.200 34.600 403.800 35.200 ;
        RECT 398.000 33.600 400.600 34.400 ;
        RECT 391.600 33.000 392.400 33.200 ;
        RECT 383.800 32.400 392.400 33.000 ;
        RECT 394.800 33.000 395.600 33.200 ;
        RECT 403.200 33.000 403.800 34.600 ;
        RECT 394.800 32.400 403.800 33.000 ;
        RECT 403.200 30.600 403.800 32.400 ;
        RECT 404.400 32.000 405.200 39.800 ;
        RECT 404.400 31.200 405.400 32.000 ;
        RECT 373.800 30.000 397.200 30.600 ;
        RECT 403.200 30.000 404.000 30.600 ;
        RECT 373.800 29.800 374.600 30.000 ;
        RECT 378.800 29.600 379.600 30.000 ;
        RECT 396.400 29.400 397.200 30.000 ;
        RECT 366.000 28.200 366.800 28.400 ;
        RECT 366.000 27.600 367.600 28.200 ;
        RECT 369.000 27.600 371.600 28.400 ;
        RECT 372.400 28.200 381.200 29.000 ;
        RECT 381.800 28.600 383.800 29.400 ;
        RECT 387.600 28.600 390.800 29.400 ;
        RECT 366.800 27.200 367.600 27.600 ;
        RECT 366.200 26.200 369.800 26.600 ;
        RECT 370.800 26.200 371.400 27.600 ;
        RECT 366.000 26.000 370.000 26.200 ;
        RECT 366.000 22.200 366.800 26.000 ;
        RECT 369.200 22.200 370.000 26.000 ;
        RECT 370.800 22.200 371.600 26.200 ;
        RECT 372.400 22.200 373.200 28.200 ;
        RECT 374.800 26.800 377.800 27.600 ;
        RECT 377.000 26.200 377.800 26.800 ;
        RECT 383.000 26.200 383.800 28.600 ;
        RECT 385.200 26.800 386.000 28.400 ;
        RECT 390.400 27.800 391.200 28.000 ;
        RECT 386.800 27.200 391.200 27.800 ;
        RECT 386.800 27.000 387.600 27.200 ;
        RECT 393.200 26.400 394.000 29.200 ;
        RECT 399.000 28.600 402.800 29.400 ;
        RECT 399.000 27.400 399.800 28.600 ;
        RECT 403.400 28.000 404.000 30.000 ;
        RECT 386.800 26.200 387.600 26.400 ;
        RECT 377.000 25.400 379.600 26.200 ;
        RECT 383.000 25.600 387.600 26.200 ;
        RECT 388.400 25.600 390.000 26.400 ;
        RECT 393.000 25.600 394.000 26.400 ;
        RECT 398.000 26.800 399.800 27.400 ;
        RECT 402.800 27.400 404.000 28.000 ;
        RECT 398.000 26.200 398.800 26.800 ;
        RECT 378.800 22.200 379.600 25.400 ;
        RECT 396.400 25.400 398.800 26.200 ;
        RECT 380.400 22.200 381.200 25.000 ;
        RECT 382.000 22.200 382.800 25.000 ;
        RECT 383.600 22.200 384.400 25.000 ;
        RECT 386.800 22.200 387.600 25.000 ;
        RECT 390.000 22.200 390.800 25.000 ;
        RECT 391.600 22.200 392.400 25.000 ;
        RECT 393.200 22.200 394.000 25.000 ;
        RECT 394.800 22.200 395.600 25.000 ;
        RECT 396.400 22.200 397.200 25.400 ;
        RECT 402.800 22.200 403.600 27.400 ;
        RECT 404.600 26.800 405.400 31.200 ;
        RECT 404.400 26.300 405.400 26.800 ;
        RECT 409.200 30.300 410.000 39.800 ;
        RECT 413.000 34.400 413.800 39.800 ;
        RECT 411.600 33.600 412.400 34.400 ;
        RECT 413.000 33.600 414.800 34.400 ;
        RECT 422.800 33.600 423.600 34.400 ;
        RECT 411.600 32.400 412.200 33.600 ;
        RECT 413.000 32.400 413.800 33.600 ;
        RECT 422.800 32.400 423.400 33.600 ;
        RECT 424.200 32.400 425.000 39.800 ;
        RECT 410.800 31.800 412.200 32.400 ;
        RECT 412.800 31.800 413.800 32.400 ;
        RECT 422.000 31.800 423.400 32.400 ;
        RECT 424.000 31.800 425.000 32.400 ;
        RECT 410.800 31.600 411.600 31.800 ;
        RECT 410.800 30.300 411.600 30.400 ;
        RECT 409.200 29.700 411.600 30.300 ;
        RECT 407.600 26.300 408.400 26.400 ;
        RECT 404.400 25.700 408.400 26.300 ;
        RECT 404.400 22.200 405.200 25.700 ;
        RECT 407.600 24.800 408.400 25.700 ;
        RECT 409.200 22.200 410.000 29.700 ;
        RECT 410.800 29.600 411.600 29.700 ;
        RECT 412.800 28.400 413.400 31.800 ;
        RECT 422.000 31.600 422.800 31.800 ;
        RECT 414.000 28.800 414.800 30.400 ;
        RECT 424.000 28.400 424.600 31.800 ;
        RECT 425.200 30.300 426.000 30.400 ;
        RECT 428.400 30.300 429.200 39.800 ;
        RECT 433.200 36.400 434.000 39.800 ;
        RECT 433.000 35.800 434.000 36.400 ;
        RECT 433.000 35.200 433.600 35.800 ;
        RECT 436.400 35.200 437.200 39.800 ;
        RECT 439.600 37.000 440.400 39.800 ;
        RECT 441.200 37.000 442.000 39.800 ;
        RECT 425.200 29.700 429.200 30.300 ;
        RECT 425.200 28.800 426.000 29.700 ;
        RECT 410.800 27.600 413.400 28.400 ;
        RECT 415.600 28.200 416.400 28.400 ;
        RECT 414.800 27.600 416.400 28.200 ;
        RECT 422.000 27.600 424.600 28.400 ;
        RECT 426.800 28.200 427.600 28.400 ;
        RECT 426.000 27.600 427.600 28.200 ;
        RECT 411.000 26.200 411.600 27.600 ;
        RECT 414.800 27.200 415.600 27.600 ;
        RECT 412.600 26.200 416.200 26.600 ;
        RECT 422.200 26.200 422.800 27.600 ;
        RECT 426.000 27.200 426.800 27.600 ;
        RECT 423.800 26.200 427.400 26.600 ;
        RECT 410.800 22.200 411.600 26.200 ;
        RECT 412.400 26.000 416.400 26.200 ;
        RECT 412.400 22.200 413.200 26.000 ;
        RECT 415.600 22.200 416.400 26.000 ;
        RECT 417.200 24.300 418.000 24.400 ;
        RECT 422.000 24.300 422.800 26.200 ;
        RECT 417.200 23.700 422.800 24.300 ;
        RECT 417.200 23.600 418.000 23.700 ;
        RECT 422.000 22.200 422.800 23.700 ;
        RECT 423.600 26.000 427.600 26.200 ;
        RECT 423.600 22.200 424.400 26.000 ;
        RECT 426.800 22.200 427.600 26.000 ;
        RECT 428.400 22.200 429.200 29.700 ;
        RECT 431.600 34.600 433.600 35.200 ;
        RECT 431.600 29.000 432.400 34.600 ;
        RECT 434.200 34.400 438.400 35.200 ;
        RECT 442.800 35.000 443.600 39.800 ;
        RECT 446.000 35.000 446.800 39.800 ;
        RECT 434.200 34.000 434.800 34.400 ;
        RECT 433.200 33.200 434.800 34.000 ;
        RECT 437.800 33.800 443.600 34.400 ;
        RECT 435.800 33.200 437.200 33.800 ;
        RECT 435.800 33.000 442.000 33.200 ;
        RECT 436.600 32.600 442.000 33.000 ;
        RECT 441.200 32.400 442.000 32.600 ;
        RECT 443.000 33.000 443.600 33.800 ;
        RECT 444.200 33.600 446.800 34.400 ;
        RECT 449.200 33.600 450.000 39.800 ;
        RECT 450.800 37.000 451.600 39.800 ;
        RECT 452.400 37.000 453.200 39.800 ;
        RECT 454.000 37.000 454.800 39.800 ;
        RECT 452.400 34.400 456.600 35.200 ;
        RECT 457.200 34.400 458.000 39.800 ;
        RECT 460.400 35.200 461.200 39.800 ;
        RECT 460.400 34.600 463.000 35.200 ;
        RECT 457.200 33.600 459.800 34.400 ;
        RECT 450.800 33.000 451.600 33.200 ;
        RECT 443.000 32.400 451.600 33.000 ;
        RECT 454.000 33.000 454.800 33.200 ;
        RECT 462.400 33.000 463.000 34.600 ;
        RECT 454.000 32.400 463.000 33.000 ;
        RECT 462.400 30.600 463.000 32.400 ;
        RECT 463.600 32.000 464.400 39.800 ;
        RECT 469.400 32.400 470.200 39.800 ;
        RECT 470.800 33.600 471.600 34.400 ;
        RECT 471.000 32.400 471.600 33.600 ;
        RECT 474.000 33.600 474.800 34.400 ;
        RECT 474.000 32.400 474.600 33.600 ;
        RECT 475.400 32.400 476.200 39.800 ;
        RECT 480.400 33.600 481.200 34.400 ;
        RECT 480.400 32.400 481.000 33.600 ;
        RECT 481.800 32.400 482.600 39.800 ;
        RECT 486.800 33.600 487.600 34.400 ;
        RECT 486.800 32.400 487.400 33.600 ;
        RECT 488.200 32.400 489.000 39.800 ;
        RECT 463.600 31.200 464.600 32.000 ;
        RECT 469.400 31.800 470.400 32.400 ;
        RECT 471.000 31.800 472.400 32.400 ;
        RECT 433.000 30.000 456.400 30.600 ;
        RECT 462.400 30.000 463.200 30.600 ;
        RECT 433.000 29.800 433.800 30.000 ;
        RECT 434.800 29.600 435.600 30.000 ;
        RECT 438.000 29.600 438.800 30.000 ;
        RECT 455.600 29.400 456.400 30.000 ;
        RECT 431.600 28.200 440.400 29.000 ;
        RECT 441.000 28.600 443.000 29.400 ;
        RECT 446.800 28.600 450.000 29.400 ;
        RECT 430.000 24.800 430.800 26.400 ;
        RECT 431.600 22.200 432.400 28.200 ;
        RECT 434.000 26.800 437.000 27.600 ;
        RECT 436.200 26.200 437.000 26.800 ;
        RECT 442.200 26.200 443.000 28.600 ;
        RECT 444.400 26.800 445.200 28.400 ;
        RECT 449.600 27.800 450.400 28.000 ;
        RECT 446.000 27.200 450.400 27.800 ;
        RECT 446.000 27.000 446.800 27.200 ;
        RECT 452.400 26.400 453.200 29.200 ;
        RECT 458.200 28.600 462.000 29.400 ;
        RECT 458.200 27.400 459.000 28.600 ;
        RECT 462.600 28.000 463.200 30.000 ;
        RECT 446.000 26.200 446.800 26.400 ;
        RECT 436.200 25.400 438.800 26.200 ;
        RECT 442.200 25.600 446.800 26.200 ;
        RECT 447.600 25.600 449.200 26.400 ;
        RECT 452.200 25.600 453.200 26.400 ;
        RECT 457.200 26.800 459.000 27.400 ;
        RECT 462.000 27.400 463.200 28.000 ;
        RECT 457.200 26.200 458.000 26.800 ;
        RECT 438.000 22.200 438.800 25.400 ;
        RECT 455.600 25.400 458.000 26.200 ;
        RECT 439.600 22.200 440.400 25.000 ;
        RECT 441.200 22.200 442.000 25.000 ;
        RECT 442.800 22.200 443.600 25.000 ;
        RECT 446.000 22.200 446.800 25.000 ;
        RECT 449.200 22.200 450.000 25.000 ;
        RECT 450.800 22.200 451.600 25.000 ;
        RECT 452.400 22.200 453.200 25.000 ;
        RECT 454.000 22.200 454.800 25.000 ;
        RECT 455.600 22.200 456.400 25.400 ;
        RECT 462.000 22.200 462.800 27.400 ;
        RECT 463.800 26.800 464.600 31.200 ;
        RECT 466.800 30.300 467.600 30.400 ;
        RECT 468.400 30.300 469.200 30.400 ;
        RECT 466.800 29.700 469.200 30.300 ;
        RECT 466.800 29.600 467.600 29.700 ;
        RECT 468.400 28.800 469.200 29.700 ;
        RECT 469.800 28.400 470.400 31.800 ;
        RECT 471.600 31.600 472.400 31.800 ;
        RECT 473.200 31.800 474.600 32.400 ;
        RECT 475.200 31.800 476.200 32.400 ;
        RECT 479.600 31.800 481.000 32.400 ;
        RECT 473.200 31.600 474.000 31.800 ;
        RECT 471.700 30.300 472.300 31.600 ;
        RECT 475.200 30.300 475.800 31.800 ;
        RECT 479.600 31.600 480.400 31.800 ;
        RECT 481.600 31.600 483.600 32.400 ;
        RECT 486.000 31.800 487.400 32.400 ;
        RECT 488.000 31.800 489.000 32.400 ;
        RECT 486.000 31.600 486.800 31.800 ;
        RECT 471.700 29.700 475.800 30.300 ;
        RECT 475.200 28.400 475.800 29.700 ;
        RECT 476.400 28.800 477.200 30.400 ;
        RECT 481.600 28.400 482.200 31.600 ;
        RECT 482.800 28.800 483.600 30.400 ;
        RECT 488.000 28.400 488.600 31.800 ;
        RECT 489.200 28.800 490.000 30.400 ;
        RECT 465.200 28.300 466.000 28.400 ;
        RECT 466.800 28.300 467.600 28.400 ;
        RECT 465.200 28.200 467.600 28.300 ;
        RECT 465.200 27.700 468.400 28.200 ;
        RECT 465.200 27.600 466.000 27.700 ;
        RECT 466.800 27.600 468.400 27.700 ;
        RECT 469.800 27.600 472.400 28.400 ;
        RECT 473.200 27.600 475.800 28.400 ;
        RECT 478.000 28.200 478.800 28.400 ;
        RECT 477.200 27.600 478.800 28.200 ;
        RECT 479.600 27.600 482.200 28.400 ;
        RECT 484.400 28.200 485.200 28.400 ;
        RECT 483.600 27.600 485.200 28.200 ;
        RECT 486.000 27.600 488.600 28.400 ;
        RECT 490.800 28.300 491.600 28.400 ;
        RECT 492.400 28.300 493.200 39.800 ;
        RECT 497.200 32.000 498.000 39.800 ;
        RECT 500.400 35.200 501.200 39.800 ;
        RECT 490.800 28.200 493.200 28.300 ;
        RECT 490.000 27.700 493.200 28.200 ;
        RECT 490.000 27.600 491.600 27.700 ;
        RECT 467.600 27.200 468.400 27.600 ;
        RECT 463.600 26.000 464.600 26.800 ;
        RECT 467.000 26.200 470.600 26.600 ;
        RECT 471.600 26.200 472.200 27.600 ;
        RECT 473.400 26.200 474.000 27.600 ;
        RECT 477.200 27.200 478.000 27.600 ;
        RECT 475.000 26.200 478.600 26.600 ;
        RECT 479.800 26.200 480.400 27.600 ;
        RECT 483.600 27.200 484.400 27.600 ;
        RECT 481.400 26.200 485.000 26.600 ;
        RECT 486.200 26.200 486.800 27.600 ;
        RECT 490.000 27.200 490.800 27.600 ;
        RECT 487.800 26.200 491.400 26.600 ;
        RECT 466.800 26.000 470.800 26.200 ;
        RECT 463.600 22.200 464.400 26.000 ;
        RECT 466.800 22.200 467.600 26.000 ;
        RECT 470.000 22.200 470.800 26.000 ;
        RECT 471.600 22.200 472.400 26.200 ;
        RECT 473.200 22.200 474.000 26.200 ;
        RECT 474.800 26.000 478.800 26.200 ;
        RECT 474.800 22.200 475.600 26.000 ;
        RECT 478.000 22.200 478.800 26.000 ;
        RECT 479.600 22.200 480.400 26.200 ;
        RECT 481.200 26.000 485.200 26.200 ;
        RECT 481.200 22.200 482.000 26.000 ;
        RECT 484.400 22.200 485.200 26.000 ;
        RECT 486.000 22.200 486.800 26.200 ;
        RECT 487.600 26.000 491.600 26.200 ;
        RECT 487.600 22.200 488.400 26.000 ;
        RECT 490.800 22.200 491.600 26.000 ;
        RECT 492.400 22.200 493.200 27.700 ;
        RECT 497.000 31.200 498.000 32.000 ;
        RECT 498.600 34.600 501.200 35.200 ;
        RECT 498.600 33.000 499.200 34.600 ;
        RECT 503.600 34.400 504.400 39.800 ;
        RECT 506.800 37.000 507.600 39.800 ;
        RECT 508.400 37.000 509.200 39.800 ;
        RECT 510.000 37.000 510.800 39.800 ;
        RECT 505.000 34.400 509.200 35.200 ;
        RECT 501.800 33.600 504.400 34.400 ;
        RECT 511.600 33.600 512.400 39.800 ;
        RECT 514.800 35.000 515.600 39.800 ;
        RECT 518.000 35.000 518.800 39.800 ;
        RECT 519.600 37.000 520.400 39.800 ;
        RECT 521.200 37.000 522.000 39.800 ;
        RECT 524.400 35.200 525.200 39.800 ;
        RECT 527.600 36.400 528.400 39.800 ;
        RECT 527.600 35.800 528.600 36.400 ;
        RECT 528.000 35.200 528.600 35.800 ;
        RECT 523.200 34.400 527.400 35.200 ;
        RECT 528.000 34.600 530.000 35.200 ;
        RECT 514.800 33.600 517.400 34.400 ;
        RECT 518.000 33.800 523.800 34.400 ;
        RECT 526.800 34.000 527.400 34.400 ;
        RECT 506.800 33.000 507.600 33.200 ;
        RECT 498.600 32.400 507.600 33.000 ;
        RECT 510.000 33.000 510.800 33.200 ;
        RECT 518.000 33.000 518.600 33.800 ;
        RECT 524.400 33.200 525.800 33.800 ;
        RECT 526.800 33.200 528.400 34.000 ;
        RECT 510.000 32.400 518.600 33.000 ;
        RECT 519.600 33.000 525.800 33.200 ;
        RECT 519.600 32.600 525.000 33.000 ;
        RECT 519.600 32.400 520.400 32.600 ;
        RECT 497.000 26.800 497.800 31.200 ;
        RECT 498.600 30.600 499.200 32.400 ;
        RECT 498.400 30.000 499.200 30.600 ;
        RECT 505.200 30.000 528.600 30.600 ;
        RECT 498.400 28.000 499.000 30.000 ;
        RECT 505.200 29.400 506.000 30.000 ;
        RECT 522.800 29.600 523.600 30.000 ;
        RECT 527.800 29.800 528.600 30.000 ;
        RECT 499.600 28.600 503.400 29.400 ;
        RECT 498.400 27.400 499.600 28.000 ;
        RECT 497.000 26.000 498.000 26.800 ;
        RECT 497.200 22.200 498.000 26.000 ;
        RECT 498.800 22.200 499.600 27.400 ;
        RECT 502.600 27.400 503.400 28.600 ;
        RECT 502.600 26.800 504.400 27.400 ;
        RECT 503.600 26.200 504.400 26.800 ;
        RECT 508.400 26.400 509.200 29.200 ;
        RECT 511.600 28.600 514.800 29.400 ;
        RECT 518.600 28.600 520.600 29.400 ;
        RECT 529.200 29.000 530.000 34.600 ;
        RECT 531.600 33.600 532.400 34.400 ;
        RECT 531.600 32.400 532.200 33.600 ;
        RECT 533.000 32.400 533.800 39.800 ;
        RECT 530.800 31.800 532.200 32.400 ;
        RECT 532.800 31.800 533.800 32.400 ;
        RECT 539.800 32.400 540.600 39.800 ;
        RECT 541.200 33.600 542.000 34.400 ;
        RECT 541.400 32.400 542.000 33.600 ;
        RECT 544.400 33.600 545.200 34.400 ;
        RECT 544.400 32.400 545.000 33.600 ;
        RECT 545.800 32.400 546.600 39.800 ;
        RECT 539.800 31.800 540.800 32.400 ;
        RECT 541.400 31.800 542.800 32.400 ;
        RECT 530.800 31.600 531.600 31.800 ;
        RECT 530.800 30.300 531.600 30.400 ;
        RECT 532.800 30.300 533.400 31.800 ;
        RECT 530.800 29.700 533.400 30.300 ;
        RECT 530.800 29.600 531.600 29.700 ;
        RECT 511.200 27.800 512.000 28.000 ;
        RECT 511.200 27.200 515.600 27.800 ;
        RECT 514.800 27.000 515.600 27.200 ;
        RECT 516.400 26.800 517.200 28.400 ;
        RECT 503.600 25.400 506.000 26.200 ;
        RECT 508.400 25.600 509.400 26.400 ;
        RECT 512.400 25.600 514.000 26.400 ;
        RECT 514.800 26.200 515.600 26.400 ;
        RECT 518.600 26.200 519.400 28.600 ;
        RECT 521.200 28.200 530.000 29.000 ;
        RECT 532.800 28.400 533.400 29.700 ;
        RECT 534.000 30.300 534.800 30.400 ;
        RECT 538.800 30.300 539.600 30.400 ;
        RECT 534.000 29.700 539.600 30.300 ;
        RECT 534.000 28.800 534.800 29.700 ;
        RECT 538.800 28.800 539.600 29.700 ;
        RECT 540.200 28.400 540.800 31.800 ;
        RECT 542.000 31.600 542.800 31.800 ;
        RECT 543.600 31.800 545.000 32.400 ;
        RECT 545.600 31.800 546.600 32.400 ;
        RECT 552.600 32.400 553.400 39.800 ;
        RECT 554.000 33.600 554.800 34.400 ;
        RECT 554.200 32.400 554.800 33.600 ;
        RECT 552.600 31.800 553.600 32.400 ;
        RECT 554.200 31.800 555.600 32.400 ;
        RECT 543.600 31.600 544.400 31.800 ;
        RECT 542.100 30.300 542.700 31.600 ;
        RECT 545.600 30.300 546.200 31.800 ;
        RECT 542.100 29.700 546.200 30.300 ;
        RECT 545.600 28.400 546.200 29.700 ;
        RECT 546.800 28.800 547.600 30.400 ;
        RECT 551.600 28.800 552.400 30.400 ;
        RECT 553.000 28.400 553.600 31.800 ;
        RECT 554.800 31.600 555.600 31.800 ;
        RECT 556.400 31.600 557.200 33.200 ;
        RECT 554.900 30.300 555.500 31.600 ;
        RECT 558.000 30.300 558.800 39.800 ;
        RECT 565.000 38.400 565.800 39.800 ;
        RECT 564.400 37.600 565.800 38.400 ;
        RECT 565.000 32.800 565.800 37.600 ;
        RECT 569.200 35.000 570.000 39.000 ;
        RECT 564.200 32.200 565.800 32.800 ;
        RECT 554.900 29.700 558.800 30.300 ;
        RECT 524.600 26.800 527.600 27.600 ;
        RECT 524.600 26.200 525.400 26.800 ;
        RECT 514.800 25.600 519.400 26.200 ;
        RECT 505.200 22.200 506.000 25.400 ;
        RECT 522.800 25.400 525.400 26.200 ;
        RECT 506.800 22.200 507.600 25.000 ;
        RECT 508.400 22.200 509.200 25.000 ;
        RECT 510.000 22.200 510.800 25.000 ;
        RECT 511.600 22.200 512.400 25.000 ;
        RECT 514.800 22.200 515.600 25.000 ;
        RECT 518.000 22.200 518.800 25.000 ;
        RECT 519.600 22.200 520.400 25.000 ;
        RECT 521.200 22.200 522.000 25.000 ;
        RECT 522.800 22.200 523.600 25.400 ;
        RECT 529.200 22.200 530.000 28.200 ;
        RECT 530.800 27.600 533.400 28.400 ;
        RECT 535.600 28.200 536.400 28.400 ;
        RECT 534.800 27.600 536.400 28.200 ;
        RECT 537.200 28.200 538.000 28.400 ;
        RECT 537.200 27.600 538.800 28.200 ;
        RECT 540.200 27.600 542.800 28.400 ;
        RECT 543.600 27.600 546.200 28.400 ;
        RECT 548.400 28.300 549.200 28.400 ;
        RECT 550.000 28.300 550.800 28.400 ;
        RECT 548.400 28.200 550.800 28.300 ;
        RECT 547.600 27.700 551.600 28.200 ;
        RECT 547.600 27.600 549.200 27.700 ;
        RECT 550.000 27.600 551.600 27.700 ;
        RECT 553.000 27.600 555.600 28.400 ;
        RECT 531.000 26.200 531.600 27.600 ;
        RECT 534.800 27.200 535.600 27.600 ;
        RECT 538.000 27.200 538.800 27.600 ;
        RECT 532.600 26.200 536.200 26.600 ;
        RECT 537.400 26.200 541.000 26.600 ;
        RECT 542.000 26.200 542.600 27.600 ;
        RECT 543.800 26.200 544.400 27.600 ;
        RECT 547.600 27.200 548.400 27.600 ;
        RECT 550.800 27.200 551.600 27.600 ;
        RECT 545.400 26.200 549.000 26.600 ;
        RECT 550.200 26.200 553.800 26.600 ;
        RECT 554.800 26.200 555.400 27.600 ;
        RECT 558.000 26.200 558.800 29.700 ;
        RECT 559.600 30.300 560.400 30.400 ;
        RECT 562.800 30.300 563.600 31.200 ;
        RECT 559.600 29.700 563.600 30.300 ;
        RECT 559.600 29.600 560.400 29.700 ;
        RECT 562.800 29.600 563.600 29.700 ;
        RECT 564.200 28.400 564.800 32.200 ;
        RECT 569.400 31.600 570.000 35.000 ;
        RECT 572.400 34.300 573.200 34.400 ;
        RECT 575.600 34.300 576.400 39.800 ;
        RECT 579.800 35.800 581.000 39.800 ;
        RECT 584.400 35.800 585.200 39.800 ;
        RECT 588.800 36.400 589.600 39.800 ;
        RECT 588.800 35.800 590.800 36.400 ;
        RECT 580.400 35.000 581.200 35.800 ;
        RECT 584.600 35.200 585.200 35.800 ;
        RECT 583.800 34.600 587.400 35.200 ;
        RECT 590.000 35.000 590.800 35.800 ;
        RECT 583.800 34.400 584.600 34.600 ;
        RECT 586.600 34.400 587.400 34.600 ;
        RECT 572.400 33.700 576.400 34.300 ;
        RECT 572.400 33.600 573.200 33.700 ;
        RECT 566.200 31.000 570.000 31.600 ;
        RECT 575.600 31.200 576.400 33.700 ;
        RECT 579.600 33.200 581.000 34.000 ;
        RECT 580.400 32.200 581.000 33.200 ;
        RECT 582.600 33.000 584.800 33.600 ;
        RECT 582.600 32.800 583.400 33.000 ;
        RECT 580.400 31.600 582.800 32.200 ;
        RECT 566.200 29.000 566.800 31.000 ;
        RECT 575.600 30.600 579.800 31.200 ;
        RECT 559.600 26.800 560.400 28.400 ;
        RECT 562.800 27.600 564.800 28.400 ;
        RECT 565.400 28.200 566.800 29.000 ;
        RECT 567.600 28.800 568.400 30.400 ;
        RECT 569.200 28.800 570.000 30.400 ;
        RECT 564.200 27.000 564.800 27.600 ;
        RECT 565.800 27.800 566.800 28.200 ;
        RECT 565.800 27.200 570.000 27.800 ;
        RECT 530.800 22.200 531.600 26.200 ;
        RECT 532.400 26.000 536.400 26.200 ;
        RECT 532.400 22.200 533.200 26.000 ;
        RECT 535.600 22.200 536.400 26.000 ;
        RECT 537.200 26.000 541.200 26.200 ;
        RECT 537.200 22.200 538.000 26.000 ;
        RECT 540.400 22.200 541.200 26.000 ;
        RECT 542.000 22.200 542.800 26.200 ;
        RECT 543.600 22.200 544.400 26.200 ;
        RECT 545.200 26.000 549.200 26.200 ;
        RECT 545.200 22.200 546.000 26.000 ;
        RECT 548.400 22.200 549.200 26.000 ;
        RECT 550.000 26.000 554.000 26.200 ;
        RECT 550.000 22.200 550.800 26.000 ;
        RECT 553.200 22.200 554.000 26.000 ;
        RECT 554.800 22.200 555.600 26.200 ;
        RECT 557.000 25.600 558.800 26.200 ;
        RECT 564.200 26.600 565.000 27.000 ;
        RECT 564.200 26.000 565.800 26.600 ;
        RECT 557.000 22.200 557.800 25.600 ;
        RECT 565.000 23.000 565.800 26.000 ;
        RECT 569.400 25.000 570.000 27.200 ;
        RECT 569.200 23.000 570.000 25.000 ;
        RECT 575.600 27.200 576.400 30.600 ;
        RECT 579.000 30.400 579.800 30.600 ;
        RECT 577.400 29.800 578.200 30.000 ;
        RECT 577.400 29.200 581.200 29.800 ;
        RECT 580.400 29.000 581.200 29.200 ;
        RECT 582.200 28.400 582.800 31.600 ;
        RECT 584.200 31.800 584.800 33.000 ;
        RECT 585.400 33.000 586.200 33.200 ;
        RECT 590.000 33.000 590.800 33.200 ;
        RECT 585.400 32.400 590.800 33.000 ;
        RECT 584.200 31.400 589.000 31.800 ;
        RECT 593.200 31.400 594.000 39.800 ;
        RECT 584.200 31.200 594.000 31.400 ;
        RECT 588.200 31.000 594.000 31.200 ;
        RECT 588.400 30.800 594.000 31.000 ;
        RECT 583.600 30.300 584.400 30.400 ;
        RECT 586.800 30.300 587.600 30.400 ;
        RECT 583.600 30.200 587.600 30.300 ;
        RECT 583.600 29.700 591.800 30.200 ;
        RECT 583.600 29.600 584.400 29.700 ;
        RECT 586.800 29.600 591.800 29.700 ;
        RECT 591.000 29.400 591.800 29.600 ;
        RECT 589.400 28.400 590.200 28.600 ;
        RECT 582.000 27.800 593.200 28.400 ;
        RECT 582.000 27.600 583.400 27.800 ;
        RECT 575.600 26.600 579.400 27.200 ;
        RECT 575.600 22.200 576.400 26.600 ;
        RECT 578.600 26.400 579.400 26.600 ;
        RECT 588.400 25.600 589.000 27.800 ;
        RECT 591.600 27.600 593.200 27.800 ;
        RECT 586.600 25.400 587.400 25.600 ;
        RECT 580.400 24.200 581.200 25.000 ;
        RECT 584.600 24.800 587.400 25.400 ;
        RECT 588.400 24.800 589.200 25.600 ;
        RECT 584.600 24.200 585.200 24.800 ;
        RECT 590.000 24.200 590.800 25.000 ;
        RECT 579.800 23.600 581.200 24.200 ;
        RECT 579.800 22.200 581.000 23.600 ;
        RECT 584.400 22.200 585.200 24.200 ;
        RECT 588.800 23.600 590.800 24.200 ;
        RECT 588.800 22.200 589.600 23.600 ;
        RECT 593.200 22.200 594.000 27.000 ;
        RECT 594.800 22.200 595.600 39.800 ;
        RECT 598.000 31.200 598.800 39.800 ;
        RECT 602.200 35.800 603.400 39.800 ;
        RECT 606.800 35.800 607.600 39.800 ;
        RECT 611.200 36.400 612.000 39.800 ;
        RECT 611.200 35.800 613.200 36.400 ;
        RECT 602.800 35.000 603.600 35.800 ;
        RECT 607.000 35.200 607.600 35.800 ;
        RECT 606.200 34.600 609.800 35.200 ;
        RECT 612.400 35.000 613.200 35.800 ;
        RECT 606.200 34.400 607.000 34.600 ;
        RECT 609.000 34.400 609.800 34.600 ;
        RECT 602.000 33.200 603.400 34.000 ;
        RECT 602.800 32.200 603.400 33.200 ;
        RECT 605.000 33.000 607.200 33.600 ;
        RECT 605.000 32.800 605.800 33.000 ;
        RECT 602.800 31.600 605.200 32.200 ;
        RECT 598.000 30.600 602.200 31.200 ;
        RECT 598.000 27.200 598.800 30.600 ;
        RECT 601.400 30.400 602.200 30.600 ;
        RECT 599.800 29.800 600.600 30.000 ;
        RECT 599.800 29.200 603.600 29.800 ;
        RECT 602.800 29.000 603.600 29.200 ;
        RECT 604.600 28.400 605.200 31.600 ;
        RECT 606.600 31.800 607.200 33.000 ;
        RECT 607.800 33.000 608.600 33.200 ;
        RECT 612.400 33.000 613.200 33.200 ;
        RECT 607.800 32.400 613.200 33.000 ;
        RECT 606.600 31.400 611.400 31.800 ;
        RECT 615.600 31.400 616.400 39.800 ;
        RECT 619.800 32.400 620.600 39.800 ;
        RECT 625.800 34.400 626.600 39.800 ;
        RECT 621.200 33.600 622.000 34.400 ;
        RECT 621.400 32.400 622.000 33.600 ;
        RECT 624.400 33.600 625.200 34.400 ;
        RECT 625.800 33.600 627.600 34.400 ;
        RECT 624.400 32.400 625.000 33.600 ;
        RECT 625.800 32.400 626.600 33.600 ;
        RECT 633.800 32.800 634.600 39.800 ;
        RECT 638.000 35.000 638.800 39.000 ;
        RECT 619.800 31.800 620.800 32.400 ;
        RECT 621.400 31.800 622.800 32.400 ;
        RECT 606.600 31.200 616.400 31.400 ;
        RECT 610.600 31.000 616.400 31.200 ;
        RECT 610.800 30.800 616.400 31.000 ;
        RECT 609.200 30.200 610.000 30.400 ;
        RECT 609.200 29.600 614.200 30.200 ;
        RECT 610.800 29.400 611.600 29.600 ;
        RECT 613.400 29.400 614.200 29.600 ;
        RECT 618.800 28.800 619.600 30.400 ;
        RECT 620.200 30.300 620.800 31.800 ;
        RECT 622.000 31.600 622.800 31.800 ;
        RECT 623.600 31.800 625.000 32.400 ;
        RECT 625.600 31.800 626.600 32.400 ;
        RECT 633.000 32.200 634.600 32.800 ;
        RECT 623.600 31.600 624.400 31.800 ;
        RECT 623.700 30.300 624.300 31.600 ;
        RECT 620.200 29.700 624.300 30.300 ;
        RECT 611.800 28.400 612.600 28.600 ;
        RECT 620.200 28.400 620.800 29.700 ;
        RECT 625.600 28.400 626.200 31.800 ;
        RECT 626.800 30.300 627.600 30.400 ;
        RECT 626.800 29.700 630.700 30.300 ;
        RECT 626.800 28.800 627.600 29.700 ;
        RECT 604.400 27.800 615.600 28.400 ;
        RECT 604.400 27.600 605.800 27.800 ;
        RECT 598.000 26.600 601.800 27.200 ;
        RECT 596.400 26.300 597.200 26.400 ;
        RECT 598.000 26.300 598.800 26.600 ;
        RECT 601.000 26.400 601.800 26.600 ;
        RECT 596.400 25.700 598.800 26.300 ;
        RECT 596.400 24.800 597.200 25.700 ;
        RECT 598.000 22.200 598.800 25.700 ;
        RECT 610.800 25.600 611.400 27.800 ;
        RECT 614.000 27.600 615.600 27.800 ;
        RECT 617.200 28.200 618.000 28.400 ;
        RECT 617.200 27.600 618.800 28.200 ;
        RECT 620.200 27.600 622.800 28.400 ;
        RECT 623.600 27.600 626.200 28.400 ;
        RECT 628.400 28.200 629.200 28.400 ;
        RECT 627.600 27.600 629.200 28.200 ;
        RECT 630.100 28.300 630.700 29.700 ;
        RECT 631.600 29.600 632.400 31.200 ;
        RECT 633.000 28.400 633.600 32.200 ;
        RECT 638.200 31.600 638.800 35.000 ;
        RECT 635.000 31.000 638.800 31.600 ;
        RECT 639.600 35.000 640.400 39.000 ;
        RECT 639.600 31.600 640.200 35.000 ;
        RECT 643.800 32.800 644.600 39.800 ;
        RECT 643.800 32.200 645.400 32.800 ;
        RECT 639.600 31.000 643.400 31.600 ;
        RECT 635.000 29.000 635.600 31.000 ;
        RECT 631.600 28.300 633.600 28.400 ;
        RECT 630.100 27.700 633.600 28.300 ;
        RECT 634.200 28.200 635.600 29.000 ;
        RECT 636.400 28.800 637.200 30.400 ;
        RECT 638.000 30.300 638.800 30.400 ;
        RECT 639.600 30.300 640.400 30.400 ;
        RECT 638.000 29.700 640.400 30.300 ;
        RECT 638.000 28.800 638.800 29.700 ;
        RECT 639.600 28.800 640.400 29.700 ;
        RECT 641.200 28.800 642.000 30.400 ;
        RECT 642.800 29.000 643.400 31.000 ;
        RECT 631.600 27.600 633.600 27.700 ;
        RECT 618.000 27.200 618.800 27.600 ;
        RECT 609.000 25.400 609.800 25.600 ;
        RECT 602.800 24.200 603.600 25.000 ;
        RECT 607.000 24.800 609.800 25.400 ;
        RECT 610.800 24.800 611.600 25.600 ;
        RECT 607.000 24.200 607.600 24.800 ;
        RECT 612.400 24.200 613.200 25.000 ;
        RECT 602.200 23.600 603.600 24.200 ;
        RECT 602.200 22.200 603.400 23.600 ;
        RECT 606.800 22.200 607.600 24.200 ;
        RECT 611.200 23.600 613.200 24.200 ;
        RECT 611.200 22.200 612.000 23.600 ;
        RECT 615.600 22.200 616.400 27.000 ;
        RECT 617.400 26.200 621.000 26.600 ;
        RECT 622.000 26.200 622.600 27.600 ;
        RECT 623.800 26.200 624.400 27.600 ;
        RECT 627.600 27.200 628.400 27.600 ;
        RECT 633.000 27.000 633.600 27.600 ;
        RECT 634.600 27.800 635.600 28.200 ;
        RECT 642.800 28.200 644.200 29.000 ;
        RECT 644.800 28.400 645.400 32.200 ;
        RECT 651.800 32.400 652.600 39.800 ;
        RECT 653.200 33.600 654.000 34.400 ;
        RECT 653.400 32.400 654.000 33.600 ;
        RECT 656.400 33.600 657.200 34.400 ;
        RECT 656.400 32.400 657.000 33.600 ;
        RECT 657.800 32.400 658.600 39.800 ;
        RECT 651.800 31.800 652.800 32.400 ;
        RECT 653.400 31.800 654.800 32.400 ;
        RECT 646.000 30.300 646.800 31.200 ;
        RECT 647.600 30.300 648.400 30.400 ;
        RECT 646.000 29.700 648.400 30.300 ;
        RECT 646.000 29.600 646.800 29.700 ;
        RECT 647.600 29.600 648.400 29.700 ;
        RECT 650.800 28.800 651.600 30.400 ;
        RECT 652.200 30.300 652.800 31.800 ;
        RECT 654.000 31.600 654.800 31.800 ;
        RECT 655.600 31.800 657.000 32.400 ;
        RECT 657.600 31.800 658.600 32.400 ;
        RECT 664.600 32.400 665.400 39.800 ;
        RECT 670.600 38.400 671.400 39.800 ;
        RECT 670.600 37.600 672.400 38.400 ;
        RECT 666.000 33.600 666.800 34.400 ;
        RECT 666.200 32.400 666.800 33.600 ;
        RECT 669.200 33.600 670.000 34.400 ;
        RECT 669.200 32.400 669.800 33.600 ;
        RECT 670.600 32.400 671.400 37.600 ;
        RECT 664.600 31.800 665.600 32.400 ;
        RECT 666.200 31.800 667.600 32.400 ;
        RECT 655.600 31.600 656.400 31.800 ;
        RECT 655.700 30.300 656.300 31.600 ;
        RECT 652.200 29.700 656.300 30.300 ;
        RECT 652.200 28.400 652.800 29.700 ;
        RECT 657.600 28.400 658.200 31.800 ;
        RECT 658.800 28.800 659.600 30.400 ;
        RECT 660.400 30.300 661.200 30.400 ;
        RECT 663.600 30.300 664.400 30.400 ;
        RECT 660.400 29.700 664.400 30.300 ;
        RECT 660.400 29.600 661.200 29.700 ;
        RECT 663.600 28.800 664.400 29.700 ;
        RECT 665.000 30.300 665.600 31.800 ;
        RECT 666.800 31.600 667.600 31.800 ;
        RECT 668.400 31.800 669.800 32.400 ;
        RECT 670.400 31.800 671.400 32.400 ;
        RECT 674.800 32.400 675.600 39.800 ;
        RECT 679.200 38.400 680.800 39.800 ;
        RECT 679.200 37.600 682.000 38.400 ;
        RECT 676.400 32.400 677.200 32.600 ;
        RECT 679.200 32.400 680.800 37.600 ;
        RECT 674.800 31.800 677.200 32.400 ;
        RECT 678.800 31.800 680.800 32.400 ;
        RECT 683.000 32.400 683.800 32.600 ;
        RECT 684.400 32.400 685.200 39.800 ;
        RECT 683.000 31.800 685.200 32.400 ;
        RECT 668.400 31.600 669.200 31.800 ;
        RECT 668.500 30.300 669.100 31.600 ;
        RECT 665.000 29.700 669.100 30.300 ;
        RECT 665.000 28.400 665.600 29.700 ;
        RECT 670.400 28.400 671.000 31.800 ;
        RECT 678.800 30.400 679.400 31.800 ;
        RECT 683.000 31.200 683.600 31.800 ;
        RECT 680.200 30.600 683.600 31.200 ;
        RECT 680.200 30.400 681.000 30.600 ;
        RECT 671.600 28.800 672.400 30.400 ;
        RECT 678.000 29.800 679.400 30.400 ;
        RECT 682.400 29.800 683.200 30.000 ;
        RECT 678.000 29.600 679.800 29.800 ;
        RECT 678.800 29.200 679.800 29.600 ;
        RECT 644.800 28.300 646.800 28.400 ;
        RECT 647.600 28.300 648.400 28.400 ;
        RECT 642.800 27.800 643.800 28.200 ;
        RECT 634.600 27.200 638.800 27.800 ;
        RECT 633.000 26.600 633.800 27.000 ;
        RECT 625.400 26.200 629.000 26.600 ;
        RECT 617.200 26.000 621.200 26.200 ;
        RECT 617.200 22.200 618.000 26.000 ;
        RECT 620.400 22.200 621.200 26.000 ;
        RECT 622.000 22.200 622.800 26.200 ;
        RECT 623.600 22.200 624.400 26.200 ;
        RECT 625.200 26.000 629.200 26.200 ;
        RECT 633.000 26.000 634.600 26.600 ;
        RECT 625.200 22.200 626.000 26.000 ;
        RECT 628.400 22.200 629.200 26.000 ;
        RECT 633.800 23.000 634.600 26.000 ;
        RECT 638.200 25.000 638.800 27.200 ;
        RECT 638.000 23.000 638.800 25.000 ;
        RECT 639.600 27.200 643.800 27.800 ;
        RECT 644.800 27.700 648.400 28.300 ;
        RECT 644.800 27.600 646.800 27.700 ;
        RECT 647.600 27.600 648.400 27.700 ;
        RECT 649.200 28.200 650.000 28.400 ;
        RECT 649.200 27.600 650.800 28.200 ;
        RECT 652.200 27.600 654.800 28.400 ;
        RECT 655.600 27.600 658.200 28.400 ;
        RECT 660.400 28.200 661.200 28.400 ;
        RECT 659.600 27.600 661.200 28.200 ;
        RECT 662.000 28.200 662.800 28.400 ;
        RECT 662.000 27.600 663.600 28.200 ;
        RECT 665.000 27.600 667.600 28.400 ;
        RECT 668.400 27.600 671.000 28.400 ;
        RECT 673.200 28.200 674.000 28.400 ;
        RECT 672.400 27.600 674.000 28.200 ;
        RECT 674.800 27.600 676.400 28.400 ;
        RECT 677.600 27.600 678.400 28.400 ;
        RECT 639.600 25.000 640.200 27.200 ;
        RECT 644.800 27.000 645.400 27.600 ;
        RECT 650.000 27.200 650.800 27.600 ;
        RECT 644.600 26.600 645.400 27.000 ;
        RECT 643.800 26.000 645.400 26.600 ;
        RECT 649.400 26.200 653.000 26.600 ;
        RECT 654.000 26.200 654.600 27.600 ;
        RECT 655.800 26.200 656.400 27.600 ;
        RECT 659.600 27.200 660.400 27.600 ;
        RECT 662.800 27.200 663.600 27.600 ;
        RECT 657.400 26.200 661.000 26.600 ;
        RECT 662.200 26.200 665.800 26.600 ;
        RECT 666.800 26.200 667.400 27.600 ;
        RECT 668.600 26.200 669.200 27.600 ;
        RECT 672.400 27.200 673.200 27.600 ;
        RECT 677.800 27.200 678.400 27.600 ;
        RECT 676.400 26.800 677.200 27.000 ;
        RECT 670.200 26.200 673.800 26.600 ;
        RECT 674.800 26.200 677.200 26.800 ;
        RECT 677.800 26.400 678.600 27.200 ;
        RECT 649.200 26.000 653.200 26.200 ;
        RECT 639.600 23.000 640.400 25.000 ;
        RECT 643.800 23.000 644.600 26.000 ;
        RECT 649.200 22.200 650.000 26.000 ;
        RECT 652.400 22.200 653.200 26.000 ;
        RECT 654.000 22.200 654.800 26.200 ;
        RECT 655.600 22.200 656.400 26.200 ;
        RECT 657.200 26.000 661.200 26.200 ;
        RECT 657.200 22.200 658.000 26.000 ;
        RECT 660.400 22.200 661.200 26.000 ;
        RECT 662.000 26.000 666.000 26.200 ;
        RECT 662.000 22.200 662.800 26.000 ;
        RECT 665.200 22.200 666.000 26.000 ;
        RECT 666.800 22.200 667.600 26.200 ;
        RECT 668.400 22.200 669.200 26.200 ;
        RECT 670.000 26.000 674.000 26.200 ;
        RECT 670.000 22.200 670.800 26.000 ;
        RECT 673.200 22.200 674.000 26.000 ;
        RECT 674.800 22.200 675.600 26.200 ;
        RECT 679.200 25.800 679.800 29.200 ;
        RECT 680.600 29.200 683.200 29.800 ;
        RECT 680.600 28.600 681.200 29.200 ;
        RECT 680.400 27.800 681.200 28.600 ;
        RECT 683.600 28.200 685.200 28.400 ;
        RECT 681.800 27.600 685.200 28.200 ;
        RECT 681.800 27.200 682.400 27.600 ;
        RECT 680.400 26.600 682.400 27.200 ;
        RECT 683.000 26.800 683.800 27.000 ;
        RECT 680.400 26.400 682.000 26.600 ;
        RECT 683.000 26.200 685.200 26.800 ;
        RECT 679.200 22.200 680.800 25.800 ;
        RECT 684.400 22.200 685.200 26.200 ;
        RECT 1.200 15.600 2.000 17.200 ;
        RECT 2.800 2.200 3.600 19.800 ;
        RECT 4.400 13.800 5.200 19.800 ;
        RECT 10.800 16.600 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 14.000 17.000 14.800 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 26.800 17.000 27.600 19.800 ;
        RECT 9.000 15.800 11.600 16.600 ;
        RECT 28.400 16.600 29.200 19.800 ;
        RECT 15.000 15.800 19.600 16.400 ;
        RECT 9.000 15.200 9.800 15.800 ;
        RECT 6.800 14.400 9.800 15.200 ;
        RECT 4.400 13.000 13.200 13.800 ;
        RECT 15.000 13.400 15.800 15.800 ;
        RECT 18.800 15.600 19.600 15.800 ;
        RECT 20.400 15.600 22.000 16.400 ;
        RECT 25.000 15.600 26.000 16.400 ;
        RECT 28.400 15.800 30.800 16.600 ;
        RECT 17.200 13.600 18.000 15.200 ;
        RECT 18.800 14.800 19.600 15.000 ;
        RECT 18.800 14.200 23.200 14.800 ;
        RECT 22.400 14.000 23.200 14.200 ;
        RECT 4.400 7.400 5.200 13.000 ;
        RECT 13.800 12.600 15.800 13.400 ;
        RECT 19.600 12.600 22.800 13.400 ;
        RECT 25.200 12.800 26.000 15.600 ;
        RECT 30.000 15.200 30.800 15.800 ;
        RECT 30.000 14.600 31.800 15.200 ;
        RECT 31.000 13.400 31.800 14.600 ;
        RECT 34.800 14.600 35.600 19.800 ;
        RECT 36.400 16.300 37.200 19.800 ;
        RECT 38.000 16.300 38.800 16.400 ;
        RECT 36.400 15.700 38.800 16.300 ;
        RECT 36.400 15.200 37.400 15.700 ;
        RECT 38.000 15.600 38.800 15.700 ;
        RECT 42.800 15.200 43.600 19.800 ;
        RECT 34.800 14.000 36.000 14.600 ;
        RECT 31.000 12.600 34.800 13.400 ;
        RECT 5.800 12.000 6.600 12.200 ;
        RECT 7.600 12.000 8.400 12.400 ;
        RECT 10.800 12.000 11.600 12.400 ;
        RECT 28.400 12.000 29.200 12.600 ;
        RECT 35.400 12.000 36.000 14.000 ;
        RECT 5.800 11.400 29.200 12.000 ;
        RECT 35.200 11.400 36.000 12.000 ;
        RECT 35.200 9.600 35.800 11.400 ;
        RECT 36.600 10.800 37.400 15.200 ;
        RECT 41.400 14.600 43.600 15.200 ;
        RECT 41.400 11.600 42.000 14.600 ;
        RECT 42.800 12.300 43.600 13.200 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 42.800 11.700 45.200 12.300 ;
        RECT 42.800 11.600 43.600 11.700 ;
        RECT 44.400 11.600 45.200 11.700 ;
        RECT 40.800 10.800 42.000 11.600 ;
        RECT 14.000 9.400 14.800 9.600 ;
        RECT 9.400 9.000 14.800 9.400 ;
        RECT 8.600 8.800 14.800 9.000 ;
        RECT 15.800 9.000 24.400 9.600 ;
        RECT 6.000 8.000 7.600 8.800 ;
        RECT 8.600 8.200 10.000 8.800 ;
        RECT 15.800 8.200 16.400 9.000 ;
        RECT 23.600 8.800 24.400 9.000 ;
        RECT 26.800 9.000 35.800 9.600 ;
        RECT 26.800 8.800 27.600 9.000 ;
        RECT 7.000 7.600 7.600 8.000 ;
        RECT 10.600 7.600 16.400 8.200 ;
        RECT 17.000 7.600 19.600 8.400 ;
        RECT 4.400 6.800 6.400 7.400 ;
        RECT 7.000 6.800 11.200 7.600 ;
        RECT 5.800 6.200 6.400 6.800 ;
        RECT 5.800 5.600 6.800 6.200 ;
        RECT 6.000 2.200 6.800 5.600 ;
        RECT 9.200 2.200 10.000 6.800 ;
        RECT 12.400 2.200 13.200 5.000 ;
        RECT 14.000 2.200 14.800 5.000 ;
        RECT 15.600 2.200 16.400 7.000 ;
        RECT 18.800 2.200 19.600 7.000 ;
        RECT 22.000 2.200 22.800 8.400 ;
        RECT 30.000 7.600 32.600 8.400 ;
        RECT 25.200 6.800 29.400 7.600 ;
        RECT 23.600 2.200 24.400 5.000 ;
        RECT 25.200 2.200 26.000 5.000 ;
        RECT 26.800 2.200 27.600 5.000 ;
        RECT 30.000 2.200 30.800 7.600 ;
        RECT 35.200 7.400 35.800 9.000 ;
        RECT 33.200 6.800 35.800 7.400 ;
        RECT 36.400 10.000 37.400 10.800 ;
        RECT 41.400 10.200 42.000 10.800 ;
        RECT 33.200 2.200 34.000 6.800 ;
        RECT 36.400 2.200 37.200 10.000 ;
        RECT 41.400 9.600 43.600 10.200 ;
        RECT 42.800 2.200 43.600 9.600 ;
        RECT 46.000 2.200 46.800 19.800 ;
        RECT 49.200 16.000 50.000 19.800 ;
        RECT 49.000 15.200 50.000 16.000 ;
        RECT 49.000 10.800 49.800 15.200 ;
        RECT 50.800 14.600 51.600 19.800 ;
        RECT 57.200 16.600 58.000 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 60.400 17.000 61.200 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 63.600 17.000 64.400 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 71.600 17.000 72.400 19.800 ;
        RECT 73.200 17.000 74.000 19.800 ;
        RECT 55.600 15.800 58.000 16.600 ;
        RECT 74.800 16.600 75.600 19.800 ;
        RECT 55.600 15.200 56.400 15.800 ;
        RECT 50.400 14.000 51.600 14.600 ;
        RECT 54.600 14.600 56.400 15.200 ;
        RECT 60.400 15.600 61.400 16.400 ;
        RECT 64.400 15.600 66.000 16.400 ;
        RECT 66.800 15.800 71.400 16.400 ;
        RECT 74.800 15.800 77.400 16.600 ;
        RECT 66.800 15.600 67.600 15.800 ;
        RECT 50.400 12.000 51.000 14.000 ;
        RECT 54.600 13.400 55.400 14.600 ;
        RECT 51.600 12.600 55.400 13.400 ;
        RECT 60.400 12.800 61.200 15.600 ;
        RECT 66.800 14.800 67.600 15.000 ;
        RECT 63.200 14.200 67.600 14.800 ;
        RECT 63.200 14.000 64.000 14.200 ;
        RECT 68.400 13.600 69.200 15.200 ;
        RECT 70.600 13.400 71.400 15.800 ;
        RECT 76.600 15.200 77.400 15.800 ;
        RECT 76.600 14.400 79.600 15.200 ;
        RECT 81.200 13.800 82.000 19.800 ;
        RECT 84.400 16.000 85.200 19.800 ;
        RECT 63.600 12.600 66.800 13.400 ;
        RECT 70.600 12.600 72.600 13.400 ;
        RECT 73.200 13.000 82.000 13.800 ;
        RECT 57.200 12.000 58.000 12.600 ;
        RECT 74.800 12.000 75.600 12.400 ;
        RECT 78.000 12.000 78.800 12.400 ;
        RECT 79.800 12.000 80.600 12.200 ;
        RECT 50.400 11.400 51.200 12.000 ;
        RECT 57.200 11.400 80.600 12.000 ;
        RECT 49.000 10.000 50.000 10.800 ;
        RECT 49.200 2.200 50.000 10.000 ;
        RECT 50.600 9.600 51.200 11.400 ;
        RECT 50.600 9.000 59.600 9.600 ;
        RECT 50.600 7.400 51.200 9.000 ;
        RECT 58.800 8.800 59.600 9.000 ;
        RECT 62.000 9.000 70.600 9.600 ;
        RECT 62.000 8.800 62.800 9.000 ;
        RECT 53.800 7.600 56.400 8.400 ;
        RECT 50.600 6.800 53.200 7.400 ;
        RECT 52.400 2.200 53.200 6.800 ;
        RECT 55.600 2.200 56.400 7.600 ;
        RECT 57.000 6.800 61.200 7.600 ;
        RECT 58.800 2.200 59.600 5.000 ;
        RECT 60.400 2.200 61.200 5.000 ;
        RECT 62.000 2.200 62.800 5.000 ;
        RECT 63.600 2.200 64.400 8.400 ;
        RECT 66.800 7.600 69.400 8.400 ;
        RECT 70.000 8.200 70.600 9.000 ;
        RECT 71.600 9.400 72.400 9.600 ;
        RECT 71.600 9.000 77.000 9.400 ;
        RECT 71.600 8.800 77.800 9.000 ;
        RECT 76.400 8.200 77.800 8.800 ;
        RECT 70.000 7.600 75.800 8.200 ;
        RECT 78.800 8.000 80.400 8.800 ;
        RECT 78.800 7.600 79.400 8.000 ;
        RECT 66.800 2.200 67.600 7.000 ;
        RECT 70.000 2.200 70.800 7.000 ;
        RECT 75.200 6.800 79.400 7.600 ;
        RECT 81.200 7.400 82.000 13.000 ;
        RECT 84.200 15.200 85.200 16.000 ;
        RECT 84.200 10.800 85.000 15.200 ;
        RECT 86.000 14.600 86.800 19.800 ;
        RECT 92.400 16.600 93.200 19.800 ;
        RECT 94.000 17.000 94.800 19.800 ;
        RECT 95.600 17.000 96.400 19.800 ;
        RECT 97.200 17.000 98.000 19.800 ;
        RECT 98.800 17.000 99.600 19.800 ;
        RECT 102.000 17.000 102.800 19.800 ;
        RECT 105.200 17.000 106.000 19.800 ;
        RECT 106.800 17.000 107.600 19.800 ;
        RECT 108.400 17.000 109.200 19.800 ;
        RECT 90.800 15.800 93.200 16.600 ;
        RECT 110.000 16.600 110.800 19.800 ;
        RECT 90.800 15.200 91.600 15.800 ;
        RECT 85.600 14.000 86.800 14.600 ;
        RECT 89.800 14.600 91.600 15.200 ;
        RECT 95.600 15.600 96.600 16.400 ;
        RECT 99.600 15.600 101.200 16.400 ;
        RECT 102.000 15.800 106.600 16.400 ;
        RECT 110.000 15.800 112.600 16.600 ;
        RECT 102.000 15.600 102.800 15.800 ;
        RECT 85.600 12.000 86.200 14.000 ;
        RECT 89.800 13.400 90.600 14.600 ;
        RECT 86.800 12.600 90.600 13.400 ;
        RECT 95.600 12.800 96.400 15.600 ;
        RECT 102.000 14.800 102.800 15.000 ;
        RECT 98.400 14.200 102.800 14.800 ;
        RECT 98.400 14.000 99.200 14.200 ;
        RECT 103.600 13.600 104.400 15.200 ;
        RECT 105.800 13.400 106.600 15.800 ;
        RECT 111.800 15.200 112.600 15.800 ;
        RECT 111.800 14.400 114.800 15.200 ;
        RECT 116.400 13.800 117.200 19.800 ;
        RECT 122.800 15.000 123.600 19.800 ;
        RECT 127.200 18.400 128.000 19.800 ;
        RECT 126.000 17.800 128.000 18.400 ;
        RECT 131.600 17.800 132.400 19.800 ;
        RECT 135.800 18.400 137.000 19.800 ;
        RECT 135.600 17.800 137.000 18.400 ;
        RECT 126.000 17.000 126.800 17.800 ;
        RECT 131.600 17.200 132.200 17.800 ;
        RECT 127.600 16.400 128.400 17.200 ;
        RECT 129.400 16.600 132.200 17.200 ;
        RECT 135.600 17.000 136.400 17.800 ;
        RECT 129.400 16.400 130.200 16.600 ;
        RECT 98.800 12.600 102.000 13.400 ;
        RECT 105.800 12.600 107.800 13.400 ;
        RECT 108.400 13.000 117.200 13.800 ;
        RECT 123.600 14.200 125.200 14.400 ;
        RECT 127.800 14.200 128.400 16.400 ;
        RECT 137.400 15.400 138.200 15.600 ;
        RECT 140.400 15.400 141.200 19.800 ;
        RECT 137.400 14.800 141.200 15.400 ;
        RECT 133.400 14.200 134.200 14.400 ;
        RECT 123.600 13.600 134.600 14.200 ;
        RECT 126.600 13.400 127.400 13.600 ;
        RECT 92.400 12.000 93.200 12.600 ;
        RECT 110.000 12.000 110.800 12.400 ;
        RECT 111.600 12.000 112.400 12.400 ;
        RECT 115.000 12.000 115.800 12.200 ;
        RECT 85.600 11.400 86.400 12.000 ;
        RECT 92.400 11.400 115.800 12.000 ;
        RECT 84.200 10.000 85.200 10.800 ;
        RECT 80.000 6.800 82.000 7.400 ;
        RECT 71.600 2.200 72.400 5.000 ;
        RECT 73.200 2.200 74.000 5.000 ;
        RECT 76.400 2.200 77.200 6.800 ;
        RECT 80.000 6.200 80.600 6.800 ;
        RECT 79.600 5.600 80.600 6.200 ;
        RECT 79.600 2.200 80.400 5.600 ;
        RECT 84.400 2.200 85.200 10.000 ;
        RECT 85.800 9.600 86.400 11.400 ;
        RECT 85.800 9.000 94.800 9.600 ;
        RECT 85.800 7.400 86.400 9.000 ;
        RECT 94.000 8.800 94.800 9.000 ;
        RECT 97.200 9.000 105.800 9.600 ;
        RECT 97.200 8.800 98.000 9.000 ;
        RECT 89.000 7.600 91.600 8.400 ;
        RECT 85.800 6.800 88.400 7.400 ;
        RECT 87.600 2.200 88.400 6.800 ;
        RECT 90.800 2.200 91.600 7.600 ;
        RECT 92.200 6.800 96.400 7.600 ;
        RECT 94.000 2.200 94.800 5.000 ;
        RECT 95.600 2.200 96.400 5.000 ;
        RECT 97.200 2.200 98.000 5.000 ;
        RECT 98.800 2.200 99.600 8.400 ;
        RECT 102.000 7.600 104.600 8.400 ;
        RECT 105.200 8.200 105.800 9.000 ;
        RECT 106.800 9.400 107.600 9.600 ;
        RECT 106.800 9.000 112.200 9.400 ;
        RECT 106.800 8.800 113.000 9.000 ;
        RECT 111.600 8.200 113.000 8.800 ;
        RECT 105.200 7.600 111.000 8.200 ;
        RECT 114.000 8.000 115.600 8.800 ;
        RECT 114.000 7.600 114.600 8.000 ;
        RECT 102.000 2.200 102.800 7.000 ;
        RECT 105.200 2.200 106.000 7.000 ;
        RECT 110.400 6.800 114.600 7.600 ;
        RECT 116.400 7.400 117.200 13.000 ;
        RECT 125.000 12.400 125.800 12.600 ;
        RECT 127.600 12.400 128.400 12.600 ;
        RECT 125.000 11.800 130.000 12.400 ;
        RECT 129.200 11.600 130.000 11.800 ;
        RECT 115.200 6.800 117.200 7.400 ;
        RECT 122.800 11.000 128.400 11.200 ;
        RECT 122.800 10.800 128.600 11.000 ;
        RECT 122.800 10.600 132.600 10.800 ;
        RECT 106.800 2.200 107.600 5.000 ;
        RECT 108.400 2.200 109.200 5.000 ;
        RECT 111.600 2.200 112.400 6.800 ;
        RECT 115.200 6.200 115.800 6.800 ;
        RECT 114.800 5.600 115.800 6.200 ;
        RECT 114.800 2.200 115.600 5.600 ;
        RECT 122.800 2.200 123.600 10.600 ;
        RECT 127.800 10.200 132.600 10.600 ;
        RECT 126.000 9.000 131.400 9.600 ;
        RECT 126.000 8.800 126.800 9.000 ;
        RECT 130.600 8.800 131.400 9.000 ;
        RECT 132.000 9.000 132.600 10.200 ;
        RECT 134.000 10.400 134.600 13.600 ;
        RECT 135.600 12.800 136.400 13.000 ;
        RECT 135.600 12.200 139.400 12.800 ;
        RECT 138.600 12.000 139.400 12.200 ;
        RECT 137.000 11.400 137.800 11.600 ;
        RECT 140.400 11.400 141.200 14.800 ;
        RECT 143.600 17.800 144.400 19.800 ;
        RECT 143.600 14.400 144.200 17.800 ;
        RECT 145.200 15.600 146.000 17.200 ;
        RECT 146.800 15.800 147.600 19.800 ;
        RECT 151.200 16.200 152.800 19.800 ;
        RECT 146.800 15.200 149.000 15.800 ;
        RECT 150.000 15.400 151.600 15.600 ;
        RECT 148.200 15.000 149.000 15.200 ;
        RECT 149.600 14.800 151.600 15.400 ;
        RECT 149.600 14.400 150.200 14.800 ;
        RECT 143.600 14.300 144.400 14.400 ;
        RECT 146.800 14.300 150.200 14.400 ;
        RECT 143.600 13.800 150.200 14.300 ;
        RECT 143.600 13.700 148.400 13.800 ;
        RECT 143.600 13.600 144.400 13.700 ;
        RECT 146.800 13.600 148.400 13.700 ;
        RECT 137.000 10.800 141.200 11.400 ;
        RECT 142.000 10.800 142.800 12.400 ;
        RECT 134.000 9.800 136.400 10.400 ;
        RECT 133.400 9.000 134.200 9.200 ;
        RECT 132.000 8.400 134.200 9.000 ;
        RECT 135.800 8.800 136.400 9.800 ;
        RECT 135.800 8.000 137.200 8.800 ;
        RECT 129.400 7.400 130.200 7.600 ;
        RECT 132.200 7.400 133.000 7.600 ;
        RECT 126.000 6.200 126.800 7.000 ;
        RECT 129.400 6.800 133.000 7.400 ;
        RECT 131.600 6.200 132.200 6.800 ;
        RECT 135.600 6.200 136.400 7.000 ;
        RECT 126.000 5.600 128.000 6.200 ;
        RECT 127.200 2.200 128.000 5.600 ;
        RECT 131.600 2.200 132.400 6.200 ;
        RECT 135.800 2.200 137.000 6.200 ;
        RECT 140.400 2.200 141.200 10.800 ;
        RECT 143.600 10.200 144.200 13.600 ;
        RECT 150.800 13.400 151.600 14.200 ;
        RECT 150.800 12.800 151.400 13.400 ;
        RECT 148.800 12.200 151.400 12.800 ;
        RECT 152.200 12.800 152.800 16.200 ;
        RECT 156.400 15.800 157.200 19.800 ;
        RECT 153.400 14.800 154.200 15.600 ;
        RECT 154.800 15.200 157.200 15.800 ;
        RECT 154.800 15.000 155.600 15.200 ;
        RECT 153.600 14.400 154.200 14.800 ;
        RECT 153.600 13.600 154.400 14.400 ;
        RECT 155.600 14.300 157.200 14.400 ;
        RECT 158.000 14.300 158.800 19.800 ;
        RECT 162.800 17.600 163.600 19.800 ;
        RECT 159.600 15.600 160.400 17.200 ;
        RECT 161.200 15.600 162.000 17.200 ;
        RECT 161.300 14.300 161.900 15.600 ;
        RECT 163.000 14.400 163.600 17.600 ;
        RECT 167.600 16.000 168.400 19.800 ;
        RECT 155.600 13.700 161.900 14.300 ;
        RECT 155.600 13.600 157.200 13.700 ;
        RECT 152.200 12.400 153.200 12.800 ;
        RECT 152.200 12.300 154.000 12.400 ;
        RECT 156.400 12.300 157.200 12.400 ;
        RECT 152.200 12.200 157.200 12.300 ;
        RECT 148.800 12.000 149.600 12.200 ;
        RECT 152.600 11.700 157.200 12.200 ;
        RECT 152.600 11.600 154.000 11.700 ;
        RECT 156.400 11.600 157.200 11.700 ;
        RECT 151.000 11.400 151.800 11.600 ;
        RECT 148.400 10.800 151.800 11.400 ;
        RECT 148.400 10.200 149.000 10.800 ;
        RECT 152.600 10.200 153.200 11.600 ;
        RECT 142.600 9.400 144.400 10.200 ;
        RECT 146.800 9.600 149.000 10.200 ;
        RECT 142.600 2.200 143.400 9.400 ;
        RECT 146.800 2.200 147.600 9.600 ;
        RECT 148.200 9.400 149.000 9.600 ;
        RECT 151.200 9.600 153.200 10.200 ;
        RECT 154.800 9.600 157.200 10.200 ;
        RECT 151.200 2.200 152.800 9.600 ;
        RECT 154.800 9.400 155.600 9.600 ;
        RECT 156.400 2.200 157.200 9.600 ;
        RECT 158.000 2.200 158.800 13.700 ;
        RECT 162.800 13.600 163.600 14.400 ;
        RECT 163.000 10.200 163.600 13.600 ;
        RECT 167.400 15.200 168.400 16.000 ;
        RECT 164.400 10.800 165.200 12.400 ;
        RECT 167.400 10.800 168.200 15.200 ;
        RECT 169.200 14.600 170.000 19.800 ;
        RECT 175.600 16.600 176.400 19.800 ;
        RECT 177.200 17.000 178.000 19.800 ;
        RECT 178.800 17.000 179.600 19.800 ;
        RECT 180.400 17.000 181.200 19.800 ;
        RECT 182.000 17.000 182.800 19.800 ;
        RECT 185.200 17.000 186.000 19.800 ;
        RECT 188.400 17.000 189.200 19.800 ;
        RECT 190.000 17.000 190.800 19.800 ;
        RECT 191.600 17.000 192.400 19.800 ;
        RECT 174.000 15.800 176.400 16.600 ;
        RECT 193.200 16.600 194.000 19.800 ;
        RECT 174.000 15.200 174.800 15.800 ;
        RECT 168.800 14.000 170.000 14.600 ;
        RECT 173.000 14.600 174.800 15.200 ;
        RECT 178.800 15.600 179.800 16.400 ;
        RECT 182.800 15.600 184.400 16.400 ;
        RECT 185.200 15.800 189.800 16.400 ;
        RECT 193.200 15.800 195.800 16.600 ;
        RECT 185.200 15.600 186.000 15.800 ;
        RECT 168.800 12.000 169.400 14.000 ;
        RECT 173.000 13.400 173.800 14.600 ;
        RECT 170.000 12.600 173.800 13.400 ;
        RECT 178.800 12.800 179.600 15.600 ;
        RECT 185.200 14.800 186.000 15.000 ;
        RECT 181.600 14.200 186.000 14.800 ;
        RECT 181.600 14.000 182.400 14.200 ;
        RECT 186.800 13.600 187.600 15.200 ;
        RECT 189.000 13.400 189.800 15.800 ;
        RECT 195.000 15.200 195.800 15.800 ;
        RECT 195.000 14.400 198.000 15.200 ;
        RECT 199.600 13.800 200.400 19.800 ;
        RECT 182.000 12.600 185.200 13.400 ;
        RECT 189.000 12.600 191.000 13.400 ;
        RECT 191.600 13.000 200.400 13.800 ;
        RECT 175.600 12.000 176.400 12.600 ;
        RECT 193.200 12.000 194.000 12.400 ;
        RECT 196.400 12.000 197.200 12.400 ;
        RECT 198.200 12.000 199.000 12.200 ;
        RECT 168.800 11.400 169.600 12.000 ;
        RECT 175.600 11.400 199.000 12.000 ;
        RECT 162.800 9.400 164.600 10.200 ;
        RECT 167.400 10.000 168.400 10.800 ;
        RECT 163.800 2.200 164.600 9.400 ;
        RECT 167.600 2.200 168.400 10.000 ;
        RECT 169.000 9.600 169.600 11.400 ;
        RECT 169.000 9.000 178.000 9.600 ;
        RECT 169.000 7.400 169.600 9.000 ;
        RECT 177.200 8.800 178.000 9.000 ;
        RECT 180.400 9.000 189.000 9.600 ;
        RECT 180.400 8.800 181.200 9.000 ;
        RECT 172.200 7.600 174.800 8.400 ;
        RECT 169.000 6.800 171.600 7.400 ;
        RECT 170.800 2.200 171.600 6.800 ;
        RECT 174.000 2.200 174.800 7.600 ;
        RECT 175.400 6.800 179.600 7.600 ;
        RECT 177.200 2.200 178.000 5.000 ;
        RECT 178.800 2.200 179.600 5.000 ;
        RECT 180.400 2.200 181.200 5.000 ;
        RECT 182.000 2.200 182.800 8.400 ;
        RECT 185.200 7.600 187.800 8.400 ;
        RECT 188.400 8.200 189.000 9.000 ;
        RECT 190.000 9.400 190.800 9.600 ;
        RECT 190.000 9.000 195.400 9.400 ;
        RECT 190.000 8.800 196.200 9.000 ;
        RECT 194.800 8.200 196.200 8.800 ;
        RECT 188.400 7.600 194.200 8.200 ;
        RECT 197.200 8.000 198.800 8.800 ;
        RECT 197.200 7.600 197.800 8.000 ;
        RECT 185.200 2.200 186.000 7.000 ;
        RECT 188.400 2.200 189.200 7.000 ;
        RECT 193.600 6.800 197.800 7.600 ;
        RECT 199.600 7.400 200.400 13.000 ;
        RECT 198.400 6.800 200.400 7.400 ;
        RECT 201.200 13.800 202.000 19.800 ;
        RECT 207.600 16.600 208.400 19.800 ;
        RECT 209.200 17.000 210.000 19.800 ;
        RECT 210.800 17.000 211.600 19.800 ;
        RECT 212.400 17.000 213.200 19.800 ;
        RECT 215.600 17.000 216.400 19.800 ;
        RECT 218.800 17.000 219.600 19.800 ;
        RECT 220.400 17.000 221.200 19.800 ;
        RECT 222.000 17.000 222.800 19.800 ;
        RECT 223.600 17.000 224.400 19.800 ;
        RECT 205.800 15.800 208.400 16.600 ;
        RECT 225.200 16.600 226.000 19.800 ;
        RECT 211.800 15.800 216.400 16.400 ;
        RECT 205.800 15.200 206.600 15.800 ;
        RECT 203.600 14.400 206.600 15.200 ;
        RECT 201.200 13.000 210.000 13.800 ;
        RECT 211.800 13.400 212.600 15.800 ;
        RECT 215.600 15.600 216.400 15.800 ;
        RECT 217.200 15.600 218.800 16.400 ;
        RECT 221.800 15.600 222.800 16.400 ;
        RECT 225.200 15.800 227.600 16.600 ;
        RECT 214.000 13.600 214.800 15.200 ;
        RECT 215.600 14.800 216.400 15.000 ;
        RECT 215.600 14.200 220.000 14.800 ;
        RECT 219.200 14.000 220.000 14.200 ;
        RECT 201.200 7.400 202.000 13.000 ;
        RECT 210.600 12.600 212.600 13.400 ;
        RECT 216.400 12.600 219.600 13.400 ;
        RECT 222.000 12.800 222.800 15.600 ;
        RECT 226.800 15.200 227.600 15.800 ;
        RECT 226.800 14.600 228.600 15.200 ;
        RECT 227.800 13.400 228.600 14.600 ;
        RECT 231.600 14.600 232.400 19.800 ;
        RECT 233.200 16.300 234.000 19.800 ;
        RECT 236.400 16.300 237.200 17.200 ;
        RECT 233.200 15.700 237.200 16.300 ;
        RECT 233.200 15.200 234.200 15.700 ;
        RECT 236.400 15.600 237.200 15.700 ;
        RECT 231.600 14.000 232.800 14.600 ;
        RECT 227.800 12.600 231.600 13.400 ;
        RECT 202.800 12.200 203.600 12.400 ;
        RECT 202.600 12.000 203.600 12.200 ;
        RECT 207.600 12.000 208.400 12.400 ;
        RECT 225.200 12.000 226.000 12.600 ;
        RECT 232.200 12.000 232.800 14.000 ;
        RECT 202.600 11.400 226.000 12.000 ;
        RECT 232.000 11.400 232.800 12.000 ;
        RECT 232.000 9.600 232.600 11.400 ;
        RECT 233.400 10.800 234.200 15.200 ;
        RECT 210.800 9.400 211.600 9.600 ;
        RECT 206.200 9.000 211.600 9.400 ;
        RECT 205.400 8.800 211.600 9.000 ;
        RECT 212.600 9.000 221.200 9.600 ;
        RECT 202.800 8.000 204.400 8.800 ;
        RECT 205.400 8.200 206.800 8.800 ;
        RECT 212.600 8.200 213.200 9.000 ;
        RECT 220.400 8.800 221.200 9.000 ;
        RECT 223.600 9.000 232.600 9.600 ;
        RECT 223.600 8.800 224.400 9.000 ;
        RECT 203.800 7.600 204.400 8.000 ;
        RECT 207.400 7.600 213.200 8.200 ;
        RECT 213.800 7.600 216.400 8.400 ;
        RECT 201.200 6.800 203.200 7.400 ;
        RECT 203.800 6.800 208.000 7.600 ;
        RECT 190.000 2.200 190.800 5.000 ;
        RECT 191.600 2.200 192.400 5.000 ;
        RECT 194.800 2.200 195.600 6.800 ;
        RECT 198.400 6.200 199.000 6.800 ;
        RECT 198.000 5.600 199.000 6.200 ;
        RECT 202.600 6.200 203.200 6.800 ;
        RECT 202.600 5.600 203.600 6.200 ;
        RECT 198.000 2.200 198.800 5.600 ;
        RECT 202.800 2.200 203.600 5.600 ;
        RECT 206.000 2.200 206.800 6.800 ;
        RECT 209.200 2.200 210.000 5.000 ;
        RECT 210.800 2.200 211.600 5.000 ;
        RECT 212.400 2.200 213.200 7.000 ;
        RECT 215.600 2.200 216.400 7.000 ;
        RECT 218.800 2.200 219.600 8.400 ;
        RECT 226.800 7.600 229.400 8.400 ;
        RECT 222.000 6.800 226.200 7.600 ;
        RECT 220.400 2.200 221.200 5.000 ;
        RECT 222.000 2.200 222.800 5.000 ;
        RECT 223.600 2.200 224.400 5.000 ;
        RECT 226.800 2.200 227.600 7.600 ;
        RECT 232.000 7.400 232.600 9.000 ;
        RECT 230.000 6.800 232.600 7.400 ;
        RECT 233.200 10.000 234.200 10.800 ;
        RECT 230.000 2.200 230.800 6.800 ;
        RECT 233.200 2.200 234.000 10.000 ;
        RECT 238.000 2.200 238.800 19.800 ;
        RECT 239.600 15.200 240.400 19.800 ;
        RECT 244.400 15.600 245.200 19.800 ;
        RECT 246.000 16.000 246.800 19.800 ;
        RECT 249.200 16.000 250.000 19.800 ;
        RECT 253.400 16.400 254.200 19.800 ;
        RECT 246.000 15.800 250.000 16.000 ;
        RECT 252.400 15.800 254.200 16.400 ;
        RECT 239.600 14.600 241.800 15.200 ;
        RECT 239.600 11.600 240.400 13.200 ;
        RECT 241.200 11.600 241.800 14.600 ;
        RECT 244.600 14.400 245.200 15.600 ;
        RECT 246.200 15.400 249.800 15.800 ;
        RECT 248.400 14.400 249.200 14.800 ;
        RECT 244.400 13.600 247.000 14.400 ;
        RECT 248.400 14.300 250.000 14.400 ;
        RECT 250.800 14.300 251.600 15.200 ;
        RECT 248.400 13.800 251.600 14.300 ;
        RECT 249.200 13.700 251.600 13.800 ;
        RECT 249.200 13.600 250.000 13.700 ;
        RECT 250.800 13.600 251.600 13.700 ;
        RECT 241.200 10.800 242.400 11.600 ;
        RECT 241.200 10.200 241.800 10.800 ;
        RECT 239.600 9.600 241.800 10.200 ;
        RECT 244.400 10.200 245.200 10.400 ;
        RECT 246.400 10.200 247.000 13.600 ;
        RECT 247.600 11.600 248.400 13.200 ;
        RECT 250.800 10.300 251.600 10.400 ;
        RECT 252.400 10.300 253.200 15.800 ;
        RECT 258.800 15.200 259.600 19.800 ;
        RECT 262.000 18.300 262.800 19.800 ;
        RECT 266.800 18.300 267.600 18.400 ;
        RECT 262.000 17.700 267.600 18.300 ;
        RECT 260.400 15.600 261.200 17.200 ;
        RECT 257.400 14.600 259.600 15.200 ;
        RECT 257.400 11.600 258.000 14.600 ;
        RECT 258.800 12.300 259.600 13.200 ;
        RECT 260.400 12.300 261.200 12.400 ;
        RECT 258.800 11.700 261.200 12.300 ;
        RECT 258.800 11.600 259.600 11.700 ;
        RECT 260.400 11.600 261.200 11.700 ;
        RECT 256.800 10.800 258.000 11.600 ;
        RECT 244.400 9.600 245.800 10.200 ;
        RECT 246.400 9.600 247.400 10.200 ;
        RECT 250.800 9.700 253.200 10.300 ;
        RECT 250.800 9.600 251.600 9.700 ;
        RECT 239.600 2.200 240.400 9.600 ;
        RECT 245.200 8.400 245.800 9.600 ;
        RECT 245.200 7.600 246.000 8.400 ;
        RECT 246.600 2.200 247.400 9.600 ;
        RECT 252.400 2.200 253.200 9.700 ;
        RECT 254.000 8.800 254.800 10.400 ;
        RECT 257.400 10.200 258.000 10.800 ;
        RECT 257.400 9.600 259.600 10.200 ;
        RECT 258.800 2.200 259.600 9.600 ;
        RECT 262.000 2.200 262.800 17.700 ;
        RECT 266.800 17.600 267.600 17.700 ;
        RECT 271.600 15.200 272.400 19.800 ;
        RECT 273.200 15.600 274.000 17.200 ;
        RECT 270.200 14.600 272.400 15.200 ;
        RECT 270.200 11.600 270.800 14.600 ;
        RECT 271.600 12.300 272.400 13.200 ;
        RECT 273.200 12.300 274.000 12.400 ;
        RECT 271.600 11.700 274.000 12.300 ;
        RECT 271.600 11.600 272.400 11.700 ;
        RECT 273.200 11.600 274.000 11.700 ;
        RECT 274.800 12.300 275.600 19.800 ;
        RECT 276.400 16.000 277.200 19.800 ;
        RECT 279.600 16.000 280.400 19.800 ;
        RECT 276.400 15.800 280.400 16.000 ;
        RECT 281.200 16.300 282.000 19.800 ;
        RECT 282.800 16.300 283.600 16.400 ;
        RECT 276.600 15.400 280.200 15.800 ;
        RECT 281.200 15.700 283.600 16.300 ;
        RECT 284.400 16.000 285.200 19.800 ;
        RECT 277.200 14.400 278.000 14.800 ;
        RECT 281.200 14.400 281.800 15.700 ;
        RECT 282.800 15.600 283.600 15.700 ;
        RECT 284.200 15.200 285.200 16.000 ;
        RECT 276.400 13.800 278.000 14.400 ;
        RECT 276.400 13.600 277.200 13.800 ;
        RECT 279.400 13.600 282.000 14.400 ;
        RECT 282.800 14.300 283.600 14.400 ;
        RECT 284.200 14.300 285.000 15.200 ;
        RECT 286.000 14.600 286.800 19.800 ;
        RECT 292.400 16.600 293.200 19.800 ;
        RECT 294.000 17.000 294.800 19.800 ;
        RECT 295.600 17.000 296.400 19.800 ;
        RECT 297.200 17.000 298.000 19.800 ;
        RECT 298.800 17.000 299.600 19.800 ;
        RECT 302.000 17.000 302.800 19.800 ;
        RECT 305.200 17.000 306.000 19.800 ;
        RECT 306.800 17.000 307.600 19.800 ;
        RECT 308.400 17.000 309.200 19.800 ;
        RECT 290.800 15.800 293.200 16.600 ;
        RECT 310.000 16.600 310.800 19.800 ;
        RECT 290.800 15.200 291.600 15.800 ;
        RECT 282.800 13.700 285.000 14.300 ;
        RECT 282.800 13.600 283.600 13.700 ;
        RECT 278.000 12.300 278.800 13.200 ;
        RECT 274.800 11.700 278.800 12.300 ;
        RECT 269.600 10.800 270.800 11.600 ;
        RECT 270.200 10.200 270.800 10.800 ;
        RECT 270.200 9.600 272.400 10.200 ;
        RECT 271.600 2.200 272.400 9.600 ;
        RECT 274.800 2.200 275.600 11.700 ;
        RECT 278.000 11.600 278.800 11.700 ;
        RECT 279.400 10.200 280.000 13.600 ;
        RECT 284.200 10.800 285.000 13.700 ;
        RECT 285.600 14.000 286.800 14.600 ;
        RECT 289.800 14.600 291.600 15.200 ;
        RECT 295.600 15.600 296.600 16.400 ;
        RECT 299.600 15.600 301.200 16.400 ;
        RECT 302.000 15.800 306.600 16.400 ;
        RECT 310.000 15.800 312.600 16.600 ;
        RECT 302.000 15.600 302.800 15.800 ;
        RECT 285.600 12.000 286.200 14.000 ;
        RECT 289.800 13.400 290.600 14.600 ;
        RECT 286.800 12.600 290.600 13.400 ;
        RECT 295.600 12.800 296.400 15.600 ;
        RECT 302.000 14.800 302.800 15.000 ;
        RECT 298.400 14.200 302.800 14.800 ;
        RECT 298.400 14.000 299.200 14.200 ;
        RECT 303.600 13.600 304.400 15.200 ;
        RECT 305.800 13.400 306.600 15.800 ;
        RECT 311.800 15.200 312.600 15.800 ;
        RECT 311.800 14.400 314.800 15.200 ;
        RECT 316.400 13.800 317.200 19.800 ;
        RECT 321.200 15.200 322.000 19.800 ;
        RECT 298.800 12.600 302.000 13.400 ;
        RECT 305.800 12.600 307.800 13.400 ;
        RECT 308.400 13.000 317.200 13.800 ;
        RECT 292.400 12.000 293.200 12.600 ;
        RECT 310.000 12.000 310.800 12.400 ;
        RECT 313.200 12.000 314.000 12.400 ;
        RECT 315.000 12.000 315.800 12.200 ;
        RECT 285.600 11.400 286.400 12.000 ;
        RECT 292.400 11.400 315.800 12.000 ;
        RECT 281.200 10.200 282.000 10.400 ;
        RECT 279.000 9.600 280.000 10.200 ;
        RECT 280.600 9.600 282.000 10.200 ;
        RECT 284.200 10.000 285.200 10.800 ;
        RECT 279.000 2.200 279.800 9.600 ;
        RECT 280.600 8.400 281.200 9.600 ;
        RECT 280.400 7.600 281.200 8.400 ;
        RECT 284.400 2.200 285.200 10.000 ;
        RECT 285.800 9.600 286.400 11.400 ;
        RECT 285.800 9.000 294.800 9.600 ;
        RECT 285.800 7.400 286.400 9.000 ;
        RECT 294.000 8.800 294.800 9.000 ;
        RECT 297.200 9.000 305.800 9.600 ;
        RECT 297.200 8.800 298.000 9.000 ;
        RECT 289.000 7.600 291.600 8.400 ;
        RECT 285.800 6.800 288.400 7.400 ;
        RECT 287.600 2.200 288.400 6.800 ;
        RECT 290.800 2.200 291.600 7.600 ;
        RECT 292.200 6.800 296.400 7.600 ;
        RECT 294.000 2.200 294.800 5.000 ;
        RECT 295.600 2.200 296.400 5.000 ;
        RECT 297.200 2.200 298.000 5.000 ;
        RECT 298.800 2.200 299.600 8.400 ;
        RECT 302.000 7.600 304.600 8.400 ;
        RECT 305.200 8.200 305.800 9.000 ;
        RECT 306.800 9.400 307.600 9.600 ;
        RECT 306.800 9.000 312.200 9.400 ;
        RECT 306.800 8.800 313.000 9.000 ;
        RECT 311.600 8.200 313.000 8.800 ;
        RECT 305.200 7.600 311.000 8.200 ;
        RECT 314.000 8.000 315.600 8.800 ;
        RECT 314.000 7.600 314.600 8.000 ;
        RECT 302.000 2.200 302.800 7.000 ;
        RECT 305.200 2.200 306.000 7.000 ;
        RECT 310.400 6.800 314.600 7.600 ;
        RECT 316.400 7.400 317.200 13.000 ;
        RECT 319.800 14.600 322.000 15.200 ;
        RECT 324.400 15.200 325.200 19.800 ;
        RECT 327.600 15.200 328.400 19.800 ;
        RECT 334.000 15.200 334.800 19.800 ;
        RECT 337.200 16.000 338.000 19.800 ;
        RECT 319.800 11.600 320.400 14.600 ;
        RECT 324.400 14.400 328.400 15.200 ;
        RECT 332.600 14.600 334.800 15.200 ;
        RECT 337.000 15.200 338.000 16.000 ;
        RECT 321.200 11.600 322.000 13.200 ;
        RECT 324.400 11.600 325.200 14.400 ;
        RECT 332.600 11.600 333.200 14.600 ;
        RECT 334.000 12.300 334.800 13.200 ;
        RECT 337.000 12.300 337.800 15.200 ;
        RECT 338.800 14.600 339.600 19.800 ;
        RECT 345.200 16.600 346.000 19.800 ;
        RECT 346.800 17.000 347.600 19.800 ;
        RECT 348.400 17.000 349.200 19.800 ;
        RECT 350.000 17.000 350.800 19.800 ;
        RECT 351.600 17.000 352.400 19.800 ;
        RECT 354.800 17.000 355.600 19.800 ;
        RECT 358.000 17.000 358.800 19.800 ;
        RECT 359.600 17.000 360.400 19.800 ;
        RECT 361.200 17.000 362.000 19.800 ;
        RECT 343.600 15.800 346.000 16.600 ;
        RECT 362.800 16.600 363.600 19.800 ;
        RECT 343.600 15.200 344.400 15.800 ;
        RECT 334.000 11.700 337.800 12.300 ;
        RECT 334.000 11.600 334.800 11.700 ;
        RECT 319.200 10.800 320.400 11.600 ;
        RECT 319.800 10.200 320.400 10.800 ;
        RECT 324.400 10.800 328.400 11.600 ;
        RECT 332.000 10.800 333.200 11.600 ;
        RECT 319.800 9.600 322.000 10.200 ;
        RECT 315.200 6.800 317.200 7.400 ;
        RECT 306.800 2.200 307.600 5.000 ;
        RECT 308.400 2.200 309.200 5.000 ;
        RECT 311.600 2.200 312.400 6.800 ;
        RECT 315.200 6.200 315.800 6.800 ;
        RECT 314.800 5.600 315.800 6.200 ;
        RECT 314.800 2.200 315.600 5.600 ;
        RECT 321.200 2.200 322.000 9.600 ;
        RECT 324.400 2.200 325.200 10.800 ;
        RECT 327.600 2.200 328.400 10.800 ;
        RECT 332.600 10.200 333.200 10.800 ;
        RECT 337.000 10.800 337.800 11.700 ;
        RECT 338.400 14.000 339.600 14.600 ;
        RECT 342.600 14.600 344.400 15.200 ;
        RECT 348.400 15.600 349.400 16.400 ;
        RECT 352.400 15.600 354.000 16.400 ;
        RECT 354.800 15.800 359.400 16.400 ;
        RECT 362.800 15.800 365.400 16.600 ;
        RECT 354.800 15.600 355.600 15.800 ;
        RECT 338.400 12.000 339.000 14.000 ;
        RECT 342.600 13.400 343.400 14.600 ;
        RECT 339.600 12.600 343.400 13.400 ;
        RECT 348.400 12.800 349.200 15.600 ;
        RECT 354.800 14.800 355.600 15.000 ;
        RECT 351.200 14.200 355.600 14.800 ;
        RECT 351.200 14.000 352.000 14.200 ;
        RECT 356.400 13.600 357.200 15.200 ;
        RECT 358.600 13.400 359.400 15.800 ;
        RECT 364.600 15.200 365.400 15.800 ;
        RECT 364.600 14.400 367.600 15.200 ;
        RECT 369.200 13.800 370.000 19.800 ;
        RECT 370.800 15.200 371.600 19.800 ;
        RECT 375.600 15.200 376.400 19.800 ;
        RECT 370.800 14.600 373.000 15.200 ;
        RECT 375.600 14.600 377.800 15.200 ;
        RECT 351.600 12.600 354.800 13.400 ;
        RECT 358.600 12.600 360.600 13.400 ;
        RECT 361.200 13.000 370.000 13.800 ;
        RECT 345.200 12.000 346.000 12.600 ;
        RECT 362.800 12.000 363.600 12.400 ;
        RECT 366.000 12.000 366.800 12.400 ;
        RECT 367.800 12.000 368.600 12.200 ;
        RECT 338.400 11.400 339.200 12.000 ;
        RECT 345.200 11.400 368.600 12.000 ;
        RECT 332.600 9.600 334.800 10.200 ;
        RECT 337.000 10.000 338.000 10.800 ;
        RECT 334.000 2.200 334.800 9.600 ;
        RECT 337.200 2.200 338.000 10.000 ;
        RECT 338.600 9.600 339.200 11.400 ;
        RECT 338.600 9.000 347.600 9.600 ;
        RECT 338.600 7.400 339.200 9.000 ;
        RECT 346.800 8.800 347.600 9.000 ;
        RECT 350.000 9.000 358.600 9.600 ;
        RECT 350.000 8.800 350.800 9.000 ;
        RECT 341.800 7.600 344.400 8.400 ;
        RECT 338.600 6.800 341.200 7.400 ;
        RECT 340.400 2.200 341.200 6.800 ;
        RECT 343.600 2.200 344.400 7.600 ;
        RECT 345.000 6.800 349.200 7.600 ;
        RECT 346.800 2.200 347.600 5.000 ;
        RECT 348.400 2.200 349.200 5.000 ;
        RECT 350.000 2.200 350.800 5.000 ;
        RECT 351.600 2.200 352.400 8.400 ;
        RECT 354.800 7.600 357.400 8.400 ;
        RECT 358.000 8.200 358.600 9.000 ;
        RECT 359.600 9.400 360.400 9.600 ;
        RECT 359.600 9.000 365.000 9.400 ;
        RECT 359.600 8.800 365.800 9.000 ;
        RECT 364.400 8.200 365.800 8.800 ;
        RECT 358.000 7.600 363.800 8.200 ;
        RECT 366.800 8.000 368.400 8.800 ;
        RECT 366.800 7.600 367.400 8.000 ;
        RECT 354.800 2.200 355.600 7.000 ;
        RECT 358.000 2.200 358.800 7.000 ;
        RECT 363.200 6.800 367.400 7.600 ;
        RECT 369.200 7.400 370.000 13.000 ;
        RECT 370.800 11.600 371.600 13.200 ;
        RECT 372.400 11.600 373.000 14.600 ;
        RECT 375.600 11.600 376.400 13.200 ;
        RECT 377.200 11.600 377.800 14.600 ;
        RECT 380.400 13.800 381.200 19.800 ;
        RECT 386.800 16.600 387.600 19.800 ;
        RECT 388.400 17.000 389.200 19.800 ;
        RECT 390.000 17.000 390.800 19.800 ;
        RECT 391.600 17.000 392.400 19.800 ;
        RECT 394.800 17.000 395.600 19.800 ;
        RECT 398.000 17.000 398.800 19.800 ;
        RECT 399.600 17.000 400.400 19.800 ;
        RECT 401.200 17.000 402.000 19.800 ;
        RECT 402.800 17.000 403.600 19.800 ;
        RECT 385.000 15.800 387.600 16.600 ;
        RECT 404.400 16.600 405.200 19.800 ;
        RECT 391.000 15.800 395.600 16.400 ;
        RECT 385.000 15.200 385.800 15.800 ;
        RECT 382.800 14.400 385.800 15.200 ;
        RECT 380.400 13.000 389.200 13.800 ;
        RECT 391.000 13.400 391.800 15.800 ;
        RECT 394.800 15.600 395.600 15.800 ;
        RECT 396.400 15.600 398.000 16.400 ;
        RECT 401.000 15.600 402.000 16.400 ;
        RECT 404.400 15.800 406.800 16.600 ;
        RECT 393.200 13.600 394.000 15.200 ;
        RECT 394.800 14.800 395.600 15.000 ;
        RECT 394.800 14.200 399.200 14.800 ;
        RECT 398.400 14.000 399.200 14.200 ;
        RECT 372.400 10.800 373.600 11.600 ;
        RECT 377.200 10.800 378.400 11.600 ;
        RECT 372.400 10.200 373.000 10.800 ;
        RECT 377.200 10.200 377.800 10.800 ;
        RECT 368.000 6.800 370.000 7.400 ;
        RECT 370.800 9.600 373.000 10.200 ;
        RECT 375.600 9.600 377.800 10.200 ;
        RECT 359.600 2.200 360.400 5.000 ;
        RECT 361.200 2.200 362.000 5.000 ;
        RECT 364.400 2.200 365.200 6.800 ;
        RECT 368.000 6.200 368.600 6.800 ;
        RECT 367.600 5.600 368.600 6.200 ;
        RECT 367.600 2.200 368.400 5.600 ;
        RECT 370.800 2.200 371.600 9.600 ;
        RECT 375.600 2.200 376.400 9.600 ;
        RECT 380.400 7.400 381.200 13.000 ;
        RECT 389.800 12.600 391.800 13.400 ;
        RECT 395.600 12.600 398.800 13.400 ;
        RECT 401.200 12.800 402.000 15.600 ;
        RECT 406.000 15.200 406.800 15.800 ;
        RECT 406.000 14.600 407.800 15.200 ;
        RECT 407.000 13.400 407.800 14.600 ;
        RECT 410.800 14.600 411.600 19.800 ;
        RECT 412.400 16.000 413.200 19.800 ;
        RECT 412.400 15.200 413.400 16.000 ;
        RECT 418.800 15.200 419.600 19.800 ;
        RECT 410.800 14.000 412.000 14.600 ;
        RECT 407.000 12.600 410.800 13.400 ;
        RECT 381.800 12.000 382.600 12.200 ;
        RECT 383.600 12.000 384.400 12.400 ;
        RECT 386.800 12.000 387.600 12.400 ;
        RECT 404.400 12.000 405.200 12.600 ;
        RECT 411.400 12.000 412.000 14.000 ;
        RECT 381.800 11.400 405.200 12.000 ;
        RECT 411.200 11.400 412.000 12.000 ;
        RECT 411.200 9.600 411.800 11.400 ;
        RECT 412.600 10.800 413.400 15.200 ;
        RECT 417.400 14.600 419.600 15.200 ;
        RECT 417.400 11.600 418.000 14.600 ;
        RECT 425.200 13.800 426.000 19.800 ;
        RECT 431.600 16.600 432.400 19.800 ;
        RECT 433.200 17.000 434.000 19.800 ;
        RECT 434.800 17.000 435.600 19.800 ;
        RECT 436.400 17.000 437.200 19.800 ;
        RECT 439.600 17.000 440.400 19.800 ;
        RECT 442.800 17.000 443.600 19.800 ;
        RECT 444.400 17.000 445.200 19.800 ;
        RECT 446.000 17.000 446.800 19.800 ;
        RECT 447.600 17.000 448.400 19.800 ;
        RECT 429.800 15.800 432.400 16.600 ;
        RECT 449.200 16.600 450.000 19.800 ;
        RECT 435.800 15.800 440.400 16.400 ;
        RECT 429.800 15.200 430.600 15.800 ;
        RECT 427.600 14.400 430.600 15.200 ;
        RECT 418.800 11.600 419.600 13.200 ;
        RECT 425.200 13.000 434.000 13.800 ;
        RECT 435.800 13.400 436.600 15.800 ;
        RECT 439.600 15.600 440.400 15.800 ;
        RECT 441.200 15.600 442.800 16.400 ;
        RECT 445.800 15.600 446.800 16.400 ;
        RECT 449.200 15.800 451.600 16.600 ;
        RECT 438.000 13.600 438.800 15.200 ;
        RECT 439.600 14.800 440.400 15.000 ;
        RECT 439.600 14.200 444.000 14.800 ;
        RECT 443.200 14.000 444.000 14.200 ;
        RECT 416.800 10.800 418.000 11.600 ;
        RECT 390.000 9.400 390.800 9.600 ;
        RECT 385.400 9.000 390.800 9.400 ;
        RECT 384.600 8.800 390.800 9.000 ;
        RECT 391.800 9.000 400.400 9.600 ;
        RECT 382.000 8.000 383.600 8.800 ;
        RECT 384.600 8.200 386.000 8.800 ;
        RECT 391.800 8.200 392.400 9.000 ;
        RECT 399.600 8.800 400.400 9.000 ;
        RECT 402.800 9.000 411.800 9.600 ;
        RECT 402.800 8.800 403.600 9.000 ;
        RECT 383.000 7.600 383.600 8.000 ;
        RECT 386.600 7.600 392.400 8.200 ;
        RECT 393.000 7.600 395.600 8.400 ;
        RECT 380.400 6.800 382.400 7.400 ;
        RECT 383.000 6.800 387.200 7.600 ;
        RECT 381.800 6.200 382.400 6.800 ;
        RECT 381.800 5.600 382.800 6.200 ;
        RECT 382.000 2.200 382.800 5.600 ;
        RECT 385.200 2.200 386.000 6.800 ;
        RECT 388.400 2.200 389.200 5.000 ;
        RECT 390.000 2.200 390.800 5.000 ;
        RECT 391.600 2.200 392.400 7.000 ;
        RECT 394.800 2.200 395.600 7.000 ;
        RECT 398.000 2.200 398.800 8.400 ;
        RECT 406.000 7.600 408.600 8.400 ;
        RECT 401.200 6.800 405.400 7.600 ;
        RECT 399.600 2.200 400.400 5.000 ;
        RECT 401.200 2.200 402.000 5.000 ;
        RECT 402.800 2.200 403.600 5.000 ;
        RECT 406.000 2.200 406.800 7.600 ;
        RECT 411.200 7.400 411.800 9.000 ;
        RECT 409.200 6.800 411.800 7.400 ;
        RECT 412.400 10.000 413.400 10.800 ;
        RECT 417.400 10.200 418.000 10.800 ;
        RECT 409.200 2.200 410.000 6.800 ;
        RECT 412.400 2.200 413.200 10.000 ;
        RECT 417.400 9.600 419.600 10.200 ;
        RECT 418.800 2.200 419.600 9.600 ;
        RECT 425.200 7.400 426.000 13.000 ;
        RECT 434.600 12.600 436.600 13.400 ;
        RECT 440.400 12.600 443.600 13.400 ;
        RECT 446.000 12.800 446.800 15.600 ;
        RECT 450.800 15.200 451.600 15.800 ;
        RECT 450.800 14.600 452.600 15.200 ;
        RECT 451.800 13.400 452.600 14.600 ;
        RECT 455.600 14.600 456.400 19.800 ;
        RECT 457.200 16.300 458.000 19.800 ;
        RECT 458.800 16.300 459.600 16.400 ;
        RECT 457.200 15.700 459.600 16.300 ;
        RECT 457.200 15.200 458.200 15.700 ;
        RECT 458.800 15.600 459.600 15.700 ;
        RECT 455.600 14.000 456.800 14.600 ;
        RECT 451.800 12.600 455.600 13.400 ;
        RECT 426.600 12.000 427.400 12.200 ;
        RECT 428.400 12.000 429.200 12.400 ;
        RECT 431.600 12.000 432.400 12.400 ;
        RECT 449.200 12.000 450.000 12.600 ;
        RECT 456.200 12.000 456.800 14.000 ;
        RECT 426.600 11.400 450.000 12.000 ;
        RECT 456.000 11.400 456.800 12.000 ;
        RECT 456.000 9.600 456.600 11.400 ;
        RECT 457.400 10.800 458.200 15.200 ;
        RECT 458.800 14.300 459.600 14.400 ;
        RECT 460.400 14.300 461.200 19.800 ;
        RECT 462.000 15.600 462.800 17.200 ;
        RECT 458.800 13.700 461.200 14.300 ;
        RECT 458.800 13.600 459.600 13.700 ;
        RECT 434.800 9.400 435.600 9.600 ;
        RECT 430.200 9.000 435.600 9.400 ;
        RECT 429.400 8.800 435.600 9.000 ;
        RECT 436.600 9.000 445.200 9.600 ;
        RECT 426.800 8.000 428.400 8.800 ;
        RECT 429.400 8.200 430.800 8.800 ;
        RECT 436.600 8.200 437.200 9.000 ;
        RECT 444.400 8.800 445.200 9.000 ;
        RECT 447.600 9.000 456.600 9.600 ;
        RECT 447.600 8.800 448.400 9.000 ;
        RECT 427.800 7.600 428.400 8.000 ;
        RECT 431.400 7.600 437.200 8.200 ;
        RECT 437.800 7.600 440.400 8.400 ;
        RECT 425.200 6.800 427.200 7.400 ;
        RECT 427.800 6.800 432.000 7.600 ;
        RECT 426.600 6.200 427.200 6.800 ;
        RECT 426.600 5.600 427.600 6.200 ;
        RECT 426.800 2.200 427.600 5.600 ;
        RECT 430.000 2.200 430.800 6.800 ;
        RECT 433.200 2.200 434.000 5.000 ;
        RECT 434.800 2.200 435.600 5.000 ;
        RECT 436.400 2.200 437.200 7.000 ;
        RECT 439.600 2.200 440.400 7.000 ;
        RECT 442.800 2.200 443.600 8.400 ;
        RECT 450.800 7.600 453.400 8.400 ;
        RECT 446.000 6.800 450.200 7.600 ;
        RECT 444.400 2.200 445.200 5.000 ;
        RECT 446.000 2.200 446.800 5.000 ;
        RECT 447.600 2.200 448.400 5.000 ;
        RECT 450.800 2.200 451.600 7.600 ;
        RECT 456.000 7.400 456.600 9.000 ;
        RECT 454.000 6.800 456.600 7.400 ;
        RECT 457.200 10.000 458.200 10.800 ;
        RECT 454.000 2.200 454.800 6.800 ;
        RECT 457.200 2.200 458.000 10.000 ;
        RECT 460.400 2.200 461.200 13.700 ;
        RECT 465.200 2.200 466.000 19.800 ;
        RECT 468.400 16.000 469.200 19.800 ;
        RECT 468.200 15.200 469.200 16.000 ;
        RECT 468.200 10.800 469.000 15.200 ;
        RECT 470.000 14.600 470.800 19.800 ;
        RECT 476.400 16.600 477.200 19.800 ;
        RECT 478.000 17.000 478.800 19.800 ;
        RECT 479.600 17.000 480.400 19.800 ;
        RECT 481.200 17.000 482.000 19.800 ;
        RECT 482.800 17.000 483.600 19.800 ;
        RECT 486.000 17.000 486.800 19.800 ;
        RECT 489.200 17.000 490.000 19.800 ;
        RECT 490.800 17.000 491.600 19.800 ;
        RECT 492.400 17.000 493.200 19.800 ;
        RECT 474.800 15.800 477.200 16.600 ;
        RECT 494.000 16.600 494.800 19.800 ;
        RECT 474.800 15.200 475.600 15.800 ;
        RECT 469.600 14.000 470.800 14.600 ;
        RECT 473.800 14.600 475.600 15.200 ;
        RECT 479.600 15.600 480.600 16.400 ;
        RECT 483.600 15.600 485.200 16.400 ;
        RECT 486.000 15.800 490.600 16.400 ;
        RECT 494.000 15.800 496.600 16.600 ;
        RECT 486.000 15.600 486.800 15.800 ;
        RECT 469.600 12.000 470.200 14.000 ;
        RECT 473.800 13.400 474.600 14.600 ;
        RECT 470.800 12.600 474.600 13.400 ;
        RECT 479.600 12.800 480.400 15.600 ;
        RECT 486.000 14.800 486.800 15.000 ;
        RECT 482.400 14.200 486.800 14.800 ;
        RECT 482.400 14.000 483.200 14.200 ;
        RECT 487.600 13.600 488.400 15.200 ;
        RECT 489.800 13.400 490.600 15.800 ;
        RECT 495.800 15.200 496.600 15.800 ;
        RECT 495.800 14.400 498.800 15.200 ;
        RECT 500.400 13.800 501.200 19.800 ;
        RECT 482.800 12.600 486.000 13.400 ;
        RECT 489.800 12.600 491.800 13.400 ;
        RECT 492.400 13.000 501.200 13.800 ;
        RECT 476.400 12.000 477.200 12.600 ;
        RECT 494.000 12.000 494.800 12.400 ;
        RECT 498.800 12.200 499.600 12.400 ;
        RECT 498.800 12.000 499.800 12.200 ;
        RECT 469.600 11.400 470.400 12.000 ;
        RECT 476.400 11.400 499.800 12.000 ;
        RECT 468.200 10.000 469.200 10.800 ;
        RECT 468.400 2.200 469.200 10.000 ;
        RECT 469.800 9.600 470.400 11.400 ;
        RECT 469.800 9.000 478.800 9.600 ;
        RECT 469.800 7.400 470.400 9.000 ;
        RECT 478.000 8.800 478.800 9.000 ;
        RECT 481.200 9.000 489.800 9.600 ;
        RECT 481.200 8.800 482.000 9.000 ;
        RECT 473.000 7.600 475.600 8.400 ;
        RECT 469.800 6.800 472.400 7.400 ;
        RECT 471.600 2.200 472.400 6.800 ;
        RECT 474.800 2.200 475.600 7.600 ;
        RECT 476.200 6.800 480.400 7.600 ;
        RECT 478.000 2.200 478.800 5.000 ;
        RECT 479.600 2.200 480.400 5.000 ;
        RECT 481.200 2.200 482.000 5.000 ;
        RECT 482.800 2.200 483.600 8.400 ;
        RECT 486.000 7.600 488.600 8.400 ;
        RECT 489.200 8.200 489.800 9.000 ;
        RECT 490.800 9.400 491.600 9.600 ;
        RECT 490.800 9.000 496.200 9.400 ;
        RECT 490.800 8.800 497.000 9.000 ;
        RECT 495.600 8.200 497.000 8.800 ;
        RECT 489.200 7.600 495.000 8.200 ;
        RECT 498.000 8.000 499.600 8.800 ;
        RECT 498.000 7.600 498.600 8.000 ;
        RECT 486.000 2.200 486.800 7.000 ;
        RECT 489.200 2.200 490.000 7.000 ;
        RECT 494.400 6.800 498.600 7.600 ;
        RECT 500.400 7.400 501.200 13.000 ;
        RECT 499.200 6.800 501.200 7.400 ;
        RECT 490.800 2.200 491.600 5.000 ;
        RECT 492.400 2.200 493.200 5.000 ;
        RECT 495.600 2.200 496.400 6.800 ;
        RECT 499.200 6.200 499.800 6.800 ;
        RECT 498.800 5.600 499.800 6.200 ;
        RECT 498.800 2.200 499.600 5.600 ;
        RECT 503.600 2.200 504.400 19.800 ;
        RECT 505.200 13.800 506.000 19.800 ;
        RECT 511.600 16.600 512.400 19.800 ;
        RECT 513.200 17.000 514.000 19.800 ;
        RECT 514.800 17.000 515.600 19.800 ;
        RECT 516.400 17.000 517.200 19.800 ;
        RECT 519.600 17.000 520.400 19.800 ;
        RECT 522.800 17.000 523.600 19.800 ;
        RECT 524.400 17.000 525.200 19.800 ;
        RECT 526.000 17.000 526.800 19.800 ;
        RECT 527.600 17.000 528.400 19.800 ;
        RECT 509.800 15.800 512.400 16.600 ;
        RECT 529.200 16.600 530.000 19.800 ;
        RECT 515.800 15.800 520.400 16.400 ;
        RECT 509.800 15.200 510.600 15.800 ;
        RECT 507.600 14.400 510.600 15.200 ;
        RECT 505.200 13.000 514.000 13.800 ;
        RECT 515.800 13.400 516.600 15.800 ;
        RECT 519.600 15.600 520.400 15.800 ;
        RECT 521.200 15.600 522.800 16.400 ;
        RECT 525.800 15.600 526.800 16.400 ;
        RECT 529.200 15.800 531.600 16.600 ;
        RECT 518.000 13.600 518.800 15.200 ;
        RECT 519.600 14.800 520.400 15.000 ;
        RECT 519.600 14.200 524.000 14.800 ;
        RECT 523.200 14.000 524.000 14.200 ;
        RECT 505.200 7.400 506.000 13.000 ;
        RECT 514.600 12.600 516.600 13.400 ;
        RECT 520.400 12.600 523.600 13.400 ;
        RECT 526.000 12.800 526.800 15.600 ;
        RECT 530.800 15.200 531.600 15.800 ;
        RECT 530.800 14.600 532.600 15.200 ;
        RECT 531.800 13.400 532.600 14.600 ;
        RECT 535.600 14.600 536.400 19.800 ;
        RECT 537.200 16.300 538.000 19.800 ;
        RECT 538.800 16.300 539.600 16.400 ;
        RECT 537.200 15.700 539.600 16.300 ;
        RECT 537.200 15.200 538.200 15.700 ;
        RECT 538.800 15.600 539.600 15.700 ;
        RECT 535.600 14.000 536.800 14.600 ;
        RECT 531.800 12.600 535.600 13.400 ;
        RECT 506.600 12.000 507.400 12.200 ;
        RECT 508.400 12.000 509.200 12.400 ;
        RECT 511.600 12.000 512.400 12.400 ;
        RECT 529.200 12.000 530.000 12.600 ;
        RECT 536.200 12.000 536.800 14.000 ;
        RECT 506.600 11.400 530.000 12.000 ;
        RECT 536.000 11.400 536.800 12.000 ;
        RECT 536.000 9.600 536.600 11.400 ;
        RECT 537.400 10.800 538.200 15.200 ;
        RECT 514.800 9.400 515.600 9.600 ;
        RECT 510.200 9.000 515.600 9.400 ;
        RECT 509.400 8.800 515.600 9.000 ;
        RECT 516.600 9.000 525.200 9.600 ;
        RECT 506.800 8.000 508.400 8.800 ;
        RECT 509.400 8.200 510.800 8.800 ;
        RECT 516.600 8.200 517.200 9.000 ;
        RECT 524.400 8.800 525.200 9.000 ;
        RECT 527.600 9.000 536.600 9.600 ;
        RECT 527.600 8.800 528.400 9.000 ;
        RECT 507.800 7.600 508.400 8.000 ;
        RECT 511.400 7.600 517.200 8.200 ;
        RECT 517.800 7.600 520.400 8.400 ;
        RECT 505.200 6.800 507.200 7.400 ;
        RECT 507.800 6.800 512.000 7.600 ;
        RECT 506.600 6.200 507.200 6.800 ;
        RECT 506.600 5.600 507.600 6.200 ;
        RECT 506.800 2.200 507.600 5.600 ;
        RECT 510.000 2.200 510.800 6.800 ;
        RECT 513.200 2.200 514.000 5.000 ;
        RECT 514.800 2.200 515.600 5.000 ;
        RECT 516.400 2.200 517.200 7.000 ;
        RECT 519.600 2.200 520.400 7.000 ;
        RECT 522.800 2.200 523.600 8.400 ;
        RECT 530.800 7.600 533.400 8.400 ;
        RECT 526.000 6.800 530.200 7.600 ;
        RECT 524.400 2.200 525.200 5.000 ;
        RECT 526.000 2.200 526.800 5.000 ;
        RECT 527.600 2.200 528.400 5.000 ;
        RECT 530.800 2.200 531.600 7.600 ;
        RECT 536.000 7.400 536.600 9.000 ;
        RECT 534.000 6.800 536.600 7.400 ;
        RECT 537.200 10.000 538.200 10.800 ;
        RECT 534.000 2.200 534.800 6.800 ;
        RECT 537.200 2.200 538.000 10.000 ;
        RECT 540.400 2.200 541.200 19.800 ;
        RECT 543.600 13.800 544.400 19.800 ;
        RECT 550.000 16.600 550.800 19.800 ;
        RECT 551.600 17.000 552.400 19.800 ;
        RECT 553.200 17.000 554.000 19.800 ;
        RECT 554.800 17.000 555.600 19.800 ;
        RECT 558.000 17.000 558.800 19.800 ;
        RECT 561.200 17.000 562.000 19.800 ;
        RECT 562.800 17.000 563.600 19.800 ;
        RECT 564.400 17.000 565.200 19.800 ;
        RECT 566.000 17.000 566.800 19.800 ;
        RECT 548.200 15.800 550.800 16.600 ;
        RECT 567.600 16.600 568.400 19.800 ;
        RECT 554.200 15.800 558.800 16.400 ;
        RECT 548.200 15.200 549.000 15.800 ;
        RECT 546.000 14.400 549.000 15.200 ;
        RECT 543.600 13.000 552.400 13.800 ;
        RECT 554.200 13.400 555.000 15.800 ;
        RECT 558.000 15.600 558.800 15.800 ;
        RECT 559.600 15.600 561.200 16.400 ;
        RECT 564.200 15.600 565.200 16.400 ;
        RECT 567.600 15.800 570.000 16.600 ;
        RECT 556.400 13.600 557.200 15.200 ;
        RECT 558.000 14.800 558.800 15.000 ;
        RECT 558.000 14.200 562.400 14.800 ;
        RECT 561.600 14.000 562.400 14.200 ;
        RECT 543.600 7.400 544.400 13.000 ;
        RECT 553.000 12.600 555.000 13.400 ;
        RECT 558.800 12.600 562.000 13.400 ;
        RECT 564.400 12.800 565.200 15.600 ;
        RECT 569.200 15.200 570.000 15.800 ;
        RECT 569.200 14.600 571.000 15.200 ;
        RECT 570.200 13.400 571.000 14.600 ;
        RECT 574.000 14.600 574.800 19.800 ;
        RECT 575.600 16.000 576.400 19.800 ;
        RECT 575.600 15.200 576.600 16.000 ;
        RECT 574.000 14.000 575.200 14.600 ;
        RECT 570.200 12.600 574.000 13.400 ;
        RECT 545.000 12.000 545.800 12.200 ;
        RECT 546.800 12.000 547.600 12.400 ;
        RECT 550.000 12.000 550.800 12.400 ;
        RECT 567.600 12.000 568.400 12.600 ;
        RECT 574.600 12.000 575.200 14.000 ;
        RECT 545.000 11.400 568.400 12.000 ;
        RECT 574.400 11.400 575.200 12.000 ;
        RECT 575.800 12.300 576.600 15.200 ;
        RECT 583.600 15.200 584.400 19.800 ;
        RECT 588.400 15.400 589.200 19.800 ;
        RECT 592.600 18.400 593.800 19.800 ;
        RECT 592.600 17.800 594.000 18.400 ;
        RECT 597.200 17.800 598.000 19.800 ;
        RECT 601.600 18.400 602.400 19.800 ;
        RECT 601.600 17.800 603.600 18.400 ;
        RECT 593.200 17.000 594.000 17.800 ;
        RECT 597.400 17.200 598.000 17.800 ;
        RECT 597.400 16.600 600.200 17.200 ;
        RECT 599.400 16.400 600.200 16.600 ;
        RECT 601.200 16.400 602.000 17.200 ;
        RECT 602.800 17.000 603.600 17.800 ;
        RECT 591.400 15.400 592.200 15.600 ;
        RECT 583.600 14.600 585.800 15.200 ;
        RECT 583.600 12.300 584.400 13.200 ;
        RECT 575.800 11.700 584.400 12.300 ;
        RECT 574.400 9.600 575.000 11.400 ;
        RECT 575.800 10.800 576.600 11.700 ;
        RECT 583.600 11.600 584.400 11.700 ;
        RECT 585.200 11.600 585.800 14.600 ;
        RECT 588.400 14.800 592.200 15.400 ;
        RECT 553.200 9.400 554.000 9.600 ;
        RECT 548.600 9.000 554.000 9.400 ;
        RECT 547.800 8.800 554.000 9.000 ;
        RECT 555.000 9.000 563.600 9.600 ;
        RECT 545.200 8.000 546.800 8.800 ;
        RECT 547.800 8.200 549.200 8.800 ;
        RECT 555.000 8.200 555.600 9.000 ;
        RECT 562.800 8.800 563.600 9.000 ;
        RECT 566.000 9.000 575.000 9.600 ;
        RECT 566.000 8.800 566.800 9.000 ;
        RECT 546.200 7.600 546.800 8.000 ;
        RECT 549.800 7.600 555.600 8.200 ;
        RECT 556.200 7.600 558.800 8.400 ;
        RECT 543.600 6.800 545.600 7.400 ;
        RECT 546.200 6.800 550.400 7.600 ;
        RECT 545.000 6.200 545.600 6.800 ;
        RECT 545.000 5.600 546.000 6.200 ;
        RECT 545.200 2.200 546.000 5.600 ;
        RECT 548.400 2.200 549.200 6.800 ;
        RECT 551.600 2.200 552.400 5.000 ;
        RECT 553.200 2.200 554.000 5.000 ;
        RECT 554.800 2.200 555.600 7.000 ;
        RECT 558.000 2.200 558.800 7.000 ;
        RECT 561.200 2.200 562.000 8.400 ;
        RECT 569.200 7.600 571.800 8.400 ;
        RECT 564.400 6.800 568.600 7.600 ;
        RECT 562.800 2.200 563.600 5.000 ;
        RECT 564.400 2.200 565.200 5.000 ;
        RECT 566.000 2.200 566.800 5.000 ;
        RECT 569.200 2.200 570.000 7.600 ;
        RECT 574.400 7.400 575.000 9.000 ;
        RECT 572.400 6.800 575.000 7.400 ;
        RECT 575.600 10.000 576.600 10.800 ;
        RECT 585.200 10.800 586.400 11.600 ;
        RECT 588.400 11.400 589.200 14.800 ;
        RECT 595.400 14.200 596.200 14.400 ;
        RECT 601.200 14.200 601.800 16.400 ;
        RECT 606.000 15.000 606.800 19.800 ;
        RECT 607.600 16.000 608.400 19.800 ;
        RECT 610.800 16.000 611.600 19.800 ;
        RECT 607.600 15.800 611.600 16.000 ;
        RECT 612.400 15.800 613.200 19.800 ;
        RECT 614.000 15.800 614.800 19.800 ;
        RECT 615.600 16.000 616.400 19.800 ;
        RECT 618.800 16.000 619.600 19.800 ;
        RECT 615.600 15.800 619.600 16.000 ;
        RECT 620.400 16.000 621.200 19.800 ;
        RECT 623.600 16.000 624.400 19.800 ;
        RECT 620.400 15.800 624.400 16.000 ;
        RECT 625.200 15.800 626.000 19.800 ;
        RECT 626.800 15.800 627.600 19.800 ;
        RECT 628.400 16.000 629.200 19.800 ;
        RECT 631.600 16.000 632.400 19.800 ;
        RECT 628.400 15.800 632.400 16.000 ;
        RECT 607.800 15.400 611.400 15.800 ;
        RECT 608.400 14.400 609.200 14.800 ;
        RECT 612.400 14.400 613.000 15.800 ;
        RECT 614.200 14.400 614.800 15.800 ;
        RECT 615.800 15.400 619.400 15.800 ;
        RECT 620.600 15.400 624.200 15.800 ;
        RECT 618.000 14.400 618.800 14.800 ;
        RECT 621.200 14.400 622.000 14.800 ;
        RECT 625.200 14.400 625.800 15.800 ;
        RECT 627.000 14.400 627.600 15.800 ;
        RECT 628.600 15.400 632.200 15.800 ;
        RECT 630.800 14.400 631.600 14.800 ;
        RECT 604.400 14.200 606.000 14.400 ;
        RECT 595.000 13.600 606.000 14.200 ;
        RECT 607.600 13.800 609.200 14.400 ;
        RECT 607.600 13.600 608.400 13.800 ;
        RECT 610.600 13.600 613.200 14.400 ;
        RECT 614.000 13.600 616.600 14.400 ;
        RECT 618.000 14.300 619.600 14.400 ;
        RECT 620.400 14.300 622.000 14.400 ;
        RECT 618.000 13.800 622.000 14.300 ;
        RECT 618.800 13.700 621.200 13.800 ;
        RECT 618.800 13.600 619.600 13.700 ;
        RECT 620.400 13.600 621.200 13.700 ;
        RECT 623.400 13.600 626.000 14.400 ;
        RECT 626.800 13.600 629.400 14.400 ;
        RECT 630.800 13.800 632.400 14.400 ;
        RECT 631.600 13.600 632.400 13.800 ;
        RECT 593.200 12.800 594.000 13.000 ;
        RECT 590.200 12.200 594.000 12.800 ;
        RECT 590.200 12.000 591.000 12.200 ;
        RECT 591.800 11.400 592.600 11.600 ;
        RECT 588.400 10.800 592.600 11.400 ;
        RECT 585.200 10.200 585.800 10.800 ;
        RECT 572.400 2.200 573.200 6.800 ;
        RECT 575.600 2.200 576.400 10.000 ;
        RECT 583.600 9.600 585.800 10.200 ;
        RECT 583.600 2.200 584.400 9.600 ;
        RECT 588.400 2.200 589.200 10.800 ;
        RECT 595.000 10.400 595.600 13.600 ;
        RECT 602.200 13.400 603.000 13.600 ;
        RECT 601.200 12.400 602.000 12.600 ;
        RECT 603.800 12.400 604.600 12.600 ;
        RECT 599.600 11.800 604.600 12.400 ;
        RECT 599.600 11.600 600.400 11.800 ;
        RECT 609.200 11.600 610.000 13.200 ;
        RECT 601.200 11.000 606.800 11.200 ;
        RECT 601.000 10.800 606.800 11.000 ;
        RECT 593.200 9.800 595.600 10.400 ;
        RECT 597.000 10.600 606.800 10.800 ;
        RECT 597.000 10.200 601.800 10.600 ;
        RECT 593.200 8.800 593.800 9.800 ;
        RECT 592.400 8.000 593.800 8.800 ;
        RECT 595.400 9.000 596.200 9.200 ;
        RECT 597.000 9.000 597.600 10.200 ;
        RECT 595.400 8.400 597.600 9.000 ;
        RECT 598.200 9.000 603.600 9.600 ;
        RECT 598.200 8.800 599.000 9.000 ;
        RECT 602.800 8.800 603.600 9.000 ;
        RECT 596.600 7.400 597.400 7.600 ;
        RECT 599.400 7.400 600.200 7.600 ;
        RECT 593.200 6.200 594.000 7.000 ;
        RECT 596.600 6.800 600.200 7.400 ;
        RECT 597.400 6.200 598.000 6.800 ;
        RECT 602.800 6.200 603.600 7.000 ;
        RECT 592.600 2.200 593.800 6.200 ;
        RECT 597.200 2.200 598.000 6.200 ;
        RECT 601.600 5.600 603.600 6.200 ;
        RECT 601.600 2.200 602.400 5.600 ;
        RECT 606.000 2.200 606.800 10.600 ;
        RECT 610.600 10.400 611.200 13.600 ;
        RECT 616.000 12.300 616.600 13.600 ;
        RECT 612.500 11.700 616.600 12.300 ;
        RECT 612.500 10.400 613.100 11.700 ;
        RECT 609.200 9.600 611.200 10.400 ;
        RECT 612.400 10.200 613.200 10.400 ;
        RECT 611.800 9.600 613.200 10.200 ;
        RECT 614.000 10.200 614.800 10.400 ;
        RECT 616.000 10.200 616.600 11.700 ;
        RECT 617.200 12.300 618.000 13.200 ;
        RECT 620.400 12.300 621.200 12.400 ;
        RECT 622.000 12.300 622.800 13.200 ;
        RECT 617.200 11.700 622.800 12.300 ;
        RECT 617.200 11.600 618.000 11.700 ;
        RECT 620.400 11.600 621.200 11.700 ;
        RECT 622.000 11.600 622.800 11.700 ;
        RECT 623.400 12.300 624.000 13.600 ;
        RECT 623.400 11.700 627.500 12.300 ;
        RECT 623.400 10.200 624.000 11.700 ;
        RECT 626.900 10.400 627.500 11.700 ;
        RECT 628.800 10.400 629.400 13.600 ;
        RECT 630.000 11.600 630.800 13.200 ;
        RECT 625.200 10.200 626.000 10.400 ;
        RECT 614.000 9.600 615.400 10.200 ;
        RECT 616.000 9.600 617.000 10.200 ;
        RECT 610.200 2.200 611.000 9.600 ;
        RECT 611.800 8.400 612.400 9.600 ;
        RECT 611.600 7.600 612.400 8.400 ;
        RECT 614.800 8.400 615.400 9.600 ;
        RECT 614.800 7.600 615.600 8.400 ;
        RECT 616.200 2.200 617.000 9.600 ;
        RECT 623.000 9.600 624.000 10.200 ;
        RECT 624.600 9.600 626.000 10.200 ;
        RECT 626.800 10.200 627.600 10.400 ;
        RECT 626.800 9.600 628.200 10.200 ;
        RECT 628.800 9.600 630.800 10.400 ;
        RECT 623.000 2.200 623.800 9.600 ;
        RECT 624.600 8.400 625.200 9.600 ;
        RECT 624.400 7.600 625.200 8.400 ;
        RECT 627.600 8.400 628.200 9.600 ;
        RECT 627.600 7.600 628.400 8.400 ;
        RECT 629.000 2.200 629.800 9.600 ;
        RECT 633.200 2.200 634.000 19.800 ;
        RECT 634.800 15.600 635.600 17.200 ;
        RECT 636.400 15.800 637.200 19.800 ;
        RECT 638.000 16.000 638.800 19.800 ;
        RECT 641.200 16.000 642.000 19.800 ;
        RECT 638.000 15.800 642.000 16.000 ;
        RECT 636.600 14.400 637.200 15.800 ;
        RECT 638.200 15.400 641.800 15.800 ;
        RECT 642.800 15.400 643.600 19.800 ;
        RECT 647.000 18.400 648.200 19.800 ;
        RECT 647.000 17.800 648.400 18.400 ;
        RECT 651.600 17.800 652.400 19.800 ;
        RECT 656.000 18.400 656.800 19.800 ;
        RECT 656.000 17.800 658.000 18.400 ;
        RECT 647.600 17.000 648.400 17.800 ;
        RECT 651.800 17.200 652.400 17.800 ;
        RECT 651.800 16.600 654.600 17.200 ;
        RECT 653.800 16.400 654.600 16.600 ;
        RECT 655.600 16.400 656.400 17.200 ;
        RECT 657.200 17.000 658.000 17.800 ;
        RECT 645.800 15.400 646.600 15.600 ;
        RECT 642.800 14.800 646.600 15.400 ;
        RECT 640.400 14.400 641.200 14.800 ;
        RECT 636.400 13.600 639.000 14.400 ;
        RECT 640.400 13.800 642.000 14.400 ;
        RECT 641.200 13.600 642.000 13.800 ;
        RECT 636.400 10.200 637.200 10.400 ;
        RECT 638.400 10.200 639.000 13.600 ;
        RECT 639.600 11.600 640.400 13.200 ;
        RECT 642.800 11.400 643.600 14.800 ;
        RECT 649.200 14.200 650.600 14.400 ;
        RECT 655.600 14.200 656.200 16.400 ;
        RECT 660.400 15.000 661.200 19.800 ;
        RECT 662.000 15.400 662.800 19.800 ;
        RECT 666.200 18.400 667.400 19.800 ;
        RECT 666.200 17.800 667.600 18.400 ;
        RECT 670.800 17.800 671.600 19.800 ;
        RECT 675.200 18.400 676.000 19.800 ;
        RECT 675.200 17.800 677.200 18.400 ;
        RECT 666.800 17.000 667.600 17.800 ;
        RECT 671.000 17.200 671.600 17.800 ;
        RECT 671.000 16.600 673.800 17.200 ;
        RECT 673.000 16.400 673.800 16.600 ;
        RECT 674.800 16.400 675.600 17.200 ;
        RECT 676.400 17.000 677.200 17.800 ;
        RECT 665.000 15.400 665.800 15.600 ;
        RECT 662.000 14.800 665.800 15.400 ;
        RECT 658.800 14.200 660.400 14.400 ;
        RECT 649.200 13.600 660.400 14.200 ;
        RECT 647.600 12.800 648.400 13.000 ;
        RECT 644.600 12.200 648.400 12.800 ;
        RECT 644.600 12.000 645.400 12.200 ;
        RECT 646.200 11.400 647.000 11.600 ;
        RECT 642.800 10.800 647.000 11.400 ;
        RECT 636.400 9.600 637.800 10.200 ;
        RECT 638.400 9.600 639.400 10.200 ;
        RECT 637.200 8.400 637.800 9.600 ;
        RECT 637.200 7.600 638.000 8.400 ;
        RECT 638.600 2.200 639.400 9.600 ;
        RECT 642.800 2.200 643.600 10.800 ;
        RECT 649.400 10.400 650.000 13.600 ;
        RECT 656.600 13.400 657.400 13.600 ;
        RECT 658.200 12.400 659.000 12.600 ;
        RECT 654.000 11.800 659.000 12.400 ;
        RECT 654.000 11.600 654.800 11.800 ;
        RECT 662.000 11.400 662.800 14.800 ;
        RECT 669.000 14.200 669.800 14.400 ;
        RECT 674.800 14.200 675.400 16.400 ;
        RECT 679.600 15.000 680.400 19.800 ;
        RECT 681.200 15.800 682.000 19.800 ;
        RECT 682.800 16.000 683.600 19.800 ;
        RECT 686.000 16.000 686.800 19.800 ;
        RECT 682.800 15.800 686.800 16.000 ;
        RECT 681.400 14.400 682.000 15.800 ;
        RECT 683.000 15.400 686.600 15.800 ;
        RECT 685.200 14.400 686.000 14.800 ;
        RECT 678.000 14.200 679.600 14.400 ;
        RECT 668.600 13.600 679.600 14.200 ;
        RECT 681.200 13.600 683.800 14.400 ;
        RECT 685.200 14.300 686.800 14.400 ;
        RECT 687.600 14.300 688.400 14.400 ;
        RECT 685.200 13.800 688.400 14.300 ;
        RECT 686.000 13.700 688.400 13.800 ;
        RECT 686.000 13.600 686.800 13.700 ;
        RECT 687.600 13.600 688.400 13.700 ;
        RECT 666.800 12.800 667.600 13.000 ;
        RECT 663.800 12.200 667.600 12.800 ;
        RECT 668.600 12.300 669.200 13.600 ;
        RECT 675.800 13.400 676.600 13.600 ;
        RECT 677.400 12.400 678.200 12.600 ;
        RECT 670.000 12.300 670.800 12.400 ;
        RECT 663.800 12.000 664.600 12.200 ;
        RECT 668.500 11.700 670.800 12.300 ;
        RECT 665.400 11.400 666.200 11.600 ;
        RECT 655.600 11.000 661.200 11.200 ;
        RECT 655.400 10.800 661.200 11.000 ;
        RECT 647.600 9.800 650.000 10.400 ;
        RECT 651.400 10.600 661.200 10.800 ;
        RECT 651.400 10.200 656.200 10.600 ;
        RECT 647.600 8.800 648.200 9.800 ;
        RECT 646.800 8.000 648.200 8.800 ;
        RECT 649.800 9.000 650.600 9.200 ;
        RECT 651.400 9.000 652.000 10.200 ;
        RECT 649.800 8.400 652.000 9.000 ;
        RECT 652.600 9.000 658.000 9.600 ;
        RECT 652.600 8.800 653.400 9.000 ;
        RECT 657.200 8.800 658.000 9.000 ;
        RECT 651.000 7.400 651.800 7.600 ;
        RECT 653.800 7.400 654.600 7.600 ;
        RECT 647.600 6.200 648.400 7.000 ;
        RECT 651.000 6.800 654.600 7.400 ;
        RECT 651.800 6.200 652.400 6.800 ;
        RECT 657.200 6.200 658.000 7.000 ;
        RECT 647.000 2.200 648.200 6.200 ;
        RECT 651.600 2.200 652.400 6.200 ;
        RECT 656.000 5.600 658.000 6.200 ;
        RECT 656.000 2.200 656.800 5.600 ;
        RECT 660.400 2.200 661.200 10.600 ;
        RECT 662.000 10.800 666.200 11.400 ;
        RECT 662.000 2.200 662.800 10.800 ;
        RECT 668.600 10.400 669.200 11.700 ;
        RECT 670.000 11.600 670.800 11.700 ;
        RECT 673.200 11.800 678.200 12.400 ;
        RECT 673.200 11.600 674.000 11.800 ;
        RECT 674.800 11.000 680.400 11.200 ;
        RECT 674.600 10.800 680.400 11.000 ;
        RECT 666.800 9.800 669.200 10.400 ;
        RECT 670.600 10.600 680.400 10.800 ;
        RECT 670.600 10.200 675.400 10.600 ;
        RECT 666.800 8.800 667.400 9.800 ;
        RECT 666.000 8.000 667.400 8.800 ;
        RECT 669.000 9.000 669.800 9.200 ;
        RECT 670.600 9.000 671.200 10.200 ;
        RECT 669.000 8.400 671.200 9.000 ;
        RECT 671.800 9.000 677.200 9.600 ;
        RECT 671.800 8.800 672.600 9.000 ;
        RECT 676.400 8.800 677.200 9.000 ;
        RECT 670.200 7.400 671.000 7.600 ;
        RECT 673.000 7.400 673.800 7.600 ;
        RECT 666.800 6.200 667.600 7.000 ;
        RECT 670.200 6.800 673.800 7.400 ;
        RECT 671.000 6.200 671.600 6.800 ;
        RECT 676.400 6.200 677.200 7.000 ;
        RECT 666.200 2.200 667.400 6.200 ;
        RECT 670.800 2.200 671.600 6.200 ;
        RECT 675.200 5.600 677.200 6.200 ;
        RECT 675.200 2.200 676.000 5.600 ;
        RECT 679.600 2.200 680.400 10.600 ;
        RECT 681.200 10.200 682.000 10.400 ;
        RECT 683.200 10.200 683.800 13.600 ;
        RECT 684.400 11.600 685.200 13.200 ;
        RECT 681.200 9.600 682.600 10.200 ;
        RECT 683.200 9.600 684.200 10.200 ;
        RECT 682.000 8.400 682.600 9.600 ;
        RECT 682.000 7.600 682.800 8.400 ;
        RECT 683.400 2.200 684.200 9.600 ;
      LAYER via1 ;
        RECT 9.200 493.000 10.000 493.800 ;
        RECT 18.800 492.600 19.600 493.400 ;
        RECT 14.000 491.600 14.800 492.400 ;
        RECT 25.200 491.600 26.000 492.400 ;
        RECT 10.800 488.800 11.600 489.600 ;
        RECT 15.600 487.600 16.400 488.400 ;
        RECT 12.400 486.200 13.200 487.000 ;
        RECT 9.200 484.200 10.000 485.000 ;
        RECT 10.800 484.200 11.600 485.000 ;
        RECT 15.600 486.200 16.400 487.000 ;
        RECT 18.800 486.200 19.600 487.000 ;
        RECT 20.400 484.200 21.200 485.000 ;
        RECT 22.000 484.200 22.800 485.000 ;
        RECT 23.600 484.200 24.400 485.000 ;
        RECT 33.200 483.600 34.000 484.400 ;
        RECT 54.000 493.000 54.800 493.800 ;
        RECT 63.600 492.600 64.400 493.400 ;
        RECT 49.200 491.600 50.000 492.400 ;
        RECT 70.000 491.600 70.800 492.400 ;
        RECT 55.600 488.800 56.400 489.600 ;
        RECT 60.400 487.600 61.200 488.400 ;
        RECT 57.200 486.200 58.000 487.000 ;
        RECT 54.000 484.200 54.800 485.000 ;
        RECT 55.600 484.200 56.400 485.000 ;
        RECT 60.400 486.200 61.200 487.000 ;
        RECT 63.600 486.200 64.400 487.000 ;
        RECT 65.200 484.200 66.000 485.000 ;
        RECT 66.800 484.200 67.600 485.000 ;
        RECT 68.400 484.200 69.200 485.000 ;
        RECT 78.000 483.600 78.800 484.400 ;
        RECT 87.600 493.600 88.400 494.400 ;
        RECT 110.000 493.600 110.800 494.400 ;
        RECT 98.800 483.600 99.600 484.400 ;
        RECT 116.400 490.200 117.200 491.000 ;
        RECT 148.400 493.600 149.200 494.400 ;
        RECT 134.000 483.600 134.800 484.400 ;
        RECT 154.800 489.600 155.600 490.400 ;
        RECT 183.600 495.600 184.400 496.400 ;
        RECT 185.200 494.200 186.000 495.000 ;
        RECT 175.600 491.600 176.400 492.400 ;
        RECT 198.000 491.600 198.800 492.400 ;
        RECT 164.400 489.600 165.200 490.400 ;
        RECT 167.600 483.600 168.400 484.400 ;
        RECT 178.800 486.800 179.600 487.600 ;
        RECT 182.000 486.200 182.800 487.000 ;
        RECT 177.200 484.200 178.000 485.000 ;
        RECT 178.800 484.200 179.600 485.000 ;
        RECT 180.400 484.200 181.200 485.000 ;
        RECT 185.200 486.200 186.000 487.000 ;
        RECT 188.400 486.200 189.200 487.000 ;
        RECT 190.000 484.200 190.800 485.000 ;
        RECT 191.600 484.200 192.400 485.000 ;
        RECT 222.000 495.600 222.800 496.400 ;
        RECT 223.600 494.200 224.400 495.000 ;
        RECT 214.000 491.600 214.800 492.400 ;
        RECT 236.400 491.600 237.200 492.400 ;
        RECT 206.000 483.600 206.800 484.400 ;
        RECT 217.200 486.800 218.000 487.600 ;
        RECT 220.400 486.200 221.200 487.000 ;
        RECT 215.600 484.200 216.400 485.000 ;
        RECT 217.200 484.200 218.000 485.000 ;
        RECT 218.800 484.200 219.600 485.000 ;
        RECT 223.600 486.200 224.400 487.000 ;
        RECT 226.800 486.200 227.600 487.000 ;
        RECT 239.600 493.600 240.400 494.400 ;
        RECT 252.400 493.600 253.200 494.400 ;
        RECT 266.800 493.000 267.600 493.800 ;
        RECT 228.400 484.200 229.200 485.000 ;
        RECT 230.000 484.200 230.800 485.000 ;
        RECT 276.400 492.600 277.200 493.400 ;
        RECT 262.000 491.600 262.800 492.400 ;
        RECT 306.800 493.000 307.600 493.800 ;
        RECT 268.400 488.800 269.200 489.600 ;
        RECT 273.200 487.600 274.000 488.400 ;
        RECT 270.000 486.200 270.800 487.000 ;
        RECT 266.800 484.200 267.600 485.000 ;
        RECT 268.400 484.200 269.200 485.000 ;
        RECT 273.200 486.200 274.000 487.000 ;
        RECT 276.400 486.200 277.200 487.000 ;
        RECT 278.000 484.200 278.800 485.000 ;
        RECT 279.600 484.200 280.400 485.000 ;
        RECT 281.200 484.200 282.000 485.000 ;
        RECT 316.400 492.600 317.200 493.400 ;
        RECT 302.000 491.600 302.800 492.400 ;
        RECT 322.800 491.600 323.600 492.400 ;
        RECT 337.200 494.800 338.000 495.600 ;
        RECT 308.400 488.800 309.200 489.600 ;
        RECT 313.200 487.600 314.000 488.400 ;
        RECT 310.000 486.200 310.800 487.000 ;
        RECT 306.800 484.200 307.600 485.000 ;
        RECT 308.400 484.200 309.200 485.000 ;
        RECT 313.200 486.200 314.000 487.000 ;
        RECT 316.400 486.200 317.200 487.000 ;
        RECT 318.000 484.200 318.800 485.000 ;
        RECT 319.600 484.200 320.400 485.000 ;
        RECT 321.200 484.200 322.000 485.000 ;
        RECT 362.800 495.600 363.600 496.400 ;
        RECT 364.400 494.200 365.200 495.000 ;
        RECT 354.800 491.600 355.600 492.400 ;
        RECT 330.800 483.600 331.600 484.400 ;
        RECT 346.800 483.600 347.600 484.400 ;
        RECT 358.000 486.800 358.800 487.600 ;
        RECT 361.200 486.200 362.000 487.000 ;
        RECT 356.400 484.200 357.200 485.000 ;
        RECT 358.000 484.200 358.800 485.000 ;
        RECT 359.600 484.200 360.400 485.000 ;
        RECT 364.400 486.200 365.200 487.000 ;
        RECT 367.600 486.200 368.400 487.000 ;
        RECT 386.800 495.600 387.600 496.400 ;
        RECT 402.800 495.600 403.600 496.400 ;
        RECT 404.400 494.200 405.200 495.000 ;
        RECT 406.000 491.600 406.800 492.400 ;
        RECT 369.200 484.200 370.000 485.000 ;
        RECT 370.800 484.200 371.600 485.000 ;
        RECT 398.000 486.800 398.800 487.600 ;
        RECT 401.200 486.200 402.000 487.000 ;
        RECT 396.400 484.200 397.200 485.000 ;
        RECT 398.000 484.200 398.800 485.000 ;
        RECT 399.600 484.200 400.400 485.000 ;
        RECT 404.400 486.200 405.200 487.000 ;
        RECT 407.600 486.200 408.400 487.000 ;
        RECT 409.200 484.200 410.000 485.000 ;
        RECT 410.800 484.200 411.600 485.000 ;
        RECT 436.400 491.600 437.200 492.400 ;
        RECT 462.000 495.600 462.800 496.400 ;
        RECT 463.600 494.200 464.400 495.000 ;
        RECT 471.600 491.600 472.400 492.400 ;
        RECT 442.800 489.600 443.600 490.400 ;
        RECT 457.200 486.800 458.000 487.600 ;
        RECT 460.400 486.200 461.200 487.000 ;
        RECT 455.600 484.200 456.400 485.000 ;
        RECT 457.200 484.200 458.000 485.000 ;
        RECT 458.800 484.200 459.600 485.000 ;
        RECT 463.600 486.200 464.400 487.000 ;
        RECT 466.800 486.200 467.600 487.000 ;
        RECT 468.400 484.200 469.200 485.000 ;
        RECT 470.000 484.200 470.800 485.000 ;
        RECT 481.200 483.600 482.000 484.400 ;
        RECT 492.200 491.600 493.000 492.400 ;
        RECT 508.400 495.600 509.200 496.400 ;
        RECT 510.000 494.200 510.800 495.000 ;
        RECT 500.400 491.600 501.200 492.400 ;
        RECT 522.800 491.600 523.600 492.400 ;
        RECT 482.800 483.600 483.600 484.400 ;
        RECT 503.600 486.800 504.400 487.600 ;
        RECT 506.800 486.200 507.600 487.000 ;
        RECT 502.000 484.200 502.800 485.000 ;
        RECT 503.600 484.200 504.400 485.000 ;
        RECT 505.200 484.200 506.000 485.000 ;
        RECT 510.000 486.200 510.800 487.000 ;
        RECT 513.200 486.200 514.000 487.000 ;
        RECT 532.400 493.600 533.200 494.400 ;
        RECT 514.800 484.200 515.600 485.000 ;
        RECT 516.400 484.200 517.200 485.000 ;
        RECT 535.600 489.600 536.400 490.400 ;
        RECT 567.600 495.600 568.400 496.400 ;
        RECT 569.200 494.200 570.000 495.000 ;
        RECT 559.600 491.600 560.400 492.400 ;
        RECT 551.600 483.600 552.400 484.400 ;
        RECT 562.800 486.800 563.600 487.600 ;
        RECT 566.000 486.200 566.800 487.000 ;
        RECT 561.200 484.200 562.000 485.000 ;
        RECT 562.800 484.200 563.600 485.000 ;
        RECT 564.400 484.200 565.200 485.000 ;
        RECT 569.200 486.200 570.000 487.000 ;
        RECT 572.400 486.200 573.200 487.000 ;
        RECT 598.000 493.000 598.800 493.800 ;
        RECT 607.600 492.600 608.400 493.400 ;
        RECT 631.600 497.600 632.400 498.400 ;
        RECT 594.800 491.600 595.600 492.400 ;
        RECT 634.800 493.600 635.600 494.400 ;
        RECT 636.400 493.600 637.200 494.400 ;
        RECT 599.600 488.800 600.400 489.600 ;
        RECT 604.400 487.600 605.200 488.400 ;
        RECT 574.000 484.200 574.800 485.000 ;
        RECT 575.600 484.200 576.400 485.000 ;
        RECT 601.200 486.200 602.000 487.000 ;
        RECT 598.000 484.200 598.800 485.000 ;
        RECT 599.600 484.200 600.400 485.000 ;
        RECT 604.400 486.200 605.200 487.000 ;
        RECT 607.600 486.200 608.400 487.000 ;
        RECT 609.200 484.200 610.000 485.000 ;
        RECT 610.800 484.200 611.600 485.000 ;
        RECT 612.400 484.200 613.200 485.000 ;
        RECT 668.400 495.600 669.200 496.400 ;
        RECT 670.000 494.200 670.800 495.000 ;
        RECT 660.400 491.600 661.200 492.400 ;
        RECT 622.000 483.600 622.800 484.400 ;
        RECT 647.600 483.600 648.400 484.400 ;
        RECT 652.400 483.600 653.200 484.400 ;
        RECT 663.600 486.800 664.400 487.600 ;
        RECT 666.800 486.200 667.600 487.000 ;
        RECT 662.000 484.200 662.800 485.000 ;
        RECT 663.600 484.200 664.400 485.000 ;
        RECT 665.200 484.200 666.000 485.000 ;
        RECT 670.000 486.200 670.800 487.000 ;
        RECT 673.200 486.200 674.000 487.000 ;
        RECT 674.800 484.200 675.600 485.000 ;
        RECT 676.400 484.200 677.200 485.000 ;
        RECT 14.000 474.400 14.800 475.200 ;
        RECT 17.200 475.000 18.000 475.800 ;
        RECT 39.600 477.600 40.400 478.400 ;
        RECT 12.400 472.400 13.200 473.200 ;
        RECT 10.800 469.600 11.600 470.400 ;
        RECT 2.800 463.600 3.600 464.400 ;
        RECT 22.000 467.600 22.800 468.400 ;
        RECT 18.800 465.600 19.600 466.400 ;
        RECT 39.600 469.600 40.400 470.400 ;
        RECT 12.400 464.200 13.200 465.000 ;
        RECT 14.000 464.200 14.800 465.000 ;
        RECT 15.600 464.200 16.400 465.000 ;
        RECT 17.200 464.200 18.000 465.000 ;
        RECT 20.400 464.200 21.200 465.000 ;
        RECT 23.600 464.200 24.400 465.000 ;
        RECT 25.200 464.200 26.000 465.000 ;
        RECT 26.800 464.200 27.600 465.000 ;
        RECT 41.200 467.600 42.000 468.400 ;
        RECT 62.000 473.600 62.800 474.400 ;
        RECT 71.600 473.600 72.400 474.400 ;
        RECT 46.000 467.600 46.800 468.400 ;
        RECT 47.600 466.200 48.400 467.000 ;
        RECT 73.200 469.600 74.000 470.400 ;
        RECT 74.800 469.600 75.600 470.400 ;
        RECT 78.000 469.600 78.800 470.400 ;
        RECT 89.200 473.600 90.000 474.400 ;
        RECT 86.000 469.600 86.800 470.400 ;
        RECT 65.200 463.600 66.000 464.400 ;
        RECT 87.600 467.600 88.400 468.400 ;
        RECT 92.400 467.600 93.200 468.400 ;
        RECT 95.600 467.600 96.400 468.400 ;
        RECT 81.200 463.600 82.000 464.400 ;
        RECT 94.000 466.200 94.800 467.000 ;
        RECT 90.800 463.600 91.600 464.400 ;
        RECT 119.600 469.600 120.400 470.400 ;
        RECT 127.600 469.600 128.400 470.400 ;
        RECT 130.800 469.600 131.600 470.400 ;
        RECT 132.400 469.600 133.200 470.400 ;
        RECT 129.200 467.600 130.000 468.400 ;
        RECT 111.600 463.600 112.400 464.400 ;
        RECT 154.800 472.400 155.600 473.200 ;
        RECT 158.000 471.000 158.800 471.800 ;
        RECT 159.600 467.600 160.400 468.400 ;
        RECT 158.000 466.200 158.800 467.000 ;
        RECT 140.400 463.600 141.200 464.400 ;
        RECT 164.400 467.600 165.200 468.400 ;
        RECT 178.800 469.600 179.600 470.400 ;
        RECT 162.800 463.600 163.600 464.400 ;
        RECT 172.400 465.600 173.200 466.400 ;
        RECT 174.000 465.600 174.800 466.400 ;
        RECT 170.800 463.600 171.600 464.400 ;
        RECT 175.600 463.600 176.400 464.400 ;
        RECT 198.000 474.400 198.800 475.200 ;
        RECT 201.200 475.000 202.000 475.800 ;
        RECT 196.400 472.400 197.200 473.200 ;
        RECT 180.400 465.600 181.200 466.400 ;
        RECT 183.600 465.600 184.400 466.400 ;
        RECT 221.800 471.800 222.600 472.600 ;
        RECT 244.400 474.400 245.200 475.200 ;
        RECT 247.600 475.000 248.400 475.800 ;
        RECT 242.800 472.400 243.600 473.200 ;
        RECT 206.000 467.600 206.800 468.400 ;
        RECT 202.800 465.600 203.600 466.400 ;
        RECT 196.400 464.200 197.200 465.000 ;
        RECT 198.000 464.200 198.800 465.000 ;
        RECT 199.600 464.200 200.400 465.000 ;
        RECT 201.200 464.200 202.000 465.000 ;
        RECT 204.400 464.200 205.200 465.000 ;
        RECT 207.600 464.200 208.400 465.000 ;
        RECT 209.200 464.200 210.000 465.000 ;
        RECT 210.800 464.200 211.600 465.000 ;
        RECT 221.800 466.200 222.600 467.000 ;
        RECT 230.000 467.600 230.800 468.400 ;
        RECT 241.200 469.600 242.000 470.400 ;
        RECT 252.400 467.600 253.200 468.400 ;
        RECT 249.200 465.600 250.000 466.400 ;
        RECT 273.200 469.600 274.000 470.400 ;
        RECT 292.400 477.600 293.200 478.400 ;
        RECT 303.600 477.600 304.400 478.400 ;
        RECT 242.800 464.200 243.600 465.000 ;
        RECT 244.400 464.200 245.200 465.000 ;
        RECT 246.000 464.200 246.800 465.000 ;
        RECT 247.600 464.200 248.400 465.000 ;
        RECT 250.800 464.200 251.600 465.000 ;
        RECT 254.000 464.200 254.800 465.000 ;
        RECT 255.600 464.200 256.400 465.000 ;
        RECT 257.200 464.200 258.000 465.000 ;
        RECT 279.600 465.600 280.400 466.400 ;
        RECT 295.600 465.600 296.400 466.400 ;
        RECT 292.400 463.600 293.200 464.400 ;
        RECT 305.200 467.600 306.000 468.400 ;
        RECT 306.800 465.600 307.600 466.400 ;
        RECT 319.600 467.600 320.400 468.400 ;
        RECT 327.600 467.600 328.400 468.400 ;
        RECT 332.400 467.600 333.200 468.400 ;
        RECT 338.800 469.600 339.600 470.400 ;
        RECT 343.600 467.600 344.400 468.400 ;
        RECT 330.800 463.600 331.600 464.400 ;
        RECT 335.600 463.600 336.400 464.400 ;
        RECT 350.000 463.600 350.800 464.400 ;
        RECT 359.600 467.600 360.400 468.400 ;
        RECT 369.200 469.600 370.000 470.400 ;
        RECT 370.800 467.600 371.600 468.400 ;
        RECT 394.800 475.000 395.600 475.800 ;
        RECT 391.600 473.600 392.400 474.400 ;
        RECT 409.200 477.600 410.000 478.400 ;
        RECT 396.400 472.400 397.200 473.200 ;
        RECT 401.200 469.600 402.000 470.400 ;
        RECT 385.200 468.200 386.000 469.000 ;
        RECT 394.800 468.600 395.600 469.400 ;
        RECT 354.800 463.600 355.600 464.400 ;
        RECT 358.000 463.600 358.800 464.400 ;
        RECT 364.400 463.600 365.200 464.400 ;
        RECT 390.000 467.600 390.800 468.400 ;
        RECT 385.200 464.200 386.000 465.000 ;
        RECT 386.800 464.200 387.600 465.000 ;
        RECT 388.400 464.200 389.200 465.000 ;
        RECT 391.600 464.200 392.400 465.000 ;
        RECT 394.800 464.200 395.600 465.000 ;
        RECT 396.400 464.200 397.200 465.000 ;
        RECT 398.000 464.200 398.800 465.000 ;
        RECT 399.600 464.200 400.400 465.000 ;
        RECT 428.400 471.600 429.200 472.400 ;
        RECT 442.800 473.600 443.600 474.400 ;
        RECT 423.600 469.600 424.400 470.400 ;
        RECT 434.800 469.600 435.600 470.400 ;
        RECT 457.200 474.400 458.000 475.200 ;
        RECT 460.400 475.000 461.200 475.800 ;
        RECT 455.600 472.400 456.400 473.200 ;
        RECT 445.800 469.600 446.600 470.400 ;
        RECT 430.000 467.600 430.800 468.400 ;
        RECT 454.000 469.600 454.800 470.400 ;
        RECT 431.600 463.600 432.400 464.400 ;
        RECT 442.800 463.600 443.600 464.400 ;
        RECT 465.200 467.600 466.000 468.400 ;
        RECT 462.000 465.600 462.800 466.400 ;
        RECT 455.600 464.200 456.400 465.000 ;
        RECT 457.200 464.200 458.000 465.000 ;
        RECT 458.800 464.200 459.600 465.000 ;
        RECT 460.400 464.200 461.200 465.000 ;
        RECT 463.600 464.200 464.400 465.000 ;
        RECT 466.800 464.200 467.600 465.000 ;
        RECT 468.400 464.200 469.200 465.000 ;
        RECT 470.000 464.200 470.800 465.000 ;
        RECT 497.200 475.000 498.000 475.800 ;
        RECT 494.000 473.600 494.800 474.400 ;
        RECT 511.600 477.600 512.400 478.400 ;
        RECT 498.800 472.400 499.600 473.200 ;
        RECT 529.200 477.600 530.000 478.400 ;
        RECT 487.600 468.200 488.400 469.000 ;
        RECT 497.200 468.600 498.000 469.400 ;
        RECT 492.400 467.600 493.200 468.400 ;
        RECT 487.600 464.200 488.400 465.000 ;
        RECT 489.200 464.200 490.000 465.000 ;
        RECT 490.800 464.200 491.600 465.000 ;
        RECT 494.000 464.200 494.800 465.000 ;
        RECT 497.200 464.200 498.000 465.000 ;
        RECT 498.800 464.200 499.600 465.000 ;
        RECT 500.400 464.200 501.200 465.000 ;
        RECT 502.000 464.200 502.800 465.000 ;
        RECT 518.000 469.600 518.800 470.400 ;
        RECT 527.600 467.600 528.400 468.400 ;
        RECT 545.200 474.400 546.000 475.200 ;
        RECT 548.400 475.000 549.200 475.800 ;
        RECT 543.600 472.400 544.400 473.200 ;
        RECT 514.800 463.600 515.600 464.400 ;
        RECT 526.000 463.600 526.800 464.400 ;
        RECT 586.800 477.600 587.600 478.400 ;
        RECT 553.200 467.600 554.000 468.400 ;
        RECT 550.000 465.600 550.800 466.400 ;
        RECT 543.600 464.200 544.400 465.000 ;
        RECT 545.200 464.200 546.000 465.000 ;
        RECT 546.800 464.200 547.600 465.000 ;
        RECT 548.400 464.200 549.200 465.000 ;
        RECT 551.600 464.200 552.400 465.000 ;
        RECT 554.800 464.200 555.600 465.000 ;
        RECT 556.400 464.200 557.200 465.000 ;
        RECT 558.000 464.200 558.800 465.000 ;
        RECT 567.600 465.600 568.400 466.400 ;
        RECT 585.200 467.600 586.000 468.400 ;
        RECT 593.200 469.600 594.000 470.400 ;
        RECT 609.200 469.600 610.000 470.400 ;
        RECT 610.800 467.600 611.600 468.400 ;
        RECT 612.400 467.600 613.200 468.400 ;
        RECT 623.600 471.800 624.400 472.600 ;
        RECT 633.200 469.600 634.000 470.400 ;
        RECT 634.800 469.600 635.600 470.400 ;
        RECT 620.400 467.600 621.200 468.400 ;
        RECT 602.800 463.600 603.600 464.400 ;
        RECT 623.600 466.200 624.400 467.000 ;
        RECT 631.600 467.600 632.400 468.400 ;
        RECT 642.800 469.600 643.600 470.400 ;
        RECT 644.400 469.600 645.200 470.400 ;
        RECT 655.600 469.600 656.400 470.400 ;
        RECT 628.400 466.400 629.200 467.200 ;
        RECT 657.200 467.600 658.000 468.400 ;
        RECT 673.200 472.400 674.000 473.200 ;
        RECT 676.400 471.000 677.200 471.800 ;
        RECT 678.000 469.600 678.800 470.400 ;
        RECT 647.600 463.600 648.400 464.400 ;
        RECT 652.400 463.600 653.200 464.400 ;
        RECT 676.400 466.200 677.200 467.000 ;
        RECT 658.800 463.600 659.600 464.400 ;
        RECT 38.000 457.600 38.800 458.400 ;
        RECT 17.200 453.600 18.000 454.400 ;
        RECT 6.000 452.200 6.800 453.000 ;
        RECT 14.000 451.800 14.800 452.600 ;
        RECT 18.800 450.200 19.600 451.000 ;
        RECT 1.200 443.600 2.000 444.400 ;
        RECT 52.400 453.600 53.200 454.400 ;
        RECT 39.600 449.600 40.400 450.400 ;
        RECT 49.200 449.600 50.000 450.400 ;
        RECT 58.800 451.600 59.600 452.400 ;
        RECT 70.000 449.600 70.800 450.400 ;
        RECT 84.400 451.800 85.200 452.600 ;
        RECT 79.600 450.200 80.400 451.000 ;
        RECT 97.200 443.600 98.000 444.400 ;
        RECT 103.600 449.600 104.400 450.400 ;
        RECT 126.000 453.600 126.800 454.400 ;
        RECT 121.200 452.200 122.000 453.000 ;
        RECT 134.000 450.200 134.800 451.000 ;
        RECT 116.400 443.600 117.200 444.400 ;
        RECT 153.200 457.600 154.000 458.400 ;
        RECT 145.200 453.600 146.000 454.400 ;
        RECT 135.600 443.600 136.400 444.400 ;
        RECT 182.000 453.600 182.800 454.400 ;
        RECT 153.200 449.600 154.000 450.400 ;
        RECT 161.200 451.600 162.000 452.400 ;
        RECT 167.600 451.600 168.400 452.400 ;
        RECT 180.400 451.800 181.200 452.600 ;
        RECT 174.000 449.600 174.800 450.400 ;
        RECT 175.600 450.200 176.400 451.000 ;
        RECT 206.000 457.600 206.800 458.400 ;
        RECT 206.000 454.800 206.800 455.600 ;
        RECT 209.200 453.600 210.000 454.400 ;
        RECT 198.000 451.600 198.800 452.400 ;
        RECT 214.000 451.600 214.800 452.400 ;
        RECT 190.000 447.600 190.800 448.400 ;
        RECT 193.200 447.600 194.000 448.400 ;
        RECT 210.800 443.600 211.600 444.400 ;
        RECT 222.000 449.600 222.800 450.400 ;
        RECT 244.400 455.600 245.200 456.400 ;
        RECT 246.000 454.200 246.800 455.000 ;
        RECT 257.200 451.600 258.000 452.400 ;
        RECT 225.200 443.600 226.000 444.400 ;
        RECT 239.600 446.800 240.400 447.600 ;
        RECT 242.800 446.200 243.600 447.000 ;
        RECT 238.000 444.200 238.800 445.000 ;
        RECT 239.600 444.200 240.400 445.000 ;
        RECT 241.200 444.200 242.000 445.000 ;
        RECT 246.000 446.200 246.800 447.000 ;
        RECT 249.200 446.200 250.000 447.000 ;
        RECT 274.800 453.000 275.600 453.800 ;
        RECT 284.400 452.600 285.200 453.400 ;
        RECT 290.800 451.600 291.600 452.400 ;
        RECT 276.400 448.800 277.200 449.600 ;
        RECT 281.200 447.600 282.000 448.400 ;
        RECT 250.800 444.200 251.600 445.000 ;
        RECT 252.400 444.200 253.200 445.000 ;
        RECT 278.000 446.200 278.800 447.000 ;
        RECT 274.800 444.200 275.600 445.000 ;
        RECT 276.400 444.200 277.200 445.000 ;
        RECT 281.200 446.200 282.000 447.000 ;
        RECT 284.400 446.200 285.200 447.000 ;
        RECT 286.000 444.200 286.800 445.000 ;
        RECT 287.600 444.200 288.400 445.000 ;
        RECT 289.200 444.200 290.000 445.000 ;
        RECT 311.600 453.600 312.400 454.400 ;
        RECT 350.000 453.600 350.800 454.400 ;
        RECT 314.800 451.600 315.600 452.400 ;
        RECT 322.800 451.600 323.600 452.400 ;
        RECT 298.800 443.600 299.600 444.400 ;
        RECT 342.000 451.600 342.800 452.400 ;
        RECT 366.000 451.600 366.800 452.400 ;
        RECT 372.400 451.600 373.200 452.400 ;
        RECT 378.800 451.600 379.600 452.400 ;
        RECT 410.800 455.600 411.600 456.400 ;
        RECT 412.400 454.200 413.200 455.000 ;
        RECT 436.400 457.600 437.200 458.400 ;
        RECT 423.600 451.600 424.400 452.400 ;
        RECT 359.600 443.600 360.400 444.400 ;
        RECT 362.800 445.600 363.600 446.400 ;
        RECT 366.000 443.600 366.800 444.400 ;
        RECT 372.400 445.600 373.200 446.400 ;
        RECT 378.800 443.600 379.600 444.400 ;
        RECT 388.400 445.600 389.200 446.400 ;
        RECT 394.800 443.600 395.600 444.400 ;
        RECT 406.000 446.800 406.800 447.600 ;
        RECT 409.200 446.200 410.000 447.000 ;
        RECT 404.400 444.200 405.200 445.000 ;
        RECT 406.000 444.200 406.800 445.000 ;
        RECT 407.600 444.200 408.400 445.000 ;
        RECT 412.400 446.200 413.200 447.000 ;
        RECT 415.600 446.200 416.400 447.000 ;
        RECT 417.200 444.200 418.000 445.000 ;
        RECT 418.800 444.200 419.600 445.000 ;
        RECT 446.000 453.000 446.800 453.800 ;
        RECT 436.400 449.600 437.200 450.400 ;
        RECT 455.600 452.600 456.400 453.400 ;
        RECT 476.400 457.600 477.200 458.400 ;
        RECT 450.800 451.600 451.600 452.400 ;
        RECT 447.600 448.800 448.400 449.600 ;
        RECT 452.400 447.600 453.200 448.400 ;
        RECT 449.200 446.200 450.000 447.000 ;
        RECT 446.000 444.200 446.800 445.000 ;
        RECT 447.600 444.200 448.400 445.000 ;
        RECT 452.400 446.200 453.200 447.000 ;
        RECT 455.600 446.200 456.400 447.000 ;
        RECT 457.200 444.200 458.000 445.000 ;
        RECT 458.800 444.200 459.600 445.000 ;
        RECT 460.400 444.200 461.200 445.000 ;
        RECT 470.000 443.600 470.800 444.400 ;
        RECT 478.000 455.600 478.800 456.400 ;
        RECT 476.400 449.600 477.200 450.400 ;
        RECT 484.400 451.600 485.200 452.400 ;
        RECT 486.000 449.600 486.800 450.400 ;
        RECT 492.400 457.600 493.200 458.400 ;
        RECT 505.200 453.000 506.000 453.800 ;
        RECT 495.600 451.600 496.400 452.400 ;
        RECT 514.800 452.600 515.600 453.400 ;
        RECT 502.000 451.600 502.800 452.400 ;
        RECT 503.600 451.600 504.400 452.400 ;
        RECT 550.000 457.600 550.800 458.400 ;
        RECT 506.800 448.800 507.600 449.600 ;
        RECT 511.600 447.600 512.400 448.400 ;
        RECT 508.400 446.200 509.200 447.000 ;
        RECT 505.200 444.200 506.000 445.000 ;
        RECT 506.800 444.200 507.600 445.000 ;
        RECT 511.600 446.200 512.400 447.000 ;
        RECT 514.800 446.200 515.600 447.000 ;
        RECT 516.400 444.200 517.200 445.000 ;
        RECT 518.000 444.200 518.800 445.000 ;
        RECT 519.600 444.200 520.400 445.000 ;
        RECT 550.000 449.600 550.800 450.400 ;
        RECT 578.800 455.600 579.600 456.400 ;
        RECT 580.400 454.200 581.200 455.000 ;
        RECT 596.400 457.600 597.200 458.400 ;
        RECT 610.800 457.600 611.600 458.400 ;
        RECT 570.800 451.600 571.600 452.400 ;
        RECT 591.600 451.600 592.400 452.400 ;
        RECT 554.800 443.600 555.600 444.400 ;
        RECT 574.000 446.800 574.800 447.600 ;
        RECT 577.200 446.200 578.000 447.000 ;
        RECT 572.400 444.200 573.200 445.000 ;
        RECT 574.000 444.200 574.800 445.000 ;
        RECT 575.600 444.200 576.400 445.000 ;
        RECT 580.400 446.200 581.200 447.000 ;
        RECT 583.600 446.200 584.400 447.000 ;
        RECT 612.400 453.600 613.200 454.400 ;
        RECT 614.000 451.600 614.800 452.400 ;
        RECT 636.400 457.600 637.200 458.400 ;
        RECT 620.400 451.600 621.200 452.400 ;
        RECT 585.200 444.200 586.000 445.000 ;
        RECT 586.800 444.200 587.600 445.000 ;
        RECT 617.200 449.600 618.000 450.400 ;
        RECT 631.600 451.600 632.400 452.400 ;
        RECT 652.400 455.600 653.200 456.400 ;
        RECT 654.000 454.200 654.800 455.000 ;
        RECT 681.200 457.600 682.000 458.400 ;
        RECT 670.000 453.600 670.800 454.400 ;
        RECT 644.400 451.600 645.200 452.400 ;
        RECT 662.000 451.600 662.800 452.400 ;
        RECT 626.800 447.600 627.600 448.400 ;
        RECT 628.400 445.600 629.200 446.400 ;
        RECT 647.600 446.800 648.400 447.600 ;
        RECT 650.800 446.200 651.600 447.000 ;
        RECT 646.000 444.200 646.800 445.000 ;
        RECT 647.600 444.200 648.400 445.000 ;
        RECT 649.200 444.200 650.000 445.000 ;
        RECT 654.000 446.200 654.800 447.000 ;
        RECT 657.200 446.200 658.000 447.000 ;
        RECT 658.800 444.200 659.600 445.000 ;
        RECT 660.400 444.200 661.200 445.000 ;
        RECT 681.200 443.600 682.000 444.400 ;
        RECT 1.200 433.600 2.000 434.400 ;
        RECT 15.600 432.400 16.400 433.200 ;
        RECT 18.800 431.000 19.600 431.800 ;
        RECT 22.000 429.600 22.800 430.400 ;
        RECT 23.600 429.600 24.400 430.400 ;
        RECT 30.000 429.600 30.800 430.400 ;
        RECT 18.800 426.200 19.600 427.000 ;
        RECT 31.600 427.600 32.400 428.400 ;
        RECT 39.600 429.600 40.400 430.400 ;
        RECT 41.200 429.600 42.000 430.400 ;
        RECT 46.000 429.600 46.800 430.400 ;
        RECT 47.600 427.600 48.400 428.400 ;
        RECT 54.000 429.600 54.800 430.400 ;
        RECT 55.600 429.600 56.400 430.400 ;
        RECT 57.200 429.600 58.000 430.400 ;
        RECT 50.800 423.600 51.600 424.400 ;
        RECT 71.600 429.600 72.400 430.400 ;
        RECT 73.200 429.600 74.000 430.400 ;
        RECT 76.400 429.600 77.200 430.400 ;
        RECT 84.400 431.600 85.200 432.400 ;
        RECT 84.400 429.600 85.200 430.400 ;
        RECT 86.000 427.600 86.800 428.400 ;
        RECT 102.000 432.400 102.800 433.200 ;
        RECT 105.200 431.000 106.000 431.800 ;
        RECT 124.400 437.600 125.200 438.400 ;
        RECT 129.200 437.600 130.000 438.400 ;
        RECT 118.000 429.600 118.800 430.400 ;
        RECT 119.600 429.600 120.400 430.400 ;
        RECT 137.200 437.600 138.000 438.400 ;
        RECT 105.200 426.200 106.000 427.000 ;
        RECT 87.600 423.600 88.400 424.400 ;
        RECT 132.400 429.600 133.200 430.400 ;
        RECT 154.800 432.400 155.600 433.200 ;
        RECT 158.000 431.000 158.800 431.800 ;
        RECT 169.200 433.600 170.000 434.400 ;
        RECT 162.800 429.600 163.600 430.400 ;
        RECT 185.200 437.600 186.000 438.400 ;
        RECT 169.200 429.600 170.000 430.400 ;
        RECT 172.400 429.600 173.200 430.400 ;
        RECT 174.000 429.600 174.800 430.400 ;
        RECT 158.000 426.200 158.800 427.000 ;
        RECT 164.400 427.600 165.200 428.400 ;
        RECT 170.800 427.600 171.600 428.400 ;
        RECT 185.200 429.600 186.000 430.400 ;
        RECT 140.400 423.600 141.200 424.400 ;
        RECT 186.800 427.600 187.600 428.400 ;
        RECT 209.200 432.400 210.000 433.200 ;
        RECT 212.400 431.000 213.200 431.800 ;
        RECT 212.400 426.200 213.200 427.000 ;
        RECT 194.800 423.600 195.600 424.400 ;
        RECT 214.000 425.600 214.800 426.400 ;
        RECT 215.600 423.600 216.400 424.400 ;
        RECT 220.400 425.600 221.200 426.400 ;
        RECT 223.600 423.600 224.400 424.400 ;
        RECT 252.400 434.400 253.200 435.200 ;
        RECT 255.600 435.000 256.400 435.800 ;
        RECT 281.200 437.600 282.000 438.400 ;
        RECT 250.800 432.400 251.600 433.200 ;
        RECT 231.600 427.600 232.400 428.400 ;
        RECT 238.000 425.600 238.800 426.400 ;
        RECT 241.200 425.600 242.000 426.400 ;
        RECT 236.400 423.600 237.200 424.400 ;
        RECT 279.600 433.600 280.400 434.400 ;
        RECT 260.400 427.600 261.200 428.400 ;
        RECT 257.200 425.600 258.000 426.400 ;
        RECT 250.800 424.200 251.600 425.000 ;
        RECT 252.400 424.200 253.200 425.000 ;
        RECT 254.000 424.200 254.800 425.000 ;
        RECT 255.600 424.200 256.400 425.000 ;
        RECT 258.800 424.200 259.600 425.000 ;
        RECT 262.000 424.200 262.800 425.000 ;
        RECT 263.600 424.200 264.400 425.000 ;
        RECT 265.200 424.200 266.000 425.000 ;
        RECT 308.400 437.600 309.200 438.400 ;
        RECT 282.800 427.600 283.600 428.400 ;
        RECT 300.400 429.600 301.200 430.400 ;
        RECT 308.400 429.600 309.200 430.400 ;
        RECT 286.000 423.600 286.800 424.400 ;
        RECT 313.200 425.600 314.000 426.400 ;
        RECT 314.800 425.600 315.600 426.400 ;
        RECT 324.400 427.600 325.200 428.400 ;
        RECT 330.800 437.600 331.600 438.400 ;
        RECT 329.200 427.600 330.000 428.400 ;
        RECT 342.000 433.600 342.800 434.400 ;
        RECT 351.600 437.600 352.400 438.400 ;
        RECT 340.400 429.600 341.200 430.400 ;
        RECT 345.200 429.600 346.000 430.400 ;
        RECT 348.400 429.600 349.200 430.400 ;
        RECT 346.800 427.600 347.600 428.400 ;
        RECT 350.000 427.600 350.800 428.400 ;
        RECT 362.800 437.600 363.600 438.400 ;
        RECT 369.200 437.600 370.000 438.400 ;
        RECT 364.400 433.600 365.200 434.400 ;
        RECT 356.400 429.600 357.200 430.400 ;
        RECT 359.600 429.600 360.400 430.400 ;
        RECT 367.600 431.600 368.400 432.400 ;
        RECT 366.000 429.600 366.800 430.400 ;
        RECT 358.000 427.600 358.800 428.400 ;
        RECT 353.200 425.600 354.000 426.400 ;
        RECT 361.200 427.600 362.000 428.400 ;
        RECT 372.400 437.600 373.200 438.400 ;
        RECT 374.000 433.600 374.800 434.400 ;
        RECT 377.200 431.600 378.000 432.400 ;
        RECT 398.000 437.600 398.800 438.400 ;
        RECT 375.600 429.600 376.400 430.400 ;
        RECT 370.800 425.600 371.600 426.400 ;
        RECT 388.400 429.600 389.200 430.400 ;
        RECT 393.200 429.600 394.000 430.400 ;
        RECT 391.600 427.600 392.400 428.400 ;
        RECT 385.200 423.600 386.000 424.400 ;
        RECT 394.800 427.600 395.600 428.400 ;
        RECT 396.400 427.600 397.200 428.400 ;
        RECT 423.600 435.000 424.400 435.800 ;
        RECT 420.400 433.600 421.200 434.400 ;
        RECT 438.000 437.600 438.800 438.400 ;
        RECT 425.200 432.400 426.000 433.200 ;
        RECT 430.000 429.600 430.800 430.400 ;
        RECT 414.000 428.200 414.800 429.000 ;
        RECT 423.600 428.600 424.400 429.400 ;
        RECT 418.800 427.600 419.600 428.400 ;
        RECT 414.000 424.200 414.800 425.000 ;
        RECT 415.600 424.200 416.400 425.000 ;
        RECT 417.200 424.200 418.000 425.000 ;
        RECT 420.400 424.200 421.200 425.000 ;
        RECT 423.600 424.200 424.400 425.000 ;
        RECT 425.200 424.200 426.000 425.000 ;
        RECT 426.800 424.200 427.600 425.000 ;
        RECT 428.400 424.200 429.200 425.000 ;
        RECT 446.000 437.600 446.800 438.400 ;
        RECT 452.400 437.600 453.200 438.400 ;
        RECT 442.800 425.600 443.600 426.400 ;
        RECT 449.200 429.600 450.000 430.400 ;
        RECT 482.800 435.000 483.600 435.800 ;
        RECT 479.600 433.600 480.400 434.400 ;
        RECT 484.400 432.400 485.200 433.200 ;
        RECT 473.200 428.200 474.000 429.000 ;
        RECT 482.800 428.600 483.600 429.400 ;
        RECT 441.200 423.600 442.000 424.400 ;
        RECT 452.400 423.600 453.200 424.400 ;
        RECT 478.000 427.600 478.800 428.400 ;
        RECT 473.200 424.200 474.000 425.000 ;
        RECT 474.800 424.200 475.600 425.000 ;
        RECT 476.400 424.200 477.200 425.000 ;
        RECT 479.600 424.200 480.400 425.000 ;
        RECT 482.800 424.200 483.600 425.000 ;
        RECT 484.400 424.200 485.200 425.000 ;
        RECT 486.000 424.200 486.800 425.000 ;
        RECT 487.600 424.200 488.400 425.000 ;
        RECT 518.000 437.600 518.800 438.400 ;
        RECT 503.600 429.600 504.400 430.400 ;
        RECT 505.200 427.600 506.000 428.400 ;
        RECT 522.800 427.600 523.600 428.400 ;
        RECT 526.000 429.600 526.800 430.400 ;
        RECT 529.200 429.600 530.000 430.400 ;
        RECT 538.800 437.600 539.600 438.400 ;
        RECT 543.600 437.600 544.400 438.400 ;
        RECT 550.000 437.600 550.800 438.400 ;
        RECT 534.000 425.600 534.800 426.400 ;
        RECT 566.000 434.400 566.800 435.200 ;
        RECT 569.200 435.000 570.000 435.800 ;
        RECT 564.400 432.400 565.200 433.200 ;
        RECT 550.000 429.600 550.800 430.400 ;
        RECT 538.800 423.600 539.600 424.400 ;
        RECT 551.600 427.600 552.400 428.400 ;
        RECT 583.600 431.600 584.400 432.400 ;
        RECT 554.800 423.600 555.600 424.400 ;
        RECT 574.000 427.600 574.800 428.400 ;
        RECT 570.800 425.600 571.600 426.400 ;
        RECT 564.400 424.200 565.200 425.000 ;
        RECT 566.000 424.200 566.800 425.000 ;
        RECT 567.600 424.200 568.400 425.000 ;
        RECT 569.200 424.200 570.000 425.000 ;
        RECT 572.400 424.200 573.200 425.000 ;
        RECT 575.600 424.200 576.400 425.000 ;
        RECT 577.200 424.200 578.000 425.000 ;
        RECT 578.800 424.200 579.600 425.000 ;
        RECT 612.400 434.400 613.200 435.200 ;
        RECT 615.600 435.000 616.400 435.800 ;
        RECT 636.400 437.600 637.200 438.400 ;
        RECT 610.800 432.400 611.600 433.200 ;
        RECT 609.200 429.600 610.000 430.400 ;
        RECT 601.200 423.600 602.000 424.400 ;
        RECT 620.400 427.600 621.200 428.400 ;
        RECT 617.200 425.600 618.000 426.400 ;
        RECT 610.800 424.200 611.600 425.000 ;
        RECT 612.400 424.200 613.200 425.000 ;
        RECT 614.000 424.200 614.800 425.000 ;
        RECT 615.600 424.200 616.400 425.000 ;
        RECT 618.800 424.200 619.600 425.000 ;
        RECT 622.000 424.200 622.800 425.000 ;
        RECT 623.600 424.200 624.400 425.000 ;
        RECT 625.200 424.200 626.000 425.000 ;
        RECT 662.000 434.400 662.800 435.200 ;
        RECT 665.200 435.000 666.000 435.800 ;
        RECT 660.400 432.400 661.200 433.200 ;
        RECT 658.800 429.600 659.600 430.400 ;
        RECT 650.800 423.600 651.600 424.400 ;
        RECT 670.000 427.600 670.800 428.400 ;
        RECT 666.800 425.600 667.600 426.400 ;
        RECT 660.400 424.200 661.200 425.000 ;
        RECT 662.000 424.200 662.800 425.000 ;
        RECT 663.600 424.200 664.400 425.000 ;
        RECT 665.200 424.200 666.000 425.000 ;
        RECT 668.400 424.200 669.200 425.000 ;
        RECT 671.600 424.200 672.400 425.000 ;
        RECT 673.200 424.200 674.000 425.000 ;
        RECT 674.800 424.200 675.600 425.000 ;
        RECT 1.200 410.200 2.000 411.000 ;
        RECT 23.600 411.600 24.400 412.400 ;
        RECT 18.800 407.600 19.600 408.400 ;
        RECT 25.200 409.600 26.000 410.400 ;
        RECT 50.800 413.600 51.600 414.400 ;
        RECT 47.600 409.600 48.400 410.400 ;
        RECT 57.200 411.600 58.000 412.400 ;
        RECT 58.800 411.600 59.600 412.400 ;
        RECT 66.800 403.600 67.600 404.400 ;
        RECT 84.400 413.600 85.200 414.400 ;
        RECT 73.200 412.200 74.000 413.000 ;
        RECT 86.000 410.200 86.800 411.000 ;
        RECT 68.400 407.600 69.200 408.400 ;
        RECT 98.800 413.600 99.600 414.400 ;
        RECT 97.200 410.200 98.000 411.000 ;
        RECT 89.200 403.600 90.000 404.400 ;
        RECT 92.400 403.600 93.200 404.400 ;
        RECT 129.200 403.600 130.000 404.400 ;
        RECT 140.400 411.600 141.200 412.400 ;
        RECT 150.000 411.600 150.800 412.400 ;
        RECT 185.200 417.600 186.000 418.400 ;
        RECT 193.200 417.600 194.000 418.400 ;
        RECT 166.000 413.600 166.800 414.400 ;
        RECT 143.600 403.600 144.400 404.400 ;
        RECT 150.000 403.600 150.800 404.400 ;
        RECT 167.600 409.600 168.400 410.400 ;
        RECT 174.000 409.600 174.800 410.400 ;
        RECT 183.600 409.600 184.400 410.400 ;
        RECT 209.200 415.600 210.000 416.400 ;
        RECT 210.800 414.200 211.600 415.000 ;
        RECT 201.200 411.600 202.000 412.400 ;
        RECT 193.200 403.600 194.000 404.400 ;
        RECT 204.400 406.800 205.200 407.600 ;
        RECT 207.600 406.200 208.400 407.000 ;
        RECT 202.800 404.200 203.600 405.000 ;
        RECT 204.400 404.200 205.200 405.000 ;
        RECT 206.000 404.200 206.800 405.000 ;
        RECT 210.800 406.200 211.600 407.000 ;
        RECT 214.000 406.200 214.800 407.000 ;
        RECT 215.600 404.200 216.400 405.000 ;
        RECT 217.200 404.200 218.000 405.000 ;
        RECT 236.400 413.600 237.200 414.400 ;
        RECT 231.600 409.600 232.400 410.400 ;
        RECT 247.600 409.600 248.400 410.400 ;
        RECT 273.200 413.000 274.000 413.800 ;
        RECT 282.800 412.600 283.600 413.400 ;
        RECT 274.800 408.800 275.600 409.600 ;
        RECT 279.600 407.600 280.400 408.400 ;
        RECT 276.400 406.200 277.200 407.000 ;
        RECT 273.200 404.200 274.000 405.000 ;
        RECT 274.800 404.200 275.600 405.000 ;
        RECT 279.600 406.200 280.400 407.000 ;
        RECT 282.800 406.200 283.600 407.000 ;
        RECT 284.400 404.200 285.200 405.000 ;
        RECT 286.000 404.200 286.800 405.000 ;
        RECT 287.600 404.200 288.400 405.000 ;
        RECT 300.400 409.600 301.200 410.400 ;
        RECT 297.200 403.600 298.000 404.400 ;
        RECT 322.800 417.600 323.600 418.400 ;
        RECT 330.800 417.600 331.600 418.400 ;
        RECT 340.400 417.600 341.200 418.400 ;
        RECT 348.400 417.600 349.200 418.400 ;
        RECT 311.600 409.600 312.400 410.400 ;
        RECT 332.400 413.600 333.200 414.400 ;
        RECT 334.000 411.600 334.800 412.400 ;
        RECT 335.600 409.600 336.400 410.400 ;
        RECT 350.000 413.600 350.800 414.400 ;
        RECT 351.600 411.600 352.400 412.400 ;
        RECT 356.400 411.600 357.200 412.400 ;
        RECT 337.200 407.600 338.000 408.400 ;
        RECT 366.000 411.600 366.800 412.400 ;
        RECT 361.200 409.600 362.000 410.400 ;
        RECT 390.000 413.600 390.800 414.400 ;
        RECT 378.800 411.600 379.600 412.400 ;
        RECT 382.000 411.600 382.800 412.400 ;
        RECT 359.600 407.600 360.400 408.400 ;
        RECT 362.800 403.600 363.600 404.400 ;
        RECT 370.800 405.600 371.600 406.400 ;
        RECT 378.800 405.600 379.600 406.400 ;
        RECT 385.200 411.600 386.000 412.400 ;
        RECT 391.600 411.600 392.400 412.400 ;
        RECT 386.800 405.600 387.600 406.400 ;
        RECT 417.200 417.600 418.000 418.400 ;
        RECT 402.800 413.600 403.600 414.400 ;
        RECT 406.000 411.600 406.800 412.400 ;
        RECT 433.200 415.600 434.000 416.400 ;
        RECT 434.800 414.200 435.600 415.000 ;
        RECT 425.200 411.600 426.000 412.400 ;
        RECT 447.600 411.600 448.400 412.400 ;
        RECT 394.800 403.600 395.600 404.400 ;
        RECT 428.400 406.800 429.200 407.600 ;
        RECT 431.600 406.200 432.400 407.000 ;
        RECT 426.800 404.200 427.600 405.000 ;
        RECT 428.400 404.200 429.200 405.000 ;
        RECT 430.000 404.200 430.800 405.000 ;
        RECT 434.800 406.200 435.600 407.000 ;
        RECT 438.000 406.200 438.800 407.000 ;
        RECT 458.800 413.000 459.600 413.800 ;
        RECT 468.400 412.600 469.200 413.400 ;
        RECT 492.400 417.600 493.200 418.400 ;
        RECT 454.000 411.600 454.800 412.400 ;
        RECT 455.600 411.600 456.400 412.400 ;
        RECT 489.200 411.600 490.000 412.400 ;
        RECT 460.400 408.800 461.200 409.600 ;
        RECT 465.200 407.600 466.000 408.400 ;
        RECT 439.600 404.200 440.400 405.000 ;
        RECT 441.200 404.200 442.000 405.000 ;
        RECT 462.000 406.200 462.800 407.000 ;
        RECT 458.800 404.200 459.600 405.000 ;
        RECT 460.400 404.200 461.200 405.000 ;
        RECT 465.200 406.200 466.000 407.000 ;
        RECT 468.400 406.200 469.200 407.000 ;
        RECT 470.000 404.200 470.800 405.000 ;
        RECT 471.600 404.200 472.400 405.000 ;
        RECT 473.200 404.200 474.000 405.000 ;
        RECT 482.800 403.600 483.600 404.400 ;
        RECT 490.800 409.600 491.600 410.400 ;
        RECT 506.800 413.600 507.600 414.400 ;
        RECT 526.000 415.600 526.800 416.400 ;
        RECT 527.600 414.200 528.400 415.000 ;
        RECT 518.000 411.600 518.800 412.400 ;
        RECT 540.400 411.600 541.200 412.400 ;
        RECT 506.800 409.600 507.600 410.400 ;
        RECT 510.000 407.600 510.800 408.400 ;
        RECT 521.200 406.800 522.000 407.600 ;
        RECT 524.400 406.200 525.200 407.000 ;
        RECT 519.600 404.200 520.400 405.000 ;
        RECT 521.200 404.200 522.000 405.000 ;
        RECT 522.800 404.200 523.600 405.000 ;
        RECT 527.600 406.200 528.400 407.000 ;
        RECT 530.800 406.200 531.600 407.000 ;
        RECT 554.800 417.600 555.600 418.400 ;
        RECT 548.400 411.600 549.200 412.400 ;
        RECT 569.200 413.600 570.000 414.400 ;
        RECT 532.400 404.200 533.200 405.000 ;
        RECT 534.000 404.200 534.800 405.000 ;
        RECT 545.200 403.600 546.000 404.400 ;
        RECT 554.800 409.600 555.600 410.400 ;
        RECT 556.400 409.600 557.200 410.400 ;
        RECT 594.800 415.600 595.600 416.400 ;
        RECT 596.400 414.200 597.200 415.000 ;
        RECT 618.800 417.600 619.600 418.400 ;
        RECT 615.600 414.800 616.400 415.600 ;
        RECT 586.800 411.600 587.600 412.400 ;
        RECT 609.200 411.600 610.000 412.400 ;
        RECT 570.800 409.600 571.600 410.400 ;
        RECT 590.000 406.800 590.800 407.600 ;
        RECT 593.200 406.200 594.000 407.000 ;
        RECT 588.400 404.200 589.200 405.000 ;
        RECT 590.000 404.200 590.800 405.000 ;
        RECT 591.600 404.200 592.400 405.000 ;
        RECT 596.400 406.200 597.200 407.000 ;
        RECT 599.600 406.200 600.400 407.000 ;
        RECT 622.000 413.600 622.800 414.400 ;
        RECT 644.400 417.600 645.200 418.400 ;
        RECT 601.200 404.200 602.000 405.000 ;
        RECT 602.800 404.200 603.600 405.000 ;
        RECT 623.600 409.600 624.400 410.400 ;
        RECT 641.200 414.800 642.000 415.600 ;
        RECT 647.600 413.600 648.400 414.400 ;
        RECT 636.400 409.600 637.200 410.400 ;
        RECT 666.800 415.600 667.600 416.400 ;
        RECT 668.400 414.200 669.200 415.000 ;
        RECT 658.800 411.600 659.600 412.400 ;
        RECT 679.600 411.600 680.400 412.400 ;
        RECT 650.800 409.600 651.600 410.400 ;
        RECT 662.000 406.800 662.800 407.600 ;
        RECT 665.200 406.200 666.000 407.000 ;
        RECT 660.400 404.200 661.200 405.000 ;
        RECT 662.000 404.200 662.800 405.000 ;
        RECT 663.600 404.200 664.400 405.000 ;
        RECT 668.400 406.200 669.200 407.000 ;
        RECT 671.600 406.200 672.400 407.000 ;
        RECT 673.200 404.200 674.000 405.000 ;
        RECT 674.800 404.200 675.600 405.000 ;
        RECT 23.600 397.600 24.400 398.400 ;
        RECT 4.400 389.600 5.200 390.400 ;
        RECT 28.400 397.600 29.200 398.400 ;
        RECT 47.600 393.600 48.400 394.400 ;
        RECT 6.000 386.200 6.800 387.000 ;
        RECT 30.000 387.600 30.800 388.400 ;
        RECT 33.200 387.600 34.000 388.400 ;
        RECT 36.400 389.600 37.200 390.400 ;
        RECT 39.600 389.600 40.400 390.400 ;
        RECT 47.600 389.600 48.400 390.400 ;
        RECT 57.200 389.600 58.000 390.400 ;
        RECT 58.800 389.600 59.600 390.400 ;
        RECT 66.800 389.600 67.600 390.400 ;
        RECT 68.400 389.600 69.200 390.400 ;
        RECT 70.000 385.600 70.800 386.400 ;
        RECT 81.200 393.600 82.000 394.400 ;
        RECT 78.000 389.600 78.800 390.400 ;
        RECT 79.600 387.600 80.400 388.400 ;
        RECT 71.600 383.600 72.400 384.400 ;
        RECT 74.800 383.600 75.600 384.400 ;
        RECT 98.800 397.600 99.600 398.400 ;
        RECT 95.600 387.600 96.400 388.400 ;
        RECT 105.200 389.600 106.000 390.400 ;
        RECT 121.200 389.600 122.000 390.400 ;
        RECT 134.000 393.600 134.800 394.400 ;
        RECT 129.200 389.600 130.000 390.400 ;
        RECT 142.000 391.600 142.800 392.400 ;
        RECT 135.600 389.600 136.400 390.400 ;
        RECT 87.600 383.600 88.400 384.400 ;
        RECT 90.800 383.600 91.600 384.400 ;
        RECT 114.800 385.600 115.600 386.400 ;
        RECT 130.800 387.600 131.600 388.400 ;
        RECT 116.400 383.600 117.200 384.400 ;
        RECT 126.000 383.600 126.800 384.400 ;
        RECT 143.600 387.600 144.400 388.400 ;
        RECT 153.200 389.600 154.000 390.400 ;
        RECT 156.400 389.600 157.200 390.400 ;
        RECT 158.000 389.600 158.800 390.400 ;
        RECT 148.400 387.600 149.200 388.400 ;
        RECT 154.800 387.600 155.600 388.400 ;
        RECT 175.600 389.600 176.400 390.400 ;
        RECT 178.800 389.600 179.600 390.400 ;
        RECT 180.400 389.600 181.200 390.400 ;
        RECT 177.200 387.600 178.000 388.400 ;
        RECT 201.200 393.600 202.000 394.400 ;
        RECT 196.400 389.600 197.200 390.400 ;
        RECT 170.800 383.600 171.600 384.400 ;
        RECT 199.600 387.600 200.400 388.400 ;
        RECT 215.600 392.400 216.400 393.200 ;
        RECT 226.800 393.600 227.600 394.400 ;
        RECT 222.200 391.800 223.000 392.600 ;
        RECT 218.800 391.000 219.600 391.800 ;
        RECT 223.400 389.800 224.200 390.600 ;
        RECT 246.000 397.600 246.800 398.400 ;
        RECT 231.600 389.600 232.400 390.400 ;
        RECT 233.200 389.600 234.000 390.400 ;
        RECT 218.800 386.200 219.600 387.000 ;
        RECT 222.200 386.200 223.000 387.000 ;
        RECT 230.000 387.600 230.800 388.400 ;
        RECT 241.200 389.600 242.000 390.400 ;
        RECT 242.800 389.600 243.600 390.400 ;
        RECT 254.000 397.600 254.800 398.400 ;
        RECT 258.800 393.600 259.600 394.400 ;
        RECT 274.800 397.600 275.600 398.400 ;
        RECT 276.400 389.600 277.200 390.400 ;
        RECT 278.000 389.600 278.800 390.400 ;
        RECT 297.200 395.000 298.000 395.800 ;
        RECT 294.000 393.600 294.800 394.400 ;
        RECT 298.800 392.400 299.600 393.200 ;
        RECT 303.600 389.600 304.400 390.400 ;
        RECT 287.600 388.200 288.400 389.000 ;
        RECT 297.200 388.600 298.000 389.400 ;
        RECT 292.400 387.600 293.200 388.400 ;
        RECT 287.600 384.200 288.400 385.000 ;
        RECT 289.200 384.200 290.000 385.000 ;
        RECT 290.800 384.200 291.600 385.000 ;
        RECT 294.000 384.200 294.800 385.000 ;
        RECT 297.200 384.200 298.000 385.000 ;
        RECT 298.800 384.200 299.600 385.000 ;
        RECT 300.400 384.200 301.200 385.000 ;
        RECT 302.000 384.200 302.800 385.000 ;
        RECT 321.200 389.600 322.000 390.400 ;
        RECT 334.000 397.600 334.800 398.400 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 311.600 383.600 312.400 384.400 ;
        RECT 324.400 385.600 325.200 386.400 ;
        RECT 343.600 393.600 344.400 394.400 ;
        RECT 334.000 389.600 334.800 390.400 ;
        RECT 340.400 389.600 341.200 390.400 ;
        RECT 329.200 387.600 330.000 388.400 ;
        RECT 335.600 387.600 336.400 388.400 ;
        RECT 337.200 383.600 338.000 384.400 ;
        RECT 351.600 389.600 352.400 390.400 ;
        RECT 356.400 387.600 357.200 388.400 ;
        RECT 351.600 383.600 352.400 384.400 ;
        RECT 375.600 397.600 376.400 398.400 ;
        RECT 382.000 397.600 382.800 398.400 ;
        RECT 377.200 393.600 378.000 394.400 ;
        RECT 374.000 391.600 374.800 392.400 ;
        RECT 372.400 387.600 373.200 388.400 ;
        RECT 380.400 387.600 381.200 388.400 ;
        RECT 402.800 395.000 403.600 395.800 ;
        RECT 399.600 393.600 400.400 394.400 ;
        RECT 404.400 392.400 405.200 393.200 ;
        RECT 417.200 393.600 418.000 394.400 ;
        RECT 393.200 388.200 394.000 389.000 ;
        RECT 402.800 388.600 403.600 389.400 ;
        RECT 398.000 387.600 398.800 388.400 ;
        RECT 393.200 384.200 394.000 385.000 ;
        RECT 394.800 384.200 395.600 385.000 ;
        RECT 396.400 384.200 397.200 385.000 ;
        RECT 399.600 384.200 400.400 385.000 ;
        RECT 402.800 384.200 403.600 385.000 ;
        RECT 404.400 384.200 405.200 385.000 ;
        RECT 406.000 384.200 406.800 385.000 ;
        RECT 407.600 384.200 408.400 385.000 ;
        RECT 426.800 389.600 427.600 390.400 ;
        RECT 436.400 387.600 437.200 388.400 ;
        RECT 439.600 389.600 440.400 390.400 ;
        RECT 442.800 389.600 443.600 390.400 ;
        RECT 460.400 394.400 461.200 395.200 ;
        RECT 463.600 395.000 464.400 395.800 ;
        RECT 458.800 392.400 459.600 393.200 ;
        RECT 457.200 389.600 458.000 390.400 ;
        RECT 449.200 383.600 450.000 384.400 ;
        RECT 468.400 387.600 469.200 388.400 ;
        RECT 465.200 385.600 466.000 386.400 ;
        RECT 458.800 384.200 459.600 385.000 ;
        RECT 460.400 384.200 461.200 385.000 ;
        RECT 462.000 384.200 462.800 385.000 ;
        RECT 463.600 384.200 464.400 385.000 ;
        RECT 466.800 384.200 467.600 385.000 ;
        RECT 470.000 384.200 470.800 385.000 ;
        RECT 471.600 384.200 472.400 385.000 ;
        RECT 473.200 384.200 474.000 385.000 ;
        RECT 482.800 387.600 483.600 388.400 ;
        RECT 487.600 393.600 488.400 394.400 ;
        RECT 494.000 397.600 494.800 398.400 ;
        RECT 500.400 393.600 501.200 394.400 ;
        RECT 490.800 387.600 491.600 388.400 ;
        RECT 521.200 397.600 522.000 398.400 ;
        RECT 508.400 389.600 509.200 390.400 ;
        RECT 530.800 393.600 531.600 394.400 ;
        RECT 514.800 389.600 515.600 390.400 ;
        RECT 521.200 389.600 522.000 390.400 ;
        RECT 503.600 387.600 504.400 388.400 ;
        RECT 510.000 387.600 510.800 388.400 ;
        RECT 516.400 387.600 517.200 388.400 ;
        RECT 522.800 387.600 523.600 388.400 ;
        RECT 529.200 389.600 530.000 390.400 ;
        RECT 526.000 383.600 526.800 384.400 ;
        RECT 537.200 389.600 538.000 390.400 ;
        RECT 545.200 391.600 546.000 392.400 ;
        RECT 554.800 389.600 555.600 390.400 ;
        RECT 534.000 387.600 534.800 388.400 ;
        RECT 546.800 387.600 547.600 388.400 ;
        RECT 548.400 386.200 549.200 387.000 ;
        RECT 564.400 387.600 565.200 388.400 ;
        RECT 567.600 397.600 568.400 398.400 ;
        RECT 575.600 393.600 576.400 394.400 ;
        RECT 569.200 385.600 570.000 386.400 ;
        RECT 583.600 397.600 584.400 398.400 ;
        RECT 606.000 397.600 606.800 398.400 ;
        RECT 604.400 393.600 605.200 394.400 ;
        RECT 583.600 389.600 584.400 390.400 ;
        RECT 607.600 393.600 608.400 394.400 ;
        RECT 578.800 387.600 579.600 388.400 ;
        RECT 585.200 387.600 586.000 388.400 ;
        RECT 588.400 387.600 589.200 388.400 ;
        RECT 586.800 386.200 587.600 387.000 ;
        RECT 610.800 391.600 611.600 392.400 ;
        RECT 609.200 389.600 610.000 390.400 ;
        RECT 614.000 389.600 614.800 390.400 ;
        RECT 622.000 387.600 622.800 388.400 ;
        RECT 638.000 392.400 638.800 393.200 ;
        RECT 641.200 391.000 642.000 391.800 ;
        RECT 646.000 389.600 646.800 390.400 ;
        RECT 666.800 395.000 667.600 395.800 ;
        RECT 663.600 393.600 664.400 394.400 ;
        RECT 681.200 397.600 682.000 398.400 ;
        RECT 668.400 392.400 669.200 393.200 ;
        RECT 641.200 386.200 642.000 387.000 ;
        RECT 647.600 387.600 648.400 388.400 ;
        RECT 657.200 388.200 658.000 389.000 ;
        RECT 666.800 388.600 667.600 389.400 ;
        RECT 623.600 383.600 624.400 384.400 ;
        RECT 642.800 383.600 643.600 384.400 ;
        RECT 662.000 387.600 662.800 388.400 ;
        RECT 657.200 384.200 658.000 385.000 ;
        RECT 658.800 384.200 659.600 385.000 ;
        RECT 660.400 384.200 661.200 385.000 ;
        RECT 663.600 384.200 664.400 385.000 ;
        RECT 666.800 384.200 667.600 385.000 ;
        RECT 668.400 384.200 669.200 385.000 ;
        RECT 670.000 384.200 670.800 385.000 ;
        RECT 671.600 384.200 672.400 385.000 ;
        RECT 18.800 377.600 19.600 378.400 ;
        RECT 22.000 377.600 22.800 378.400 ;
        RECT 1.200 370.200 2.000 371.000 ;
        RECT 57.200 375.600 58.000 376.400 ;
        RECT 28.400 369.600 29.200 370.400 ;
        RECT 38.000 371.600 38.800 372.400 ;
        RECT 47.600 371.600 48.400 372.400 ;
        RECT 62.000 367.600 62.800 368.400 ;
        RECT 66.800 365.600 67.600 366.400 ;
        RECT 71.600 363.600 72.400 364.400 ;
        RECT 78.000 369.600 78.800 370.400 ;
        RECT 129.200 377.600 130.000 378.400 ;
        RECT 94.000 369.600 94.800 370.400 ;
        RECT 86.000 363.600 86.800 364.400 ;
        RECT 100.400 369.600 101.200 370.400 ;
        RECT 138.800 373.600 139.600 374.400 ;
        RECT 132.400 371.600 133.200 372.400 ;
        RECT 114.800 365.600 115.600 366.400 ;
        RECT 122.800 365.600 123.600 366.400 ;
        RECT 150.000 377.600 150.800 378.400 ;
        RECT 143.600 363.600 144.400 364.400 ;
        RECT 162.800 373.600 163.600 374.400 ;
        RECT 154.800 372.200 155.600 373.000 ;
        RECT 177.200 375.600 178.000 376.400 ;
        RECT 167.600 370.200 168.400 371.000 ;
        RECT 188.400 373.000 189.200 373.800 ;
        RECT 198.000 372.600 198.800 373.400 ;
        RECT 183.600 371.600 184.400 372.400 ;
        RECT 204.400 371.600 205.200 372.400 ;
        RECT 190.000 368.800 190.800 369.600 ;
        RECT 194.800 367.600 195.600 368.400 ;
        RECT 191.600 366.200 192.400 367.000 ;
        RECT 188.400 364.200 189.200 365.000 ;
        RECT 190.000 364.200 190.800 365.000 ;
        RECT 194.800 366.200 195.600 367.000 ;
        RECT 198.000 366.200 198.800 367.000 ;
        RECT 199.600 364.200 200.400 365.000 ;
        RECT 201.200 364.200 202.000 365.000 ;
        RECT 202.800 364.200 203.600 365.000 ;
        RECT 234.800 375.600 235.600 376.400 ;
        RECT 212.400 363.600 213.200 364.400 ;
        RECT 233.200 369.600 234.000 370.400 ;
        RECT 230.000 363.600 230.800 364.400 ;
        RECT 246.000 373.000 246.800 373.800 ;
        RECT 255.600 372.600 256.400 373.400 ;
        RECT 241.200 371.600 242.000 372.400 ;
        RECT 247.600 368.800 248.400 369.600 ;
        RECT 252.400 367.600 253.200 368.400 ;
        RECT 249.200 366.200 250.000 367.000 ;
        RECT 246.000 364.200 246.800 365.000 ;
        RECT 247.600 364.200 248.400 365.000 ;
        RECT 252.400 366.200 253.200 367.000 ;
        RECT 255.600 366.200 256.400 367.000 ;
        RECT 257.200 364.200 258.000 365.000 ;
        RECT 258.800 364.200 259.600 365.000 ;
        RECT 260.400 364.200 261.200 365.000 ;
        RECT 290.800 373.600 291.600 374.400 ;
        RECT 313.200 377.600 314.000 378.400 ;
        RECT 302.000 363.600 302.800 364.400 ;
        RECT 319.600 373.600 320.400 374.400 ;
        RECT 314.800 371.600 315.600 372.400 ;
        RECT 332.400 377.600 333.200 378.400 ;
        RECT 313.200 369.600 314.000 370.400 ;
        RECT 342.000 375.600 342.800 376.400 ;
        RECT 335.600 371.600 336.400 372.400 ;
        RECT 346.800 371.600 347.600 372.400 ;
        RECT 353.200 371.600 354.000 372.400 ;
        RECT 362.800 377.600 363.600 378.400 ;
        RECT 359.600 371.600 360.400 372.400 ;
        RECT 366.000 371.600 366.800 372.400 ;
        RECT 358.000 369.600 358.800 370.400 ;
        RECT 348.400 365.600 349.200 366.400 ;
        RECT 407.600 377.600 408.400 378.400 ;
        RECT 377.200 371.600 378.000 372.400 ;
        RECT 382.000 371.600 382.800 372.400 ;
        RECT 375.600 365.600 376.400 366.400 ;
        RECT 393.200 365.600 394.000 366.400 ;
        RECT 401.200 363.600 402.000 364.400 ;
        RECT 433.200 375.600 434.000 376.400 ;
        RECT 434.800 374.200 435.600 375.000 ;
        RECT 425.200 371.600 426.000 372.400 ;
        RECT 446.000 371.600 446.800 372.400 ;
        RECT 417.200 365.600 418.000 366.400 ;
        RECT 428.400 366.800 429.200 367.600 ;
        RECT 431.600 366.200 432.400 367.000 ;
        RECT 426.800 364.200 427.600 365.000 ;
        RECT 428.400 364.200 429.200 365.000 ;
        RECT 430.000 364.200 430.800 365.000 ;
        RECT 434.800 366.200 435.600 367.000 ;
        RECT 438.000 366.200 438.800 367.000 ;
        RECT 458.800 373.000 459.600 373.800 ;
        RECT 468.400 372.600 469.200 373.400 ;
        RECT 455.600 371.600 456.400 372.400 ;
        RECT 516.400 377.600 517.200 378.400 ;
        RECT 486.000 373.600 486.800 374.400 ;
        RECT 460.400 368.800 461.200 369.600 ;
        RECT 465.200 367.600 466.000 368.400 ;
        RECT 439.600 364.200 440.400 365.000 ;
        RECT 441.200 364.200 442.000 365.000 ;
        RECT 462.000 366.200 462.800 367.000 ;
        RECT 458.800 364.200 459.600 365.000 ;
        RECT 460.400 364.200 461.200 365.000 ;
        RECT 465.200 366.200 466.000 367.000 ;
        RECT 468.400 366.200 469.200 367.000 ;
        RECT 470.000 364.200 470.800 365.000 ;
        RECT 471.600 364.200 472.400 365.000 ;
        RECT 473.200 364.200 474.000 365.000 ;
        RECT 482.800 369.600 483.600 370.400 ;
        RECT 527.600 377.600 528.400 378.400 ;
        RECT 497.200 363.600 498.000 364.400 ;
        RECT 503.600 369.600 504.400 370.400 ;
        RECT 508.400 369.600 509.200 370.400 ;
        RECT 526.000 369.600 526.800 370.400 ;
        RECT 554.800 372.200 555.600 373.000 ;
        RECT 562.800 371.800 563.600 372.600 ;
        RECT 538.800 363.600 539.600 364.400 ;
        RECT 567.600 370.200 568.400 371.000 ;
        RECT 550.000 363.600 550.800 364.400 ;
        RECT 582.000 373.600 582.800 374.400 ;
        RECT 599.600 375.600 600.400 376.400 ;
        RECT 572.400 369.600 573.200 370.400 ;
        RECT 604.400 377.600 605.200 378.400 ;
        RECT 602.800 371.600 603.600 372.400 ;
        RECT 607.600 371.600 608.400 372.400 ;
        RECT 609.200 369.600 610.000 370.400 ;
        RECT 636.400 377.600 637.200 378.400 ;
        RECT 625.200 369.600 626.000 370.400 ;
        RECT 633.200 371.600 634.000 372.400 ;
        RECT 646.000 369.600 646.800 370.400 ;
        RECT 650.800 371.600 651.600 372.400 ;
        RECT 670.000 375.600 670.800 376.400 ;
        RECT 671.600 374.200 672.400 375.000 ;
        RECT 681.200 371.600 682.000 372.400 ;
        RECT 644.400 363.600 645.200 364.400 ;
        RECT 650.800 363.600 651.600 364.400 ;
        RECT 654.000 363.600 654.800 364.400 ;
        RECT 665.200 366.800 666.000 367.600 ;
        RECT 668.400 366.200 669.200 367.000 ;
        RECT 663.600 364.200 664.400 365.000 ;
        RECT 665.200 364.200 666.000 365.000 ;
        RECT 666.800 364.200 667.600 365.000 ;
        RECT 671.600 366.200 672.400 367.000 ;
        RECT 674.800 366.200 675.600 367.000 ;
        RECT 676.400 364.200 677.200 365.000 ;
        RECT 678.000 364.200 678.800 365.000 ;
        RECT 18.800 357.600 19.600 358.400 ;
        RECT 23.600 351.600 24.400 352.400 ;
        RECT 7.600 349.600 8.400 350.400 ;
        RECT 1.200 346.200 2.000 347.000 ;
        RECT 23.600 349.600 24.400 350.400 ;
        RECT 30.000 349.600 30.800 350.400 ;
        RECT 34.800 349.600 35.600 350.400 ;
        RECT 42.800 349.600 43.600 350.400 ;
        RECT 57.200 357.600 58.000 358.400 ;
        RECT 25.200 347.600 26.000 348.400 ;
        RECT 31.600 347.600 32.400 348.400 ;
        RECT 44.400 347.600 45.200 348.400 ;
        RECT 52.400 349.600 53.200 350.400 ;
        RECT 54.000 349.600 54.800 350.400 ;
        RECT 39.600 343.600 40.400 344.400 ;
        RECT 55.600 347.600 56.400 348.400 ;
        RECT 63.600 349.600 64.400 350.400 ;
        RECT 66.800 349.600 67.600 350.400 ;
        RECT 68.400 349.600 69.200 350.400 ;
        RECT 73.200 349.600 74.000 350.400 ;
        RECT 78.000 349.600 78.800 350.400 ;
        RECT 92.400 357.600 93.200 358.400 ;
        RECT 86.000 349.600 86.800 350.400 ;
        RECT 92.400 349.600 93.200 350.400 ;
        RECT 74.800 347.600 75.600 348.400 ;
        RECT 87.600 347.600 88.400 348.400 ;
        RECT 100.400 349.600 101.200 350.400 ;
        RECT 103.600 349.600 104.400 350.400 ;
        RECT 114.800 349.600 115.600 350.400 ;
        RECT 119.600 349.600 120.400 350.400 ;
        RECT 121.200 349.600 122.000 350.400 ;
        RECT 70.000 343.600 70.800 344.400 ;
        RECT 81.200 343.600 82.000 344.400 ;
        RECT 97.200 343.600 98.000 344.400 ;
        RECT 129.200 345.600 130.000 346.400 ;
        RECT 135.600 349.600 136.400 350.400 ;
        RECT 142.000 349.600 142.800 350.400 ;
        RECT 146.800 349.600 147.600 350.400 ;
        RECT 154.800 351.600 155.600 352.400 ;
        RECT 161.200 349.600 162.000 350.400 ;
        RECT 167.600 349.600 168.400 350.400 ;
        RECT 188.400 355.000 189.200 355.800 ;
        RECT 185.200 353.600 186.000 354.400 ;
        RECT 190.000 352.400 190.800 353.200 ;
        RECT 207.600 351.800 208.400 352.600 ;
        RECT 137.200 347.600 138.000 348.400 ;
        RECT 140.400 347.600 141.200 348.400 ;
        RECT 143.600 347.600 144.400 348.400 ;
        RECT 156.400 347.600 157.200 348.400 ;
        RECT 159.600 347.600 160.400 348.400 ;
        RECT 162.800 347.600 163.600 348.400 ;
        RECT 169.200 347.600 170.000 348.400 ;
        RECT 178.800 348.200 179.600 349.000 ;
        RECT 188.400 348.600 189.200 349.400 ;
        RECT 150.000 343.600 150.800 344.400 ;
        RECT 183.600 347.600 184.400 348.400 ;
        RECT 178.800 344.200 179.600 345.000 ;
        RECT 180.400 344.200 181.200 345.000 ;
        RECT 182.000 344.200 182.800 345.000 ;
        RECT 185.200 344.200 186.000 345.000 ;
        RECT 188.400 344.200 189.200 345.000 ;
        RECT 190.000 344.200 190.800 345.000 ;
        RECT 191.600 344.200 192.400 345.000 ;
        RECT 193.200 344.200 194.000 345.000 ;
        RECT 228.400 357.600 229.200 358.400 ;
        RECT 220.400 349.600 221.200 350.400 ;
        RECT 207.600 346.200 208.400 347.000 ;
        RECT 212.400 346.400 213.200 347.200 ;
        RECT 223.600 345.600 224.400 346.400 ;
        RECT 231.600 349.600 232.400 350.400 ;
        RECT 238.000 347.600 238.800 348.400 ;
        RECT 258.800 355.000 259.600 355.800 ;
        RECT 255.600 353.600 256.400 354.400 ;
        RECT 260.400 352.400 261.200 353.200 ;
        RECT 273.200 353.600 274.000 354.400 ;
        RECT 249.200 348.200 250.000 349.000 ;
        RECT 258.800 348.600 259.600 349.400 ;
        RECT 254.000 347.600 254.800 348.400 ;
        RECT 249.200 344.200 250.000 345.000 ;
        RECT 250.800 344.200 251.600 345.000 ;
        RECT 252.400 344.200 253.200 345.000 ;
        RECT 255.600 344.200 256.400 345.000 ;
        RECT 258.800 344.200 259.600 345.000 ;
        RECT 260.400 344.200 261.200 345.000 ;
        RECT 262.000 344.200 262.800 345.000 ;
        RECT 263.600 344.200 264.400 345.000 ;
        RECT 292.400 357.600 293.200 358.400 ;
        RECT 298.800 347.600 299.600 348.400 ;
        RECT 297.200 345.600 298.000 346.400 ;
        RECT 306.800 357.600 307.600 358.400 ;
        RECT 313.200 357.600 314.000 358.400 ;
        RECT 311.600 353.600 312.400 354.400 ;
        RECT 306.800 349.600 307.600 350.400 ;
        RECT 314.800 351.600 315.600 352.400 ;
        RECT 329.200 357.600 330.000 358.400 ;
        RECT 337.200 353.600 338.000 354.400 ;
        RECT 342.000 357.600 342.800 358.400 ;
        RECT 343.600 353.600 344.400 354.400 ;
        RECT 340.400 351.600 341.200 352.400 ;
        RECT 313.200 349.600 314.000 350.400 ;
        RECT 348.400 355.600 349.200 356.400 ;
        RECT 358.000 357.600 358.800 358.400 ;
        RECT 356.400 353.600 357.200 354.400 ;
        RECT 308.400 347.600 309.200 348.400 ;
        RECT 302.000 343.600 302.800 344.400 ;
        RECT 359.600 351.600 360.400 352.400 ;
        RECT 358.000 349.600 358.800 350.400 ;
        RECT 364.400 347.600 365.200 348.400 ;
        RECT 375.600 353.600 376.400 354.400 ;
        RECT 380.400 357.600 381.200 358.400 ;
        RECT 382.000 353.600 382.800 354.400 ;
        RECT 378.800 351.600 379.600 352.400 ;
        RECT 369.200 347.600 370.000 348.400 ;
        RECT 398.000 354.400 398.800 355.200 ;
        RECT 401.200 355.000 402.000 355.800 ;
        RECT 396.400 352.400 397.200 353.200 ;
        RECT 433.200 357.600 434.000 358.400 ;
        RECT 406.000 347.600 406.800 348.400 ;
        RECT 402.800 345.600 403.600 346.400 ;
        RECT 428.400 349.600 429.200 350.400 ;
        RECT 396.400 344.200 397.200 345.000 ;
        RECT 398.000 344.200 398.800 345.000 ;
        RECT 399.600 344.200 400.400 345.000 ;
        RECT 401.200 344.200 402.000 345.000 ;
        RECT 404.400 344.200 405.200 345.000 ;
        RECT 407.600 344.200 408.400 345.000 ;
        RECT 409.200 344.200 410.000 345.000 ;
        RECT 410.800 344.200 411.600 345.000 ;
        RECT 426.800 347.600 427.600 348.400 ;
        RECT 430.000 347.600 430.800 348.400 ;
        RECT 431.600 347.600 432.400 348.400 ;
        RECT 449.200 354.400 450.000 355.200 ;
        RECT 452.400 355.000 453.200 355.800 ;
        RECT 447.600 352.400 448.400 353.200 ;
        RECT 438.000 343.600 438.800 344.400 ;
        RECT 457.200 347.600 458.000 348.400 ;
        RECT 454.000 345.600 454.800 346.400 ;
        RECT 447.600 344.200 448.400 345.000 ;
        RECT 449.200 344.200 450.000 345.000 ;
        RECT 450.800 344.200 451.600 345.000 ;
        RECT 452.400 344.200 453.200 345.000 ;
        RECT 455.600 344.200 456.400 345.000 ;
        RECT 458.800 344.200 459.600 345.000 ;
        RECT 460.400 344.200 461.200 345.000 ;
        RECT 462.000 344.200 462.800 345.000 ;
        RECT 471.600 347.600 472.400 348.400 ;
        RECT 474.800 353.600 475.600 354.400 ;
        RECT 478.000 349.600 478.800 350.400 ;
        RECT 497.200 352.400 498.000 353.200 ;
        RECT 500.400 351.000 501.200 351.800 ;
        RECT 519.600 355.600 520.400 356.400 ;
        RECT 516.400 353.600 517.200 354.400 ;
        RECT 503.600 347.600 504.400 348.400 ;
        RECT 481.200 343.600 482.000 344.400 ;
        RECT 500.400 346.200 501.200 347.000 ;
        RECT 482.800 343.600 483.600 344.400 ;
        RECT 502.000 346.200 502.800 347.000 ;
        RECT 521.200 345.600 522.000 346.400 ;
        RECT 527.600 349.600 528.400 350.400 ;
        RECT 530.800 349.600 531.600 350.400 ;
        RECT 532.400 349.600 533.200 350.400 ;
        RECT 529.200 347.600 530.000 348.400 ;
        RECT 542.000 349.600 542.800 350.400 ;
        RECT 548.400 349.600 549.200 350.400 ;
        RECT 556.400 349.600 557.200 350.400 ;
        RECT 522.800 343.600 523.600 344.400 ;
        RECT 577.200 357.600 578.000 358.400 ;
        RECT 561.200 345.600 562.000 346.400 ;
        RECT 566.000 347.600 566.800 348.400 ;
        RECT 578.800 349.600 579.600 350.400 ;
        RECT 580.400 349.600 581.200 350.400 ;
        RECT 606.000 351.600 606.800 352.400 ;
        RECT 588.400 349.600 589.200 350.400 ;
        RECT 590.000 349.600 590.800 350.400 ;
        RECT 591.600 346.200 592.400 347.000 ;
        RECT 612.400 349.600 613.200 350.400 ;
        RECT 614.000 349.600 614.800 350.400 ;
        RECT 620.400 349.600 621.200 350.400 ;
        RECT 623.600 349.600 624.400 350.400 ;
        RECT 625.200 349.600 626.000 350.400 ;
        RECT 622.000 347.600 622.800 348.400 ;
        RECT 634.800 349.600 635.600 350.400 ;
        RECT 642.800 349.600 643.600 350.400 ;
        RECT 609.200 343.600 610.000 344.400 ;
        RECT 641.200 347.600 642.000 348.400 ;
        RECT 665.200 352.400 666.000 353.200 ;
        RECT 668.400 351.000 669.200 351.800 ;
        RECT 649.200 345.600 650.000 346.400 ;
        RECT 668.400 346.200 669.200 347.000 ;
        RECT 650.800 343.600 651.600 344.400 ;
        RECT 673.200 345.600 674.000 346.400 ;
        RECT 678.000 345.600 678.800 346.400 ;
        RECT 679.600 345.600 680.400 346.400 ;
        RECT 671.600 343.600 672.400 344.400 ;
        RECT 676.400 343.600 677.200 344.400 ;
        RECT 1.200 330.200 2.000 331.000 ;
        RECT 60.400 337.600 61.200 338.400 ;
        RECT 65.200 337.600 66.000 338.400 ;
        RECT 34.800 331.600 35.600 332.400 ;
        RECT 23.600 327.600 24.400 328.400 ;
        RECT 47.600 331.800 48.400 332.600 ;
        RECT 42.800 330.200 43.600 331.000 ;
        RECT 90.800 337.600 91.600 338.400 ;
        RECT 70.000 333.600 70.800 334.400 ;
        RECT 127.600 337.600 128.400 338.400 ;
        RECT 65.200 329.600 66.000 330.400 ;
        RECT 73.200 330.200 74.000 331.000 ;
        RECT 118.000 333.600 118.800 334.400 ;
        RECT 90.800 323.600 91.600 324.400 ;
        RECT 97.200 329.600 98.000 330.400 ;
        RECT 114.800 331.800 115.600 332.600 ;
        RECT 103.600 329.600 104.400 330.400 ;
        RECT 110.000 330.200 110.800 331.000 ;
        RECT 132.400 329.600 133.200 330.400 ;
        RECT 145.200 334.800 146.000 335.600 ;
        RECT 158.000 337.600 158.800 338.400 ;
        RECT 185.200 335.600 186.000 336.400 ;
        RECT 186.800 334.200 187.600 335.000 ;
        RECT 204.400 337.600 205.200 338.400 ;
        RECT 198.000 331.600 198.800 332.400 ;
        RECT 180.400 326.800 181.200 327.600 ;
        RECT 183.600 326.200 184.400 327.000 ;
        RECT 178.800 324.200 179.600 325.000 ;
        RECT 180.400 324.200 181.200 325.000 ;
        RECT 182.000 324.200 182.800 325.000 ;
        RECT 186.800 326.200 187.600 327.000 ;
        RECT 190.000 326.200 190.800 327.000 ;
        RECT 217.200 333.600 218.000 334.400 ;
        RECT 191.600 324.200 192.400 325.000 ;
        RECT 193.200 324.200 194.000 325.000 ;
        RECT 212.400 329.600 213.200 330.400 ;
        RECT 225.200 331.600 226.000 332.400 ;
        RECT 247.600 335.600 248.400 336.400 ;
        RECT 249.200 334.200 250.000 335.000 ;
        RECT 239.600 331.600 240.400 332.400 ;
        RECT 242.800 326.800 243.600 327.600 ;
        RECT 246.000 326.200 246.800 327.000 ;
        RECT 241.200 324.200 242.000 325.000 ;
        RECT 242.800 324.200 243.600 325.000 ;
        RECT 244.400 324.200 245.200 325.000 ;
        RECT 249.200 326.200 250.000 327.000 ;
        RECT 252.400 326.200 253.200 327.000 ;
        RECT 278.000 333.000 278.800 333.800 ;
        RECT 287.600 332.600 288.400 333.400 ;
        RECT 319.600 337.600 320.400 338.400 ;
        RECT 294.000 331.600 294.800 332.400 ;
        RECT 279.600 328.800 280.400 329.600 ;
        RECT 284.400 327.600 285.200 328.400 ;
        RECT 254.000 324.200 254.800 325.000 ;
        RECT 255.600 324.200 256.400 325.000 ;
        RECT 281.200 326.200 282.000 327.000 ;
        RECT 278.000 324.200 278.800 325.000 ;
        RECT 279.600 324.200 280.400 325.000 ;
        RECT 284.400 326.200 285.200 327.000 ;
        RECT 287.600 326.200 288.400 327.000 ;
        RECT 289.200 324.200 290.000 325.000 ;
        RECT 290.800 324.200 291.600 325.000 ;
        RECT 292.400 324.200 293.200 325.000 ;
        RECT 302.000 323.600 302.800 324.400 ;
        RECT 318.000 329.600 318.800 330.400 ;
        RECT 327.600 333.600 328.400 334.400 ;
        RECT 343.600 333.600 344.400 334.400 ;
        RECT 359.600 335.600 360.400 336.400 ;
        RECT 378.800 337.600 379.600 338.400 ;
        RECT 351.600 333.600 352.400 334.400 ;
        RECT 356.400 333.600 357.200 334.400 ;
        RECT 322.800 331.600 323.600 332.400 ;
        RECT 329.200 331.600 330.000 332.400 ;
        RECT 330.800 331.600 331.600 332.400 ;
        RECT 337.200 331.600 338.000 332.400 ;
        RECT 338.800 331.600 339.600 332.400 ;
        RECT 345.200 331.600 346.000 332.400 ;
        RECT 346.800 331.600 347.600 332.400 ;
        RECT 353.200 331.600 354.000 332.400 ;
        RECT 361.200 331.600 362.000 332.400 ;
        RECT 324.400 327.600 325.200 328.400 ;
        RECT 340.400 323.600 341.200 324.400 ;
        RECT 372.400 333.600 373.200 334.400 ;
        RECT 367.600 331.600 368.400 332.400 ;
        RECT 374.000 331.600 374.800 332.400 ;
        RECT 366.000 329.600 366.800 330.400 ;
        RECT 369.200 325.600 370.000 326.400 ;
        RECT 378.800 329.600 379.600 330.400 ;
        RECT 380.400 329.600 381.200 330.400 ;
        RECT 390.000 333.600 390.800 334.400 ;
        RECT 391.600 331.600 392.400 332.400 ;
        RECT 393.200 329.600 394.000 330.400 ;
        RECT 399.600 333.600 400.400 334.400 ;
        RECT 407.600 333.600 408.400 334.400 ;
        RECT 404.400 331.600 405.200 332.400 ;
        RECT 415.600 329.600 416.400 330.400 ;
        RECT 426.800 329.600 427.600 330.400 ;
        RECT 452.400 335.600 453.200 336.400 ;
        RECT 454.000 334.200 454.800 335.000 ;
        RECT 463.600 331.600 464.400 332.400 ;
        RECT 433.200 329.600 434.000 330.400 ;
        RECT 436.400 329.600 437.200 330.400 ;
        RECT 447.600 326.800 448.400 327.600 ;
        RECT 450.800 326.200 451.600 327.000 ;
        RECT 446.000 324.200 446.800 325.000 ;
        RECT 447.600 324.200 448.400 325.000 ;
        RECT 449.200 324.200 450.000 325.000 ;
        RECT 454.000 326.200 454.800 327.000 ;
        RECT 457.200 326.200 458.000 327.000 ;
        RECT 458.800 324.200 459.600 325.000 ;
        RECT 460.400 324.200 461.200 325.000 ;
        RECT 490.800 337.600 491.600 338.400 ;
        RECT 510.000 337.600 510.800 338.400 ;
        RECT 478.000 329.600 478.800 330.400 ;
        RECT 487.600 329.600 488.400 330.400 ;
        RECT 502.000 333.600 502.800 334.400 ;
        RECT 519.600 335.600 520.400 336.400 ;
        RECT 524.400 333.600 525.200 334.400 ;
        RECT 545.200 333.600 546.000 334.400 ;
        RECT 559.600 337.600 560.400 338.400 ;
        RECT 556.400 333.600 557.200 334.400 ;
        RECT 526.000 329.600 526.800 330.400 ;
        RECT 535.600 323.600 536.400 324.400 ;
        RECT 545.200 329.600 546.000 330.400 ;
        RECT 569.200 333.600 570.000 334.400 ;
        RECT 609.200 337.600 610.000 338.400 ;
        RECT 564.400 332.200 565.200 333.000 ;
        RECT 558.000 329.600 558.800 330.400 ;
        RECT 572.400 331.800 573.200 332.600 ;
        RECT 586.800 331.600 587.600 332.400 ;
        RECT 577.200 330.200 578.000 331.000 ;
        RECT 588.400 329.600 589.200 330.400 ;
        RECT 625.200 333.600 626.000 334.400 ;
        RECT 634.800 335.600 635.600 336.400 ;
        RECT 642.800 337.600 643.600 338.400 ;
        RECT 631.600 331.600 632.400 332.400 ;
        RECT 687.600 337.600 688.400 338.400 ;
        RECT 644.400 331.600 645.200 332.400 ;
        RECT 671.600 333.600 672.400 334.400 ;
        RECT 652.400 329.600 653.200 330.400 ;
        RECT 674.800 331.800 675.600 332.600 ;
        RECT 670.000 330.200 670.800 331.000 ;
        RECT 666.800 327.600 667.600 328.400 ;
        RECT 18.800 315.000 19.600 315.800 ;
        RECT 15.600 313.600 16.400 314.400 ;
        RECT 20.400 312.400 21.200 313.200 ;
        RECT 33.200 313.600 34.000 314.400 ;
        RECT 25.200 309.600 26.000 310.400 ;
        RECT 9.200 308.200 10.000 309.000 ;
        RECT 18.800 308.600 19.600 309.400 ;
        RECT 14.000 307.600 14.800 308.400 ;
        RECT 9.200 304.200 10.000 305.000 ;
        RECT 10.800 304.200 11.600 305.000 ;
        RECT 12.400 304.200 13.200 305.000 ;
        RECT 15.600 304.200 16.400 305.000 ;
        RECT 18.800 304.200 19.600 305.000 ;
        RECT 20.400 304.200 21.200 305.000 ;
        RECT 22.000 304.200 22.800 305.000 ;
        RECT 23.600 304.200 24.400 305.000 ;
        RECT 46.000 309.600 46.800 310.400 ;
        RECT 50.800 305.600 51.600 306.400 ;
        RECT 55.600 307.600 56.400 308.400 ;
        RECT 57.200 307.600 58.000 308.400 ;
        RECT 79.600 315.000 80.400 315.800 ;
        RECT 76.400 313.600 77.200 314.400 ;
        RECT 94.000 317.600 94.800 318.400 ;
        RECT 81.200 312.400 82.000 313.200 ;
        RECT 97.200 317.600 98.000 318.400 ;
        RECT 86.000 309.600 86.800 310.400 ;
        RECT 70.000 308.200 70.800 309.000 ;
        RECT 79.600 308.600 80.400 309.400 ;
        RECT 54.000 303.600 54.800 304.400 ;
        RECT 74.800 307.600 75.600 308.400 ;
        RECT 70.000 304.200 70.800 305.000 ;
        RECT 71.600 304.200 72.400 305.000 ;
        RECT 73.200 304.200 74.000 305.000 ;
        RECT 76.400 304.200 77.200 305.000 ;
        RECT 79.600 304.200 80.400 305.000 ;
        RECT 81.200 304.200 82.000 305.000 ;
        RECT 82.800 304.200 83.600 305.000 ;
        RECT 84.400 304.200 85.200 305.000 ;
        RECT 102.000 317.600 102.800 318.400 ;
        RECT 103.600 313.600 104.400 314.400 ;
        RECT 100.400 311.600 101.200 312.400 ;
        RECT 129.200 315.000 130.000 315.800 ;
        RECT 126.000 313.600 126.800 314.400 ;
        RECT 130.800 312.400 131.600 313.200 ;
        RECT 154.800 317.600 155.600 318.400 ;
        RECT 135.600 309.600 136.400 310.400 ;
        RECT 119.600 308.200 120.400 309.000 ;
        RECT 129.200 308.600 130.000 309.400 ;
        RECT 98.800 305.600 99.600 306.400 ;
        RECT 124.400 307.600 125.200 308.400 ;
        RECT 119.600 304.200 120.400 305.000 ;
        RECT 121.200 304.200 122.000 305.000 ;
        RECT 122.800 304.200 123.600 305.000 ;
        RECT 126.000 304.200 126.800 305.000 ;
        RECT 129.200 304.200 130.000 305.000 ;
        RECT 130.800 304.200 131.600 305.000 ;
        RECT 132.400 304.200 133.200 305.000 ;
        RECT 134.000 304.200 134.800 305.000 ;
        RECT 150.000 309.600 150.800 310.400 ;
        RECT 151.600 307.600 152.400 308.400 ;
        RECT 159.600 317.600 160.400 318.400 ;
        RECT 156.400 307.600 157.200 308.400 ;
        RECT 146.800 303.600 147.600 304.400 ;
        RECT 158.000 305.600 158.800 306.400 ;
        RECT 169.200 315.600 170.000 316.400 ;
        RECT 180.400 314.400 181.200 315.200 ;
        RECT 183.600 315.000 184.400 315.800 ;
        RECT 178.800 312.400 179.600 313.200 ;
        RECT 166.000 309.600 166.800 310.400 ;
        RECT 162.800 303.600 163.600 304.400 ;
        RECT 177.200 309.600 178.000 310.400 ;
        RECT 188.400 307.600 189.200 308.400 ;
        RECT 185.200 305.600 186.000 306.400 ;
        RECT 178.800 304.200 179.600 305.000 ;
        RECT 180.400 304.200 181.200 305.000 ;
        RECT 182.000 304.200 182.800 305.000 ;
        RECT 183.600 304.200 184.400 305.000 ;
        RECT 186.800 304.200 187.600 305.000 ;
        RECT 190.000 304.200 190.800 305.000 ;
        RECT 191.600 304.200 192.400 305.000 ;
        RECT 193.200 304.200 194.000 305.000 ;
        RECT 202.800 307.600 203.600 308.400 ;
        RECT 215.600 309.600 216.400 310.400 ;
        RECT 217.200 307.600 218.000 308.400 ;
        RECT 222.000 309.600 222.800 310.400 ;
        RECT 218.800 303.600 219.600 304.400 ;
        RECT 234.800 317.600 235.600 318.400 ;
        RECT 231.600 303.600 232.400 304.400 ;
        RECT 244.400 309.600 245.200 310.400 ;
        RECT 271.600 315.000 272.400 315.800 ;
        RECT 268.400 313.600 269.200 314.400 ;
        RECT 273.200 312.400 274.000 313.200 ;
        RECT 286.000 313.600 286.800 314.400 ;
        RECT 290.800 317.600 291.600 318.400 ;
        RECT 241.200 307.600 242.000 308.400 ;
        RECT 246.000 307.600 246.800 308.400 ;
        RECT 262.000 308.200 262.800 309.000 ;
        RECT 271.600 308.600 272.400 309.400 ;
        RECT 266.800 307.600 267.600 308.400 ;
        RECT 262.000 304.200 262.800 305.000 ;
        RECT 263.600 304.200 264.400 305.000 ;
        RECT 265.200 304.200 266.000 305.000 ;
        RECT 268.400 304.200 269.200 305.000 ;
        RECT 271.600 304.200 272.400 305.000 ;
        RECT 273.200 304.200 274.000 305.000 ;
        RECT 274.800 304.200 275.600 305.000 ;
        RECT 276.400 304.200 277.200 305.000 ;
        RECT 295.600 317.600 296.400 318.400 ;
        RECT 300.400 309.600 301.200 310.400 ;
        RECT 297.200 307.600 298.000 308.400 ;
        RECT 313.200 317.600 314.000 318.400 ;
        RECT 321.200 315.600 322.000 316.400 ;
        RECT 314.800 313.600 315.600 314.400 ;
        RECT 308.400 307.600 309.200 308.400 ;
        RECT 306.800 305.600 307.600 306.400 ;
        RECT 318.000 311.600 318.800 312.400 ;
        RECT 316.400 309.600 317.200 310.400 ;
        RECT 334.000 313.600 334.800 314.400 ;
        RECT 322.800 307.600 323.600 308.400 ;
        RECT 330.800 311.600 331.600 312.400 ;
        RECT 342.000 309.600 342.800 310.400 ;
        RECT 343.600 307.600 344.400 308.400 ;
        RECT 369.200 317.600 370.000 318.400 ;
        RECT 358.000 309.600 358.800 310.400 ;
        RECT 362.800 309.600 363.600 310.400 ;
        RECT 380.400 314.400 381.200 315.200 ;
        RECT 383.600 315.000 384.400 315.800 ;
        RECT 378.800 312.400 379.600 313.200 ;
        RECT 345.200 303.600 346.000 304.400 ;
        RECT 358.000 305.600 358.800 306.400 ;
        RECT 388.400 307.600 389.200 308.400 ;
        RECT 385.200 305.600 386.000 306.400 ;
        RECT 378.800 304.200 379.600 305.000 ;
        RECT 380.400 304.200 381.200 305.000 ;
        RECT 382.000 304.200 382.800 305.000 ;
        RECT 383.600 304.200 384.400 305.000 ;
        RECT 386.800 304.200 387.600 305.000 ;
        RECT 390.000 304.200 390.800 305.000 ;
        RECT 391.600 304.200 392.400 305.000 ;
        RECT 393.200 304.200 394.000 305.000 ;
        RECT 425.200 315.000 426.000 315.800 ;
        RECT 422.000 313.600 422.800 314.400 ;
        RECT 439.600 317.600 440.400 318.400 ;
        RECT 426.800 312.400 427.600 313.200 ;
        RECT 431.600 309.600 432.400 310.400 ;
        RECT 415.600 308.200 416.400 309.000 ;
        RECT 425.200 308.600 426.000 309.400 ;
        RECT 420.400 307.600 421.200 308.400 ;
        RECT 415.600 304.200 416.400 305.000 ;
        RECT 417.200 304.200 418.000 305.000 ;
        RECT 418.800 304.200 419.600 305.000 ;
        RECT 422.000 304.200 422.800 305.000 ;
        RECT 425.200 304.200 426.000 305.000 ;
        RECT 426.800 304.200 427.600 305.000 ;
        RECT 428.400 304.200 429.200 305.000 ;
        RECT 430.000 304.200 430.800 305.000 ;
        RECT 466.800 317.600 467.600 318.400 ;
        RECT 452.400 309.600 453.200 310.400 ;
        RECT 444.400 307.600 445.200 308.400 ;
        RECT 447.600 307.600 448.400 308.400 ;
        RECT 439.600 303.600 440.400 304.400 ;
        RECT 446.000 306.200 446.800 307.000 ;
        RECT 465.200 305.600 466.000 306.400 ;
        RECT 470.000 309.600 470.800 310.400 ;
        RECT 481.200 309.600 482.000 310.400 ;
        RECT 482.800 309.600 483.600 310.400 ;
        RECT 486.000 309.600 486.800 310.400 ;
        RECT 505.200 317.600 506.000 318.400 ;
        RECT 494.000 309.600 494.800 310.400 ;
        RECT 500.400 309.600 501.200 310.400 ;
        RECT 479.600 305.600 480.400 306.400 ;
        RECT 495.600 307.600 496.400 308.400 ;
        RECT 498.800 307.600 499.600 308.400 ;
        RECT 502.000 307.600 502.800 308.400 ;
        RECT 503.600 305.600 504.400 306.400 ;
        RECT 516.400 313.600 517.200 314.400 ;
        RECT 511.600 307.600 512.400 308.400 ;
        RECT 529.200 309.600 530.000 310.400 ;
        RECT 532.400 309.600 533.200 310.400 ;
        RECT 546.800 317.600 547.600 318.400 ;
        RECT 553.200 317.600 554.000 318.400 ;
        RECT 538.800 309.600 539.600 310.400 ;
        RECT 526.000 303.600 526.800 304.400 ;
        RECT 553.200 309.600 554.000 310.400 ;
        RECT 558.000 309.600 558.800 310.400 ;
        RECT 554.800 307.600 555.600 308.400 ;
        RECT 559.600 307.600 560.400 308.400 ;
        RECT 594.800 313.600 595.600 314.400 ;
        RECT 583.600 309.600 584.400 310.400 ;
        RECT 578.800 307.600 579.600 308.400 ;
        RECT 570.800 305.600 571.600 306.400 ;
        RECT 577.200 306.200 578.000 307.000 ;
        RECT 598.000 309.600 598.800 310.400 ;
        RECT 606.000 309.600 606.800 310.400 ;
        RECT 609.200 309.600 610.000 310.400 ;
        RECT 610.800 309.600 611.600 310.400 ;
        RECT 607.600 307.600 608.400 308.400 ;
        RECT 602.800 303.600 603.600 304.400 ;
        RECT 633.200 317.600 634.000 318.400 ;
        RECT 625.200 307.600 626.000 308.400 ;
        RECT 633.200 309.600 634.000 310.400 ;
        RECT 634.800 307.600 635.600 308.400 ;
        RECT 642.800 309.600 643.600 310.400 ;
        RECT 639.600 307.600 640.400 308.400 ;
        RECT 622.000 303.600 622.800 304.400 ;
        RECT 641.200 305.600 642.000 306.400 ;
        RECT 652.400 309.600 653.200 310.400 ;
        RECT 654.000 309.600 654.800 310.400 ;
        RECT 657.200 309.600 658.000 310.400 ;
        RECT 686.000 313.600 686.800 314.400 ;
        RECT 665.200 309.600 666.000 310.400 ;
        RECT 644.400 305.600 645.200 306.400 ;
        RECT 650.800 305.600 651.600 306.400 ;
        RECT 666.800 307.600 667.600 308.400 ;
        RECT 668.400 306.200 669.200 307.000 ;
        RECT 23.600 293.600 24.400 294.400 ;
        RECT 49.200 297.600 50.000 298.400 ;
        RECT 55.600 297.600 56.400 298.400 ;
        RECT 33.200 289.600 34.000 290.400 ;
        RECT 38.000 283.600 38.800 284.400 ;
        RECT 47.600 289.600 48.400 290.400 ;
        RECT 70.000 293.000 70.800 293.800 ;
        RECT 79.600 292.600 80.400 293.400 ;
        RECT 110.000 297.600 110.800 298.400 ;
        RECT 86.000 291.600 86.800 292.400 ;
        RECT 71.600 288.800 72.400 289.600 ;
        RECT 76.400 287.600 77.200 288.400 ;
        RECT 73.200 286.200 74.000 287.000 ;
        RECT 70.000 284.200 70.800 285.000 ;
        RECT 71.600 284.200 72.400 285.000 ;
        RECT 76.400 286.200 77.200 287.000 ;
        RECT 79.600 286.200 80.400 287.000 ;
        RECT 81.200 284.200 82.000 285.000 ;
        RECT 82.800 284.200 83.600 285.000 ;
        RECT 84.400 284.200 85.200 285.000 ;
        RECT 94.000 289.600 94.800 290.400 ;
        RECT 97.200 289.600 98.000 290.400 ;
        RECT 108.400 289.600 109.200 290.400 ;
        RECT 126.000 293.000 126.800 293.800 ;
        RECT 135.600 292.600 136.400 293.400 ;
        RECT 142.000 291.600 142.800 292.400 ;
        RECT 127.600 288.800 128.400 289.600 ;
        RECT 132.400 287.600 133.200 288.400 ;
        RECT 129.200 286.200 130.000 287.000 ;
        RECT 126.000 284.200 126.800 285.000 ;
        RECT 127.600 284.200 128.400 285.000 ;
        RECT 132.400 286.200 133.200 287.000 ;
        RECT 135.600 286.200 136.400 287.000 ;
        RECT 137.200 284.200 138.000 285.000 ;
        RECT 138.800 284.200 139.600 285.000 ;
        RECT 140.400 284.200 141.200 285.000 ;
        RECT 153.200 289.600 154.000 290.400 ;
        RECT 150.000 287.600 150.800 288.400 ;
        RECT 172.400 293.000 173.200 293.800 ;
        RECT 182.000 292.600 182.800 293.400 ;
        RECT 170.800 291.600 171.600 292.400 ;
        RECT 202.800 293.600 203.600 294.400 ;
        RECT 174.000 288.800 174.800 289.600 ;
        RECT 178.800 287.600 179.600 288.400 ;
        RECT 175.600 286.200 176.400 287.000 ;
        RECT 172.400 284.200 173.200 285.000 ;
        RECT 174.000 284.200 174.800 285.000 ;
        RECT 178.800 286.200 179.600 287.000 ;
        RECT 182.000 286.200 182.800 287.000 ;
        RECT 183.600 284.200 184.400 285.000 ;
        RECT 185.200 284.200 186.000 285.000 ;
        RECT 186.800 284.200 187.600 285.000 ;
        RECT 196.400 289.600 197.200 290.400 ;
        RECT 214.000 293.000 214.800 293.800 ;
        RECT 204.400 289.600 205.200 290.400 ;
        RECT 223.600 292.600 224.400 293.400 ;
        RECT 218.800 291.600 219.600 292.400 ;
        RECT 215.600 288.800 216.400 289.600 ;
        RECT 220.400 287.600 221.200 288.400 ;
        RECT 217.200 286.200 218.000 287.000 ;
        RECT 214.000 284.200 214.800 285.000 ;
        RECT 215.600 284.200 216.400 285.000 ;
        RECT 220.400 286.200 221.200 287.000 ;
        RECT 223.600 286.200 224.400 287.000 ;
        RECT 225.200 284.200 226.000 285.000 ;
        RECT 226.800 284.200 227.600 285.000 ;
        RECT 228.400 284.200 229.200 285.000 ;
        RECT 250.800 295.600 251.600 296.400 ;
        RECT 242.800 283.600 243.600 284.400 ;
        RECT 247.600 289.600 248.400 290.400 ;
        RECT 266.800 293.000 267.600 293.800 ;
        RECT 252.400 289.600 253.200 290.400 ;
        RECT 276.400 292.600 277.200 293.400 ;
        RECT 290.800 297.600 291.600 298.400 ;
        RECT 282.800 291.600 283.600 292.400 ;
        RECT 268.400 288.800 269.200 289.600 ;
        RECT 273.200 287.600 274.000 288.400 ;
        RECT 270.000 286.200 270.800 287.000 ;
        RECT 266.800 284.200 267.600 285.000 ;
        RECT 268.400 284.200 269.200 285.000 ;
        RECT 273.200 286.200 274.000 287.000 ;
        RECT 276.400 286.200 277.200 287.000 ;
        RECT 278.000 284.200 278.800 285.000 ;
        RECT 279.600 284.200 280.400 285.000 ;
        RECT 281.200 284.200 282.000 285.000 ;
        RECT 330.800 297.600 331.600 298.400 ;
        RECT 308.400 291.600 309.200 292.400 ;
        RECT 314.800 291.600 315.600 292.400 ;
        RECT 321.200 291.600 322.000 292.400 ;
        RECT 295.600 283.600 296.400 284.400 ;
        RECT 324.400 289.600 325.200 290.400 ;
        RECT 308.400 283.600 309.200 284.400 ;
        RECT 314.800 283.600 315.600 284.400 ;
        RECT 321.200 285.600 322.000 286.400 ;
        RECT 359.600 295.600 360.400 296.400 ;
        RECT 369.200 297.600 370.000 298.400 ;
        RECT 364.400 295.600 365.200 296.400 ;
        RECT 345.200 291.600 346.000 292.400 ;
        RECT 356.400 291.600 357.200 292.400 ;
        RECT 326.000 283.600 326.800 284.400 ;
        RECT 337.200 283.600 338.000 284.400 ;
        RECT 350.000 283.600 350.800 284.400 ;
        RECT 385.200 295.600 386.000 296.400 ;
        RECT 386.800 294.200 387.600 295.000 ;
        RECT 407.600 297.600 408.400 298.400 ;
        RECT 394.800 291.600 395.600 292.400 ;
        RECT 380.400 286.800 381.200 287.600 ;
        RECT 383.600 286.200 384.400 287.000 ;
        RECT 378.800 284.200 379.600 285.000 ;
        RECT 380.400 284.200 381.200 285.000 ;
        RECT 382.000 284.200 382.800 285.000 ;
        RECT 386.800 286.200 387.600 287.000 ;
        RECT 390.000 286.200 390.800 287.000 ;
        RECT 391.600 284.200 392.400 285.000 ;
        RECT 393.200 284.200 394.000 285.000 ;
        RECT 428.400 293.000 429.200 293.800 ;
        RECT 438.000 292.600 438.800 293.400 ;
        RECT 452.400 297.600 453.200 298.400 ;
        RECT 426.800 291.600 427.600 292.400 ;
        RECT 433.200 291.600 434.000 292.400 ;
        RECT 430.000 288.800 430.800 289.600 ;
        RECT 434.800 287.600 435.600 288.400 ;
        RECT 431.600 286.200 432.400 287.000 ;
        RECT 428.400 284.200 429.200 285.000 ;
        RECT 430.000 284.200 430.800 285.000 ;
        RECT 434.800 286.200 435.600 287.000 ;
        RECT 438.000 286.200 438.800 287.000 ;
        RECT 439.600 284.200 440.400 285.000 ;
        RECT 441.200 284.200 442.000 285.000 ;
        RECT 442.800 284.200 443.600 285.000 ;
        RECT 476.400 295.600 477.200 296.400 ;
        RECT 487.600 297.600 488.400 298.400 ;
        RECT 473.200 291.600 474.000 292.400 ;
        RECT 470.000 289.600 470.800 290.400 ;
        RECT 486.000 293.600 486.800 294.400 ;
        RECT 508.400 297.600 509.200 298.400 ;
        RECT 500.400 293.600 501.200 294.400 ;
        RECT 492.400 292.200 493.200 293.000 ;
        RECT 486.000 289.600 486.800 290.400 ;
        RECT 505.200 290.200 506.000 291.000 ;
        RECT 511.600 291.600 512.400 292.400 ;
        RECT 542.000 297.600 542.800 298.400 ;
        RECT 514.800 283.600 515.600 284.400 ;
        RECT 530.800 289.600 531.600 290.400 ;
        RECT 538.800 291.600 539.600 292.400 ;
        RECT 558.000 290.200 558.800 291.000 ;
        RECT 554.800 283.600 555.600 284.400 ;
        RECT 614.000 297.600 614.800 298.400 ;
        RECT 588.400 291.600 589.200 292.400 ;
        RECT 586.800 287.600 587.600 288.400 ;
        RECT 598.000 291.600 598.800 292.400 ;
        RECT 631.600 295.600 632.400 296.400 ;
        RECT 639.600 297.600 640.400 298.400 ;
        RECT 626.800 289.600 627.600 290.400 ;
        RECT 649.200 297.600 650.000 298.400 ;
        RECT 650.800 297.600 651.600 298.400 ;
        RECT 641.200 291.600 642.000 292.400 ;
        RECT 681.200 297.600 682.000 298.400 ;
        RECT 666.800 293.600 667.600 294.400 ;
        RECT 670.000 293.600 670.800 294.400 ;
        RECT 655.600 292.200 656.400 293.000 ;
        RECT 668.400 290.200 669.200 291.000 ;
        RECT 18.800 275.000 19.600 275.800 ;
        RECT 15.600 273.600 16.400 274.400 ;
        RECT 33.200 277.600 34.000 278.400 ;
        RECT 20.400 272.400 21.200 273.200 ;
        RECT 25.200 269.600 26.000 270.400 ;
        RECT 9.200 268.200 10.000 269.000 ;
        RECT 18.800 268.600 19.600 269.400 ;
        RECT 14.000 267.600 14.800 268.400 ;
        RECT 9.200 264.200 10.000 265.000 ;
        RECT 10.800 264.200 11.600 265.000 ;
        RECT 12.400 264.200 13.200 265.000 ;
        RECT 15.600 264.200 16.400 265.000 ;
        RECT 18.800 264.200 19.600 265.000 ;
        RECT 20.400 264.200 21.200 265.000 ;
        RECT 22.000 264.200 22.800 265.000 ;
        RECT 23.600 264.200 24.400 265.000 ;
        RECT 54.000 269.600 54.800 270.400 ;
        RECT 68.400 277.600 69.200 278.400 ;
        RECT 55.600 267.600 56.400 268.400 ;
        RECT 50.800 263.600 51.600 264.400 ;
        RECT 57.200 265.600 58.000 266.400 ;
        RECT 79.600 274.400 80.400 275.200 ;
        RECT 82.800 275.000 83.600 275.800 ;
        RECT 102.000 277.600 102.800 278.400 ;
        RECT 78.000 272.400 78.800 273.200 ;
        RECT 76.400 269.600 77.200 270.400 ;
        RECT 65.200 263.600 66.000 264.400 ;
        RECT 87.600 267.600 88.400 268.400 ;
        RECT 84.400 265.600 85.200 266.400 ;
        RECT 78.000 264.200 78.800 265.000 ;
        RECT 79.600 264.200 80.400 265.000 ;
        RECT 81.200 264.200 82.000 265.000 ;
        RECT 82.800 264.200 83.600 265.000 ;
        RECT 86.000 264.200 86.800 265.000 ;
        RECT 89.200 264.200 90.000 265.000 ;
        RECT 90.800 264.200 91.600 265.000 ;
        RECT 92.400 264.200 93.200 265.000 ;
        RECT 105.200 277.600 106.000 278.400 ;
        RECT 103.600 265.600 104.400 266.400 ;
        RECT 119.600 277.600 120.400 278.400 ;
        RECT 132.400 277.600 133.200 278.400 ;
        RECT 111.600 267.600 112.400 268.400 ;
        RECT 106.800 265.600 107.600 266.400 ;
        RECT 137.200 273.600 138.000 274.400 ;
        RECT 148.400 274.400 149.200 275.200 ;
        RECT 151.600 275.000 152.400 275.800 ;
        RECT 146.800 272.400 147.600 273.200 ;
        RECT 134.000 265.600 134.800 266.400 ;
        RECT 156.400 267.600 157.200 268.400 ;
        RECT 153.200 265.600 154.000 266.400 ;
        RECT 146.800 264.200 147.600 265.000 ;
        RECT 148.400 264.200 149.200 265.000 ;
        RECT 150.000 264.200 150.800 265.000 ;
        RECT 151.600 264.200 152.400 265.000 ;
        RECT 154.800 264.200 155.600 265.000 ;
        RECT 158.000 264.200 158.800 265.000 ;
        RECT 159.600 264.200 160.400 265.000 ;
        RECT 161.200 264.200 162.000 265.000 ;
        RECT 190.000 277.600 190.800 278.400 ;
        RECT 178.800 269.600 179.600 270.400 ;
        RECT 180.400 267.600 181.200 268.400 ;
        RECT 201.200 274.400 202.000 275.200 ;
        RECT 204.400 275.000 205.200 275.800 ;
        RECT 199.600 272.400 200.400 273.200 ;
        RECT 183.600 263.600 184.400 264.400 ;
        RECT 230.000 277.600 230.800 278.400 ;
        RECT 209.200 267.600 210.000 268.400 ;
        RECT 206.000 265.600 206.800 266.400 ;
        RECT 199.600 264.200 200.400 265.000 ;
        RECT 201.200 264.200 202.000 265.000 ;
        RECT 202.800 264.200 203.600 265.000 ;
        RECT 204.400 264.200 205.200 265.000 ;
        RECT 207.600 264.200 208.400 265.000 ;
        RECT 210.800 264.200 211.600 265.000 ;
        RECT 212.400 264.200 213.200 265.000 ;
        RECT 214.000 264.200 214.800 265.000 ;
        RECT 241.200 274.400 242.000 275.200 ;
        RECT 244.400 275.000 245.200 275.800 ;
        RECT 239.600 272.400 240.400 273.200 ;
        RECT 238.000 269.600 238.800 270.400 ;
        RECT 230.000 263.600 230.800 264.400 ;
        RECT 276.400 273.600 277.200 274.400 ;
        RECT 249.200 267.600 250.000 268.400 ;
        RECT 246.000 265.600 246.800 266.400 ;
        RECT 239.600 264.200 240.400 265.000 ;
        RECT 241.200 264.200 242.000 265.000 ;
        RECT 242.800 264.200 243.600 265.000 ;
        RECT 244.400 264.200 245.200 265.000 ;
        RECT 247.600 264.200 248.400 265.000 ;
        RECT 250.800 264.200 251.600 265.000 ;
        RECT 252.400 264.200 253.200 265.000 ;
        RECT 254.000 264.200 254.800 265.000 ;
        RECT 284.400 271.600 285.200 272.400 ;
        RECT 278.000 269.600 278.800 270.400 ;
        RECT 284.400 269.600 285.200 270.400 ;
        RECT 311.600 275.000 312.400 275.800 ;
        RECT 308.400 273.600 309.200 274.400 ;
        RECT 313.200 272.400 314.000 273.200 ;
        RECT 286.000 267.600 286.800 268.400 ;
        RECT 302.000 268.200 302.800 269.000 ;
        RECT 311.600 268.600 312.400 269.400 ;
        RECT 306.800 267.600 307.600 268.400 ;
        RECT 326.200 267.600 327.000 268.400 ;
        RECT 302.000 264.200 302.800 265.000 ;
        RECT 303.600 264.200 304.400 265.000 ;
        RECT 305.200 264.200 306.000 265.000 ;
        RECT 308.400 264.200 309.200 265.000 ;
        RECT 311.600 264.200 312.400 265.000 ;
        RECT 313.200 264.200 314.000 265.000 ;
        RECT 314.800 264.200 315.600 265.000 ;
        RECT 316.400 264.200 317.200 265.000 ;
        RECT 334.000 275.600 334.800 276.400 ;
        RECT 332.400 263.600 333.200 264.400 ;
        RECT 335.600 267.600 336.400 268.400 ;
        RECT 350.000 269.600 350.800 270.400 ;
        RECT 358.000 269.600 358.800 270.400 ;
        RECT 346.800 263.600 347.600 264.400 ;
        RECT 354.800 265.600 355.600 266.400 ;
        RECT 370.800 265.600 371.600 266.400 ;
        RECT 378.800 277.600 379.600 278.400 ;
        RECT 377.200 271.600 378.000 272.400 ;
        RECT 394.800 277.600 395.600 278.400 ;
        RECT 406.000 273.600 406.800 274.400 ;
        RECT 388.400 269.600 389.200 270.400 ;
        RECT 398.000 269.600 398.800 270.400 ;
        RECT 385.200 263.600 386.000 264.400 ;
        RECT 409.200 269.600 410.000 270.400 ;
        RECT 410.800 269.600 411.600 270.400 ;
        RECT 401.200 263.600 402.000 264.400 ;
        RECT 414.000 263.600 414.800 264.400 ;
        RECT 444.400 275.000 445.200 275.800 ;
        RECT 441.200 273.600 442.000 274.400 ;
        RECT 446.000 272.400 446.800 273.200 ;
        RECT 463.600 277.600 464.400 278.400 ;
        RECT 450.800 269.600 451.600 270.400 ;
        RECT 434.800 268.200 435.600 269.000 ;
        RECT 444.400 268.600 445.200 269.400 ;
        RECT 425.200 265.600 426.000 266.400 ;
        RECT 439.600 267.600 440.400 268.400 ;
        RECT 434.800 264.200 435.600 265.000 ;
        RECT 436.400 264.200 437.200 265.000 ;
        RECT 438.000 264.200 438.800 265.000 ;
        RECT 441.200 264.200 442.000 265.000 ;
        RECT 444.400 264.200 445.200 265.000 ;
        RECT 446.000 264.200 446.800 265.000 ;
        RECT 447.600 264.200 448.400 265.000 ;
        RECT 449.200 264.200 450.000 265.000 ;
        RECT 462.000 265.600 462.800 266.400 ;
        RECT 482.800 275.000 483.600 275.800 ;
        RECT 479.600 273.600 480.400 274.400 ;
        RECT 484.400 272.400 485.200 273.200 ;
        RECT 502.000 277.600 502.800 278.400 ;
        RECT 473.200 268.200 474.000 269.000 ;
        RECT 482.800 268.600 483.600 269.400 ;
        RECT 478.000 267.600 478.800 268.400 ;
        RECT 473.200 264.200 474.000 265.000 ;
        RECT 474.800 264.200 475.600 265.000 ;
        RECT 476.400 264.200 477.200 265.000 ;
        RECT 479.600 264.200 480.400 265.000 ;
        RECT 482.800 264.200 483.600 265.000 ;
        RECT 484.400 264.200 485.200 265.000 ;
        RECT 486.000 264.200 486.800 265.000 ;
        RECT 487.600 264.200 488.400 265.000 ;
        RECT 497.200 263.600 498.000 264.400 ;
        RECT 503.600 277.600 504.400 278.400 ;
        RECT 529.200 277.600 530.000 278.400 ;
        RECT 524.400 269.600 525.200 270.400 ;
        RECT 529.200 267.600 530.000 268.400 ;
        RECT 505.200 265.600 506.000 266.400 ;
        RECT 532.400 269.600 533.200 270.400 ;
        RECT 535.600 269.600 536.400 270.400 ;
        RECT 558.000 277.600 558.800 278.400 ;
        RECT 561.200 277.600 562.000 278.400 ;
        RECT 542.000 267.600 542.800 268.400 ;
        RECT 521.200 263.600 522.000 264.400 ;
        RECT 540.400 266.200 541.200 267.000 ;
        RECT 583.600 275.600 584.400 276.400 ;
        RECT 562.800 267.600 563.600 268.400 ;
        RECT 570.800 269.600 571.600 270.400 ;
        RECT 572.400 269.600 573.200 270.400 ;
        RECT 591.600 271.600 592.400 272.400 ;
        RECT 585.200 269.600 586.000 270.400 ;
        RECT 586.800 269.600 587.600 270.400 ;
        RECT 598.000 269.600 598.800 270.400 ;
        RECT 593.200 267.600 594.000 268.400 ;
        RECT 599.600 267.600 600.400 268.400 ;
        RECT 609.200 269.600 610.000 270.400 ;
        RECT 620.400 277.600 621.200 278.400 ;
        RECT 617.200 269.600 618.000 270.400 ;
        RECT 594.800 263.600 595.600 264.400 ;
        RECT 618.800 267.600 619.600 268.400 ;
        RECT 614.000 263.600 614.800 264.400 ;
        RECT 625.200 277.600 626.000 278.400 ;
        RECT 622.000 265.600 622.800 266.400 ;
        RECT 628.400 269.600 629.200 270.400 ;
        RECT 630.000 269.600 630.800 270.400 ;
        RECT 626.800 267.600 627.600 268.400 ;
        RECT 639.600 269.600 640.400 270.400 ;
        RECT 646.000 269.600 646.800 270.400 ;
        RECT 654.000 271.600 654.800 272.400 ;
        RECT 666.800 275.600 667.600 276.400 ;
        RECT 663.600 273.600 664.400 274.400 ;
        RECT 641.200 267.600 642.000 268.400 ;
        RECT 657.200 269.600 658.000 270.400 ;
        RECT 658.800 269.600 659.600 270.400 ;
        RECT 663.600 269.600 664.400 270.400 ;
        RECT 665.200 267.600 666.000 268.400 ;
        RECT 681.200 272.400 682.000 273.200 ;
        RECT 684.400 271.000 685.200 271.800 ;
        RECT 684.400 266.200 685.200 267.000 ;
        RECT 12.400 257.600 13.200 258.400 ;
        RECT 31.600 255.600 32.400 256.400 ;
        RECT 33.200 254.200 34.000 255.000 ;
        RECT 23.600 251.600 24.400 252.400 ;
        RECT 44.400 251.600 45.200 252.400 ;
        RECT 26.800 246.800 27.600 247.600 ;
        RECT 30.000 246.200 30.800 247.000 ;
        RECT 25.200 244.200 26.000 245.000 ;
        RECT 26.800 244.200 27.600 245.000 ;
        RECT 28.400 244.200 29.200 245.000 ;
        RECT 33.200 246.200 34.000 247.000 ;
        RECT 36.400 246.200 37.200 247.000 ;
        RECT 66.800 255.600 67.600 256.400 ;
        RECT 68.400 254.200 69.200 255.000 ;
        RECT 58.800 251.600 59.600 252.400 ;
        RECT 76.400 251.600 77.200 252.400 ;
        RECT 50.800 249.600 51.600 250.400 ;
        RECT 38.000 244.200 38.800 245.000 ;
        RECT 39.600 244.200 40.400 245.000 ;
        RECT 62.000 246.800 62.800 247.600 ;
        RECT 65.200 246.200 66.000 247.000 ;
        RECT 60.400 244.200 61.200 245.000 ;
        RECT 62.000 244.200 62.800 245.000 ;
        RECT 63.600 244.200 64.400 245.000 ;
        RECT 68.400 246.200 69.200 247.000 ;
        RECT 71.600 246.200 72.400 247.000 ;
        RECT 73.200 244.200 74.000 245.000 ;
        RECT 74.800 244.200 75.600 245.000 ;
        RECT 89.200 257.600 90.000 258.400 ;
        RECT 105.200 255.600 106.000 256.400 ;
        RECT 106.800 254.200 107.600 255.000 ;
        RECT 129.200 257.600 130.000 258.400 ;
        RECT 118.000 251.600 118.800 252.400 ;
        RECT 84.400 243.600 85.200 244.400 ;
        RECT 100.400 246.800 101.200 247.600 ;
        RECT 103.600 246.200 104.400 247.000 ;
        RECT 98.800 244.200 99.600 245.000 ;
        RECT 100.400 244.200 101.200 245.000 ;
        RECT 102.000 244.200 102.800 245.000 ;
        RECT 106.800 246.200 107.600 247.000 ;
        RECT 110.000 246.200 110.800 247.000 ;
        RECT 142.000 253.600 142.800 254.400 ;
        RECT 111.600 244.200 112.400 245.000 ;
        RECT 113.200 244.200 114.000 245.000 ;
        RECT 153.200 243.600 154.000 244.400 ;
        RECT 183.600 253.600 184.400 254.400 ;
        RECT 193.200 253.000 194.000 253.800 ;
        RECT 202.800 252.600 203.600 253.400 ;
        RECT 217.200 257.600 218.000 258.400 ;
        RECT 186.800 251.600 187.600 252.400 ;
        RECT 209.200 251.600 210.000 252.400 ;
        RECT 194.800 248.800 195.600 249.600 ;
        RECT 199.600 247.600 200.400 248.400 ;
        RECT 196.400 246.200 197.200 247.000 ;
        RECT 193.200 244.200 194.000 245.000 ;
        RECT 194.800 244.200 195.600 245.000 ;
        RECT 199.600 246.200 200.400 247.000 ;
        RECT 202.800 246.200 203.600 247.000 ;
        RECT 204.400 244.200 205.200 245.000 ;
        RECT 206.000 244.200 206.800 245.000 ;
        RECT 207.600 244.200 208.400 245.000 ;
        RECT 225.200 257.600 226.000 258.400 ;
        RECT 241.200 255.600 242.000 256.400 ;
        RECT 242.800 254.200 243.600 255.000 ;
        RECT 244.400 251.600 245.200 252.400 ;
        RECT 222.000 243.600 222.800 244.400 ;
        RECT 236.400 246.800 237.200 247.600 ;
        RECT 239.600 246.200 240.400 247.000 ;
        RECT 234.800 244.200 235.600 245.000 ;
        RECT 236.400 244.200 237.200 245.000 ;
        RECT 238.000 244.200 238.800 245.000 ;
        RECT 242.800 246.200 243.600 247.000 ;
        RECT 246.000 246.200 246.800 247.000 ;
        RECT 274.800 257.600 275.600 258.400 ;
        RECT 247.600 244.200 248.400 245.000 ;
        RECT 249.200 244.200 250.000 245.000 ;
        RECT 270.000 253.600 270.800 254.400 ;
        RECT 290.800 255.600 291.600 256.400 ;
        RECT 292.400 254.200 293.200 255.000 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 302.000 251.600 302.800 252.400 ;
        RECT 271.600 249.600 272.400 250.400 ;
        RECT 286.000 246.800 286.800 247.600 ;
        RECT 289.200 246.200 290.000 247.000 ;
        RECT 284.400 244.200 285.200 245.000 ;
        RECT 286.000 244.200 286.800 245.000 ;
        RECT 287.600 244.200 288.400 245.000 ;
        RECT 292.400 246.200 293.200 247.000 ;
        RECT 295.600 246.200 296.400 247.000 ;
        RECT 324.400 249.600 325.200 250.400 ;
        RECT 297.200 244.200 298.000 245.000 ;
        RECT 298.800 244.200 299.600 245.000 ;
        RECT 310.000 243.600 310.800 244.400 ;
        RECT 316.400 243.600 317.200 244.400 ;
        RECT 340.400 253.600 341.200 254.400 ;
        RECT 353.200 253.600 354.000 254.400 ;
        RECT 367.600 253.600 368.400 254.400 ;
        RECT 338.800 249.600 339.600 250.400 ;
        RECT 337.200 243.600 338.000 244.400 ;
        RECT 358.000 249.600 358.800 250.400 ;
        RECT 372.400 249.600 373.200 250.400 ;
        RECT 378.800 249.600 379.600 250.400 ;
        RECT 383.600 251.600 384.400 252.400 ;
        RECT 391.600 249.600 392.400 250.400 ;
        RECT 370.800 243.600 371.600 244.400 ;
        RECT 386.800 243.600 387.600 244.400 ;
        RECT 390.000 245.600 390.800 246.400 ;
        RECT 402.800 257.600 403.600 258.400 ;
        RECT 406.000 257.600 406.800 258.400 ;
        RECT 402.800 243.600 403.600 244.400 ;
        RECT 431.600 253.000 432.400 253.800 ;
        RECT 441.200 252.600 442.000 253.400 ;
        RECT 455.600 257.600 456.400 258.400 ;
        RECT 463.600 257.600 464.400 258.400 ;
        RECT 426.800 251.600 427.600 252.400 ;
        RECT 433.200 248.800 434.000 249.600 ;
        RECT 438.000 247.600 438.800 248.400 ;
        RECT 414.000 245.600 414.800 246.400 ;
        RECT 434.800 246.200 435.600 247.000 ;
        RECT 431.600 244.200 432.400 245.000 ;
        RECT 433.200 244.200 434.000 245.000 ;
        RECT 438.000 246.200 438.800 247.000 ;
        RECT 441.200 246.200 442.000 247.000 ;
        RECT 442.800 244.200 443.600 245.000 ;
        RECT 444.400 244.200 445.200 245.000 ;
        RECT 446.000 244.200 446.800 245.000 ;
        RECT 471.600 253.600 472.400 254.400 ;
        RECT 484.400 253.600 485.200 254.400 ;
        RECT 519.600 253.000 520.400 253.800 ;
        RECT 529.200 252.600 530.000 253.400 ;
        RECT 543.600 255.600 544.400 256.400 ;
        RECT 546.800 257.600 547.600 258.400 ;
        RECT 514.800 251.600 515.600 252.400 ;
        RECT 521.200 248.800 522.000 249.600 ;
        RECT 526.000 247.600 526.800 248.400 ;
        RECT 522.800 246.200 523.600 247.000 ;
        RECT 519.600 244.200 520.400 245.000 ;
        RECT 521.200 244.200 522.000 245.000 ;
        RECT 526.000 246.200 526.800 247.000 ;
        RECT 529.200 246.200 530.000 247.000 ;
        RECT 530.800 244.200 531.600 245.000 ;
        RECT 532.400 244.200 533.200 245.000 ;
        RECT 534.000 244.200 534.800 245.000 ;
        RECT 601.200 257.600 602.000 258.400 ;
        RECT 551.600 252.200 552.400 253.000 ;
        RECT 564.400 250.200 565.200 251.000 ;
        RECT 588.400 251.800 589.200 252.600 ;
        RECT 583.600 250.200 584.400 251.000 ;
        RECT 602.800 257.600 603.600 258.400 ;
        RECT 622.000 257.600 622.800 258.400 ;
        RECT 618.800 253.600 619.600 254.400 ;
        RECT 607.600 252.200 608.400 253.000 ;
        RECT 687.600 257.600 688.400 258.400 ;
        RECT 626.800 252.200 627.600 253.000 ;
        RECT 620.400 250.200 621.200 251.000 ;
        RECT 639.600 250.200 640.400 251.000 ;
        RECT 671.600 253.600 672.400 254.400 ;
        RECT 655.600 251.600 656.400 252.400 ;
        RECT 657.200 251.600 658.000 252.400 ;
        RECT 644.400 247.600 645.200 248.400 ;
        RECT 674.800 251.800 675.600 252.600 ;
        RECT 668.400 249.600 669.200 250.400 ;
        RECT 670.000 250.200 670.800 251.000 ;
        RECT 20.400 237.600 21.200 238.400 ;
        RECT 2.800 223.600 3.600 224.400 ;
        RECT 18.800 225.600 19.600 226.400 ;
        RECT 34.800 234.400 35.600 235.200 ;
        RECT 38.000 235.000 38.800 235.800 ;
        RECT 33.200 232.400 34.000 233.200 ;
        RECT 23.600 225.600 24.400 226.400 ;
        RECT 42.800 227.600 43.600 228.400 ;
        RECT 39.600 225.600 40.400 226.400 ;
        RECT 82.800 237.600 83.600 238.400 ;
        RECT 33.200 224.200 34.000 225.000 ;
        RECT 34.800 224.200 35.600 225.000 ;
        RECT 36.400 224.200 37.200 225.000 ;
        RECT 38.000 224.200 38.800 225.000 ;
        RECT 41.200 224.200 42.000 225.000 ;
        RECT 44.400 224.200 45.200 225.000 ;
        RECT 46.000 224.200 46.800 225.000 ;
        RECT 47.600 224.200 48.400 225.000 ;
        RECT 63.600 229.600 64.400 230.400 ;
        RECT 65.200 229.600 66.000 230.400 ;
        RECT 66.800 225.600 67.600 226.400 ;
        RECT 78.000 229.600 78.800 230.400 ;
        RECT 79.600 229.600 80.400 230.400 ;
        RECT 105.200 235.000 106.000 235.800 ;
        RECT 102.000 233.600 102.800 234.400 ;
        RECT 119.600 237.600 120.400 238.400 ;
        RECT 106.800 232.400 107.600 233.200 ;
        RECT 140.400 237.600 141.200 238.400 ;
        RECT 111.600 229.600 112.400 230.400 ;
        RECT 73.200 223.600 74.000 224.400 ;
        RECT 95.600 228.200 96.400 229.000 ;
        RECT 105.200 228.600 106.000 229.400 ;
        RECT 100.400 227.600 101.200 228.400 ;
        RECT 95.600 224.200 96.400 225.000 ;
        RECT 97.200 224.200 98.000 225.000 ;
        RECT 98.800 224.200 99.600 225.000 ;
        RECT 102.000 224.200 102.800 225.000 ;
        RECT 105.200 224.200 106.000 225.000 ;
        RECT 106.800 224.200 107.600 225.000 ;
        RECT 108.400 224.200 109.200 225.000 ;
        RECT 110.000 224.200 110.800 225.000 ;
        RECT 151.600 234.400 152.400 235.200 ;
        RECT 154.800 235.000 155.600 235.800 ;
        RECT 150.000 232.400 150.800 233.200 ;
        RECT 130.800 225.600 131.600 226.400 ;
        RECT 148.400 229.600 149.200 230.400 ;
        RECT 134.000 223.600 134.800 224.400 ;
        RECT 159.600 227.600 160.400 228.400 ;
        RECT 156.400 225.600 157.200 226.400 ;
        RECT 150.000 224.200 150.800 225.000 ;
        RECT 151.600 224.200 152.400 225.000 ;
        RECT 153.200 224.200 154.000 225.000 ;
        RECT 154.800 224.200 155.600 225.000 ;
        RECT 158.000 224.200 158.800 225.000 ;
        RECT 161.200 224.200 162.000 225.000 ;
        RECT 162.800 224.200 163.600 225.000 ;
        RECT 164.400 224.200 165.200 225.000 ;
        RECT 174.000 225.600 174.800 226.400 ;
        RECT 199.600 234.400 200.400 235.200 ;
        RECT 202.800 235.000 203.600 235.800 ;
        RECT 226.800 237.600 227.600 238.400 ;
        RECT 198.000 232.400 198.800 233.200 ;
        RECT 183.600 229.600 184.400 230.400 ;
        RECT 185.200 229.600 186.000 230.400 ;
        RECT 188.400 223.600 189.200 224.400 ;
        RECT 207.600 227.600 208.400 228.400 ;
        RECT 204.400 225.600 205.200 226.400 ;
        RECT 198.000 224.200 198.800 225.000 ;
        RECT 199.600 224.200 200.400 225.000 ;
        RECT 201.200 224.200 202.000 225.000 ;
        RECT 202.800 224.200 203.600 225.000 ;
        RECT 206.000 224.200 206.800 225.000 ;
        RECT 209.200 224.200 210.000 225.000 ;
        RECT 210.800 224.200 211.600 225.000 ;
        RECT 212.400 224.200 213.200 225.000 ;
        RECT 228.400 229.600 229.200 230.400 ;
        RECT 230.000 229.600 230.800 230.400 ;
        RECT 234.800 229.600 235.600 230.400 ;
        RECT 255.600 235.000 256.400 235.800 ;
        RECT 252.400 233.600 253.200 234.400 ;
        RECT 257.200 232.400 258.000 233.200 ;
        RECT 262.000 229.600 262.800 230.400 ;
        RECT 236.400 227.600 237.200 228.400 ;
        RECT 246.000 228.200 246.800 229.000 ;
        RECT 255.600 228.600 256.400 229.400 ;
        RECT 250.800 227.600 251.600 228.400 ;
        RECT 270.200 229.600 271.000 230.400 ;
        RECT 246.000 224.200 246.800 225.000 ;
        RECT 247.600 224.200 248.400 225.000 ;
        RECT 249.200 224.200 250.000 225.000 ;
        RECT 252.400 224.200 253.200 225.000 ;
        RECT 255.600 224.200 256.400 225.000 ;
        RECT 257.200 224.200 258.000 225.000 ;
        RECT 258.800 224.200 259.600 225.000 ;
        RECT 260.400 224.200 261.200 225.000 ;
        RECT 284.400 237.600 285.200 238.400 ;
        RECT 282.800 225.600 283.600 226.400 ;
        RECT 287.600 227.600 288.400 228.400 ;
        RECT 286.000 225.600 286.800 226.400 ;
        RECT 290.800 227.600 291.600 228.400 ;
        RECT 300.400 227.600 301.200 228.400 ;
        RECT 306.800 229.600 307.600 230.400 ;
        RECT 313.200 229.600 314.000 230.400 ;
        RECT 335.600 235.000 336.400 235.800 ;
        RECT 332.400 233.600 333.200 234.400 ;
        RECT 337.200 232.400 338.000 233.200 ;
        RECT 354.800 237.600 355.600 238.400 ;
        RECT 294.000 223.600 294.800 224.400 ;
        RECT 295.600 223.600 296.400 224.400 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 326.000 228.200 326.800 229.000 ;
        RECT 335.600 228.600 336.400 229.400 ;
        RECT 310.000 223.600 310.800 224.400 ;
        RECT 330.800 227.600 331.600 228.400 ;
        RECT 326.000 224.200 326.800 225.000 ;
        RECT 327.600 224.200 328.400 225.000 ;
        RECT 329.200 224.200 330.000 225.000 ;
        RECT 332.400 224.200 333.200 225.000 ;
        RECT 335.600 224.200 336.400 225.000 ;
        RECT 337.200 224.200 338.000 225.000 ;
        RECT 338.800 224.200 339.600 225.000 ;
        RECT 340.400 224.200 341.200 225.000 ;
        RECT 353.200 227.600 354.000 228.400 ;
        RECT 356.400 227.600 357.200 228.400 ;
        RECT 374.000 237.600 374.800 238.400 ;
        RECT 383.600 237.600 384.400 238.400 ;
        RECT 375.600 233.600 376.400 234.400 ;
        RECT 382.000 233.600 382.800 234.400 ;
        RECT 364.400 229.600 365.200 230.400 ;
        RECT 366.000 227.600 366.800 228.400 ;
        RECT 378.800 231.600 379.600 232.400 ;
        RECT 377.200 229.600 378.000 230.400 ;
        RECT 385.200 231.600 386.000 232.400 ;
        RECT 383.600 229.600 384.400 230.400 ;
        RECT 404.400 235.000 405.200 235.800 ;
        RECT 401.200 233.600 402.000 234.400 ;
        RECT 406.000 232.400 406.800 233.200 ;
        RECT 410.800 229.600 411.600 230.400 ;
        RECT 394.800 228.200 395.600 229.000 ;
        RECT 404.400 228.600 405.200 229.400 ;
        RECT 359.600 223.600 360.400 224.400 ;
        RECT 399.600 227.600 400.400 228.400 ;
        RECT 394.800 224.200 395.600 225.000 ;
        RECT 396.400 224.200 397.200 225.000 ;
        RECT 398.000 224.200 398.800 225.000 ;
        RECT 401.200 224.200 402.000 225.000 ;
        RECT 404.400 224.200 405.200 225.000 ;
        RECT 406.000 224.200 406.800 225.000 ;
        RECT 407.600 224.200 408.400 225.000 ;
        RECT 409.200 224.200 410.000 225.000 ;
        RECT 428.400 229.600 429.200 230.400 ;
        RECT 450.800 237.600 451.600 238.400 ;
        RECT 436.400 225.600 437.200 226.400 ;
        RECT 471.600 235.000 472.400 235.800 ;
        RECT 468.400 233.600 469.200 234.400 ;
        RECT 473.200 232.400 474.000 233.200 ;
        RECT 478.000 229.600 478.800 230.400 ;
        RECT 462.000 228.200 462.800 229.000 ;
        RECT 471.600 228.600 472.400 229.400 ;
        RECT 450.800 223.600 451.600 224.400 ;
        RECT 466.800 227.600 467.600 228.400 ;
        RECT 462.000 224.200 462.800 225.000 ;
        RECT 463.600 224.200 464.400 225.000 ;
        RECT 465.200 224.200 466.000 225.000 ;
        RECT 468.400 224.200 469.200 225.000 ;
        RECT 471.600 224.200 472.400 225.000 ;
        RECT 473.200 224.200 474.000 225.000 ;
        RECT 474.800 224.200 475.600 225.000 ;
        RECT 476.400 224.200 477.200 225.000 ;
        RECT 489.200 229.600 490.000 230.400 ;
        RECT 490.800 229.600 491.600 230.400 ;
        RECT 486.000 223.600 486.800 224.400 ;
        RECT 519.600 235.000 520.400 235.800 ;
        RECT 516.400 233.600 517.200 234.400 ;
        RECT 521.200 232.400 522.000 233.200 ;
        RECT 510.000 228.200 510.800 229.000 ;
        RECT 519.600 228.600 520.400 229.400 ;
        RECT 500.400 225.600 501.200 226.400 ;
        RECT 514.800 227.600 515.600 228.400 ;
        RECT 510.000 224.200 510.800 225.000 ;
        RECT 511.600 224.200 512.400 225.000 ;
        RECT 513.200 224.200 514.000 225.000 ;
        RECT 516.400 224.200 517.200 225.000 ;
        RECT 519.600 224.200 520.400 225.000 ;
        RECT 521.200 224.200 522.000 225.000 ;
        RECT 522.800 224.200 523.600 225.000 ;
        RECT 524.400 224.200 525.200 225.000 ;
        RECT 534.000 225.600 534.800 226.400 ;
        RECT 538.800 225.600 539.600 226.400 ;
        RECT 537.200 223.600 538.000 224.400 ;
        RECT 546.800 225.600 547.600 226.400 ;
        RECT 553.200 229.600 554.000 230.400 ;
        RECT 558.000 229.600 558.800 230.400 ;
        RECT 545.200 223.600 546.000 224.400 ;
        RECT 548.400 223.600 549.200 224.400 ;
        RECT 559.600 227.600 560.400 228.400 ;
        RECT 561.200 227.600 562.000 228.400 ;
        RECT 588.400 234.400 589.200 235.200 ;
        RECT 591.600 235.000 592.400 235.800 ;
        RECT 610.800 237.600 611.600 238.400 ;
        RECT 586.800 232.400 587.600 233.200 ;
        RECT 569.200 227.600 570.000 228.400 ;
        RECT 585.200 229.600 586.000 230.400 ;
        RECT 596.400 227.600 597.200 228.400 ;
        RECT 593.200 225.600 594.000 226.400 ;
        RECT 586.800 224.200 587.600 225.000 ;
        RECT 588.400 224.200 589.200 225.000 ;
        RECT 590.000 224.200 590.800 225.000 ;
        RECT 591.600 224.200 592.400 225.000 ;
        RECT 594.800 224.200 595.600 225.000 ;
        RECT 598.000 224.200 598.800 225.000 ;
        RECT 599.600 224.200 600.400 225.000 ;
        RECT 601.200 224.200 602.000 225.000 ;
        RECT 625.200 232.400 626.000 233.200 ;
        RECT 628.400 231.000 629.200 231.800 ;
        RECT 647.600 235.000 648.400 235.800 ;
        RECT 644.400 233.600 645.200 234.400 ;
        RECT 649.200 232.400 650.000 233.200 ;
        RECT 666.800 237.600 667.600 238.400 ;
        RECT 638.000 228.200 638.800 229.000 ;
        RECT 647.600 228.600 648.400 229.400 ;
        RECT 628.400 226.200 629.200 227.000 ;
        RECT 642.800 227.600 643.600 228.400 ;
        RECT 638.000 224.200 638.800 225.000 ;
        RECT 639.600 224.200 640.400 225.000 ;
        RECT 641.200 224.200 642.000 225.000 ;
        RECT 644.400 224.200 645.200 225.000 ;
        RECT 647.600 224.200 648.400 225.000 ;
        RECT 649.200 224.200 650.000 225.000 ;
        RECT 650.800 224.200 651.600 225.000 ;
        RECT 652.400 224.200 653.200 225.000 ;
        RECT 662.000 223.600 662.800 224.400 ;
        RECT 674.800 229.600 675.600 230.400 ;
        RECT 668.400 226.200 669.200 227.000 ;
        RECT 686.000 223.600 686.800 224.400 ;
        RECT 9.200 213.600 10.000 214.400 ;
        RECT 18.800 213.000 19.600 213.800 ;
        RECT 9.200 209.600 10.000 210.400 ;
        RECT 28.400 212.600 29.200 213.400 ;
        RECT 62.000 217.600 62.800 218.400 ;
        RECT 23.600 211.600 24.400 212.400 ;
        RECT 58.800 213.600 59.600 214.400 ;
        RECT 20.400 208.800 21.200 209.600 ;
        RECT 25.200 207.600 26.000 208.400 ;
        RECT 22.000 206.200 22.800 207.000 ;
        RECT 18.800 204.200 19.600 205.000 ;
        RECT 20.400 204.200 21.200 205.000 ;
        RECT 25.200 206.200 26.000 207.000 ;
        RECT 28.400 206.200 29.200 207.000 ;
        RECT 30.000 204.200 30.800 205.000 ;
        RECT 31.600 204.200 32.400 205.000 ;
        RECT 33.200 204.200 34.000 205.000 ;
        RECT 42.800 203.600 43.600 204.400 ;
        RECT 47.600 203.600 48.400 204.400 ;
        RECT 78.000 215.600 78.800 216.400 ;
        RECT 79.600 214.200 80.400 215.000 ;
        RECT 95.600 213.600 96.400 214.400 ;
        RECT 108.400 213.600 109.200 214.400 ;
        RECT 70.000 211.600 70.800 212.400 ;
        RECT 90.800 211.600 91.600 212.400 ;
        RECT 62.000 203.600 62.800 204.400 ;
        RECT 73.200 206.800 74.000 207.600 ;
        RECT 76.400 206.200 77.200 207.000 ;
        RECT 71.600 204.200 72.400 205.000 ;
        RECT 73.200 204.200 74.000 205.000 ;
        RECT 74.800 204.200 75.600 205.000 ;
        RECT 79.600 206.200 80.400 207.000 ;
        RECT 82.800 206.200 83.600 207.000 ;
        RECT 84.400 204.200 85.200 205.000 ;
        RECT 86.000 204.200 86.800 205.000 ;
        RECT 106.800 203.600 107.600 204.400 ;
        RECT 119.600 217.600 120.400 218.400 ;
        RECT 135.600 215.600 136.400 216.400 ;
        RECT 137.200 214.200 138.000 215.000 ;
        RECT 154.800 217.600 155.600 218.400 ;
        RECT 148.400 211.600 149.200 212.400 ;
        RECT 130.800 206.800 131.600 207.600 ;
        RECT 134.000 206.200 134.800 207.000 ;
        RECT 129.200 204.200 130.000 205.000 ;
        RECT 130.800 204.200 131.600 205.000 ;
        RECT 132.400 204.200 133.200 205.000 ;
        RECT 137.200 206.200 138.000 207.000 ;
        RECT 140.400 206.200 141.200 207.000 ;
        RECT 170.800 215.600 171.600 216.400 ;
        RECT 172.400 214.200 173.200 215.000 ;
        RECT 183.600 211.600 184.400 212.400 ;
        RECT 142.000 204.200 142.800 205.000 ;
        RECT 143.600 204.200 144.400 205.000 ;
        RECT 166.000 206.800 166.800 207.600 ;
        RECT 169.200 206.200 170.000 207.000 ;
        RECT 164.400 204.200 165.200 205.000 ;
        RECT 166.000 204.200 166.800 205.000 ;
        RECT 167.600 204.200 168.400 205.000 ;
        RECT 172.400 206.200 173.200 207.000 ;
        RECT 175.600 206.200 176.400 207.000 ;
        RECT 196.400 213.000 197.200 213.800 ;
        RECT 206.000 212.600 206.800 213.400 ;
        RECT 190.000 211.600 190.800 212.400 ;
        RECT 212.400 211.600 213.200 212.400 ;
        RECT 198.000 208.800 198.800 209.600 ;
        RECT 202.800 207.600 203.600 208.400 ;
        RECT 177.200 204.200 178.000 205.000 ;
        RECT 178.800 204.200 179.600 205.000 ;
        RECT 199.600 206.200 200.400 207.000 ;
        RECT 196.400 204.200 197.200 205.000 ;
        RECT 198.000 204.200 198.800 205.000 ;
        RECT 202.800 206.200 203.600 207.000 ;
        RECT 206.000 206.200 206.800 207.000 ;
        RECT 207.600 204.200 208.400 205.000 ;
        RECT 209.200 204.200 210.000 205.000 ;
        RECT 210.800 204.200 211.600 205.000 ;
        RECT 226.800 211.600 227.600 212.400 ;
        RECT 231.600 213.600 232.400 214.400 ;
        RECT 233.200 211.600 234.000 212.400 ;
        RECT 220.400 203.600 221.200 204.400 ;
        RECT 238.000 209.600 238.800 210.400 ;
        RECT 242.800 211.600 243.600 212.400 ;
        RECT 249.200 211.600 250.000 212.400 ;
        RECT 255.600 211.600 256.400 212.400 ;
        RECT 252.400 203.600 253.200 204.400 ;
        RECT 257.200 209.600 258.000 210.400 ;
        RECT 273.200 213.000 274.000 213.800 ;
        RECT 282.800 212.600 283.600 213.400 ;
        RECT 313.200 217.600 314.000 218.400 ;
        RECT 270.000 211.600 270.800 212.400 ;
        RECT 274.800 208.800 275.600 209.600 ;
        RECT 279.600 207.600 280.400 208.400 ;
        RECT 276.400 206.200 277.200 207.000 ;
        RECT 273.200 204.200 274.000 205.000 ;
        RECT 274.800 204.200 275.600 205.000 ;
        RECT 279.600 206.200 280.400 207.000 ;
        RECT 282.800 206.200 283.600 207.000 ;
        RECT 284.400 204.200 285.200 205.000 ;
        RECT 286.000 204.200 286.800 205.000 ;
        RECT 287.600 204.200 288.400 205.000 ;
        RECT 303.600 209.600 304.400 210.400 ;
        RECT 318.000 217.600 318.800 218.400 ;
        RECT 324.400 217.600 325.200 218.400 ;
        RECT 324.400 203.600 325.200 204.400 ;
        RECT 334.000 209.600 334.800 210.400 ;
        RECT 330.800 203.600 331.600 204.400 ;
        RECT 338.800 209.600 339.600 210.400 ;
        RECT 348.400 209.600 349.200 210.400 ;
        RECT 350.000 209.600 350.800 210.400 ;
        RECT 372.400 215.600 373.200 216.400 ;
        RECT 374.000 214.200 374.800 215.000 ;
        RECT 385.200 211.600 386.000 212.400 ;
        RECT 367.600 206.800 368.400 207.600 ;
        RECT 370.800 206.200 371.600 207.000 ;
        RECT 366.000 204.200 366.800 205.000 ;
        RECT 367.600 204.200 368.400 205.000 ;
        RECT 369.200 204.200 370.000 205.000 ;
        RECT 374.000 206.200 374.800 207.000 ;
        RECT 377.200 206.200 378.000 207.000 ;
        RECT 391.600 213.600 392.400 214.400 ;
        RECT 415.600 213.000 416.400 213.800 ;
        RECT 378.800 204.200 379.600 205.000 ;
        RECT 380.400 204.200 381.200 205.000 ;
        RECT 401.200 209.600 402.000 210.400 ;
        RECT 425.200 212.600 426.000 213.400 ;
        RECT 410.800 211.600 411.600 212.400 ;
        RECT 417.200 208.800 418.000 209.600 ;
        RECT 422.000 207.600 422.800 208.400 ;
        RECT 418.800 206.200 419.600 207.000 ;
        RECT 415.600 204.200 416.400 205.000 ;
        RECT 417.200 204.200 418.000 205.000 ;
        RECT 422.000 206.200 422.800 207.000 ;
        RECT 425.200 206.200 426.000 207.000 ;
        RECT 426.800 204.200 427.600 205.000 ;
        RECT 428.400 204.200 429.200 205.000 ;
        RECT 430.000 204.200 430.800 205.000 ;
        RECT 439.600 203.600 440.400 204.400 ;
        RECT 450.600 211.600 451.400 212.400 ;
        RECT 466.800 215.600 467.600 216.400 ;
        RECT 468.400 214.200 469.200 215.000 ;
        RECT 446.000 203.600 446.800 204.400 ;
        RECT 462.000 206.800 462.800 207.600 ;
        RECT 465.200 206.200 466.000 207.000 ;
        RECT 460.400 204.200 461.200 205.000 ;
        RECT 462.000 204.200 462.800 205.000 ;
        RECT 463.600 204.200 464.400 205.000 ;
        RECT 468.400 206.200 469.200 207.000 ;
        RECT 471.600 206.200 472.400 207.000 ;
        RECT 473.200 204.200 474.000 205.000 ;
        RECT 474.800 204.200 475.600 205.000 ;
        RECT 495.600 213.000 496.400 213.800 ;
        RECT 505.200 212.600 506.000 213.400 ;
        RECT 527.600 217.600 528.400 218.400 ;
        RECT 489.200 211.600 490.000 212.400 ;
        RECT 500.400 211.600 501.200 212.400 ;
        RECT 511.600 211.600 512.400 212.400 ;
        RECT 497.200 208.800 498.000 209.600 ;
        RECT 502.000 207.600 502.800 208.400 ;
        RECT 486.000 203.600 486.800 204.400 ;
        RECT 498.800 206.200 499.600 207.000 ;
        RECT 495.600 204.200 496.400 205.000 ;
        RECT 497.200 204.200 498.000 205.000 ;
        RECT 502.000 206.200 502.800 207.000 ;
        RECT 505.200 206.200 506.000 207.000 ;
        RECT 506.800 204.200 507.600 205.000 ;
        RECT 508.400 204.200 509.200 205.000 ;
        RECT 510.000 204.200 510.800 205.000 ;
        RECT 519.600 203.600 520.400 204.400 ;
        RECT 527.600 209.600 528.400 210.400 ;
        RECT 529.200 209.600 530.000 210.400 ;
        RECT 545.200 211.600 546.000 212.400 ;
        RECT 554.800 209.600 555.600 210.400 ;
        RECT 561.200 211.600 562.000 212.400 ;
        RECT 586.800 217.600 587.600 218.400 ;
        RECT 566.000 211.600 566.800 212.400 ;
        RECT 577.200 213.600 578.000 214.400 ;
        RECT 590.000 213.600 590.800 214.400 ;
        RECT 598.000 211.600 598.800 212.400 ;
        RECT 607.600 211.600 608.400 212.400 ;
        RECT 612.200 211.600 613.000 212.400 ;
        RECT 628.400 215.600 629.200 216.400 ;
        RECT 630.000 214.200 630.800 215.000 ;
        RECT 649.200 214.800 650.000 215.600 ;
        RECT 620.400 211.600 621.200 212.400 ;
        RECT 642.800 211.600 643.600 212.400 ;
        RECT 623.600 206.800 624.400 207.600 ;
        RECT 626.800 206.200 627.600 207.000 ;
        RECT 622.000 204.200 622.800 205.000 ;
        RECT 623.600 204.200 624.400 205.000 ;
        RECT 625.200 204.200 626.000 205.000 ;
        RECT 630.000 206.200 630.800 207.000 ;
        RECT 633.200 206.200 634.000 207.000 ;
        RECT 668.400 217.600 669.200 218.400 ;
        RECT 655.600 213.600 656.400 214.400 ;
        RECT 671.600 213.600 672.400 214.400 ;
        RECT 634.800 204.200 635.600 205.000 ;
        RECT 636.400 204.200 637.200 205.000 ;
        RECT 682.800 203.600 683.600 204.400 ;
        RECT 14.000 197.600 14.800 198.400 ;
        RECT 6.000 189.600 6.800 190.400 ;
        RECT 14.000 189.600 14.800 190.400 ;
        RECT 34.800 195.000 35.600 195.800 ;
        RECT 31.600 193.600 32.400 194.400 ;
        RECT 49.200 195.600 50.000 196.400 ;
        RECT 36.400 192.400 37.200 193.200 ;
        RECT 9.200 185.600 10.000 186.400 ;
        RECT 15.600 187.600 16.400 188.400 ;
        RECT 25.200 188.200 26.000 189.000 ;
        RECT 34.800 188.600 35.600 189.400 ;
        RECT 30.000 187.600 30.800 188.400 ;
        RECT 25.200 184.200 26.000 185.000 ;
        RECT 26.800 184.200 27.600 185.000 ;
        RECT 28.400 184.200 29.200 185.000 ;
        RECT 31.600 184.200 32.400 185.000 ;
        RECT 34.800 184.200 35.600 185.000 ;
        RECT 36.400 184.200 37.200 185.000 ;
        RECT 38.000 184.200 38.800 185.000 ;
        RECT 39.600 184.200 40.400 185.000 ;
        RECT 55.600 189.600 56.400 190.400 ;
        RECT 58.800 185.600 59.600 186.400 ;
        RECT 68.400 193.600 69.200 194.400 ;
        RECT 71.600 191.600 72.400 192.400 ;
        RECT 65.200 187.600 66.000 188.400 ;
        RECT 63.600 183.600 64.400 184.400 ;
        RECT 70.000 185.600 70.800 186.400 ;
        RECT 76.400 189.600 77.200 190.400 ;
        RECT 82.800 189.600 83.600 190.400 ;
        RECT 105.200 193.600 106.000 194.400 ;
        RECT 78.000 187.600 78.800 188.400 ;
        RECT 84.400 187.600 85.200 188.400 ;
        RECT 87.600 187.600 88.400 188.400 ;
        RECT 86.000 186.200 86.800 187.000 ;
        RECT 73.200 183.600 74.000 184.400 ;
        RECT 79.600 183.600 80.400 184.400 ;
        RECT 118.000 189.600 118.800 190.400 ;
        RECT 108.400 187.600 109.200 188.400 ;
        RECT 119.600 187.600 120.400 188.400 ;
        RECT 122.800 187.600 123.600 188.400 ;
        RECT 121.200 186.200 122.000 187.000 ;
        RECT 103.600 183.600 104.400 184.400 ;
        RECT 114.800 183.600 115.600 184.400 ;
        RECT 138.800 183.600 139.600 184.400 ;
        RECT 140.400 191.600 141.200 192.400 ;
        RECT 142.000 185.600 142.800 186.400 ;
        RECT 143.600 186.200 144.400 187.000 ;
        RECT 169.200 189.600 170.000 190.400 ;
        RECT 164.400 187.600 165.200 188.400 ;
        RECT 161.200 183.600 162.000 184.400 ;
        RECT 162.800 186.200 163.600 187.000 ;
        RECT 194.800 194.400 195.600 195.200 ;
        RECT 198.000 195.000 198.800 195.800 ;
        RECT 193.200 192.400 194.000 193.200 ;
        RECT 180.400 183.600 181.200 184.400 ;
        RECT 183.600 183.600 184.400 184.400 ;
        RECT 202.800 187.600 203.600 188.400 ;
        RECT 199.600 185.600 200.400 186.400 ;
        RECT 193.200 184.200 194.000 185.000 ;
        RECT 194.800 184.200 195.600 185.000 ;
        RECT 196.400 184.200 197.200 185.000 ;
        RECT 198.000 184.200 198.800 185.000 ;
        RECT 201.200 184.200 202.000 185.000 ;
        RECT 204.400 184.200 205.200 185.000 ;
        RECT 206.000 184.200 206.800 185.000 ;
        RECT 207.600 184.200 208.400 185.000 ;
        RECT 241.200 194.400 242.000 195.200 ;
        RECT 244.400 195.000 245.200 195.800 ;
        RECT 239.600 192.400 240.400 193.200 ;
        RECT 229.800 187.600 230.600 188.400 ;
        RECT 220.400 185.600 221.200 186.400 ;
        RECT 223.600 185.600 224.400 186.400 ;
        RECT 238.000 189.600 238.800 190.400 ;
        RECT 249.200 187.600 250.000 188.400 ;
        RECT 246.000 185.600 246.800 186.400 ;
        RECT 239.600 184.200 240.400 185.000 ;
        RECT 241.200 184.200 242.000 185.000 ;
        RECT 242.800 184.200 243.600 185.000 ;
        RECT 244.400 184.200 245.200 185.000 ;
        RECT 247.600 184.200 248.400 185.000 ;
        RECT 250.800 184.200 251.600 185.000 ;
        RECT 252.400 184.200 253.200 185.000 ;
        RECT 254.000 184.200 254.800 185.000 ;
        RECT 281.200 194.400 282.000 195.200 ;
        RECT 284.400 195.000 285.200 195.800 ;
        RECT 303.600 197.600 304.400 198.400 ;
        RECT 279.600 192.400 280.400 193.200 ;
        RECT 278.000 189.600 278.800 190.400 ;
        RECT 270.000 183.600 270.800 184.400 ;
        RECT 289.200 187.600 290.000 188.400 ;
        RECT 286.000 185.600 286.800 186.400 ;
        RECT 279.600 184.200 280.400 185.000 ;
        RECT 281.200 184.200 282.000 185.000 ;
        RECT 282.800 184.200 283.600 185.000 ;
        RECT 284.400 184.200 285.200 185.000 ;
        RECT 287.600 184.200 288.400 185.000 ;
        RECT 290.800 184.200 291.600 185.000 ;
        RECT 292.400 184.200 293.200 185.000 ;
        RECT 294.000 184.200 294.800 185.000 ;
        RECT 324.400 195.000 325.200 195.800 ;
        RECT 321.200 193.600 322.000 194.400 ;
        RECT 326.000 192.400 326.800 193.200 ;
        RECT 314.800 188.200 315.600 189.000 ;
        RECT 324.400 188.600 325.200 189.400 ;
        RECT 305.200 185.600 306.000 186.400 ;
        RECT 319.600 187.600 320.400 188.400 ;
        RECT 339.000 187.600 339.800 188.400 ;
        RECT 314.800 184.200 315.600 185.000 ;
        RECT 316.400 184.200 317.200 185.000 ;
        RECT 318.000 184.200 318.800 185.000 ;
        RECT 321.200 184.200 322.000 185.000 ;
        RECT 324.400 184.200 325.200 185.000 ;
        RECT 326.000 184.200 326.800 185.000 ;
        RECT 327.600 184.200 328.400 185.000 ;
        RECT 329.200 184.200 330.000 185.000 ;
        RECT 350.000 187.600 350.800 188.400 ;
        RECT 370.800 195.600 371.600 196.400 ;
        RECT 369.200 187.600 370.000 188.400 ;
        RECT 353.200 183.600 354.000 184.400 ;
        RECT 356.400 185.600 357.200 186.400 ;
        RECT 372.400 187.600 373.200 188.400 ;
        RECT 383.600 189.600 384.400 190.400 ;
        RECT 396.400 197.600 397.200 198.400 ;
        RECT 402.800 197.600 403.600 198.400 ;
        RECT 398.000 193.600 398.800 194.400 ;
        RECT 404.400 193.600 405.200 194.400 ;
        RECT 401.200 191.600 402.000 192.400 ;
        RECT 388.400 187.600 389.200 188.400 ;
        RECT 428.400 197.600 429.200 198.400 ;
        RECT 393.200 187.600 394.000 188.400 ;
        RECT 439.600 194.400 440.400 195.200 ;
        RECT 442.800 195.000 443.600 195.800 ;
        RECT 438.000 192.400 438.800 193.200 ;
        RECT 380.400 183.600 381.200 184.400 ;
        RECT 383.600 183.600 384.400 184.400 ;
        RECT 409.200 183.600 410.000 184.400 ;
        RECT 447.600 187.600 448.400 188.400 ;
        RECT 444.400 185.600 445.200 186.400 ;
        RECT 465.200 189.600 466.000 190.400 ;
        RECT 438.000 184.200 438.800 185.000 ;
        RECT 439.600 184.200 440.400 185.000 ;
        RECT 441.200 184.200 442.000 185.000 ;
        RECT 442.800 184.200 443.600 185.000 ;
        RECT 446.000 184.200 446.800 185.000 ;
        RECT 449.200 184.200 450.000 185.000 ;
        RECT 450.800 184.200 451.600 185.000 ;
        RECT 452.400 184.200 453.200 185.000 ;
        RECT 466.800 187.600 467.600 188.400 ;
        RECT 482.800 189.600 483.600 190.400 ;
        RECT 484.400 189.600 485.200 190.400 ;
        RECT 506.800 197.600 507.600 198.400 ;
        RECT 462.000 183.600 462.800 184.400 ;
        RECT 470.000 185.600 470.800 186.400 ;
        RECT 526.000 197.600 526.800 198.400 ;
        RECT 529.000 191.800 529.800 192.600 ;
        RECT 494.000 185.600 494.800 186.400 ;
        RECT 506.800 183.600 507.600 184.400 ;
        RECT 516.400 185.600 517.200 186.400 ;
        RECT 513.200 183.600 514.000 184.400 ;
        RECT 545.200 189.600 546.000 190.400 ;
        RECT 522.800 185.600 523.600 186.400 ;
        RECT 521.200 183.600 522.000 184.400 ;
        RECT 529.000 186.200 529.800 187.000 ;
        RECT 537.200 187.600 538.000 188.400 ;
        RECT 540.400 187.600 541.200 188.400 ;
        RECT 538.800 186.200 539.600 187.000 ;
        RECT 559.600 189.600 560.400 190.400 ;
        RECT 561.200 189.600 562.000 190.400 ;
        RECT 567.600 189.600 568.400 190.400 ;
        RECT 575.600 189.600 576.400 190.400 ;
        RECT 577.200 189.600 578.000 190.400 ;
        RECT 569.200 187.600 570.000 188.400 ;
        RECT 586.800 189.600 587.600 190.400 ;
        RECT 588.400 189.600 589.200 190.400 ;
        RECT 594.800 189.600 595.600 190.400 ;
        RECT 556.400 183.600 557.200 184.400 ;
        RECT 596.400 187.600 597.200 188.400 ;
        RECT 612.400 192.400 613.200 193.200 ;
        RECT 615.600 191.000 616.400 191.800 ;
        RECT 618.800 189.600 619.600 190.400 ;
        RECT 620.400 189.600 621.200 190.400 ;
        RECT 625.200 189.600 626.000 190.400 ;
        RECT 639.600 193.600 640.400 194.400 ;
        RECT 615.600 186.200 616.400 187.000 ;
        RECT 636.400 189.600 637.200 190.400 ;
        RECT 638.000 189.600 638.800 190.400 ;
        RECT 598.000 183.600 598.800 184.400 ;
        RECT 654.000 192.400 654.800 193.200 ;
        RECT 657.200 191.000 658.000 191.800 ;
        RECT 657.200 186.200 658.000 187.000 ;
        RECT 658.800 185.600 659.600 186.400 ;
        RECT 679.600 191.800 680.400 192.600 ;
        RECT 670.000 185.600 670.800 186.400 ;
        RECT 676.400 187.600 677.200 188.400 ;
        RECT 679.600 186.200 680.400 187.000 ;
        RECT 671.600 183.600 672.400 184.400 ;
        RECT 687.600 187.600 688.400 188.400 ;
        RECT 684.400 186.400 685.200 187.200 ;
        RECT 9.200 173.000 10.000 173.800 ;
        RECT 18.800 172.600 19.600 173.400 ;
        RECT 14.000 171.600 14.800 172.400 ;
        RECT 25.200 171.600 26.000 172.400 ;
        RECT 57.200 177.600 58.000 178.400 ;
        RECT 41.200 171.800 42.000 172.600 ;
        RECT 10.800 168.800 11.600 169.600 ;
        RECT 15.600 167.600 16.400 168.400 ;
        RECT 12.400 166.200 13.200 167.000 ;
        RECT 9.200 164.200 10.000 165.000 ;
        RECT 10.800 164.200 11.600 165.000 ;
        RECT 15.600 166.200 16.400 167.000 ;
        RECT 18.800 166.200 19.600 167.000 ;
        RECT 20.400 164.200 21.200 165.000 ;
        RECT 22.000 164.200 22.800 165.000 ;
        RECT 23.600 164.200 24.400 165.000 ;
        RECT 36.400 170.200 37.200 171.000 ;
        RECT 33.200 167.600 34.000 168.400 ;
        RECT 54.000 163.600 54.800 164.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 65.200 169.600 66.000 170.400 ;
        RECT 84.400 173.000 85.200 173.800 ;
        RECT 94.000 172.600 94.800 173.400 ;
        RECT 79.600 171.600 80.400 172.400 ;
        RECT 86.000 168.800 86.800 169.600 ;
        RECT 90.800 167.600 91.600 168.400 ;
        RECT 87.600 166.200 88.400 167.000 ;
        RECT 84.400 164.200 85.200 165.000 ;
        RECT 86.000 164.200 86.800 165.000 ;
        RECT 90.800 166.200 91.600 167.000 ;
        RECT 94.000 166.200 94.800 167.000 ;
        RECT 95.600 164.200 96.400 165.000 ;
        RECT 97.200 164.200 98.000 165.000 ;
        RECT 98.800 164.200 99.600 165.000 ;
        RECT 108.400 169.600 109.200 170.400 ;
        RECT 130.800 177.600 131.600 178.400 ;
        RECT 121.200 167.600 122.000 168.400 ;
        RECT 162.800 173.600 163.600 174.400 ;
        RECT 127.600 163.600 128.400 164.400 ;
        RECT 143.600 171.600 144.400 172.400 ;
        RECT 146.800 171.600 147.600 172.400 ;
        RECT 148.400 169.600 149.200 170.400 ;
        RECT 188.400 177.600 189.200 178.400 ;
        RECT 154.800 167.600 155.600 168.400 ;
        RECT 174.000 171.600 174.800 172.400 ;
        RECT 182.000 169.600 182.800 170.400 ;
        RECT 212.400 177.600 213.200 178.400 ;
        RECT 209.200 171.600 210.000 172.400 ;
        RECT 217.200 177.600 218.000 178.400 ;
        RECT 214.000 173.600 214.800 174.400 ;
        RECT 215.600 171.600 216.400 172.400 ;
        RECT 202.800 167.600 203.600 168.400 ;
        RECT 196.400 163.600 197.200 164.400 ;
        RECT 238.000 175.600 238.800 176.400 ;
        RECT 239.600 174.200 240.400 175.000 ;
        RECT 230.000 171.600 230.800 172.400 ;
        RECT 250.800 171.600 251.600 172.400 ;
        RECT 233.200 166.800 234.000 167.600 ;
        RECT 236.400 166.200 237.200 167.000 ;
        RECT 231.600 164.200 232.400 165.000 ;
        RECT 233.200 164.200 234.000 165.000 ;
        RECT 234.800 164.200 235.600 165.000 ;
        RECT 239.600 166.200 240.400 167.000 ;
        RECT 242.800 166.200 243.600 167.000 ;
        RECT 262.000 177.600 262.800 178.400 ;
        RECT 255.600 171.600 256.400 172.400 ;
        RECT 263.600 173.600 264.400 174.400 ;
        RECT 279.600 173.000 280.400 173.800 ;
        RECT 265.200 171.600 266.000 172.400 ;
        RECT 244.400 164.200 245.200 165.000 ;
        RECT 246.000 164.200 246.800 165.000 ;
        RECT 289.200 172.600 290.000 173.400 ;
        RECT 274.800 171.600 275.600 172.400 ;
        RECT 295.600 171.600 296.400 172.400 ;
        RECT 314.800 175.600 315.600 176.400 ;
        RECT 281.200 168.800 282.000 169.600 ;
        RECT 286.000 167.600 286.800 168.400 ;
        RECT 282.800 166.200 283.600 167.000 ;
        RECT 279.600 164.200 280.400 165.000 ;
        RECT 281.200 164.200 282.000 165.000 ;
        RECT 286.000 166.200 286.800 167.000 ;
        RECT 289.200 166.200 290.000 167.000 ;
        RECT 290.800 164.200 291.600 165.000 ;
        RECT 292.400 164.200 293.200 165.000 ;
        RECT 294.000 164.200 294.800 165.000 ;
        RECT 303.600 163.600 304.400 164.400 ;
        RECT 313.200 169.600 314.000 170.400 ;
        RECT 332.400 173.000 333.200 173.800 ;
        RECT 321.200 171.600 322.000 172.400 ;
        RECT 322.800 169.600 323.600 170.400 ;
        RECT 342.000 172.600 342.800 173.400 ;
        RECT 361.200 177.600 362.000 178.400 ;
        RECT 329.200 171.600 330.000 172.400 ;
        RECT 334.000 168.800 334.800 169.600 ;
        RECT 338.800 167.600 339.600 168.400 ;
        RECT 335.600 166.200 336.400 167.000 ;
        RECT 332.400 164.200 333.200 165.000 ;
        RECT 334.000 164.200 334.800 165.000 ;
        RECT 338.800 166.200 339.600 167.000 ;
        RECT 342.000 166.200 342.800 167.000 ;
        RECT 343.600 164.200 344.400 165.000 ;
        RECT 345.200 164.200 346.000 165.000 ;
        RECT 346.800 164.200 347.600 165.000 ;
        RECT 356.400 169.600 357.200 170.400 ;
        RECT 377.200 175.600 378.000 176.400 ;
        RECT 378.800 174.200 379.600 175.000 ;
        RECT 407.600 177.600 408.400 178.400 ;
        RECT 417.200 177.600 418.000 178.400 ;
        RECT 380.400 171.600 381.200 172.400 ;
        RECT 372.400 166.800 373.200 167.600 ;
        RECT 375.600 166.200 376.400 167.000 ;
        RECT 370.800 164.200 371.600 165.000 ;
        RECT 372.400 164.200 373.200 165.000 ;
        RECT 374.000 164.200 374.800 165.000 ;
        RECT 378.800 166.200 379.600 167.000 ;
        RECT 382.000 166.200 382.800 167.000 ;
        RECT 401.200 171.600 402.000 172.400 ;
        RECT 383.600 164.200 384.400 165.000 ;
        RECT 385.200 164.200 386.000 165.000 ;
        RECT 433.200 175.600 434.000 176.400 ;
        RECT 434.800 174.200 435.600 175.000 ;
        RECT 425.200 171.600 426.000 172.400 ;
        RECT 447.600 171.600 448.400 172.400 ;
        RECT 428.400 166.800 429.200 167.600 ;
        RECT 431.600 166.200 432.400 167.000 ;
        RECT 426.800 164.200 427.600 165.000 ;
        RECT 428.400 164.200 429.200 165.000 ;
        RECT 430.000 164.200 430.800 165.000 ;
        RECT 434.800 166.200 435.600 167.000 ;
        RECT 438.000 166.200 438.800 167.000 ;
        RECT 439.600 164.200 440.400 165.000 ;
        RECT 441.200 164.200 442.000 165.000 ;
        RECT 454.000 169.600 454.800 170.400 ;
        RECT 458.800 169.600 459.600 170.400 ;
        RECT 457.200 163.600 458.000 164.400 ;
        RECT 489.200 163.600 490.000 164.400 ;
        RECT 500.400 173.600 501.200 174.400 ;
        RECT 513.200 173.000 514.000 173.800 ;
        RECT 503.600 171.600 504.400 172.400 ;
        RECT 497.200 163.600 498.000 164.400 ;
        RECT 522.800 172.600 523.600 173.400 ;
        RECT 508.400 171.600 509.200 172.400 ;
        RECT 514.800 168.800 515.600 169.600 ;
        RECT 519.600 167.600 520.400 168.400 ;
        RECT 516.400 166.200 517.200 167.000 ;
        RECT 513.200 164.200 514.000 165.000 ;
        RECT 514.800 164.200 515.600 165.000 ;
        RECT 519.600 166.200 520.400 167.000 ;
        RECT 522.800 166.200 523.600 167.000 ;
        RECT 524.400 164.200 525.200 165.000 ;
        RECT 526.000 164.200 526.800 165.000 ;
        RECT 527.600 164.200 528.400 165.000 ;
        RECT 542.000 175.600 542.800 176.400 ;
        RECT 550.000 177.600 550.800 178.400 ;
        RECT 545.200 171.600 546.000 172.400 ;
        RECT 537.200 163.600 538.000 164.400 ;
        RECT 542.000 163.600 542.800 164.400 ;
        RECT 577.200 177.600 578.000 178.400 ;
        RECT 553.200 163.600 554.000 164.400 ;
        RECT 574.000 171.600 574.800 172.400 ;
        RECT 566.000 169.600 566.800 170.400 ;
        RECT 591.600 177.600 592.400 178.400 ;
        RECT 564.400 163.600 565.200 164.400 ;
        RECT 607.600 173.600 608.400 174.400 ;
        RECT 596.400 172.200 597.200 173.000 ;
        RECT 604.400 171.800 605.200 172.600 ;
        RECT 609.200 170.200 610.000 171.000 ;
        RECT 610.800 163.600 611.600 164.400 ;
        RECT 618.800 169.600 619.600 170.400 ;
        RECT 623.600 167.600 624.400 168.400 ;
        RECT 633.200 171.600 634.000 172.400 ;
        RECT 636.400 169.600 637.200 170.400 ;
        RECT 650.800 177.600 651.600 178.400 ;
        RECT 655.600 177.600 656.400 178.400 ;
        RECT 646.000 171.600 646.800 172.400 ;
        RECT 644.400 163.600 645.200 164.400 ;
        RECT 671.600 175.600 672.400 176.400 ;
        RECT 673.200 174.200 674.000 175.000 ;
        RECT 674.800 171.600 675.600 172.400 ;
        RECT 666.800 166.800 667.600 167.600 ;
        RECT 670.000 166.200 670.800 167.000 ;
        RECT 665.200 164.200 666.000 165.000 ;
        RECT 666.800 164.200 667.600 165.000 ;
        RECT 668.400 164.200 669.200 165.000 ;
        RECT 673.200 166.200 674.000 167.000 ;
        RECT 676.400 166.200 677.200 167.000 ;
        RECT 678.000 164.200 678.800 165.000 ;
        RECT 679.600 164.200 680.400 165.000 ;
        RECT 6.000 149.600 6.800 150.400 ;
        RECT 39.600 157.600 40.400 158.400 ;
        RECT 14.000 149.600 14.800 150.400 ;
        RECT 18.800 147.600 19.600 148.400 ;
        RECT 2.800 145.600 3.600 146.400 ;
        RECT 22.000 149.600 22.800 150.400 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 31.600 149.600 32.400 150.400 ;
        RECT 39.600 149.600 40.400 150.400 ;
        RECT 25.200 143.600 26.000 144.400 ;
        RECT 41.200 147.600 42.000 148.400 ;
        RECT 49.200 149.600 50.000 150.400 ;
        RECT 50.800 149.600 51.600 150.400 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 58.800 149.600 59.600 150.400 ;
        RECT 60.400 149.600 61.200 150.400 ;
        RECT 63.600 149.600 64.400 150.400 ;
        RECT 90.800 157.600 91.600 158.400 ;
        RECT 71.600 149.600 72.400 150.400 ;
        RECT 66.800 147.600 67.600 148.400 ;
        RECT 73.200 147.600 74.000 148.400 ;
        RECT 79.600 149.600 80.400 150.400 ;
        RECT 82.800 149.600 83.600 150.400 ;
        RECT 94.000 153.600 94.800 154.400 ;
        RECT 90.800 149.600 91.600 150.400 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 108.400 152.400 109.200 153.200 ;
        RECT 111.600 151.000 112.400 151.800 ;
        RECT 118.000 149.600 118.800 150.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 137.200 157.600 138.000 158.400 ;
        RECT 130.800 149.600 131.600 150.400 ;
        RECT 111.600 146.200 112.400 147.000 ;
        RECT 140.400 149.600 141.200 150.400 ;
        RECT 142.000 149.600 142.800 150.400 ;
        RECT 151.600 149.600 152.400 150.400 ;
        RECT 159.600 149.600 160.400 150.400 ;
        RECT 146.800 147.600 147.600 148.400 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 161.200 147.600 162.000 148.400 ;
        RECT 164.400 147.600 165.200 148.400 ;
        RECT 162.800 146.200 163.600 147.000 ;
        RECT 182.000 145.600 182.800 146.400 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 186.800 149.600 187.600 150.400 ;
        RECT 194.800 149.600 195.600 150.400 ;
        RECT 196.400 149.600 197.200 150.400 ;
        RECT 183.600 143.600 184.400 144.400 ;
        RECT 206.000 149.600 206.800 150.400 ;
        RECT 217.200 153.600 218.000 154.400 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 215.600 147.600 216.400 148.400 ;
        RECT 231.600 152.400 232.400 153.200 ;
        RECT 234.800 151.000 235.600 151.800 ;
        RECT 241.200 157.600 242.000 158.400 ;
        RECT 236.400 149.600 237.200 150.400 ;
        RECT 238.000 149.600 238.800 150.400 ;
        RECT 246.000 149.600 246.800 150.400 ;
        RECT 247.600 149.600 248.400 150.400 ;
        RECT 257.400 151.800 258.200 152.600 ;
        RECT 258.600 149.800 259.400 150.600 ;
        RECT 234.800 146.200 235.600 147.000 ;
        RECT 289.200 155.000 290.000 155.800 ;
        RECT 286.000 153.600 286.800 154.400 ;
        RECT 290.800 152.400 291.600 153.200 ;
        RECT 274.800 151.600 275.600 152.400 ;
        RECT 311.600 153.600 312.400 154.400 ;
        RECT 257.400 146.200 258.200 147.000 ;
        RECT 265.200 147.600 266.000 148.400 ;
        RECT 279.600 148.200 280.400 149.000 ;
        RECT 289.200 148.600 290.000 149.400 ;
        RECT 284.400 147.600 285.200 148.400 ;
        RECT 330.800 155.000 331.600 155.800 ;
        RECT 327.600 153.600 328.400 154.400 ;
        RECT 332.400 152.400 333.200 153.200 ;
        RECT 345.200 153.600 346.000 154.400 ;
        RECT 337.200 149.600 338.000 150.400 ;
        RECT 303.800 147.600 304.600 148.400 ;
        RECT 321.200 148.200 322.000 149.000 ;
        RECT 330.800 148.600 331.600 149.400 ;
        RECT 279.600 144.200 280.400 145.000 ;
        RECT 281.200 144.200 282.000 145.000 ;
        RECT 282.800 144.200 283.600 145.000 ;
        RECT 286.000 144.200 286.800 145.000 ;
        RECT 289.200 144.200 290.000 145.000 ;
        RECT 290.800 144.200 291.600 145.000 ;
        RECT 292.400 144.200 293.200 145.000 ;
        RECT 294.000 144.200 294.800 145.000 ;
        RECT 311.600 143.600 312.400 144.400 ;
        RECT 326.000 147.600 326.800 148.400 ;
        RECT 321.200 144.200 322.000 145.000 ;
        RECT 322.800 144.200 323.600 145.000 ;
        RECT 324.400 144.200 325.200 145.000 ;
        RECT 327.600 144.200 328.400 145.000 ;
        RECT 330.800 144.200 331.600 145.000 ;
        RECT 332.400 144.200 333.200 145.000 ;
        RECT 334.000 144.200 334.800 145.000 ;
        RECT 335.600 144.200 336.400 145.000 ;
        RECT 361.200 154.400 362.000 155.200 ;
        RECT 364.400 155.000 365.200 155.800 ;
        RECT 359.600 152.400 360.400 153.200 ;
        RECT 358.000 149.600 358.800 150.400 ;
        RECT 369.200 147.600 370.000 148.400 ;
        RECT 366.000 145.600 366.800 146.400 ;
        RECT 359.600 144.200 360.400 145.000 ;
        RECT 361.200 144.200 362.000 145.000 ;
        RECT 362.800 144.200 363.600 145.000 ;
        RECT 364.400 144.200 365.200 145.000 ;
        RECT 367.600 144.200 368.400 145.000 ;
        RECT 370.800 144.200 371.600 145.000 ;
        RECT 372.400 144.200 373.200 145.000 ;
        RECT 374.000 144.200 374.800 145.000 ;
        RECT 401.200 155.000 402.000 155.800 ;
        RECT 398.000 153.600 398.800 154.400 ;
        RECT 402.800 152.400 403.600 153.200 ;
        RECT 407.600 149.600 408.400 150.400 ;
        RECT 391.600 148.200 392.400 149.000 ;
        RECT 401.200 148.600 402.000 149.400 ;
        RECT 396.400 147.600 397.200 148.400 ;
        RECT 391.600 144.200 392.400 145.000 ;
        RECT 393.200 144.200 394.000 145.000 ;
        RECT 394.800 144.200 395.600 145.000 ;
        RECT 398.000 144.200 398.800 145.000 ;
        RECT 401.200 144.200 402.000 145.000 ;
        RECT 402.800 144.200 403.600 145.000 ;
        RECT 404.400 144.200 405.200 145.000 ;
        RECT 406.000 144.200 406.800 145.000 ;
        RECT 415.600 145.600 416.400 146.400 ;
        RECT 428.400 149.600 429.200 150.400 ;
        RECT 425.200 145.600 426.000 146.400 ;
        RECT 455.600 155.000 456.400 155.800 ;
        RECT 452.400 153.600 453.200 154.400 ;
        RECT 457.200 152.400 458.000 153.200 ;
        RECT 473.200 157.600 474.000 158.400 ;
        RECT 462.000 149.600 462.800 150.400 ;
        RECT 446.000 148.200 446.800 149.000 ;
        RECT 455.600 148.600 456.400 149.400 ;
        RECT 450.800 147.600 451.600 148.400 ;
        RECT 446.000 144.200 446.800 145.000 ;
        RECT 447.600 144.200 448.400 145.000 ;
        RECT 449.200 144.200 450.000 145.000 ;
        RECT 452.400 144.200 453.200 145.000 ;
        RECT 455.600 144.200 456.400 145.000 ;
        RECT 457.200 144.200 458.000 145.000 ;
        RECT 458.800 144.200 459.600 145.000 ;
        RECT 460.400 144.200 461.200 145.000 ;
        RECT 470.000 145.600 470.800 146.400 ;
        RECT 494.000 155.000 494.800 155.800 ;
        RECT 490.800 153.600 491.600 154.400 ;
        RECT 508.400 157.600 509.200 158.400 ;
        RECT 495.600 152.400 496.400 153.200 ;
        RECT 484.400 148.200 485.200 149.000 ;
        RECT 494.000 148.600 494.800 149.400 ;
        RECT 474.800 145.600 475.600 146.400 ;
        RECT 489.200 147.600 490.000 148.400 ;
        RECT 484.400 144.200 485.200 145.000 ;
        RECT 486.000 144.200 486.800 145.000 ;
        RECT 487.600 144.200 488.400 145.000 ;
        RECT 490.800 144.200 491.600 145.000 ;
        RECT 494.000 144.200 494.800 145.000 ;
        RECT 495.600 144.200 496.400 145.000 ;
        RECT 497.200 144.200 498.000 145.000 ;
        RECT 498.800 144.200 499.600 145.000 ;
        RECT 518.000 157.600 518.800 158.400 ;
        RECT 518.000 149.600 518.800 150.400 ;
        RECT 522.800 149.600 523.600 150.400 ;
        RECT 540.400 157.600 541.200 158.400 ;
        RECT 530.800 149.600 531.600 150.400 ;
        RECT 519.600 147.600 520.400 148.400 ;
        RECT 532.400 147.600 533.200 148.400 ;
        RECT 526.000 143.600 526.800 144.400 ;
        RECT 534.000 145.600 534.800 146.400 ;
        RECT 538.800 145.600 539.600 146.400 ;
        RECT 535.600 143.600 536.400 144.400 ;
        RECT 550.000 147.600 550.800 148.400 ;
        RECT 546.800 143.600 547.600 144.400 ;
        RECT 548.400 145.600 549.200 146.400 ;
        RECT 558.000 157.600 558.800 158.400 ;
        RECT 561.200 149.600 562.000 150.400 ;
        RECT 577.200 149.600 578.000 150.400 ;
        RECT 582.000 149.600 582.800 150.400 ;
        RECT 590.000 149.600 590.800 150.400 ;
        RECT 593.200 149.600 594.000 150.400 ;
        RECT 594.800 149.600 595.600 150.400 ;
        RECT 567.600 147.600 568.400 148.400 ;
        RECT 578.800 147.600 579.600 148.400 ;
        RECT 591.600 147.600 592.400 148.400 ;
        RECT 617.200 157.600 618.000 158.400 ;
        RECT 586.800 143.600 587.600 144.400 ;
        RECT 610.800 149.600 611.600 150.400 ;
        RECT 623.600 153.600 624.400 154.400 ;
        RECT 631.600 157.600 632.400 158.400 ;
        RECT 620.400 149.600 621.200 150.400 ;
        RECT 626.800 151.600 627.600 152.400 ;
        RECT 638.000 157.600 638.800 158.400 ;
        RECT 641.200 155.600 642.000 156.400 ;
        RECT 625.200 149.600 626.000 150.400 ;
        RECT 606.000 143.600 606.800 144.400 ;
        RECT 614.000 143.600 614.800 144.400 ;
        RECT 617.200 143.600 618.000 144.400 ;
        RECT 631.600 143.600 632.400 144.400 ;
        RECT 638.000 143.600 638.800 144.400 ;
        RECT 644.400 149.600 645.200 150.400 ;
        RECT 646.000 149.600 646.800 150.400 ;
        RECT 654.000 149.600 654.800 150.400 ;
        RECT 655.600 149.600 656.400 150.400 ;
        RECT 670.000 153.600 670.800 154.400 ;
        RECT 642.800 145.600 643.600 146.400 ;
        RECT 684.400 152.400 685.200 153.200 ;
        RECT 687.600 151.000 688.400 151.800 ;
        RECT 682.800 145.600 683.600 146.400 ;
        RECT 687.600 146.200 688.400 147.000 ;
        RECT 26.800 137.600 27.600 138.400 ;
        RECT 1.200 130.200 2.000 131.000 ;
        RECT 50.800 137.600 51.600 138.400 ;
        RECT 23.600 129.600 24.400 130.400 ;
        RECT 33.200 130.200 34.000 131.000 ;
        RECT 18.800 123.600 19.600 124.400 ;
        RECT 47.600 127.600 48.400 128.400 ;
        RECT 57.200 129.600 58.000 130.400 ;
        RECT 66.800 131.600 67.600 132.400 ;
        RECT 92.400 131.600 93.200 132.400 ;
        RECT 108.400 133.600 109.200 134.400 ;
        RECT 159.600 137.600 160.400 138.400 ;
        RECT 95.600 123.600 96.400 124.400 ;
        RECT 121.200 129.600 122.000 130.400 ;
        RECT 126.000 123.600 126.800 124.400 ;
        RECT 134.000 123.600 134.800 124.400 ;
        RECT 167.600 137.600 168.400 138.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 146.800 129.600 147.600 130.400 ;
        RECT 159.600 129.600 160.400 130.400 ;
        RECT 172.400 133.600 173.200 134.400 ;
        RECT 178.800 133.600 179.600 134.400 ;
        RECT 174.000 131.600 174.800 132.400 ;
        RECT 183.600 129.600 184.400 130.400 ;
        RECT 191.600 129.600 192.400 130.400 ;
        RECT 218.800 135.600 219.600 136.400 ;
        RECT 220.400 134.200 221.200 135.000 ;
        RECT 230.000 131.600 230.800 132.400 ;
        RECT 199.600 129.600 200.400 130.400 ;
        RECT 202.800 123.600 203.600 124.400 ;
        RECT 214.000 126.800 214.800 127.600 ;
        RECT 217.200 126.200 218.000 127.000 ;
        RECT 212.400 124.200 213.200 125.000 ;
        RECT 214.000 124.200 214.800 125.000 ;
        RECT 215.600 124.200 216.400 125.000 ;
        RECT 220.400 126.200 221.200 127.000 ;
        RECT 223.600 126.200 224.400 127.000 ;
        RECT 242.800 137.600 243.600 138.400 ;
        RECT 239.600 131.600 240.400 132.400 ;
        RECT 268.400 137.600 269.200 138.400 ;
        RECT 274.800 135.600 275.600 136.400 ;
        RECT 246.000 133.600 246.800 134.400 ;
        RECT 249.200 131.600 250.000 132.400 ;
        RECT 225.200 124.200 226.000 125.000 ;
        RECT 226.800 124.200 227.600 125.000 ;
        RECT 236.400 123.600 237.200 124.400 ;
        RECT 250.800 123.600 251.600 124.400 ;
        RECT 303.600 137.600 304.400 138.400 ;
        RECT 271.600 131.600 272.400 132.400 ;
        RECT 279.600 129.600 280.400 130.400 ;
        RECT 290.800 129.600 291.600 130.400 ;
        RECT 300.400 129.600 301.200 130.400 ;
        RECT 302.000 129.600 302.800 130.400 ;
        RECT 324.400 135.600 325.200 136.400 ;
        RECT 326.000 134.200 326.800 135.000 ;
        RECT 337.200 131.600 338.000 132.400 ;
        RECT 308.400 129.600 309.200 130.400 ;
        RECT 319.600 126.800 320.400 127.600 ;
        RECT 322.800 126.200 323.600 127.000 ;
        RECT 318.000 124.200 318.800 125.000 ;
        RECT 319.600 124.200 320.400 125.000 ;
        RECT 321.200 124.200 322.000 125.000 ;
        RECT 326.000 126.200 326.800 127.000 ;
        RECT 329.200 126.200 330.000 127.000 ;
        RECT 342.000 131.600 342.800 132.400 ;
        RECT 359.600 133.000 360.400 133.800 ;
        RECT 350.000 131.600 350.800 132.400 ;
        RECT 330.800 124.200 331.600 125.000 ;
        RECT 332.400 124.200 333.200 125.000 ;
        RECT 369.200 132.600 370.000 133.400 ;
        RECT 375.600 131.600 376.400 132.400 ;
        RECT 361.200 128.800 362.000 129.600 ;
        RECT 366.000 127.600 366.800 128.400 ;
        RECT 350.000 123.600 350.800 124.400 ;
        RECT 362.800 126.200 363.600 127.000 ;
        RECT 359.600 124.200 360.400 125.000 ;
        RECT 361.200 124.200 362.000 125.000 ;
        RECT 366.000 126.200 366.800 127.000 ;
        RECT 369.200 126.200 370.000 127.000 ;
        RECT 370.800 124.200 371.600 125.000 ;
        RECT 372.400 124.200 373.200 125.000 ;
        RECT 374.000 124.200 374.800 125.000 ;
        RECT 394.800 137.600 395.600 138.400 ;
        RECT 391.600 131.600 392.400 132.400 ;
        RECT 410.800 135.600 411.600 136.400 ;
        RECT 412.400 134.200 413.200 135.000 ;
        RECT 402.800 131.600 403.600 132.400 ;
        RECT 423.600 131.600 424.400 132.400 ;
        RECT 383.600 123.600 384.400 124.400 ;
        RECT 388.400 123.600 389.200 124.400 ;
        RECT 406.000 126.800 406.800 127.600 ;
        RECT 409.200 126.200 410.000 127.000 ;
        RECT 404.400 124.200 405.200 125.000 ;
        RECT 406.000 124.200 406.800 125.000 ;
        RECT 407.600 124.200 408.400 125.000 ;
        RECT 412.400 126.200 413.200 127.000 ;
        RECT 415.600 126.200 416.400 127.000 ;
        RECT 417.200 124.200 418.000 125.000 ;
        RECT 418.800 124.200 419.600 125.000 ;
        RECT 449.200 133.000 450.000 133.800 ;
        RECT 458.800 132.600 459.600 133.400 ;
        RECT 473.200 137.600 474.000 138.400 ;
        RECT 444.400 131.600 445.200 132.400 ;
        RECT 450.800 128.800 451.600 129.600 ;
        RECT 455.600 127.600 456.400 128.400 ;
        RECT 439.600 123.600 440.400 124.400 ;
        RECT 452.400 126.200 453.200 127.000 ;
        RECT 449.200 124.200 450.000 125.000 ;
        RECT 450.800 124.200 451.600 125.000 ;
        RECT 455.600 126.200 456.400 127.000 ;
        RECT 458.800 126.200 459.600 127.000 ;
        RECT 460.400 124.200 461.200 125.000 ;
        RECT 462.000 124.200 462.800 125.000 ;
        RECT 463.600 124.200 464.400 125.000 ;
        RECT 484.400 133.000 485.200 133.800 ;
        RECT 494.000 132.600 494.800 133.400 ;
        RECT 508.400 137.600 509.200 138.400 ;
        RECT 511.600 137.600 512.400 138.400 ;
        RECT 500.400 131.600 501.200 132.400 ;
        RECT 486.000 128.800 486.800 129.600 ;
        RECT 490.800 127.600 491.600 128.400 ;
        RECT 473.200 123.600 474.000 124.400 ;
        RECT 487.600 126.200 488.400 127.000 ;
        RECT 484.400 124.200 485.200 125.000 ;
        RECT 486.000 124.200 486.800 125.000 ;
        RECT 490.800 126.200 491.600 127.000 ;
        RECT 494.000 126.200 494.800 127.000 ;
        RECT 495.600 124.200 496.400 125.000 ;
        RECT 497.200 124.200 498.000 125.000 ;
        RECT 498.800 124.200 499.600 125.000 ;
        RECT 534.000 133.600 534.800 134.400 ;
        RECT 522.800 132.200 523.600 133.000 ;
        RECT 530.800 131.800 531.600 132.600 ;
        RECT 535.600 130.200 536.400 131.000 ;
        RECT 546.800 131.600 547.600 132.400 ;
        RECT 518.000 127.600 518.800 128.400 ;
        RECT 559.600 131.600 560.400 132.400 ;
        RECT 561.200 130.200 562.000 131.000 ;
        RECT 585.200 129.600 586.000 130.400 ;
        RECT 596.400 137.600 597.200 138.400 ;
        RECT 625.200 137.600 626.000 138.400 ;
        RECT 593.200 131.600 594.000 132.400 ;
        RECT 609.200 131.600 610.000 132.400 ;
        RECT 617.200 133.600 618.000 134.400 ;
        RECT 641.200 133.600 642.000 134.400 ;
        RECT 630.000 132.200 630.800 133.000 ;
        RECT 617.200 129.600 618.000 130.400 ;
        RECT 642.800 130.200 643.600 131.000 ;
        RECT 670.000 137.600 670.800 138.400 ;
        RECT 644.400 127.600 645.200 128.400 ;
        RECT 654.000 131.600 654.800 132.400 ;
        RECT 674.800 132.200 675.600 133.000 ;
        RECT 652.400 123.600 653.200 124.400 ;
        RECT 668.400 129.600 669.200 130.400 ;
        RECT 687.600 130.200 688.400 131.000 ;
        RECT 1.200 106.200 2.000 107.000 ;
        RECT 25.200 109.600 26.000 110.400 ;
        RECT 26.800 109.600 27.600 110.400 ;
        RECT 28.400 109.600 29.200 110.400 ;
        RECT 46.000 117.600 46.800 118.400 ;
        RECT 18.800 103.600 19.600 104.400 ;
        RECT 22.000 103.600 22.800 104.400 ;
        RECT 66.800 113.600 67.600 114.400 ;
        RECT 55.600 109.600 56.400 110.400 ;
        RECT 73.200 117.600 74.000 118.400 ;
        RECT 50.800 107.600 51.600 108.400 ;
        RECT 49.200 106.200 50.000 107.000 ;
        RECT 46.000 103.600 46.800 104.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 70.000 109.600 70.800 110.400 ;
        RECT 78.000 105.600 78.800 106.400 ;
        RECT 98.800 117.600 99.600 118.400 ;
        RECT 87.600 109.600 88.400 110.400 ;
        RECT 79.600 103.600 80.400 104.400 ;
        RECT 81.200 106.200 82.000 107.000 ;
        RECT 102.000 109.600 102.800 110.400 ;
        RECT 111.600 107.600 112.400 108.400 ;
        RECT 124.400 107.600 125.200 108.400 ;
        RECT 130.800 109.600 131.600 110.400 ;
        RECT 138.800 109.600 139.600 110.400 ;
        RECT 142.000 109.600 142.800 110.400 ;
        RECT 143.600 109.600 144.400 110.400 ;
        RECT 146.800 109.600 147.600 110.400 ;
        RECT 169.200 117.600 170.000 118.400 ;
        RECT 153.200 107.600 154.000 108.400 ;
        RECT 134.000 105.600 134.800 106.400 ;
        RECT 151.600 106.200 152.400 107.000 ;
        RECT 175.600 109.600 176.400 110.400 ;
        RECT 199.600 117.600 200.400 118.400 ;
        RECT 193.200 111.600 194.000 112.400 ;
        RECT 193.200 109.600 194.000 110.400 ;
        RECT 199.600 109.600 200.400 110.400 ;
        RECT 218.800 117.600 219.600 118.400 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 186.800 105.600 187.600 106.400 ;
        RECT 194.800 107.600 195.600 108.400 ;
        RECT 201.200 107.600 202.000 108.400 ;
        RECT 202.800 105.600 203.600 106.400 ;
        RECT 204.400 103.600 205.200 104.400 ;
        RECT 210.800 107.600 211.600 108.400 ;
        RECT 212.400 105.600 213.200 106.400 ;
        RECT 223.600 117.600 224.400 118.400 ;
        RECT 217.200 107.600 218.000 108.400 ;
        RECT 220.400 105.600 221.200 106.400 ;
        RECT 225.200 105.600 226.000 106.400 ;
        RECT 241.200 109.600 242.000 110.400 ;
        RECT 252.400 109.600 253.200 110.400 ;
        RECT 268.400 113.600 269.200 114.400 ;
        RECT 279.600 114.400 280.400 115.200 ;
        RECT 282.800 115.000 283.600 115.800 ;
        RECT 278.000 112.400 278.800 113.200 ;
        RECT 249.200 103.600 250.000 104.400 ;
        RECT 287.600 107.600 288.400 108.400 ;
        RECT 284.400 105.600 285.200 106.400 ;
        RECT 278.000 104.200 278.800 105.000 ;
        RECT 279.600 104.200 280.400 105.000 ;
        RECT 281.200 104.200 282.000 105.000 ;
        RECT 282.800 104.200 283.600 105.000 ;
        RECT 286.000 104.200 286.800 105.000 ;
        RECT 289.200 104.200 290.000 105.000 ;
        RECT 290.800 104.200 291.600 105.000 ;
        RECT 292.400 104.200 293.200 105.000 ;
        RECT 308.400 109.600 309.200 110.400 ;
        RECT 311.600 107.600 312.400 108.400 ;
        RECT 313.200 117.600 314.000 118.400 ;
        RECT 318.000 109.600 318.800 110.400 ;
        RECT 314.800 105.600 315.600 106.400 ;
        RECT 329.200 113.600 330.000 114.400 ;
        RECT 340.400 114.400 341.200 115.200 ;
        RECT 343.600 115.000 344.400 115.800 ;
        RECT 364.400 117.600 365.200 118.400 ;
        RECT 338.800 112.400 339.600 113.200 ;
        RECT 337.200 109.600 338.000 110.400 ;
        RECT 348.400 107.600 349.200 108.400 ;
        RECT 345.200 105.600 346.000 106.400 ;
        RECT 338.800 104.200 339.600 105.000 ;
        RECT 340.400 104.200 341.200 105.000 ;
        RECT 342.000 104.200 342.800 105.000 ;
        RECT 343.600 104.200 344.400 105.000 ;
        RECT 346.800 104.200 347.600 105.000 ;
        RECT 350.000 104.200 350.800 105.000 ;
        RECT 351.600 104.200 352.400 105.000 ;
        RECT 353.200 104.200 354.000 105.000 ;
        RECT 375.600 114.400 376.400 115.200 ;
        RECT 378.800 115.000 379.600 115.800 ;
        RECT 374.000 112.400 374.800 113.200 ;
        RECT 372.400 109.600 373.200 110.400 ;
        RECT 364.400 103.600 365.200 104.400 ;
        RECT 383.600 107.600 384.400 108.400 ;
        RECT 380.400 105.600 381.200 106.400 ;
        RECT 374.000 104.200 374.800 105.000 ;
        RECT 375.600 104.200 376.400 105.000 ;
        RECT 377.200 104.200 378.000 105.000 ;
        RECT 378.800 104.200 379.600 105.000 ;
        RECT 382.000 104.200 382.800 105.000 ;
        RECT 385.200 104.200 386.000 105.000 ;
        RECT 386.800 104.200 387.600 105.000 ;
        RECT 388.400 104.200 389.200 105.000 ;
        RECT 409.200 117.600 410.000 118.400 ;
        RECT 404.400 109.600 405.200 110.400 ;
        RECT 398.000 107.600 398.800 108.400 ;
        RECT 402.800 107.600 403.600 108.400 ;
        RECT 399.600 105.600 400.400 106.400 ;
        RECT 406.000 107.600 406.800 108.400 ;
        RECT 407.600 107.600 408.400 108.400 ;
        RECT 425.200 115.600 426.000 116.400 ;
        RECT 436.400 114.400 437.200 115.200 ;
        RECT 439.600 115.000 440.400 115.800 ;
        RECT 434.800 112.400 435.600 113.200 ;
        RECT 415.600 109.600 416.400 110.400 ;
        RECT 417.200 107.600 418.000 108.400 ;
        RECT 433.200 109.600 434.000 110.400 ;
        RECT 412.400 103.600 413.200 104.400 ;
        RECT 444.400 107.600 445.200 108.400 ;
        RECT 441.200 105.600 442.000 106.400 ;
        RECT 434.800 104.200 435.600 105.000 ;
        RECT 436.400 104.200 437.200 105.000 ;
        RECT 438.000 104.200 438.800 105.000 ;
        RECT 439.600 104.200 440.400 105.000 ;
        RECT 442.800 104.200 443.600 105.000 ;
        RECT 446.000 104.200 446.800 105.000 ;
        RECT 447.600 104.200 448.400 105.000 ;
        RECT 449.200 104.200 450.000 105.000 ;
        RECT 463.600 109.600 464.400 110.400 ;
        RECT 466.800 109.600 467.600 110.400 ;
        RECT 470.000 107.600 470.800 108.400 ;
        RECT 471.600 107.600 472.400 108.400 ;
        RECT 476.400 107.600 477.200 108.400 ;
        RECT 482.800 115.600 483.600 116.400 ;
        RECT 494.000 114.400 494.800 115.200 ;
        RECT 497.200 115.000 498.000 115.800 ;
        RECT 492.400 112.400 493.200 113.200 ;
        RECT 490.800 109.600 491.600 110.400 ;
        RECT 474.800 103.600 475.600 104.400 ;
        RECT 502.000 107.600 502.800 108.400 ;
        RECT 498.800 105.600 499.600 106.400 ;
        RECT 526.000 113.600 526.800 114.400 ;
        RECT 492.400 104.200 493.200 105.000 ;
        RECT 494.000 104.200 494.800 105.000 ;
        RECT 495.600 104.200 496.400 105.000 ;
        RECT 497.200 104.200 498.000 105.000 ;
        RECT 500.400 104.200 501.200 105.000 ;
        RECT 503.600 104.200 504.400 105.000 ;
        RECT 505.200 104.200 506.000 105.000 ;
        RECT 506.800 104.200 507.600 105.000 ;
        RECT 521.200 109.600 522.000 110.400 ;
        RECT 526.000 109.600 526.800 110.400 ;
        RECT 551.600 111.600 552.400 112.400 ;
        RECT 527.600 107.600 528.400 108.400 ;
        RECT 546.800 109.600 547.600 110.400 ;
        RECT 548.400 107.600 549.200 108.400 ;
        RECT 550.000 107.600 550.800 108.400 ;
        RECT 577.200 117.600 578.000 118.400 ;
        RECT 561.200 109.600 562.000 110.400 ;
        RECT 562.800 109.600 563.600 110.400 ;
        RECT 586.800 117.600 587.600 118.400 ;
        RECT 567.600 103.600 568.400 104.400 ;
        RECT 586.800 109.600 587.600 110.400 ;
        RECT 582.000 105.600 582.800 106.400 ;
        RECT 588.400 107.600 589.200 108.400 ;
        RECT 599.600 107.600 600.400 108.400 ;
        RECT 604.400 115.600 605.200 116.400 ;
        RECT 618.800 112.400 619.600 113.200 ;
        RECT 622.000 111.000 622.800 111.800 ;
        RECT 625.200 109.600 626.000 110.400 ;
        RECT 636.400 109.600 637.200 110.400 ;
        RECT 638.000 109.600 638.800 110.400 ;
        RECT 601.200 103.600 602.000 104.400 ;
        RECT 622.000 106.200 622.800 107.000 ;
        RECT 634.800 107.600 635.600 108.400 ;
        RECT 660.400 117.600 661.200 118.400 ;
        RECT 647.600 105.600 648.400 106.400 ;
        RECT 657.200 109.600 658.000 110.400 ;
        RECT 674.800 109.600 675.600 110.400 ;
        RECT 679.600 109.600 680.400 110.400 ;
        RECT 681.200 109.600 682.000 110.400 ;
        RECT 654.000 103.600 654.800 104.400 ;
        RECT 678.000 103.600 678.800 104.400 ;
        RECT 1.200 97.600 2.000 98.400 ;
        RECT 34.800 97.600 35.600 98.400 ;
        RECT 9.200 91.600 10.000 92.400 ;
        RECT 71.600 97.600 72.400 98.400 ;
        RECT 26.800 85.600 27.600 86.400 ;
        RECT 34.800 89.600 35.600 90.400 ;
        RECT 41.200 89.600 42.000 90.400 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 52.400 87.600 53.200 88.400 ;
        RECT 70.000 91.600 70.800 92.400 ;
        RECT 87.600 93.600 88.400 94.400 ;
        RECT 76.400 92.200 77.200 93.000 ;
        RECT 92.400 91.600 93.200 92.400 ;
        RECT 121.200 97.600 122.000 98.400 ;
        RECT 89.200 90.200 90.000 91.000 ;
        RECT 126.000 91.600 126.800 92.400 ;
        RECT 97.200 87.600 98.000 88.400 ;
        RECT 110.000 83.600 110.800 84.400 ;
        RECT 174.000 97.600 174.800 98.400 ;
        RECT 177.200 97.600 178.000 98.400 ;
        RECT 146.800 91.600 147.600 92.400 ;
        RECT 129.200 83.600 130.000 84.400 ;
        RECT 138.800 89.600 139.600 90.400 ;
        RECT 143.600 89.600 144.400 90.400 ;
        RECT 156.400 91.800 157.200 92.600 ;
        RECT 151.600 90.200 152.400 91.000 ;
        RECT 148.400 87.600 149.200 88.400 ;
        RECT 169.200 83.600 170.000 84.400 ;
        RECT 193.200 95.600 194.000 96.400 ;
        RECT 194.800 94.200 195.600 95.000 ;
        RECT 214.000 97.600 214.800 98.400 ;
        RECT 223.600 97.600 224.400 98.400 ;
        RECT 206.000 91.600 206.800 92.400 ;
        RECT 174.000 89.600 174.800 90.400 ;
        RECT 188.400 86.800 189.200 87.600 ;
        RECT 191.600 86.200 192.400 87.000 ;
        RECT 186.800 84.200 187.600 85.000 ;
        RECT 188.400 84.200 189.200 85.000 ;
        RECT 190.000 84.200 190.800 85.000 ;
        RECT 194.800 86.200 195.600 87.000 ;
        RECT 198.000 86.200 198.800 87.000 ;
        RECT 199.600 84.200 200.400 85.000 ;
        RECT 201.200 84.200 202.000 85.000 ;
        RECT 220.400 89.600 221.200 90.400 ;
        RECT 230.000 97.600 230.800 98.400 ;
        RECT 225.200 93.600 226.000 94.400 ;
        RECT 255.600 97.600 256.400 98.400 ;
        RECT 238.000 94.800 238.800 95.600 ;
        RECT 271.600 95.600 272.400 96.400 ;
        RECT 273.200 94.200 274.000 95.000 ;
        RECT 292.400 97.600 293.200 98.400 ;
        RECT 263.600 91.600 264.400 92.400 ;
        RECT 238.000 83.600 238.800 84.400 ;
        RECT 266.800 86.800 267.600 87.600 ;
        RECT 270.000 86.200 270.800 87.000 ;
        RECT 265.200 84.200 266.000 85.000 ;
        RECT 266.800 84.200 267.600 85.000 ;
        RECT 268.400 84.200 269.200 85.000 ;
        RECT 273.200 86.200 274.000 87.000 ;
        RECT 276.400 86.200 277.200 87.000 ;
        RECT 278.000 84.200 278.800 85.000 ;
        RECT 279.600 84.200 280.400 85.000 ;
        RECT 324.400 95.600 325.200 96.400 ;
        RECT 326.000 94.200 326.800 95.000 ;
        RECT 316.400 91.600 317.200 92.400 ;
        RECT 337.200 91.600 338.000 92.400 ;
        RECT 305.200 89.600 306.000 90.400 ;
        RECT 308.400 89.600 309.200 90.400 ;
        RECT 319.600 86.800 320.400 87.600 ;
        RECT 322.800 86.200 323.600 87.000 ;
        RECT 318.000 84.200 318.800 85.000 ;
        RECT 319.600 84.200 320.400 85.000 ;
        RECT 321.200 84.200 322.000 85.000 ;
        RECT 326.000 86.200 326.800 87.000 ;
        RECT 329.200 86.200 330.000 87.000 ;
        RECT 330.800 84.200 331.600 85.000 ;
        RECT 332.400 84.200 333.200 85.000 ;
        RECT 353.200 93.000 354.000 93.800 ;
        RECT 362.800 92.600 363.600 93.400 ;
        RECT 369.200 91.600 370.000 92.400 ;
        RECT 390.000 95.600 390.800 96.400 ;
        RECT 354.800 88.800 355.600 89.600 ;
        RECT 359.600 87.600 360.400 88.400 ;
        RECT 343.600 83.600 344.400 84.400 ;
        RECT 356.400 86.200 357.200 87.000 ;
        RECT 353.200 84.200 354.000 85.000 ;
        RECT 354.800 84.200 355.600 85.000 ;
        RECT 359.600 86.200 360.400 87.000 ;
        RECT 362.800 86.200 363.600 87.000 ;
        RECT 364.400 84.200 365.200 85.000 ;
        RECT 366.000 84.200 366.800 85.000 ;
        RECT 367.600 84.200 368.400 85.000 ;
        RECT 377.200 83.600 378.000 84.400 ;
        RECT 390.000 89.600 390.800 90.400 ;
        RECT 425.200 95.600 426.000 96.400 ;
        RECT 426.800 94.200 427.600 95.000 ;
        RECT 465.200 97.600 466.000 98.400 ;
        RECT 438.000 91.600 438.800 92.400 ;
        RECT 401.200 89.600 402.000 90.400 ;
        RECT 409.200 89.600 410.000 90.400 ;
        RECT 399.600 83.600 400.400 84.400 ;
        RECT 420.400 86.800 421.200 87.600 ;
        RECT 423.600 86.200 424.400 87.000 ;
        RECT 418.800 84.200 419.600 85.000 ;
        RECT 420.400 84.200 421.200 85.000 ;
        RECT 422.000 84.200 422.800 85.000 ;
        RECT 426.800 86.200 427.600 87.000 ;
        RECT 430.000 86.200 430.800 87.000 ;
        RECT 431.600 84.200 432.400 85.000 ;
        RECT 433.200 84.200 434.000 85.000 ;
        RECT 446.000 89.600 446.800 90.400 ;
        RECT 484.400 95.600 485.200 96.400 ;
        RECT 486.000 94.200 486.800 95.000 ;
        RECT 506.800 97.600 507.600 98.400 ;
        RECT 476.400 91.600 477.200 92.400 ;
        RECT 495.600 91.600 496.400 92.400 ;
        RECT 457.200 83.600 458.000 84.400 ;
        RECT 465.200 87.600 466.000 88.400 ;
        RECT 479.600 86.800 480.400 87.600 ;
        RECT 482.800 86.200 483.600 87.000 ;
        RECT 478.000 84.200 478.800 85.000 ;
        RECT 479.600 84.200 480.400 85.000 ;
        RECT 481.200 84.200 482.000 85.000 ;
        RECT 486.000 86.200 486.800 87.000 ;
        RECT 489.200 86.200 490.000 87.000 ;
        RECT 490.800 84.200 491.600 85.000 ;
        RECT 492.400 84.200 493.200 85.000 ;
        RECT 506.800 89.600 507.600 90.400 ;
        RECT 527.600 97.600 528.400 98.400 ;
        RECT 526.000 89.600 526.800 90.400 ;
        RECT 583.600 97.600 584.400 98.400 ;
        RECT 567.600 91.600 568.400 92.400 ;
        RECT 556.400 83.600 557.200 84.400 ;
        RECT 570.800 83.600 571.600 84.400 ;
        RECT 612.400 97.600 613.200 98.400 ;
        RECT 599.600 93.600 600.400 94.400 ;
        RECT 588.400 92.200 589.200 93.000 ;
        RECT 596.400 91.800 597.200 92.600 ;
        RECT 650.800 97.600 651.600 98.400 ;
        RECT 601.200 90.200 602.000 91.000 ;
        RECT 609.200 91.600 610.000 92.400 ;
        RECT 641.200 91.600 642.000 92.400 ;
        RECT 642.800 89.600 643.600 90.400 ;
        RECT 687.600 97.600 688.400 98.400 ;
        RECT 655.600 92.200 656.400 93.000 ;
        RECT 663.600 91.800 664.400 92.600 ;
        RECT 668.400 90.200 669.200 91.000 ;
        RECT 670.000 90.200 670.800 91.000 ;
        RECT 18.800 73.600 19.600 74.400 ;
        RECT 1.200 66.200 2.000 67.000 ;
        RECT 30.000 69.600 30.800 70.400 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 34.800 69.600 35.600 70.400 ;
        RECT 46.000 71.600 46.800 72.400 ;
        RECT 6.000 65.600 6.800 66.400 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 26.800 65.600 27.600 66.400 ;
        RECT 47.600 67.600 48.400 68.400 ;
        RECT 55.600 69.600 56.400 70.400 ;
        RECT 86.000 77.600 86.800 78.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 66.800 69.600 67.600 70.400 ;
        RECT 70.000 67.600 70.800 68.400 ;
        RECT 68.400 66.200 69.200 67.000 ;
        RECT 87.600 65.600 88.400 66.400 ;
        RECT 90.800 67.600 91.600 68.400 ;
        RECT 102.000 69.600 102.800 70.400 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 95.600 66.200 96.400 67.000 ;
        RECT 89.200 63.600 90.000 64.400 ;
        RECT 94.000 63.600 94.800 64.400 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 127.600 69.600 128.400 70.400 ;
        RECT 124.400 67.600 125.200 68.400 ;
        RECT 145.200 73.600 146.000 74.400 ;
        RECT 137.200 69.600 138.000 70.400 ;
        RECT 142.000 71.600 142.800 72.400 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 156.400 69.600 157.200 70.400 ;
        RECT 162.800 69.600 163.600 70.400 ;
        RECT 113.200 63.600 114.000 64.400 ;
        RECT 132.400 65.600 133.200 66.400 ;
        RECT 153.200 65.600 154.000 66.400 ;
        RECT 186.800 77.600 187.600 78.400 ;
        RECT 159.600 63.600 160.400 64.400 ;
        RECT 180.400 67.600 181.200 68.400 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 194.800 71.800 195.600 72.600 ;
        RECT 177.200 63.600 178.000 64.400 ;
        RECT 191.600 65.600 192.400 66.400 ;
        RECT 194.800 66.200 195.600 67.000 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 199.600 66.400 200.400 67.200 ;
        RECT 223.600 69.600 224.400 70.400 ;
        RECT 215.600 63.600 216.400 64.400 ;
        RECT 220.400 63.600 221.200 64.400 ;
        RECT 230.000 69.600 230.800 70.400 ;
        RECT 226.800 65.600 227.600 66.400 ;
        RECT 254.000 75.000 254.800 75.800 ;
        RECT 250.800 73.600 251.600 74.400 ;
        RECT 268.400 77.600 269.200 78.400 ;
        RECT 255.600 72.400 256.400 73.200 ;
        RECT 278.000 77.600 278.800 78.400 ;
        RECT 260.400 69.600 261.200 70.400 ;
        RECT 234.800 67.600 235.600 68.400 ;
        RECT 244.400 68.200 245.200 69.000 ;
        RECT 254.000 68.600 254.800 69.400 ;
        RECT 249.200 67.600 250.000 68.400 ;
        RECT 244.400 64.200 245.200 65.000 ;
        RECT 246.000 64.200 246.800 65.000 ;
        RECT 247.600 64.200 248.400 65.000 ;
        RECT 250.800 64.200 251.600 65.000 ;
        RECT 254.000 64.200 254.800 65.000 ;
        RECT 255.600 64.200 256.400 65.000 ;
        RECT 257.200 64.200 258.000 65.000 ;
        RECT 258.800 64.200 259.600 65.000 ;
        RECT 300.400 73.600 301.200 74.400 ;
        RECT 297.200 69.600 298.000 70.400 ;
        RECT 298.800 69.600 299.600 70.400 ;
        RECT 319.600 75.000 320.400 75.800 ;
        RECT 316.400 73.600 317.200 74.400 ;
        RECT 321.200 72.400 322.000 73.200 ;
        RECT 334.000 73.600 334.800 74.400 ;
        RECT 294.000 67.600 294.800 68.400 ;
        RECT 310.000 68.200 310.800 69.000 ;
        RECT 319.600 68.600 320.400 69.400 ;
        RECT 292.400 65.600 293.200 66.400 ;
        RECT 314.800 67.600 315.600 68.400 ;
        RECT 310.000 64.200 310.800 65.000 ;
        RECT 311.600 64.200 312.400 65.000 ;
        RECT 313.200 64.200 314.000 65.000 ;
        RECT 316.400 64.200 317.200 65.000 ;
        RECT 319.600 64.200 320.400 65.000 ;
        RECT 321.200 64.200 322.000 65.000 ;
        RECT 322.800 64.200 323.600 65.000 ;
        RECT 324.400 64.200 325.200 65.000 ;
        RECT 354.800 75.000 355.600 75.800 ;
        RECT 351.600 73.600 352.400 74.400 ;
        RECT 356.400 72.400 357.200 73.200 ;
        RECT 345.200 68.200 346.000 69.000 ;
        RECT 354.800 68.600 355.600 69.400 ;
        RECT 350.000 67.600 350.800 68.400 ;
        RECT 345.200 64.200 346.000 65.000 ;
        RECT 346.800 64.200 347.600 65.000 ;
        RECT 348.400 64.200 349.200 65.000 ;
        RECT 351.600 64.200 352.400 65.000 ;
        RECT 354.800 64.200 355.600 65.000 ;
        RECT 356.400 64.200 357.200 65.000 ;
        RECT 358.000 64.200 358.800 65.000 ;
        RECT 359.600 64.200 360.400 65.000 ;
        RECT 383.600 77.600 384.400 78.400 ;
        RECT 369.200 63.600 370.000 64.400 ;
        RECT 386.800 65.600 387.600 66.400 ;
        RECT 401.200 67.600 402.000 68.400 ;
        RECT 394.800 63.600 395.600 64.400 ;
        RECT 423.600 74.400 424.400 75.200 ;
        RECT 426.800 75.000 427.600 75.800 ;
        RECT 422.000 72.400 422.800 73.200 ;
        RECT 431.600 67.600 432.400 68.400 ;
        RECT 428.400 65.600 429.200 66.400 ;
        RECT 422.000 64.200 422.800 65.000 ;
        RECT 423.600 64.200 424.400 65.000 ;
        RECT 425.200 64.200 426.000 65.000 ;
        RECT 426.800 64.200 427.600 65.000 ;
        RECT 430.000 64.200 430.800 65.000 ;
        RECT 433.200 64.200 434.000 65.000 ;
        RECT 434.800 64.200 435.600 65.000 ;
        RECT 436.400 64.200 437.200 65.000 ;
        RECT 462.000 77.600 462.800 78.400 ;
        RECT 454.000 69.600 454.800 70.400 ;
        RECT 449.200 67.600 450.000 68.400 ;
        RECT 482.800 75.000 483.600 75.800 ;
        RECT 479.600 73.600 480.400 74.400 ;
        RECT 484.400 72.400 485.200 73.200 ;
        RECT 473.200 68.200 474.000 69.000 ;
        RECT 482.800 68.600 483.600 69.400 ;
        RECT 450.800 63.600 451.600 64.400 ;
        RECT 478.000 67.600 478.800 68.400 ;
        RECT 473.200 64.200 474.000 65.000 ;
        RECT 474.800 64.200 475.600 65.000 ;
        RECT 476.400 64.200 477.200 65.000 ;
        RECT 479.600 64.200 480.400 65.000 ;
        RECT 482.800 64.200 483.600 65.000 ;
        RECT 484.400 64.200 485.200 65.000 ;
        RECT 486.000 64.200 486.800 65.000 ;
        RECT 487.600 64.200 488.400 65.000 ;
        RECT 497.200 65.600 498.000 66.400 ;
        RECT 508.400 69.600 509.200 70.400 ;
        RECT 516.400 69.600 517.200 70.400 ;
        RECT 502.000 65.600 502.800 66.400 ;
        RECT 503.600 65.600 504.400 66.400 ;
        RECT 518.000 67.600 518.800 68.400 ;
        RECT 553.200 77.600 554.000 78.400 ;
        RECT 554.800 73.600 555.600 74.400 ;
        RECT 521.200 63.600 522.000 64.400 ;
        RECT 534.000 66.200 534.800 67.000 ;
        RECT 558.000 71.600 558.800 72.400 ;
        RECT 580.400 75.600 581.200 76.400 ;
        RECT 590.000 77.600 590.800 78.400 ;
        RECT 556.400 69.600 557.200 70.400 ;
        RECT 561.200 69.600 562.000 70.400 ;
        RECT 569.200 71.600 570.000 72.400 ;
        RECT 585.200 73.600 586.000 74.400 ;
        RECT 580.400 69.600 581.200 70.400 ;
        RECT 588.400 71.600 589.200 72.400 ;
        RECT 586.800 69.600 587.600 70.400 ;
        RECT 551.600 63.600 552.400 64.400 ;
        RECT 570.800 67.600 571.600 68.400 ;
        RECT 582.000 67.600 582.800 68.400 ;
        RECT 604.400 72.400 605.200 73.200 ;
        RECT 612.400 77.600 613.200 78.400 ;
        RECT 610.800 73.600 611.600 74.400 ;
        RECT 623.600 73.600 624.400 74.400 ;
        RECT 607.600 71.000 608.400 71.800 ;
        RECT 614.000 71.600 614.800 72.400 ;
        RECT 612.400 69.600 613.200 70.400 ;
        RECT 626.800 71.600 627.600 72.400 ;
        RECT 625.200 69.600 626.000 70.400 ;
        RECT 628.400 69.600 629.200 70.400 ;
        RECT 630.000 69.600 630.800 70.400 ;
        RECT 607.600 66.200 608.400 67.000 ;
        RECT 644.400 73.600 645.200 74.400 ;
        RECT 639.600 69.600 640.400 70.400 ;
        RECT 634.800 67.600 635.600 68.400 ;
        RECT 658.800 72.400 659.600 73.200 ;
        RECT 666.800 77.600 667.600 78.400 ;
        RECT 670.000 77.600 670.800 78.400 ;
        RECT 662.000 71.000 662.800 71.800 ;
        RECT 666.800 69.600 667.600 70.400 ;
        RECT 662.000 66.200 662.800 67.000 ;
        RECT 668.400 67.600 669.200 68.400 ;
        RECT 684.400 75.600 685.200 76.400 ;
        RECT 671.600 65.600 672.400 66.400 ;
        RECT 18.800 57.600 19.600 58.400 ;
        RECT 34.800 57.600 35.600 58.400 ;
        RECT 1.200 50.200 2.000 51.000 ;
        RECT 25.200 49.600 26.000 50.400 ;
        RECT 44.400 51.600 45.200 52.400 ;
        RECT 82.800 57.600 83.600 58.400 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 70.000 51.800 70.800 52.600 ;
        RECT 57.200 49.600 58.000 50.400 ;
        RECT 65.200 50.200 66.000 51.000 ;
        RECT 87.600 49.600 88.400 50.400 ;
        RECT 89.200 49.600 90.000 50.400 ;
        RECT 122.800 57.600 123.600 58.400 ;
        RECT 90.800 43.600 91.600 44.400 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 105.200 51.600 106.000 52.400 ;
        RECT 148.400 57.600 149.200 58.400 ;
        RECT 98.800 43.600 99.600 44.400 ;
        RECT 127.600 51.600 128.400 52.400 ;
        RECT 122.800 49.600 123.600 50.400 ;
        RECT 129.200 49.600 130.000 50.400 ;
        RECT 135.600 49.600 136.400 50.400 ;
        RECT 143.600 51.600 144.400 52.400 ;
        RECT 167.600 57.600 168.400 58.400 ;
        RECT 151.600 51.600 152.400 52.400 ;
        RECT 167.600 49.600 168.400 50.400 ;
        RECT 193.200 55.600 194.000 56.400 ;
        RECT 194.800 54.200 195.600 55.000 ;
        RECT 212.400 57.600 213.200 58.400 ;
        RECT 206.000 51.600 206.800 52.400 ;
        RECT 170.800 45.600 171.600 46.400 ;
        RECT 188.400 46.800 189.200 47.600 ;
        RECT 191.600 46.200 192.400 47.000 ;
        RECT 186.800 44.200 187.600 45.000 ;
        RECT 188.400 44.200 189.200 45.000 ;
        RECT 190.000 44.200 190.800 45.000 ;
        RECT 194.800 46.200 195.600 47.000 ;
        RECT 198.000 46.200 198.800 47.000 ;
        RECT 225.200 53.000 226.000 53.800 ;
        RECT 199.600 44.200 200.400 45.000 ;
        RECT 201.200 44.200 202.000 45.000 ;
        RECT 212.400 45.600 213.200 46.400 ;
        RECT 234.800 52.600 235.600 53.400 ;
        RECT 252.400 57.600 253.200 58.400 ;
        RECT 218.800 51.600 219.600 52.400 ;
        RECT 220.400 51.600 221.200 52.400 ;
        RECT 226.800 48.800 227.600 49.600 ;
        RECT 231.600 47.600 232.400 48.400 ;
        RECT 228.400 46.200 229.200 47.000 ;
        RECT 225.200 44.200 226.000 45.000 ;
        RECT 226.800 44.200 227.600 45.000 ;
        RECT 231.600 46.200 232.400 47.000 ;
        RECT 234.800 46.200 235.600 47.000 ;
        RECT 236.400 44.200 237.200 45.000 ;
        RECT 238.000 44.200 238.800 45.000 ;
        RECT 239.600 44.200 240.400 45.000 ;
        RECT 271.600 53.000 272.400 53.800 ;
        RECT 281.200 52.600 282.000 53.400 ;
        RECT 266.800 51.600 267.600 52.400 ;
        RECT 287.600 51.600 288.400 52.400 ;
        RECT 273.200 48.800 274.000 49.600 ;
        RECT 278.000 47.600 278.800 48.400 ;
        RECT 274.800 46.200 275.600 47.000 ;
        RECT 271.600 44.200 272.400 45.000 ;
        RECT 273.200 44.200 274.000 45.000 ;
        RECT 278.000 46.200 278.800 47.000 ;
        RECT 281.200 46.200 282.000 47.000 ;
        RECT 282.800 44.200 283.600 45.000 ;
        RECT 284.400 44.200 285.200 45.000 ;
        RECT 286.000 44.200 286.800 45.000 ;
        RECT 295.600 49.600 296.400 50.400 ;
        RECT 298.800 49.600 299.600 50.400 ;
        RECT 332.400 55.600 333.200 56.400 ;
        RECT 334.000 54.200 334.800 55.000 ;
        RECT 343.600 51.600 344.400 52.400 ;
        RECT 311.600 43.600 312.400 44.400 ;
        RECT 327.600 46.800 328.400 47.600 ;
        RECT 330.800 46.200 331.600 47.000 ;
        RECT 326.000 44.200 326.800 45.000 ;
        RECT 327.600 44.200 328.400 45.000 ;
        RECT 329.200 44.200 330.000 45.000 ;
        RECT 334.000 46.200 334.800 47.000 ;
        RECT 337.200 46.200 338.000 47.000 ;
        RECT 359.600 57.600 360.400 58.400 ;
        RECT 338.800 44.200 339.600 45.000 ;
        RECT 340.400 44.200 341.200 45.000 ;
        RECT 375.600 55.600 376.400 56.400 ;
        RECT 377.200 54.200 378.000 55.000 ;
        RECT 399.600 57.600 400.400 58.400 ;
        RECT 367.600 51.600 368.400 52.400 ;
        RECT 378.800 51.600 379.600 52.400 ;
        RECT 359.600 43.600 360.400 44.400 ;
        RECT 370.800 46.800 371.600 47.600 ;
        RECT 374.000 46.200 374.800 47.000 ;
        RECT 369.200 44.200 370.000 45.000 ;
        RECT 370.800 44.200 371.600 45.000 ;
        RECT 372.400 44.200 373.200 45.000 ;
        RECT 377.200 46.200 378.000 47.000 ;
        RECT 380.400 46.200 381.200 47.000 ;
        RECT 382.000 44.200 382.800 45.000 ;
        RECT 383.600 44.200 384.400 45.000 ;
        RECT 415.600 55.600 416.400 56.400 ;
        RECT 417.200 54.200 418.000 55.000 ;
        RECT 428.400 51.600 429.200 52.400 ;
        RECT 394.800 43.600 395.600 44.400 ;
        RECT 410.800 46.800 411.600 47.600 ;
        RECT 414.000 46.200 414.800 47.000 ;
        RECT 409.200 44.200 410.000 45.000 ;
        RECT 410.800 44.200 411.600 45.000 ;
        RECT 412.400 44.200 413.200 45.000 ;
        RECT 417.200 46.200 418.000 47.000 ;
        RECT 420.400 46.200 421.200 47.000 ;
        RECT 452.400 57.600 453.200 58.400 ;
        RECT 422.000 44.200 422.800 45.000 ;
        RECT 423.600 44.200 424.400 45.000 ;
        RECT 447.600 43.600 448.400 44.400 ;
        RECT 466.800 53.000 467.600 53.800 ;
        RECT 476.400 52.600 477.200 53.400 ;
        RECT 490.800 57.600 491.600 58.400 ;
        RECT 462.000 51.600 462.800 52.400 ;
        RECT 468.400 48.800 469.200 49.600 ;
        RECT 473.200 47.600 474.000 48.400 ;
        RECT 470.000 46.200 470.800 47.000 ;
        RECT 466.800 44.200 467.600 45.000 ;
        RECT 468.400 44.200 469.200 45.000 ;
        RECT 473.200 46.200 474.000 47.000 ;
        RECT 476.400 46.200 477.200 47.000 ;
        RECT 478.000 44.200 478.800 45.000 ;
        RECT 479.600 44.200 480.400 45.000 ;
        RECT 481.200 44.200 482.000 45.000 ;
        RECT 519.600 55.600 520.400 56.400 ;
        RECT 535.600 57.600 536.400 58.400 ;
        RECT 522.800 51.600 523.600 52.400 ;
        RECT 514.800 43.600 515.600 44.400 ;
        RECT 561.200 57.600 562.000 58.400 ;
        RECT 580.400 57.600 581.200 58.400 ;
        RECT 534.000 49.600 534.800 50.400 ;
        RECT 554.800 51.600 555.600 52.400 ;
        RECT 556.400 49.600 557.200 50.400 ;
        RECT 580.400 54.800 581.200 55.600 ;
        RECT 561.200 49.600 562.000 50.400 ;
        RECT 583.600 53.600 584.400 54.400 ;
        RECT 566.000 43.600 566.800 44.400 ;
        RECT 585.200 49.600 586.000 50.400 ;
        RECT 599.600 57.600 600.400 58.400 ;
        RECT 591.600 51.600 592.400 52.400 ;
        RECT 604.400 52.200 605.200 53.000 ;
        RECT 612.400 51.800 613.200 52.600 ;
        RECT 617.200 50.200 618.000 51.000 ;
        RECT 625.200 51.600 626.000 52.400 ;
        RECT 633.200 51.600 634.000 52.400 ;
        RECT 682.800 57.600 683.600 58.400 ;
        RECT 630.000 43.600 630.800 44.400 ;
        RECT 641.200 51.600 642.000 52.400 ;
        RECT 658.800 51.600 659.600 52.400 ;
        RECT 647.600 47.600 648.400 48.400 ;
        RECT 639.600 43.600 640.400 44.400 ;
        RECT 673.200 53.600 674.000 54.400 ;
        RECT 662.000 43.600 662.800 44.400 ;
        RECT 681.200 49.600 682.000 50.400 ;
        RECT 18.800 35.000 19.600 35.800 ;
        RECT 15.600 33.600 16.400 34.400 ;
        RECT 33.200 37.600 34.000 38.400 ;
        RECT 20.400 32.400 21.200 33.200 ;
        RECT 9.200 28.200 10.000 29.000 ;
        RECT 18.800 28.600 19.600 29.400 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 9.200 24.200 10.000 25.000 ;
        RECT 10.800 24.200 11.600 25.000 ;
        RECT 12.400 24.200 13.200 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 18.800 24.200 19.600 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 22.000 24.200 22.800 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 66.800 37.600 67.600 38.400 ;
        RECT 60.400 29.600 61.200 30.400 ;
        RECT 90.800 37.600 91.600 38.400 ;
        RECT 103.600 35.600 104.400 36.400 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 110.000 31.600 110.800 32.400 ;
        RECT 135.600 37.600 136.400 38.400 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 110.000 29.600 110.800 30.400 ;
        RECT 145.200 37.600 146.000 38.400 ;
        RECT 63.600 23.600 64.400 24.400 ;
        RECT 98.800 27.600 99.600 28.400 ;
        RECT 105.200 27.600 106.000 28.400 ;
        RECT 111.600 27.600 112.400 28.400 ;
        RECT 118.000 26.200 118.800 27.000 ;
        RECT 90.800 23.600 91.600 24.400 ;
        RECT 94.000 23.600 94.800 24.400 ;
        RECT 172.400 37.600 173.200 38.400 ;
        RECT 146.800 27.600 147.600 28.400 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 154.800 26.200 155.600 27.000 ;
        RECT 188.200 31.800 189.000 32.600 ;
        RECT 174.000 25.600 174.800 26.400 ;
        RECT 210.800 34.400 211.600 35.200 ;
        RECT 214.000 35.000 214.800 35.800 ;
        RECT 209.200 32.400 210.000 33.200 ;
        RECT 180.400 25.600 181.200 26.400 ;
        RECT 182.000 25.600 182.800 26.400 ;
        RECT 178.800 23.600 179.600 24.400 ;
        RECT 188.200 26.200 189.000 27.000 ;
        RECT 196.400 27.600 197.200 28.400 ;
        RECT 207.600 29.600 208.400 30.400 ;
        RECT 218.800 27.600 219.600 28.400 ;
        RECT 215.600 25.600 216.400 26.400 ;
        RECT 209.200 24.200 210.000 25.000 ;
        RECT 210.800 24.200 211.600 25.000 ;
        RECT 212.400 24.200 213.200 25.000 ;
        RECT 214.000 24.200 214.800 25.000 ;
        RECT 217.200 24.200 218.000 25.000 ;
        RECT 220.400 24.200 221.200 25.000 ;
        RECT 222.000 24.200 222.800 25.000 ;
        RECT 223.600 24.200 224.400 25.000 ;
        RECT 250.800 35.000 251.600 35.800 ;
        RECT 247.600 33.600 248.400 34.400 ;
        RECT 252.400 32.400 253.200 33.200 ;
        RECT 257.200 29.600 258.000 30.400 ;
        RECT 241.200 28.200 242.000 29.000 ;
        RECT 250.800 28.600 251.600 29.400 ;
        RECT 246.000 27.600 246.800 28.400 ;
        RECT 241.200 24.200 242.000 25.000 ;
        RECT 242.800 24.200 243.600 25.000 ;
        RECT 244.400 24.200 245.200 25.000 ;
        RECT 247.600 24.200 248.400 25.000 ;
        RECT 250.800 24.200 251.600 25.000 ;
        RECT 252.400 24.200 253.200 25.000 ;
        RECT 254.000 24.200 254.800 25.000 ;
        RECT 255.600 24.200 256.400 25.000 ;
        RECT 276.400 29.600 277.200 30.400 ;
        RECT 284.400 27.600 285.200 28.400 ;
        RECT 265.200 23.600 266.000 24.400 ;
        RECT 290.800 37.600 291.600 38.400 ;
        RECT 305.200 29.600 306.000 30.400 ;
        RECT 290.800 23.600 291.600 24.400 ;
        RECT 308.400 25.600 309.200 26.400 ;
        RECT 326.000 34.400 326.800 35.200 ;
        RECT 329.200 35.000 330.000 35.800 ;
        RECT 324.400 32.400 325.200 33.200 ;
        RECT 322.800 29.600 323.600 30.400 ;
        RECT 314.800 23.600 315.600 24.400 ;
        RECT 334.000 27.600 334.800 28.400 ;
        RECT 330.800 25.600 331.600 26.400 ;
        RECT 324.400 24.200 325.200 25.000 ;
        RECT 326.000 24.200 326.800 25.000 ;
        RECT 327.600 24.200 328.400 25.000 ;
        RECT 329.200 24.200 330.000 25.000 ;
        RECT 332.400 24.200 333.200 25.000 ;
        RECT 335.600 24.200 336.400 25.000 ;
        RECT 337.200 24.200 338.000 25.000 ;
        RECT 338.800 24.200 339.600 25.000 ;
        RECT 362.800 25.600 363.600 26.400 ;
        RECT 359.600 23.600 360.400 24.400 ;
        RECT 390.000 35.000 390.800 35.800 ;
        RECT 386.800 33.600 387.600 34.400 ;
        RECT 391.600 32.400 392.400 33.200 ;
        RECT 369.200 27.600 370.000 28.400 ;
        RECT 380.400 28.200 381.200 29.000 ;
        RECT 390.000 28.600 390.800 29.400 ;
        RECT 385.200 27.600 386.000 28.400 ;
        RECT 380.400 24.200 381.200 25.000 ;
        RECT 382.000 24.200 382.800 25.000 ;
        RECT 383.600 24.200 384.400 25.000 ;
        RECT 386.800 24.200 387.600 25.000 ;
        RECT 390.000 24.200 390.800 25.000 ;
        RECT 391.600 24.200 392.400 25.000 ;
        RECT 393.200 24.200 394.000 25.000 ;
        RECT 394.800 24.200 395.600 25.000 ;
        RECT 414.000 33.600 414.800 34.400 ;
        RECT 404.400 23.600 405.200 24.400 ;
        RECT 414.000 29.600 414.800 30.400 ;
        RECT 415.600 27.600 416.400 28.400 ;
        RECT 426.800 27.600 427.600 28.400 ;
        RECT 449.200 35.000 450.000 35.800 ;
        RECT 446.000 33.600 446.800 34.400 ;
        RECT 463.600 37.600 464.400 38.400 ;
        RECT 450.800 32.400 451.600 33.200 ;
        RECT 455.600 29.600 456.400 30.400 ;
        RECT 439.600 28.200 440.400 29.000 ;
        RECT 449.200 28.600 450.000 29.400 ;
        RECT 430.000 25.600 430.800 26.400 ;
        RECT 444.400 27.600 445.200 28.400 ;
        RECT 439.600 24.200 440.400 25.000 ;
        RECT 441.200 24.200 442.000 25.000 ;
        RECT 442.800 24.200 443.600 25.000 ;
        RECT 446.000 24.200 446.800 25.000 ;
        RECT 449.200 24.200 450.000 25.000 ;
        RECT 450.800 24.200 451.600 25.000 ;
        RECT 452.400 24.200 453.200 25.000 ;
        RECT 454.000 24.200 454.800 25.000 ;
        RECT 482.800 31.600 483.600 32.400 ;
        RECT 476.400 29.600 477.200 30.400 ;
        RECT 482.800 29.600 483.600 30.400 ;
        RECT 489.200 29.600 490.000 30.400 ;
        RECT 470.000 27.600 470.800 28.400 ;
        RECT 478.000 27.600 478.800 28.400 ;
        RECT 484.400 27.600 485.200 28.400 ;
        RECT 487.600 27.600 488.400 28.400 ;
        RECT 497.200 37.600 498.000 38.400 ;
        RECT 508.400 34.400 509.200 35.200 ;
        RECT 511.600 35.000 512.400 35.800 ;
        RECT 506.800 32.400 507.600 33.200 ;
        RECT 505.200 29.600 506.000 30.400 ;
        RECT 516.400 27.600 517.200 28.400 ;
        RECT 513.200 25.600 514.000 26.400 ;
        RECT 534.000 29.600 534.800 30.400 ;
        RECT 546.800 29.600 547.600 30.400 ;
        RECT 551.600 29.600 552.400 30.400 ;
        RECT 506.800 24.200 507.600 25.000 ;
        RECT 508.400 24.200 509.200 25.000 ;
        RECT 510.000 24.200 510.800 25.000 ;
        RECT 511.600 24.200 512.400 25.000 ;
        RECT 514.800 24.200 515.600 25.000 ;
        RECT 518.000 24.200 518.800 25.000 ;
        RECT 519.600 24.200 520.400 25.000 ;
        RECT 521.200 24.200 522.000 25.000 ;
        RECT 535.600 27.600 536.400 28.400 ;
        RECT 540.400 27.600 541.200 28.400 ;
        RECT 559.600 27.600 560.400 28.400 ;
        RECT 567.600 29.600 568.400 30.400 ;
        RECT 569.200 29.600 570.000 30.400 ;
        RECT 554.800 23.600 555.600 24.400 ;
        RECT 590.000 32.400 590.800 33.200 ;
        RECT 593.200 31.000 594.000 31.800 ;
        RECT 594.800 37.600 595.600 38.400 ;
        RECT 593.200 26.200 594.000 27.000 ;
        RECT 598.000 33.600 598.800 34.400 ;
        RECT 612.400 32.400 613.200 33.200 ;
        RECT 626.800 33.600 627.600 34.400 ;
        RECT 615.600 31.000 616.400 31.800 ;
        RECT 618.800 29.600 619.600 30.400 ;
        RECT 615.600 26.200 616.400 27.000 ;
        RECT 628.400 27.600 629.200 28.400 ;
        RECT 636.400 29.600 637.200 30.400 ;
        RECT 638.000 29.600 638.800 30.400 ;
        RECT 641.200 29.600 642.000 30.400 ;
        RECT 650.800 29.600 651.600 30.400 ;
        RECT 671.600 37.600 672.400 38.400 ;
        RECT 658.800 29.600 659.600 30.400 ;
        RECT 681.200 37.600 682.000 38.400 ;
        RECT 676.400 31.800 677.200 32.600 ;
        RECT 671.600 29.600 672.400 30.400 ;
        RECT 660.400 27.600 661.200 28.400 ;
        RECT 673.200 27.600 674.000 28.400 ;
        RECT 676.400 26.200 677.200 27.000 ;
        RECT 655.600 23.600 656.400 24.400 ;
        RECT 684.400 27.600 685.200 28.400 ;
        RECT 681.200 26.400 682.000 27.200 ;
        RECT 2.800 13.600 3.600 14.400 ;
        RECT 12.400 13.000 13.200 13.800 ;
        RECT 22.000 12.600 22.800 13.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 28.400 11.600 29.200 12.400 ;
        RECT 46.000 17.600 46.800 18.400 ;
        RECT 14.000 8.800 14.800 9.600 ;
        RECT 18.800 7.600 19.600 8.400 ;
        RECT 15.600 6.200 16.400 7.000 ;
        RECT 12.400 4.200 13.200 5.000 ;
        RECT 14.000 4.200 14.800 5.000 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 22.000 6.200 22.800 7.000 ;
        RECT 23.600 4.200 24.400 5.000 ;
        RECT 25.200 4.200 26.000 5.000 ;
        RECT 26.800 4.200 27.600 5.000 ;
        RECT 49.200 17.600 50.000 18.400 ;
        RECT 65.200 15.600 66.000 16.400 ;
        RECT 66.800 14.200 67.600 15.000 ;
        RECT 57.200 11.600 58.000 12.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 60.400 6.800 61.200 7.600 ;
        RECT 63.600 6.200 64.400 7.000 ;
        RECT 58.800 4.200 59.600 5.000 ;
        RECT 60.400 4.200 61.200 5.000 ;
        RECT 62.000 4.200 62.800 5.000 ;
        RECT 66.800 6.200 67.600 7.000 ;
        RECT 70.000 6.200 70.800 7.000 ;
        RECT 84.200 13.600 85.000 14.400 ;
        RECT 100.400 15.600 101.200 16.400 ;
        RECT 102.000 14.200 102.800 15.000 ;
        RECT 140.400 17.600 141.200 18.400 ;
        RECT 124.400 13.600 125.200 14.400 ;
        RECT 92.400 11.600 93.200 12.400 ;
        RECT 111.600 11.600 112.400 12.400 ;
        RECT 71.600 4.200 72.400 5.000 ;
        RECT 73.200 4.200 74.000 5.000 ;
        RECT 95.600 6.800 96.400 7.600 ;
        RECT 98.800 6.200 99.600 7.000 ;
        RECT 94.000 4.200 94.800 5.000 ;
        RECT 95.600 4.200 96.400 5.000 ;
        RECT 97.200 4.200 98.000 5.000 ;
        RECT 102.000 6.200 102.800 7.000 ;
        RECT 105.200 6.200 106.000 7.000 ;
        RECT 127.600 11.800 128.400 12.600 ;
        RECT 122.800 10.200 123.600 11.000 ;
        RECT 106.800 4.200 107.600 5.000 ;
        RECT 108.400 4.200 109.200 5.000 ;
        RECT 150.000 14.800 150.800 15.600 ;
        RECT 142.000 11.600 142.800 12.400 ;
        RECT 167.600 15.600 168.400 16.400 ;
        RECT 164.400 11.600 165.200 12.400 ;
        RECT 183.600 15.600 184.400 16.400 ;
        RECT 185.200 14.200 186.000 15.000 ;
        RECT 196.400 11.600 197.200 12.400 ;
        RECT 178.800 6.800 179.600 7.600 ;
        RECT 182.000 6.200 182.800 7.000 ;
        RECT 177.200 4.200 178.000 5.000 ;
        RECT 178.800 4.200 179.600 5.000 ;
        RECT 180.400 4.200 181.200 5.000 ;
        RECT 185.200 6.200 186.000 7.000 ;
        RECT 188.400 6.200 189.200 7.000 ;
        RECT 209.200 13.000 210.000 13.800 ;
        RECT 218.800 12.600 219.600 13.400 ;
        RECT 202.800 11.600 203.600 12.400 ;
        RECT 225.200 11.600 226.000 12.400 ;
        RECT 210.800 8.800 211.600 9.600 ;
        RECT 215.600 7.600 216.400 8.400 ;
        RECT 190.000 4.200 190.800 5.000 ;
        RECT 191.600 4.200 192.400 5.000 ;
        RECT 212.400 6.200 213.200 7.000 ;
        RECT 209.200 4.200 210.000 5.000 ;
        RECT 210.800 4.200 211.600 5.000 ;
        RECT 215.600 6.200 216.400 7.000 ;
        RECT 218.800 6.200 219.600 7.000 ;
        RECT 220.400 4.200 221.200 5.000 ;
        RECT 222.000 4.200 222.800 5.000 ;
        RECT 223.600 4.200 224.400 5.000 ;
        RECT 238.000 11.600 238.800 12.400 ;
        RECT 254.000 9.600 254.800 10.400 ;
        RECT 300.400 15.600 301.200 16.400 ;
        RECT 302.000 14.200 302.800 15.000 ;
        RECT 292.400 11.600 293.200 12.400 ;
        RECT 313.200 11.600 314.000 12.400 ;
        RECT 281.200 9.600 282.000 10.400 ;
        RECT 295.600 6.800 296.400 7.600 ;
        RECT 298.800 6.200 299.600 7.000 ;
        RECT 294.000 4.200 294.800 5.000 ;
        RECT 295.600 4.200 296.400 5.000 ;
        RECT 297.200 4.200 298.000 5.000 ;
        RECT 302.000 6.200 302.800 7.000 ;
        RECT 305.200 6.200 306.000 7.000 ;
        RECT 324.400 17.600 325.200 18.400 ;
        RECT 337.200 17.600 338.000 18.400 ;
        RECT 306.800 4.200 307.600 5.000 ;
        RECT 308.400 4.200 309.200 5.000 ;
        RECT 353.200 15.600 354.000 16.400 ;
        RECT 354.800 14.200 355.600 15.000 ;
        RECT 366.000 11.600 366.800 12.400 ;
        RECT 348.400 6.800 349.200 7.600 ;
        RECT 351.600 6.200 352.400 7.000 ;
        RECT 346.800 4.200 347.600 5.000 ;
        RECT 348.400 4.200 349.200 5.000 ;
        RECT 350.000 4.200 350.800 5.000 ;
        RECT 354.800 6.200 355.600 7.000 ;
        RECT 358.000 6.200 358.800 7.000 ;
        RECT 388.400 13.000 389.200 13.800 ;
        RECT 359.600 4.200 360.400 5.000 ;
        RECT 361.200 4.200 362.000 5.000 ;
        RECT 398.000 12.600 398.800 13.400 ;
        RECT 383.600 11.600 384.400 12.400 ;
        RECT 404.400 11.600 405.200 12.400 ;
        RECT 412.600 13.600 413.400 14.400 ;
        RECT 433.200 13.000 434.000 13.800 ;
        RECT 390.000 8.800 390.800 9.600 ;
        RECT 394.800 7.600 395.600 8.400 ;
        RECT 391.600 6.200 392.400 7.000 ;
        RECT 388.400 4.200 389.200 5.000 ;
        RECT 390.000 4.200 390.800 5.000 ;
        RECT 394.800 6.200 395.600 7.000 ;
        RECT 398.000 6.200 398.800 7.000 ;
        RECT 399.600 4.200 400.400 5.000 ;
        RECT 401.200 4.200 402.000 5.000 ;
        RECT 402.800 4.200 403.600 5.000 ;
        RECT 442.800 12.600 443.600 13.400 ;
        RECT 428.400 11.600 429.200 12.400 ;
        RECT 449.200 11.600 450.000 12.400 ;
        RECT 465.200 17.600 466.000 18.400 ;
        RECT 434.800 8.800 435.600 9.600 ;
        RECT 439.600 7.600 440.400 8.400 ;
        RECT 436.400 6.200 437.200 7.000 ;
        RECT 433.200 4.200 434.000 5.000 ;
        RECT 434.800 4.200 435.600 5.000 ;
        RECT 439.600 6.200 440.400 7.000 ;
        RECT 442.800 6.200 443.600 7.000 ;
        RECT 444.400 4.200 445.200 5.000 ;
        RECT 446.000 4.200 446.800 5.000 ;
        RECT 447.600 4.200 448.400 5.000 ;
        RECT 468.400 17.600 469.200 18.400 ;
        RECT 484.400 15.600 485.200 16.400 ;
        RECT 486.000 14.200 486.800 15.000 ;
        RECT 476.400 11.600 477.200 12.400 ;
        RECT 498.800 11.600 499.600 12.400 ;
        RECT 479.600 6.800 480.400 7.600 ;
        RECT 482.800 6.200 483.600 7.000 ;
        RECT 478.000 4.200 478.800 5.000 ;
        RECT 479.600 4.200 480.400 5.000 ;
        RECT 481.200 4.200 482.000 5.000 ;
        RECT 486.000 6.200 486.800 7.000 ;
        RECT 489.200 6.200 490.000 7.000 ;
        RECT 503.600 17.600 504.400 18.400 ;
        RECT 490.800 4.200 491.600 5.000 ;
        RECT 492.400 4.200 493.200 5.000 ;
        RECT 513.200 13.000 514.000 13.800 ;
        RECT 522.800 12.600 523.600 13.400 ;
        RECT 540.400 17.600 541.200 18.400 ;
        RECT 508.400 11.600 509.200 12.400 ;
        RECT 529.200 11.600 530.000 12.400 ;
        RECT 514.800 8.800 515.600 9.600 ;
        RECT 519.600 7.600 520.400 8.400 ;
        RECT 516.400 6.200 517.200 7.000 ;
        RECT 513.200 4.200 514.000 5.000 ;
        RECT 514.800 4.200 515.600 5.000 ;
        RECT 519.600 6.200 520.400 7.000 ;
        RECT 522.800 6.200 523.600 7.000 ;
        RECT 524.400 4.200 525.200 5.000 ;
        RECT 526.000 4.200 526.800 5.000 ;
        RECT 527.600 4.200 528.400 5.000 ;
        RECT 551.600 13.000 552.400 13.800 ;
        RECT 561.200 12.600 562.000 13.400 ;
        RECT 575.600 17.600 576.400 18.400 ;
        RECT 546.800 11.600 547.600 12.400 ;
        RECT 588.400 17.600 589.200 18.400 ;
        RECT 553.200 8.800 554.000 9.600 ;
        RECT 558.000 7.600 558.800 8.400 ;
        RECT 554.800 6.200 555.600 7.000 ;
        RECT 551.600 4.200 552.400 5.000 ;
        RECT 553.200 4.200 554.000 5.000 ;
        RECT 558.000 6.200 558.800 7.000 ;
        RECT 561.200 6.200 562.000 7.000 ;
        RECT 562.800 4.200 563.600 5.000 ;
        RECT 564.400 4.200 565.200 5.000 ;
        RECT 566.000 4.200 566.800 5.000 ;
        RECT 633.200 17.600 634.000 18.400 ;
        RECT 604.400 13.600 605.200 14.400 ;
        RECT 593.200 12.200 594.000 13.000 ;
        RECT 601.200 11.800 602.000 12.600 ;
        RECT 606.000 10.200 606.800 11.000 ;
        RECT 625.200 9.600 626.000 10.400 ;
        RECT 630.000 9.600 630.800 10.400 ;
        RECT 636.400 17.600 637.200 18.400 ;
        RECT 642.800 17.600 643.600 18.400 ;
        RECT 662.000 17.600 662.800 18.400 ;
        RECT 658.800 13.600 659.600 14.400 ;
        RECT 647.600 12.200 648.400 13.000 ;
        RECT 681.200 17.600 682.000 18.400 ;
        RECT 666.800 12.200 667.600 13.000 ;
        RECT 660.400 10.200 661.200 11.000 ;
        RECT 679.600 10.200 680.400 11.000 ;
      LAYER metal2 ;
        RECT 9.200 484.200 10.000 497.800 ;
        RECT 10.800 484.200 11.600 497.800 ;
        RECT 12.400 486.200 13.200 497.800 ;
        RECT 14.000 493.600 14.800 494.400 ;
        RECT 14.000 491.600 14.800 492.400 ;
        RECT 14.100 482.400 14.700 491.600 ;
        RECT 15.600 486.200 16.400 497.800 ;
        RECT 17.200 495.600 18.000 496.400 ;
        RECT 17.300 484.300 17.900 495.600 ;
        RECT 18.800 486.200 19.600 497.800 ;
        RECT 17.300 483.700 19.500 484.300 ;
        RECT 20.400 484.200 21.200 497.800 ;
        RECT 22.000 484.200 22.800 497.800 ;
        RECT 23.600 484.200 24.400 497.800 ;
        RECT 34.800 493.600 35.600 494.400 ;
        RECT 25.200 491.600 26.000 492.400 ;
        RECT 41.200 491.600 42.000 492.400 ;
        RECT 49.200 491.600 50.000 492.400 ;
        RECT 41.300 490.400 41.900 491.600 ;
        RECT 36.400 489.600 37.200 490.400 ;
        RECT 39.600 489.600 40.400 490.400 ;
        RECT 41.200 489.600 42.000 490.400 ;
        RECT 10.800 481.600 11.600 482.400 ;
        RECT 14.000 481.600 14.800 482.400 ;
        RECT 10.900 470.400 11.500 481.600 ;
        RECT 10.800 469.600 11.600 470.400 ;
        RECT 2.800 463.600 3.600 464.400 ;
        RECT 2.900 448.400 3.500 463.600 ;
        RECT 2.800 447.600 3.600 448.400 ;
        RECT 1.200 443.600 2.000 444.400 ;
        RECT 1.200 433.600 2.000 434.400 ;
        RECT 1.300 432.400 1.900 433.600 ;
        RECT 1.200 431.600 2.000 432.400 ;
        RECT 1.200 410.200 2.000 415.800 ;
        RECT 2.900 404.300 3.500 447.600 ;
        RECT 6.000 446.200 6.800 457.800 ;
        RECT 6.000 424.200 6.800 435.800 ;
        RECT 4.400 406.200 5.200 417.800 ;
        RECT 7.600 411.600 8.400 412.400 ;
        RECT 2.900 403.700 5.100 404.300 ;
        RECT 1.200 370.200 2.000 375.800 ;
        RECT 1.200 346.200 2.000 351.800 ;
        RECT 1.200 330.200 2.000 335.800 ;
        RECT 2.900 292.400 3.500 403.700 ;
        RECT 4.500 390.400 5.100 403.700 ;
        RECT 4.400 389.600 5.200 390.400 ;
        RECT 6.000 386.200 6.800 391.800 ;
        RECT 9.200 384.200 10.000 395.800 ;
        RECT 4.400 366.200 5.200 377.800 ;
        RECT 7.600 371.600 8.400 372.400 ;
        RECT 4.400 344.200 5.200 355.800 ;
        RECT 7.600 349.600 8.400 350.400 ;
        RECT 7.700 348.400 8.300 349.600 ;
        RECT 7.600 347.600 8.400 348.400 ;
        RECT 4.400 326.200 5.200 337.800 ;
        RECT 7.600 331.600 8.400 332.400 ;
        RECT 10.900 330.400 11.500 469.600 ;
        RECT 12.400 464.200 13.200 477.800 ;
        RECT 14.000 464.200 14.800 477.800 ;
        RECT 15.600 464.200 16.400 477.800 ;
        RECT 17.200 464.200 18.000 475.800 ;
        RECT 18.900 466.400 19.500 483.700 ;
        RECT 33.200 483.600 34.000 484.400 ;
        RECT 18.800 465.600 19.600 466.400 ;
        RECT 18.900 460.400 19.500 465.600 ;
        RECT 20.400 464.200 21.200 475.800 ;
        RECT 22.000 467.600 22.800 468.400 ;
        RECT 23.600 464.200 24.400 475.800 ;
        RECT 25.200 464.200 26.000 477.800 ;
        RECT 26.800 464.200 27.600 477.800 ;
        RECT 33.300 472.400 33.900 483.600 ;
        RECT 39.700 478.400 40.300 489.600 ;
        RECT 54.000 484.200 54.800 497.800 ;
        RECT 55.600 484.200 56.400 497.800 ;
        RECT 57.200 486.200 58.000 497.800 ;
        RECT 58.800 493.600 59.600 494.400 ;
        RECT 60.400 486.200 61.200 497.800 ;
        RECT 62.000 495.600 62.800 496.400 ;
        RECT 39.600 477.600 40.400 478.400 ;
        RECT 39.600 475.600 40.400 476.400 ;
        RECT 33.200 471.600 34.000 472.400 ;
        RECT 36.400 471.600 37.200 472.400 ;
        RECT 39.700 470.400 40.300 475.600 ;
        RECT 42.800 471.600 43.600 472.400 ;
        RECT 39.600 469.600 40.400 470.400 ;
        RECT 38.000 467.600 38.800 468.400 ;
        RECT 18.800 460.300 19.600 460.400 ;
        RECT 17.300 459.700 19.600 460.300 ;
        RECT 14.000 451.800 14.800 452.600 ;
        RECT 14.100 450.400 14.700 451.800 ;
        RECT 14.000 449.600 14.800 450.400 ;
        RECT 15.600 446.200 16.400 457.800 ;
        RECT 17.300 454.400 17.900 459.700 ;
        RECT 18.800 459.600 19.600 459.700 ;
        RECT 38.100 458.400 38.700 467.600 ;
        RECT 38.000 457.600 38.800 458.400 ;
        RECT 17.200 453.600 18.000 454.400 ;
        RECT 14.000 429.400 14.800 430.400 ;
        RECT 15.600 424.200 16.400 435.800 ;
        RECT 17.300 428.400 17.900 453.600 ;
        RECT 18.800 450.200 19.600 455.800 ;
        RECT 20.400 453.600 21.200 454.400 ;
        RECT 31.600 453.600 32.400 454.400 ;
        RECT 34.800 453.600 35.600 454.400 ;
        RECT 20.500 446.400 21.100 453.600 ;
        RECT 22.000 452.300 22.800 452.400 ;
        RECT 22.000 451.700 24.300 452.300 ;
        RECT 22.000 451.600 22.800 451.700 ;
        RECT 22.000 449.600 22.800 450.400 ;
        RECT 20.400 445.600 21.200 446.400 ;
        RECT 17.200 427.600 18.000 428.400 ;
        RECT 18.800 426.200 19.600 431.800 ;
        RECT 20.500 428.400 21.100 445.600 ;
        RECT 23.700 442.400 24.300 451.700 ;
        RECT 30.000 451.600 30.800 452.400 ;
        RECT 26.800 449.600 27.600 450.400 ;
        RECT 26.900 444.400 27.500 449.600 ;
        RECT 26.800 443.600 27.600 444.400 ;
        RECT 23.600 441.600 24.400 442.400 ;
        RECT 26.800 431.600 27.600 432.400 ;
        RECT 30.100 430.400 30.700 451.600 ;
        RECT 31.700 450.400 32.300 453.600 ;
        RECT 34.900 452.400 35.500 453.600 ;
        RECT 34.800 451.600 35.600 452.400 ;
        RECT 39.700 450.400 40.300 469.600 ;
        RECT 41.200 467.600 42.000 468.400 ;
        RECT 46.000 467.600 46.800 468.400 ;
        RECT 41.300 450.400 41.900 467.600 ;
        RECT 42.800 463.600 43.600 464.400 ;
        RECT 42.900 456.400 43.500 463.600 ;
        RECT 42.800 455.600 43.600 456.400 ;
        RECT 46.100 454.400 46.700 467.600 ;
        RECT 47.600 466.200 48.400 471.800 ;
        RECT 50.800 464.200 51.600 475.800 ;
        RECT 52.400 469.400 53.200 470.200 ;
        RECT 52.500 454.400 53.100 469.400 ;
        RECT 55.600 467.600 56.400 468.400 ;
        RECT 55.700 460.400 56.300 467.600 ;
        RECT 58.800 463.600 59.600 464.400 ;
        RECT 60.400 464.200 61.200 475.800 ;
        RECT 62.100 474.400 62.700 495.600 ;
        RECT 63.600 486.200 64.400 497.800 ;
        RECT 65.200 484.200 66.000 497.800 ;
        RECT 66.800 484.200 67.600 497.800 ;
        RECT 68.400 484.200 69.200 497.800 ;
        RECT 86.000 495.600 86.800 496.400 ;
        RECT 86.100 492.400 86.700 495.600 ;
        RECT 87.600 493.600 88.400 494.400 ;
        RECT 95.600 493.600 96.400 494.400 ;
        RECT 110.000 493.600 110.800 494.400 ;
        RECT 70.000 491.600 70.800 492.400 ;
        RECT 86.000 491.600 86.800 492.400 ;
        RECT 94.000 491.600 94.800 492.400 ;
        RECT 70.100 486.400 70.700 491.600 ;
        RECT 86.100 490.400 86.700 491.600 ;
        RECT 94.100 490.400 94.700 491.600 ;
        RECT 86.000 489.600 86.800 490.400 ;
        RECT 90.800 490.300 91.600 490.400 ;
        RECT 89.300 489.700 91.600 490.300 ;
        RECT 87.600 487.600 88.400 488.400 ;
        RECT 70.000 485.600 70.800 486.400 ;
        RECT 78.000 483.600 78.800 484.400 ;
        RECT 62.000 473.600 62.800 474.400 ;
        RECT 71.600 473.600 72.400 474.400 ;
        RECT 78.000 473.600 78.800 474.400 ;
        RECT 84.400 473.600 85.200 474.400 ;
        RECT 68.400 471.600 69.200 472.400 ;
        RECT 68.500 470.400 69.100 471.600 ;
        RECT 78.100 470.400 78.700 473.600 ;
        RECT 82.800 471.600 83.600 472.400 ;
        RECT 82.900 470.400 83.500 471.600 ;
        RECT 68.400 469.600 69.200 470.400 ;
        RECT 73.200 469.600 74.000 470.400 ;
        RECT 74.800 469.600 75.600 470.400 ;
        RECT 78.000 469.600 78.800 470.400 ;
        RECT 82.800 469.600 83.600 470.400 ;
        RECT 68.500 464.400 69.100 469.600 ;
        RECT 71.600 465.600 72.400 466.400 ;
        RECT 65.200 464.300 66.000 464.400 ;
        RECT 63.700 463.700 66.000 464.300 ;
        RECT 55.600 459.600 56.400 460.400 ;
        RECT 42.800 453.600 43.600 454.400 ;
        RECT 46.000 454.300 46.800 454.400 ;
        RECT 46.000 453.700 48.300 454.300 ;
        RECT 46.000 453.600 46.800 453.700 ;
        RECT 42.900 450.400 43.500 453.600 ;
        RECT 44.400 451.600 45.200 452.400 ;
        RECT 31.600 449.600 32.400 450.400 ;
        RECT 39.600 449.600 40.400 450.400 ;
        RECT 41.200 449.600 42.000 450.400 ;
        RECT 42.800 449.600 43.600 450.400 ;
        RECT 22.000 429.600 22.800 430.400 ;
        RECT 23.600 429.600 24.400 430.400 ;
        RECT 30.000 429.600 30.800 430.400 ;
        RECT 20.400 427.600 21.200 428.400 ;
        RECT 12.400 411.600 13.200 412.400 ;
        RECT 12.500 388.400 13.100 411.600 ;
        RECT 14.000 406.200 14.800 417.800 ;
        RECT 20.500 414.400 21.100 427.600 ;
        RECT 22.100 416.400 22.700 429.600 ;
        RECT 31.700 428.400 32.300 449.600 ;
        RECT 39.700 448.400 40.300 449.600 ;
        RECT 39.600 447.600 40.400 448.400 ;
        RECT 39.600 443.600 40.400 444.400 ;
        RECT 36.400 441.600 37.200 442.400 ;
        RECT 36.500 438.400 37.100 441.600 ;
        RECT 36.400 437.600 37.200 438.400 ;
        RECT 39.700 430.400 40.300 443.600 ;
        RECT 41.200 437.600 42.000 438.400 ;
        RECT 41.300 430.400 41.900 437.600 ;
        RECT 42.800 435.600 43.600 436.400 ;
        RECT 42.900 432.400 43.500 435.600 ;
        RECT 44.500 434.400 45.100 451.600 ;
        RECT 44.400 433.600 45.200 434.400 ;
        RECT 42.800 431.600 43.600 432.400 ;
        RECT 34.800 429.600 35.600 430.400 ;
        RECT 39.600 429.600 40.400 430.400 ;
        RECT 41.200 429.600 42.000 430.400 ;
        RECT 42.800 429.600 43.600 430.400 ;
        RECT 31.600 427.600 32.400 428.400 ;
        RECT 31.700 416.400 32.300 427.600 ;
        RECT 34.800 417.600 35.600 418.400 ;
        RECT 22.000 415.600 22.800 416.400 ;
        RECT 31.600 415.600 32.400 416.400 ;
        RECT 20.400 413.600 21.200 414.400 ;
        RECT 22.000 413.600 22.800 414.400 ;
        RECT 26.800 413.600 27.600 414.400 ;
        RECT 18.800 409.600 19.600 410.400 ;
        RECT 18.900 408.400 19.500 409.600 ;
        RECT 18.800 407.600 19.600 408.400 ;
        RECT 20.500 402.400 21.100 413.600 ;
        RECT 22.100 412.400 22.700 413.600 ;
        RECT 34.900 412.400 35.500 417.600 ;
        RECT 22.000 411.600 22.800 412.400 ;
        RECT 23.600 411.600 24.400 412.400 ;
        RECT 26.800 411.600 27.600 412.400 ;
        RECT 33.200 411.600 34.000 412.400 ;
        RECT 34.800 411.600 35.600 412.400 ;
        RECT 36.400 411.600 37.200 412.400 ;
        RECT 26.900 410.400 27.500 411.600 ;
        RECT 25.200 409.600 26.000 410.400 ;
        RECT 26.800 409.600 27.600 410.400 ;
        RECT 25.300 408.400 25.900 409.600 ;
        RECT 25.200 407.600 26.000 408.400 ;
        RECT 20.400 401.600 21.200 402.400 ;
        RECT 23.600 397.600 24.400 398.400 ;
        RECT 14.000 393.600 14.800 394.400 ;
        RECT 14.100 390.400 14.700 393.600 ;
        RECT 14.000 389.600 14.800 390.400 ;
        RECT 12.400 387.600 13.200 388.400 ;
        RECT 12.500 372.400 13.100 387.600 ;
        RECT 18.800 384.200 19.600 395.800 ;
        RECT 20.400 391.600 21.200 392.400 ;
        RECT 25.200 392.300 26.000 392.400 ;
        RECT 26.900 392.300 27.500 409.600 ;
        RECT 28.400 407.600 29.200 408.400 ;
        RECT 28.500 398.400 29.100 407.600 ;
        RECT 33.300 402.300 33.900 411.600 ;
        RECT 33.300 401.700 35.500 402.300 ;
        RECT 28.400 397.600 29.200 398.400 ;
        RECT 25.200 391.700 27.500 392.300 ;
        RECT 25.200 391.600 26.000 391.700 ;
        RECT 12.400 371.600 13.200 372.400 ;
        RECT 12.500 350.400 13.100 371.600 ;
        RECT 14.000 366.200 14.800 377.800 ;
        RECT 18.800 377.600 19.600 378.400 ;
        RECT 18.900 374.400 19.500 377.600 ;
        RECT 20.500 376.400 21.100 391.600 ;
        RECT 25.200 389.600 26.000 390.400 ;
        RECT 33.200 389.600 34.000 390.400 ;
        RECT 23.600 381.600 24.400 382.400 ;
        RECT 22.000 379.600 22.800 380.400 ;
        RECT 22.100 378.400 22.700 379.600 ;
        RECT 22.000 377.600 22.800 378.400 ;
        RECT 20.400 375.600 21.200 376.400 ;
        RECT 23.700 374.400 24.300 381.600 ;
        RECT 18.800 373.600 19.600 374.400 ;
        RECT 23.600 373.600 24.400 374.400 ;
        RECT 18.800 359.600 19.600 360.400 ;
        RECT 18.900 358.400 19.500 359.600 ;
        RECT 18.800 357.600 19.600 358.400 ;
        RECT 12.400 349.600 13.200 350.400 ;
        RECT 12.500 332.400 13.100 349.600 ;
        RECT 14.000 344.200 14.800 355.800 ;
        RECT 23.700 354.300 24.300 373.600 ;
        RECT 25.300 372.400 25.900 389.600 ;
        RECT 33.300 388.400 33.900 389.600 ;
        RECT 30.000 387.600 30.800 388.400 ;
        RECT 33.200 387.600 34.000 388.400 ;
        RECT 30.100 382.400 30.700 387.600 ;
        RECT 30.000 381.600 30.800 382.400 ;
        RECT 33.200 375.600 34.000 376.400 ;
        RECT 28.400 373.600 29.200 374.400 ;
        RECT 30.000 373.600 30.800 374.400 ;
        RECT 25.200 371.600 26.000 372.400 ;
        RECT 25.300 356.400 25.900 371.600 ;
        RECT 28.500 370.400 29.100 373.600 ;
        RECT 30.100 372.400 30.700 373.600 ;
        RECT 33.300 372.400 33.900 375.600 ;
        RECT 34.900 372.400 35.500 401.700 ;
        RECT 36.500 396.400 37.100 411.600 ;
        RECT 39.700 408.400 40.300 429.600 ;
        RECT 42.800 415.600 43.600 416.400 ;
        RECT 42.900 414.400 43.500 415.600 ;
        RECT 42.800 413.600 43.600 414.400 ;
        RECT 44.500 412.400 45.100 433.600 ;
        RECT 46.000 429.600 46.800 430.400 ;
        RECT 46.100 424.400 46.700 429.600 ;
        RECT 47.700 428.400 48.300 453.700 ;
        RECT 52.400 453.600 53.200 454.400 ;
        RECT 55.600 453.600 56.400 454.400 ;
        RECT 49.200 449.600 50.000 450.400 ;
        RECT 55.700 446.400 56.300 453.600 ;
        RECT 58.900 452.400 59.500 463.600 ;
        RECT 63.700 452.400 64.300 463.700 ;
        RECT 65.200 463.600 66.000 463.700 ;
        RECT 68.400 463.600 69.200 464.400 ;
        RECT 71.700 454.400 72.300 465.600 ;
        RECT 71.600 453.600 72.400 454.400 ;
        RECT 58.800 451.600 59.600 452.400 ;
        RECT 63.600 451.600 64.400 452.400 ;
        RECT 65.200 451.600 66.000 452.400 ;
        RECT 66.800 451.600 67.600 452.400 ;
        RECT 70.000 452.300 70.800 452.400 ;
        RECT 68.500 451.700 70.800 452.300 ;
        RECT 55.600 445.600 56.400 446.400 ;
        RECT 55.600 435.600 56.400 436.400 ;
        RECT 55.700 430.400 56.300 435.600 ;
        RECT 54.000 429.600 54.800 430.400 ;
        RECT 55.600 429.600 56.400 430.400 ;
        RECT 57.200 429.600 58.000 430.400 ;
        RECT 47.600 427.600 48.400 428.400 ;
        RECT 46.000 423.600 46.800 424.400 ;
        RECT 50.800 423.600 51.600 424.400 ;
        RECT 50.900 416.400 51.500 423.600 ;
        RECT 50.800 415.600 51.600 416.400 ;
        RECT 50.800 413.600 51.600 414.400 ;
        RECT 44.400 411.600 45.200 412.400 ;
        RECT 52.400 411.600 53.200 412.400 ;
        RECT 47.600 409.600 48.400 410.400 ;
        RECT 39.600 407.600 40.400 408.400 ;
        RECT 47.700 406.400 48.300 409.600 ;
        RECT 47.600 405.600 48.400 406.400 ;
        RECT 54.100 404.400 54.700 429.600 ;
        RECT 55.700 418.400 56.300 429.600 ;
        RECT 58.900 428.300 59.500 451.600 ;
        RECT 63.700 450.400 64.300 451.600 ;
        RECT 63.600 449.600 64.400 450.400 ;
        RECT 65.300 438.400 65.900 451.600 ;
        RECT 66.900 450.400 67.500 451.600 ;
        RECT 66.800 449.600 67.600 450.400 ;
        RECT 68.500 438.400 69.100 451.700 ;
        RECT 70.000 451.600 70.800 451.700 ;
        RECT 70.000 449.600 70.800 450.400 ;
        RECT 71.700 446.400 72.300 453.600 ;
        RECT 73.200 451.600 74.000 452.400 ;
        RECT 73.200 449.600 74.000 450.400 ;
        RECT 71.600 445.600 72.400 446.400 ;
        RECT 73.300 444.400 73.900 449.600 ;
        RECT 73.200 444.300 74.000 444.400 ;
        RECT 71.700 443.700 74.000 444.300 ;
        RECT 65.200 437.600 66.000 438.400 ;
        RECT 68.400 437.600 69.200 438.400 ;
        RECT 70.000 437.600 70.800 438.400 ;
        RECT 66.800 431.600 67.600 432.400 ;
        RECT 66.900 430.400 67.500 431.600 ;
        RECT 63.600 429.600 64.400 430.400 ;
        RECT 65.200 429.600 66.000 430.400 ;
        RECT 66.800 429.600 67.600 430.400 ;
        RECT 57.300 427.700 59.500 428.300 ;
        RECT 55.600 417.600 56.400 418.400 ;
        RECT 55.600 413.600 56.400 414.400 ;
        RECT 54.000 403.600 54.800 404.400 ;
        RECT 55.700 402.400 56.300 413.600 ;
        RECT 57.300 412.400 57.900 427.700 ;
        RECT 63.700 426.400 64.300 429.600 ;
        RECT 65.300 428.400 65.900 429.600 ;
        RECT 65.200 427.600 66.000 428.400 ;
        RECT 63.600 425.600 64.400 426.400 ;
        RECT 65.200 419.600 66.000 420.400 ;
        RECT 65.300 416.400 65.900 419.600 ;
        RECT 65.200 415.600 66.000 416.400 ;
        RECT 57.200 411.600 58.000 412.400 ;
        RECT 58.800 411.600 59.600 412.400 ;
        RECT 62.000 411.600 62.800 412.400 ;
        RECT 63.600 411.600 64.400 412.400 ;
        RECT 68.400 411.600 69.200 412.400 ;
        RECT 57.300 410.400 57.900 411.600 ;
        RECT 57.200 409.600 58.000 410.400 ;
        RECT 62.100 406.400 62.700 411.600 ;
        RECT 63.700 410.400 64.300 411.600 ;
        RECT 63.600 409.600 64.400 410.400 ;
        RECT 65.200 409.600 66.000 410.400 ;
        RECT 62.000 405.600 62.800 406.400 ;
        RECT 50.800 401.600 51.600 402.400 ;
        RECT 55.600 401.600 56.400 402.400 ;
        RECT 42.800 397.600 43.600 398.400 ;
        RECT 36.400 395.600 37.200 396.400 ;
        RECT 36.500 390.400 37.100 395.600 ;
        RECT 42.900 392.400 43.500 397.600 ;
        RECT 47.600 393.600 48.400 394.400 ;
        RECT 42.800 391.600 43.600 392.400 ;
        RECT 49.200 391.600 50.000 392.400 ;
        RECT 49.300 390.400 49.900 391.600 ;
        RECT 36.400 389.600 37.200 390.400 ;
        RECT 39.600 389.600 40.400 390.400 ;
        RECT 47.600 389.600 48.400 390.400 ;
        RECT 49.200 389.600 50.000 390.400 ;
        RECT 38.000 387.600 38.800 388.400 ;
        RECT 49.300 384.400 49.900 389.600 ;
        RECT 50.900 388.400 51.500 401.600 ;
        RECT 63.600 399.600 64.400 400.400 ;
        RECT 63.700 398.400 64.300 399.600 ;
        RECT 63.600 397.600 64.400 398.400 ;
        RECT 52.400 389.600 53.200 390.400 ;
        RECT 57.200 389.600 58.000 390.400 ;
        RECT 58.800 389.600 59.600 390.400 ;
        RECT 60.400 389.600 61.200 390.400 ;
        RECT 52.500 388.400 53.100 389.600 ;
        RECT 57.300 388.400 57.900 389.600 ;
        RECT 60.500 388.400 61.100 389.600 ;
        RECT 50.800 387.600 51.600 388.400 ;
        RECT 52.400 387.600 53.200 388.400 ;
        RECT 57.200 387.600 58.000 388.400 ;
        RECT 60.400 387.600 61.200 388.400 ;
        RECT 49.200 383.600 50.000 384.400 ;
        RECT 47.600 377.600 48.400 378.400 ;
        RECT 54.000 377.600 54.800 378.400 ;
        RECT 46.000 375.600 46.800 376.400 ;
        RECT 46.100 374.400 46.700 375.600 ;
        RECT 36.400 373.600 37.200 374.400 ;
        RECT 46.000 373.600 46.800 374.400 ;
        RECT 30.000 371.600 30.800 372.400 ;
        RECT 33.200 371.600 34.000 372.400 ;
        RECT 34.800 371.600 35.600 372.400 ;
        RECT 28.400 369.600 29.200 370.400 ;
        RECT 25.200 355.600 26.000 356.400 ;
        RECT 34.800 355.600 35.600 356.400 ;
        RECT 23.700 353.700 25.900 354.300 ;
        RECT 23.600 351.600 24.400 352.400 ;
        RECT 23.600 349.600 24.400 350.400 ;
        RECT 12.400 331.600 13.200 332.400 ;
        RECT 12.500 330.400 13.100 331.600 ;
        RECT 7.600 329.600 8.400 330.400 ;
        RECT 10.800 329.600 11.600 330.400 ;
        RECT 12.400 329.600 13.200 330.400 ;
        RECT 7.700 310.400 8.300 329.600 ;
        RECT 14.000 326.200 14.800 337.800 ;
        RECT 23.700 332.400 24.300 349.600 ;
        RECT 25.300 348.400 25.900 353.700 ;
        RECT 30.000 353.600 30.800 354.400 ;
        RECT 26.800 351.600 27.600 352.400 ;
        RECT 30.100 350.400 30.700 353.600 ;
        RECT 34.900 350.400 35.500 355.600 ;
        RECT 30.000 349.600 30.800 350.400 ;
        RECT 34.800 349.600 35.600 350.400 ;
        RECT 25.200 347.600 26.000 348.400 ;
        RECT 26.800 347.600 27.600 348.400 ;
        RECT 31.600 347.600 32.400 348.400 ;
        RECT 33.200 347.600 34.000 348.400 ;
        RECT 34.800 347.600 35.600 348.400 ;
        RECT 25.300 346.400 25.900 347.600 ;
        RECT 25.200 345.600 26.000 346.400 ;
        RECT 25.300 334.400 25.900 345.600 ;
        RECT 31.700 344.400 32.300 347.600 ;
        RECT 33.300 346.400 33.900 347.600 ;
        RECT 33.200 345.600 34.000 346.400 ;
        RECT 31.600 343.600 32.400 344.400 ;
        RECT 31.700 334.400 32.300 343.600 ;
        RECT 25.200 333.600 26.000 334.400 ;
        RECT 31.600 333.600 32.400 334.400 ;
        RECT 33.200 333.600 34.000 334.400 ;
        RECT 33.300 332.400 33.900 333.600 ;
        RECT 34.900 332.400 35.500 347.600 ;
        RECT 36.500 344.400 37.100 373.600 ;
        RECT 47.700 372.400 48.300 377.600 ;
        RECT 52.400 373.600 53.200 374.400 ;
        RECT 52.500 372.400 53.100 373.600 ;
        RECT 54.100 372.400 54.700 377.600 ;
        RECT 55.600 375.600 56.400 376.400 ;
        RECT 57.200 375.600 58.000 376.400 ;
        RECT 38.000 371.600 38.800 372.400 ;
        RECT 42.800 371.600 43.600 372.400 ;
        RECT 44.400 371.600 45.200 372.400 ;
        RECT 47.600 371.600 48.400 372.400 ;
        RECT 52.400 371.600 53.200 372.400 ;
        RECT 54.000 371.600 54.800 372.400 ;
        RECT 38.100 358.400 38.700 371.600 ;
        RECT 42.900 370.400 43.500 371.600 ;
        RECT 42.800 369.600 43.600 370.400 ;
        RECT 39.600 363.600 40.400 364.400 ;
        RECT 38.000 357.600 38.800 358.400 ;
        RECT 39.700 354.400 40.300 363.600 ;
        RECT 42.900 360.400 43.500 369.600 ;
        RECT 42.800 359.600 43.600 360.400 ;
        RECT 46.000 357.600 46.800 358.400 ;
        RECT 39.600 353.600 40.400 354.400 ;
        RECT 38.000 351.600 38.800 352.400 ;
        RECT 46.100 350.400 46.700 357.600 ;
        RECT 54.100 350.400 54.700 371.600 ;
        RECT 55.700 370.400 56.300 375.600 ;
        RECT 55.600 369.600 56.400 370.400 ;
        RECT 58.800 370.300 59.600 370.400 ;
        RECT 57.300 369.700 59.600 370.300 ;
        RECT 57.300 358.400 57.900 369.700 ;
        RECT 58.800 369.600 59.600 369.700 ;
        RECT 57.200 357.600 58.000 358.400 ;
        RECT 58.800 355.600 59.600 356.400 ;
        RECT 58.900 352.400 59.500 355.600 ;
        RECT 58.800 351.600 59.600 352.400 ;
        RECT 42.800 349.600 43.600 350.400 ;
        RECT 46.000 349.600 46.800 350.400 ;
        RECT 47.600 349.600 48.400 350.400 ;
        RECT 52.400 349.600 53.200 350.400 ;
        RECT 54.000 349.600 54.800 350.400 ;
        RECT 55.600 349.600 56.400 350.400 ;
        RECT 47.700 348.400 48.300 349.600 ;
        RECT 44.400 347.600 45.200 348.400 ;
        RECT 47.600 347.600 48.400 348.400 ;
        RECT 44.500 344.400 45.100 347.600 ;
        RECT 36.400 343.600 37.200 344.400 ;
        RECT 39.600 343.600 40.400 344.400 ;
        RECT 44.400 343.600 45.200 344.400 ;
        RECT 39.700 334.400 40.300 343.600 ;
        RECT 54.100 338.400 54.700 349.600 ;
        RECT 55.700 348.400 56.300 349.600 ;
        RECT 55.600 347.600 56.400 348.400 ;
        RECT 55.700 340.400 56.300 347.600 ;
        RECT 55.600 339.600 56.400 340.400 ;
        RECT 41.200 337.600 42.000 338.400 ;
        RECT 39.600 333.600 40.400 334.400 ;
        RECT 41.300 332.400 41.900 337.600 ;
        RECT 23.600 331.600 24.400 332.400 ;
        RECT 25.200 331.600 26.000 332.400 ;
        RECT 30.000 331.600 30.800 332.400 ;
        RECT 31.600 331.600 32.400 332.400 ;
        RECT 33.200 331.600 34.000 332.400 ;
        RECT 34.800 331.600 35.600 332.400 ;
        RECT 39.600 331.600 40.400 332.400 ;
        RECT 41.200 331.600 42.000 332.400 ;
        RECT 20.400 329.600 21.200 330.400 ;
        RECT 26.800 329.600 27.600 330.400 ;
        RECT 26.900 328.400 27.500 329.600 ;
        RECT 23.600 327.600 24.400 328.400 ;
        RECT 26.800 327.600 27.600 328.400 ;
        RECT 7.600 309.600 8.400 310.400 ;
        RECT 9.200 304.200 10.000 317.800 ;
        RECT 10.800 304.200 11.600 317.800 ;
        RECT 12.400 304.200 13.200 315.800 ;
        RECT 14.000 307.600 14.800 308.400 ;
        RECT 15.600 304.200 16.400 315.800 ;
        RECT 17.200 305.600 18.000 306.400 ;
        RECT 18.800 304.200 19.600 315.800 ;
        RECT 20.400 304.200 21.200 317.800 ;
        RECT 22.000 304.200 22.800 317.800 ;
        RECT 23.600 304.200 24.400 317.800 ;
        RECT 25.200 309.600 26.000 310.400 ;
        RECT 28.400 309.600 29.200 310.400 ;
        RECT 23.600 301.600 24.400 302.400 ;
        RECT 15.600 295.600 16.400 296.400 ;
        RECT 15.700 294.400 16.300 295.600 ;
        RECT 23.700 294.400 24.300 301.600 ;
        RECT 15.600 293.600 16.400 294.400 ;
        RECT 20.400 293.600 21.200 294.400 ;
        RECT 23.600 293.600 24.400 294.400 ;
        RECT 2.800 291.600 3.600 292.400 ;
        RECT 6.000 291.600 6.800 292.400 ;
        RECT 14.000 291.600 14.800 292.400 ;
        RECT 6.100 290.400 6.700 291.600 ;
        RECT 6.000 289.600 6.800 290.400 ;
        RECT 10.800 289.600 11.600 290.400 ;
        RECT 10.900 288.400 11.500 289.600 ;
        RECT 10.800 287.600 11.600 288.400 ;
        RECT 17.200 287.600 18.000 288.400 ;
        RECT 6.000 283.600 6.800 284.400 ;
        RECT 6.100 268.400 6.700 283.600 ;
        RECT 17.300 278.400 17.900 287.600 ;
        RECT 6.000 267.600 6.800 268.400 ;
        RECT 9.200 264.200 10.000 277.800 ;
        RECT 10.800 264.200 11.600 277.800 ;
        RECT 17.200 277.600 18.000 278.400 ;
        RECT 12.400 264.200 13.200 275.800 ;
        RECT 14.000 267.600 14.800 268.400 ;
        RECT 15.600 264.200 16.400 275.800 ;
        RECT 17.200 265.600 18.000 266.400 ;
        RECT 18.800 264.200 19.600 275.800 ;
        RECT 20.400 264.200 21.200 277.800 ;
        RECT 22.000 264.200 22.800 277.800 ;
        RECT 23.600 264.200 24.400 277.800 ;
        RECT 25.300 270.400 25.900 309.600 ;
        RECT 28.500 296.400 29.100 309.600 ;
        RECT 31.700 302.400 32.300 331.600 ;
        RECT 39.700 330.400 40.300 331.600 ;
        RECT 39.600 329.600 40.400 330.400 ;
        RECT 42.800 330.200 43.600 335.800 ;
        RECT 34.800 327.600 35.600 328.400 ;
        RECT 33.200 313.600 34.000 314.400 ;
        RECT 33.300 312.400 33.900 313.600 ;
        RECT 33.200 311.600 34.000 312.400 ;
        RECT 34.900 310.400 35.500 327.600 ;
        RECT 46.000 326.200 46.800 337.800 ;
        RECT 54.000 337.600 54.800 338.400 ;
        RECT 49.200 335.600 50.000 336.400 ;
        RECT 47.600 333.600 48.400 334.400 ;
        RECT 47.700 332.600 48.300 333.600 ;
        RECT 47.600 331.800 48.400 332.600 ;
        RECT 38.000 315.600 38.800 316.400 ;
        RECT 46.000 315.600 46.800 316.400 ;
        RECT 34.800 309.600 35.600 310.400 ;
        RECT 36.400 309.600 37.200 310.400 ;
        RECT 31.600 301.600 32.400 302.400 ;
        RECT 28.400 295.600 29.200 296.400 ;
        RECT 28.500 294.400 29.100 295.600 ;
        RECT 26.800 293.600 27.600 294.400 ;
        RECT 28.400 293.600 29.200 294.400 ;
        RECT 34.900 292.400 35.500 309.600 ;
        RECT 36.500 308.400 37.100 309.600 ;
        RECT 36.400 307.600 37.200 308.400 ;
        RECT 38.100 292.400 38.700 315.600 ;
        RECT 41.200 311.600 42.000 312.400 ;
        RECT 46.100 310.400 46.700 315.600 ;
        RECT 46.000 309.600 46.800 310.400 ;
        RECT 42.800 307.600 43.600 308.400 ;
        RECT 49.300 298.400 49.900 335.600 ;
        RECT 54.000 333.600 54.800 334.400 ;
        RECT 54.100 332.400 54.700 333.600 ;
        RECT 54.000 331.600 54.800 332.400 ;
        RECT 55.600 326.200 56.400 337.800 ;
        RECT 58.900 330.400 59.500 351.600 ;
        RECT 60.500 350.300 61.100 387.600 ;
        RECT 65.300 378.400 65.900 409.600 ;
        RECT 68.500 408.400 69.100 411.600 ;
        RECT 68.400 407.600 69.200 408.400 ;
        RECT 66.800 403.600 67.600 404.400 ;
        RECT 66.900 400.400 67.500 403.600 ;
        RECT 66.800 399.600 67.600 400.400 ;
        RECT 66.800 389.600 67.600 390.400 ;
        RECT 68.400 390.300 69.200 390.400 ;
        RECT 70.100 390.300 70.700 437.600 ;
        RECT 71.700 430.400 72.300 443.700 ;
        RECT 73.200 443.600 74.000 443.700 ;
        RECT 71.600 429.600 72.400 430.400 ;
        RECT 73.200 430.300 74.000 430.400 ;
        RECT 74.900 430.300 75.500 469.600 ;
        RECT 76.400 467.600 77.200 468.400 ;
        RECT 76.500 466.400 77.100 467.600 ;
        RECT 82.900 466.400 83.500 469.600 ;
        RECT 76.400 465.600 77.200 466.400 ;
        RECT 82.800 465.600 83.600 466.400 ;
        RECT 81.200 463.600 82.000 464.400 ;
        RECT 84.500 460.400 85.100 473.600 ;
        RECT 86.000 469.600 86.800 470.400 ;
        RECT 86.100 462.400 86.700 469.600 ;
        RECT 87.700 468.400 88.300 487.600 ;
        RECT 89.300 484.400 89.900 489.700 ;
        RECT 90.800 489.600 91.600 489.700 ;
        RECT 94.000 489.600 94.800 490.400 ;
        RECT 89.200 483.600 90.000 484.400 ;
        RECT 89.300 474.400 89.900 483.600 ;
        RECT 94.100 476.400 94.700 489.600 ;
        RECT 95.700 488.400 96.300 493.600 ;
        RECT 116.400 490.200 117.200 495.800 ;
        RECT 95.600 487.600 96.400 488.400 ;
        RECT 119.600 486.200 120.400 497.800 ;
        RECT 124.400 491.600 125.200 492.400 ;
        RECT 127.600 492.300 128.400 492.400 ;
        RECT 126.100 491.700 128.400 492.300 ;
        RECT 98.800 483.600 99.600 484.400 ;
        RECT 122.800 483.600 123.600 484.400 ;
        RECT 94.000 475.600 94.800 476.400 ;
        RECT 89.200 473.600 90.000 474.400 ;
        RECT 87.600 467.600 88.400 468.400 ;
        RECT 92.400 467.600 93.200 468.400 ;
        RECT 86.000 461.600 86.800 462.400 ;
        RECT 84.400 459.600 85.200 460.400 ;
        RECT 78.000 455.600 78.800 456.400 ;
        RECT 78.100 454.400 78.700 455.600 ;
        RECT 78.000 453.600 78.800 454.400 ;
        RECT 76.400 451.600 77.200 452.400 ;
        RECT 76.500 434.400 77.100 451.600 ;
        RECT 76.400 433.600 77.200 434.400 ;
        RECT 76.500 430.400 77.100 433.600 ;
        RECT 73.200 429.700 75.500 430.300 ;
        RECT 73.200 429.600 74.000 429.700 ;
        RECT 76.400 429.600 77.200 430.400 ;
        RECT 73.300 422.400 73.900 429.600 ;
        RECT 78.100 428.400 78.700 453.600 ;
        RECT 79.600 450.200 80.400 455.800 ;
        RECT 82.800 446.200 83.600 457.800 ;
        RECT 84.500 456.400 85.100 459.600 ;
        RECT 87.700 456.400 88.300 467.600 ;
        RECT 94.000 466.200 94.800 471.800 ;
        RECT 95.600 467.600 96.400 468.400 ;
        RECT 90.800 463.600 91.600 464.400 ;
        RECT 84.400 455.600 85.200 456.400 ;
        RECT 87.600 455.600 88.400 456.400 ;
        RECT 86.000 453.600 86.800 454.400 ;
        RECT 84.400 451.800 85.200 452.600 ;
        RECT 84.500 450.400 85.100 451.800 ;
        RECT 84.400 449.600 85.200 450.400 ;
        RECT 86.100 446.400 86.700 453.600 ;
        RECT 86.000 445.600 86.800 446.400 ;
        RECT 79.600 431.600 80.400 432.400 ;
        RECT 84.400 431.600 85.200 432.400 ;
        RECT 74.800 427.600 75.600 428.400 ;
        RECT 78.000 427.600 78.800 428.400 ;
        RECT 79.700 426.400 80.300 431.600 ;
        RECT 84.400 429.600 85.200 430.400 ;
        RECT 86.100 428.400 86.700 445.600 ;
        RECT 86.000 427.600 86.800 428.400 ;
        RECT 79.600 425.600 80.400 426.400 ;
        RECT 87.600 425.600 88.400 426.400 ;
        RECT 87.700 424.400 88.300 425.600 ;
        RECT 87.600 423.600 88.400 424.400 ;
        RECT 73.200 421.600 74.000 422.400 ;
        RECT 73.200 406.200 74.000 417.800 ;
        RECT 79.600 413.600 80.400 414.400 ;
        RECT 79.700 412.400 80.300 413.600 ;
        RECT 79.600 411.600 80.400 412.400 ;
        RECT 79.600 405.600 80.400 406.400 ;
        RECT 82.800 406.200 83.600 417.800 ;
        RECT 87.700 416.400 88.300 423.600 ;
        RECT 90.900 420.400 91.500 463.600 ;
        RECT 92.400 446.200 93.200 457.800 ;
        RECT 92.400 424.200 93.200 435.800 ;
        RECT 95.700 430.400 96.300 467.600 ;
        RECT 97.200 464.200 98.000 475.800 ;
        RECT 98.900 474.400 99.500 483.600 ;
        RECT 98.800 473.600 99.600 474.400 ;
        RECT 98.800 469.400 99.600 470.200 ;
        RECT 105.200 469.600 106.000 470.400 ;
        RECT 98.900 464.400 99.500 469.400 ;
        RECT 98.800 463.600 99.600 464.400 ;
        RECT 106.800 464.200 107.600 475.800 ;
        RECT 122.900 472.400 123.500 483.600 ;
        RECT 122.800 471.600 123.600 472.400 ;
        RECT 119.600 469.600 120.400 470.400 ;
        RECT 118.000 467.600 118.800 468.400 ;
        RECT 111.600 465.600 112.400 466.400 ;
        RECT 111.700 464.400 112.300 465.600 ;
        RECT 111.600 463.600 112.400 464.400 ;
        RECT 100.400 461.600 101.200 462.400 ;
        RECT 98.800 455.600 99.600 456.400 ;
        RECT 98.900 454.400 99.500 455.600 ;
        RECT 98.800 453.600 99.600 454.400 ;
        RECT 100.500 452.400 101.100 461.600 ;
        RECT 110.000 453.600 110.800 454.400 ;
        RECT 100.400 451.600 101.200 452.400 ;
        RECT 106.800 451.600 107.600 452.400 ;
        RECT 108.400 451.600 109.200 452.400 ;
        RECT 97.200 443.600 98.000 444.400 ;
        RECT 95.600 429.600 96.400 430.400 ;
        RECT 90.800 419.600 91.600 420.400 ;
        RECT 97.300 418.400 97.900 443.600 ;
        RECT 98.800 431.600 99.600 432.400 ;
        RECT 98.900 430.400 99.500 431.600 ;
        RECT 98.800 429.600 99.600 430.400 ;
        RECT 98.800 427.600 99.600 428.400 ;
        RECT 90.800 417.600 91.600 418.400 ;
        RECT 97.200 417.600 98.000 418.400 ;
        RECT 84.400 413.600 85.200 414.400 ;
        RECT 86.000 410.200 86.800 415.800 ;
        RECT 87.600 415.600 88.400 416.400 ;
        RECT 90.900 410.400 91.500 417.600 ;
        RECT 92.400 411.600 93.200 412.400 ;
        RECT 90.800 409.600 91.600 410.400 ;
        RECT 97.200 410.200 98.000 415.800 ;
        RECT 98.900 414.400 99.500 427.600 ;
        RECT 100.500 420.400 101.100 451.600 ;
        RECT 103.600 449.600 104.400 450.400 ;
        RECT 103.700 444.400 104.300 449.600 ;
        RECT 103.600 443.600 104.400 444.400 ;
        RECT 102.000 424.200 102.800 435.800 ;
        RECT 105.200 426.200 106.000 431.800 ;
        RECT 106.800 429.600 107.600 430.400 ;
        RECT 100.400 419.600 101.200 420.400 ;
        RECT 98.800 413.600 99.600 414.400 ;
        RECT 94.000 407.600 94.800 408.400 ;
        RECT 100.400 406.200 101.200 417.800 ;
        RECT 103.600 413.600 104.400 414.400 ;
        RECT 103.700 412.400 104.300 413.600 ;
        RECT 103.600 411.600 104.400 412.400 ;
        RECT 78.000 403.600 78.800 404.400 ;
        RECT 78.100 392.400 78.700 403.600 ;
        RECT 78.000 391.600 78.800 392.400 ;
        RECT 78.100 390.400 78.700 391.600 ;
        RECT 68.400 389.700 70.700 390.300 ;
        RECT 68.400 389.600 69.200 389.700 ;
        RECT 78.000 389.600 78.800 390.400 ;
        RECT 66.900 386.400 67.500 389.600 ;
        RECT 66.800 385.600 67.600 386.400 ;
        RECT 65.200 377.600 66.000 378.400 ;
        RECT 66.900 376.400 67.500 385.600 ;
        RECT 63.600 375.600 64.400 376.400 ;
        RECT 66.800 375.600 67.600 376.400 ;
        RECT 63.700 374.400 64.300 375.600 ;
        RECT 63.600 373.600 64.400 374.400 ;
        RECT 65.200 373.600 66.000 374.400 ;
        RECT 68.500 372.400 69.100 389.600 ;
        RECT 79.700 388.400 80.300 405.600 ;
        RECT 89.200 403.600 90.000 404.400 ;
        RECT 92.400 403.600 93.200 404.400 ;
        RECT 89.300 396.400 89.900 403.600 ;
        RECT 89.200 395.600 90.000 396.400 ;
        RECT 81.200 393.600 82.000 394.400 ;
        RECT 82.800 391.600 83.600 392.400 ;
        RECT 84.400 391.600 85.200 392.400 ;
        RECT 90.800 392.300 91.600 392.400 ;
        RECT 92.500 392.300 93.100 403.600 ;
        RECT 98.800 401.600 99.600 402.400 ;
        RECT 98.900 398.400 99.500 401.600 ;
        RECT 102.000 399.600 102.800 400.400 ;
        RECT 98.800 397.600 99.600 398.400 ;
        RECT 95.600 395.600 96.400 396.400 ;
        RECT 90.800 391.700 93.100 392.300 ;
        RECT 90.800 391.600 91.600 391.700 ;
        RECT 82.900 390.400 83.500 391.600 ;
        RECT 84.500 390.400 85.100 391.600 ;
        RECT 82.800 390.300 83.600 390.400 ;
        RECT 81.300 389.700 83.600 390.300 ;
        RECT 70.000 387.600 70.800 388.400 ;
        RECT 79.600 387.600 80.400 388.400 ;
        RECT 70.100 386.400 70.700 387.600 ;
        RECT 70.000 385.600 70.800 386.400 ;
        RECT 71.600 383.600 72.400 384.400 ;
        RECT 74.800 383.600 75.600 384.400 ;
        RECT 79.600 383.600 80.400 384.400 ;
        RECT 70.000 375.600 70.800 376.400 ;
        RECT 70.000 373.600 70.800 374.400 ;
        RECT 71.700 374.300 72.300 383.600 ;
        RECT 74.900 382.400 75.500 383.600 ;
        RECT 74.800 381.600 75.600 382.400 ;
        RECT 79.700 376.400 80.300 383.600 ;
        RECT 79.600 375.600 80.400 376.400 ;
        RECT 81.300 374.400 81.900 389.700 ;
        RECT 82.800 389.600 83.600 389.700 ;
        RECT 84.400 389.600 85.200 390.400 ;
        RECT 95.700 388.400 96.300 395.600 ;
        RECT 97.200 389.600 98.000 390.400 ;
        RECT 87.600 387.600 88.400 388.400 ;
        RECT 95.600 387.600 96.400 388.400 ;
        RECT 87.700 384.400 88.300 387.600 ;
        RECT 97.300 386.400 97.900 389.600 ;
        RECT 102.100 388.300 102.700 399.600 ;
        RECT 103.600 395.600 104.400 396.400 ;
        RECT 103.700 390.400 104.300 395.600 ;
        RECT 103.600 389.600 104.400 390.400 ;
        RECT 105.200 389.600 106.000 390.400 ;
        RECT 103.600 388.300 104.400 388.400 ;
        RECT 102.100 387.700 104.400 388.300 ;
        RECT 103.600 387.600 104.400 387.700 ;
        RECT 97.200 385.600 98.000 386.400 ;
        RECT 87.600 383.600 88.400 384.400 ;
        RECT 90.800 383.600 91.600 384.400 ;
        RECT 82.800 375.600 83.600 376.400 ;
        RECT 73.200 374.300 74.000 374.400 ;
        RECT 71.700 373.700 74.000 374.300 ;
        RECT 73.200 373.600 74.000 373.700 ;
        RECT 81.200 373.600 82.000 374.400 ;
        RECT 62.000 371.600 62.800 372.400 ;
        RECT 68.400 371.600 69.200 372.400 ;
        RECT 62.100 370.400 62.700 371.600 ;
        RECT 70.100 370.400 70.700 373.600 ;
        RECT 82.900 372.400 83.500 375.600 ;
        RECT 73.200 371.600 74.000 372.400 ;
        RECT 79.600 371.600 80.400 372.400 ;
        RECT 82.800 371.600 83.600 372.400 ;
        RECT 73.300 370.400 73.900 371.600 ;
        RECT 62.000 369.600 62.800 370.400 ;
        RECT 70.000 369.600 70.800 370.400 ;
        RECT 73.200 369.600 74.000 370.400 ;
        RECT 78.000 369.600 78.800 370.400 ;
        RECT 62.000 367.600 62.800 368.400 ;
        RECT 66.800 365.600 67.600 366.400 ;
        RECT 70.100 356.400 70.700 369.600 ;
        RECT 71.600 363.600 72.400 364.400 ;
        RECT 70.000 355.600 70.800 356.400 ;
        RECT 68.400 353.600 69.200 354.400 ;
        RECT 65.200 351.600 66.000 352.400 ;
        RECT 62.000 350.300 62.800 350.400 ;
        RECT 60.500 349.700 62.800 350.300 ;
        RECT 62.000 349.600 62.800 349.700 ;
        RECT 63.600 349.600 64.400 350.400 ;
        RECT 62.100 348.400 62.700 349.600 ;
        RECT 62.000 347.600 62.800 348.400 ;
        RECT 60.400 339.600 61.200 340.400 ;
        RECT 60.500 338.400 61.100 339.600 ;
        RECT 65.300 338.400 65.900 351.600 ;
        RECT 68.500 350.400 69.100 353.600 ;
        RECT 71.700 352.400 72.300 363.600 ;
        RECT 70.000 351.600 70.800 352.400 ;
        RECT 71.600 351.600 72.400 352.400 ;
        RECT 73.300 350.400 73.900 369.600 ;
        RECT 78.100 366.400 78.700 369.600 ;
        RECT 79.600 367.600 80.400 368.400 ;
        RECT 78.000 365.600 78.800 366.400 ;
        RECT 74.800 351.600 75.600 352.400 ;
        RECT 66.800 349.600 67.600 350.400 ;
        RECT 68.400 349.600 69.200 350.400 ;
        RECT 73.200 349.600 74.000 350.400 ;
        RECT 66.900 342.400 67.500 349.600 ;
        RECT 73.300 348.400 73.900 349.600 ;
        RECT 74.900 348.400 75.500 351.600 ;
        RECT 78.000 349.600 78.800 350.400 ;
        RECT 73.200 347.600 74.000 348.400 ;
        RECT 74.800 347.600 75.600 348.400 ;
        RECT 76.400 347.600 77.200 348.400 ;
        RECT 71.600 345.600 72.400 346.400 ;
        RECT 70.000 343.600 70.800 344.400 ;
        RECT 66.800 341.600 67.600 342.400 ;
        RECT 60.400 337.600 61.200 338.400 ;
        RECT 65.200 337.600 66.000 338.400 ;
        RECT 70.100 336.400 70.700 343.600 ;
        RECT 71.700 336.400 72.300 345.600 ;
        RECT 76.500 344.400 77.100 347.600 ;
        RECT 76.400 343.600 77.200 344.400 ;
        RECT 70.000 335.600 70.800 336.400 ;
        RECT 71.600 335.600 72.400 336.400 ;
        RECT 62.000 333.600 62.800 334.400 ;
        RECT 70.000 333.600 70.800 334.400 ;
        RECT 71.600 333.600 72.400 334.400 ;
        RECT 62.100 332.400 62.700 333.600 ;
        RECT 62.000 331.600 62.800 332.400 ;
        RECT 58.800 329.600 59.600 330.400 ;
        RECT 65.200 329.600 66.000 330.400 ;
        RECT 70.100 328.400 70.700 333.600 ;
        RECT 73.200 330.200 74.000 335.800 ;
        RECT 70.000 327.600 70.800 328.400 ;
        RECT 76.400 326.200 77.200 337.800 ;
        RECT 79.700 334.400 80.300 367.600 ;
        RECT 86.000 363.600 86.800 364.400 ;
        RECT 82.800 351.600 83.600 352.400 ;
        RECT 81.200 343.600 82.000 344.400 ;
        RECT 79.600 333.600 80.400 334.400 ;
        RECT 81.300 332.400 81.900 343.600 ;
        RECT 82.900 342.400 83.500 351.600 ;
        RECT 86.100 350.400 86.700 363.600 ;
        RECT 86.000 349.600 86.800 350.400 ;
        RECT 87.700 348.400 88.300 383.600 ;
        RECT 89.200 374.300 90.000 374.400 ;
        RECT 90.900 374.300 91.500 383.600 ;
        RECT 95.600 379.600 96.400 380.400 ;
        RECT 95.700 374.400 96.300 379.600 ;
        RECT 89.200 373.700 91.500 374.300 ;
        RECT 89.200 373.600 90.000 373.700 ;
        RECT 95.600 373.600 96.400 374.400 ;
        RECT 97.300 372.400 97.900 385.600 ;
        RECT 90.800 371.600 91.600 372.400 ;
        RECT 95.600 371.600 96.400 372.400 ;
        RECT 97.200 371.600 98.000 372.400 ;
        RECT 103.600 371.600 104.400 372.400 ;
        RECT 94.000 369.600 94.800 370.400 ;
        RECT 94.100 366.400 94.700 369.600 ;
        RECT 94.000 365.600 94.800 366.400 ;
        RECT 90.800 363.600 91.600 364.400 ;
        RECT 94.000 363.600 94.800 364.400 ;
        RECT 89.200 351.600 90.000 352.400 ;
        RECT 87.600 347.600 88.400 348.400 ;
        RECT 87.700 346.400 88.300 347.600 ;
        RECT 87.600 345.600 88.400 346.400 ;
        RECT 82.800 341.600 83.600 342.400 ;
        RECT 82.900 338.400 83.500 341.600 ;
        RECT 82.800 337.600 83.600 338.400 ;
        RECT 81.200 331.600 82.000 332.400 ;
        RECT 84.400 331.600 85.200 332.400 ;
        RECT 84.500 330.400 85.100 331.600 ;
        RECT 84.400 329.600 85.200 330.400 ;
        RECT 86.000 326.200 86.800 337.800 ;
        RECT 66.800 323.600 67.600 324.400 ;
        RECT 66.900 316.400 67.500 323.600 ;
        RECT 66.800 315.600 67.600 316.400 ;
        RECT 60.400 313.600 61.200 314.400 ;
        RECT 60.500 312.400 61.100 313.600 ;
        RECT 50.800 311.600 51.600 312.400 ;
        RECT 60.400 311.600 61.200 312.400 ;
        RECT 50.900 306.400 51.500 311.600 ;
        RECT 55.600 307.600 56.400 308.400 ;
        RECT 57.200 307.600 58.000 308.400 ;
        RECT 60.400 307.600 61.200 308.400 ;
        RECT 50.800 305.600 51.600 306.400 ;
        RECT 55.600 305.600 56.400 306.400 ;
        RECT 54.000 303.600 54.800 304.400 ;
        RECT 49.200 297.600 50.000 298.400 ;
        RECT 42.800 295.600 43.600 296.400 ;
        RECT 54.100 296.300 54.700 303.600 ;
        RECT 55.700 298.400 56.300 305.600 ;
        RECT 55.600 297.600 56.400 298.400 ;
        RECT 54.100 295.700 56.300 296.300 ;
        RECT 42.900 292.400 43.500 295.600 ;
        RECT 44.400 293.600 45.200 294.400 ;
        RECT 54.000 293.600 54.800 294.400 ;
        RECT 26.800 291.600 27.600 292.400 ;
        RECT 30.000 291.600 30.800 292.400 ;
        RECT 34.800 291.600 35.600 292.400 ;
        RECT 38.000 291.600 38.800 292.400 ;
        RECT 42.800 291.600 43.600 292.400 ;
        RECT 47.600 291.600 48.400 292.400 ;
        RECT 52.400 291.600 53.200 292.400 ;
        RECT 25.200 269.600 26.000 270.400 ;
        RECT 20.400 261.600 21.200 262.400 ;
        RECT 25.300 262.300 25.900 269.600 ;
        RECT 26.900 262.400 27.500 291.600 ;
        RECT 38.100 290.400 38.700 291.600 ;
        RECT 33.200 289.600 34.000 290.400 ;
        RECT 38.000 289.600 38.800 290.400 ;
        RECT 33.300 288.400 33.900 289.600 ;
        RECT 42.900 288.400 43.500 291.600 ;
        RECT 47.700 290.400 48.300 291.600 ;
        RECT 47.600 289.600 48.400 290.400 ;
        RECT 33.200 287.600 34.000 288.400 ;
        RECT 42.800 287.600 43.600 288.400 ;
        RECT 38.000 283.600 38.800 284.400 ;
        RECT 33.200 277.600 34.000 278.400 ;
        RECT 38.100 270.400 38.700 283.600 ;
        RECT 47.700 278.400 48.300 289.600 ;
        RECT 52.500 288.400 53.100 291.600 ;
        RECT 55.700 290.400 56.300 295.700 ;
        RECT 55.600 289.600 56.400 290.400 ;
        RECT 52.400 287.600 53.200 288.400 ;
        RECT 47.600 277.600 48.400 278.400 ;
        RECT 50.800 271.600 51.600 272.400 ;
        RECT 38.000 269.600 38.800 270.400 ;
        RECT 36.400 267.600 37.200 268.400 ;
        RECT 49.200 267.600 50.000 268.400 ;
        RECT 36.500 266.400 37.100 267.600 ;
        RECT 36.400 265.600 37.200 266.400 ;
        RECT 31.600 263.600 32.400 264.400 ;
        RECT 23.700 261.700 25.900 262.300 ;
        RECT 12.400 259.600 13.200 260.400 ;
        RECT 12.500 258.400 13.100 259.600 ;
        RECT 12.400 257.600 13.200 258.400 ;
        RECT 10.800 255.600 11.600 256.400 ;
        RECT 14.000 255.600 14.800 256.400 ;
        RECT 10.900 252.400 11.500 255.600 ;
        RECT 4.400 251.600 5.200 252.400 ;
        RECT 10.800 251.600 11.600 252.400 ;
        RECT 4.500 250.400 5.100 251.600 ;
        RECT 4.400 249.600 5.200 250.400 ;
        RECT 20.500 238.400 21.100 261.600 ;
        RECT 23.700 252.400 24.300 261.700 ;
        RECT 26.800 261.600 27.600 262.400 ;
        RECT 23.600 251.600 24.400 252.400 ;
        RECT 25.200 244.200 26.000 257.800 ;
        RECT 26.800 244.200 27.600 257.800 ;
        RECT 28.400 244.200 29.200 257.800 ;
        RECT 30.000 246.200 30.800 257.800 ;
        RECT 31.700 256.400 32.300 263.600 ;
        RECT 31.600 255.600 32.400 256.400 ;
        RECT 33.200 246.200 34.000 257.800 ;
        RECT 34.800 253.600 35.600 254.400 ;
        RECT 36.400 246.200 37.200 257.800 ;
        RECT 38.000 244.200 38.800 257.800 ;
        RECT 39.600 244.200 40.400 257.800 ;
        RECT 44.400 251.600 45.200 252.400 ;
        RECT 20.400 237.600 21.200 238.400 ;
        RECT 18.800 229.600 19.600 230.400 ;
        RECT 14.000 227.600 14.800 228.400 ;
        RECT 2.800 223.600 3.600 224.400 ;
        RECT 2.900 218.400 3.500 223.600 ;
        RECT 2.800 217.600 3.600 218.400 ;
        RECT 14.100 216.400 14.700 227.600 ;
        RECT 18.800 225.600 19.600 226.400 ;
        RECT 23.600 225.600 24.400 226.400 ;
        RECT 33.200 224.200 34.000 237.800 ;
        RECT 34.800 224.200 35.600 237.800 ;
        RECT 36.400 224.200 37.200 237.800 ;
        RECT 38.000 224.200 38.800 235.800 ;
        RECT 39.600 225.600 40.400 226.400 ;
        RECT 39.700 218.400 40.300 225.600 ;
        RECT 41.200 224.200 42.000 235.800 ;
        RECT 42.800 227.600 43.600 228.400 ;
        RECT 44.400 224.200 45.200 235.800 ;
        RECT 46.000 224.200 46.800 237.800 ;
        RECT 47.600 224.200 48.400 237.800 ;
        RECT 14.000 215.600 14.800 216.400 ;
        RECT 9.200 213.600 10.000 214.400 ;
        RECT 6.000 211.600 6.800 212.400 ;
        RECT 6.100 190.400 6.700 211.600 ;
        RECT 9.200 209.600 10.000 210.400 ;
        RECT 9.300 202.400 9.900 209.600 ;
        RECT 10.800 203.600 11.600 204.400 ;
        RECT 18.800 204.200 19.600 217.800 ;
        RECT 20.400 204.200 21.200 217.800 ;
        RECT 22.000 206.200 22.800 217.800 ;
        RECT 23.600 213.600 24.400 214.400 ;
        RECT 23.600 211.600 24.400 212.400 ;
        RECT 9.200 201.600 10.000 202.400 ;
        RECT 10.900 192.400 11.500 203.600 ;
        RECT 14.000 201.600 14.800 202.400 ;
        RECT 14.100 198.400 14.700 201.600 ;
        RECT 14.000 197.600 14.800 198.400 ;
        RECT 9.200 191.600 10.000 192.400 ;
        RECT 10.800 191.600 11.600 192.400 ;
        RECT 23.700 190.400 24.300 211.600 ;
        RECT 25.200 206.200 26.000 217.800 ;
        RECT 26.800 217.600 27.600 218.400 ;
        RECT 39.600 218.300 40.400 218.400 ;
        RECT 26.900 216.400 27.500 217.600 ;
        RECT 26.800 215.600 27.600 216.400 ;
        RECT 28.400 206.200 29.200 217.800 ;
        RECT 30.000 204.200 30.800 217.800 ;
        RECT 31.600 204.200 32.400 217.800 ;
        RECT 33.200 204.200 34.000 217.800 ;
        RECT 39.600 217.700 41.900 218.300 ;
        RECT 39.600 217.600 40.400 217.700 ;
        RECT 6.000 189.600 6.800 190.400 ;
        RECT 7.600 189.600 8.400 190.400 ;
        RECT 14.000 189.600 14.800 190.400 ;
        RECT 23.600 189.600 24.400 190.400 ;
        RECT 6.000 173.600 6.800 174.400 ;
        RECT 6.100 158.400 6.700 173.600 ;
        RECT 6.000 157.600 6.800 158.400 ;
        RECT 2.800 151.600 3.600 152.400 ;
        RECT 2.900 146.400 3.500 151.600 ;
        RECT 6.000 150.300 6.800 150.400 ;
        RECT 7.700 150.300 8.300 189.600 ;
        RECT 9.200 185.600 10.000 186.400 ;
        RECT 14.100 184.400 14.700 189.600 ;
        RECT 15.600 187.600 16.400 188.400 ;
        RECT 14.000 183.600 14.800 184.400 ;
        RECT 23.700 182.300 24.300 189.600 ;
        RECT 25.200 184.200 26.000 197.800 ;
        RECT 26.800 184.200 27.600 197.800 ;
        RECT 28.400 184.200 29.200 195.800 ;
        RECT 30.000 187.600 30.800 188.400 ;
        RECT 30.100 186.400 30.700 187.600 ;
        RECT 30.000 185.600 30.800 186.400 ;
        RECT 31.600 184.200 32.400 195.800 ;
        RECT 33.200 185.600 34.000 186.400 ;
        RECT 23.700 181.700 25.900 182.300 ;
        RECT 9.200 164.200 10.000 177.800 ;
        RECT 10.800 164.200 11.600 177.800 ;
        RECT 12.400 166.200 13.200 177.800 ;
        RECT 14.000 173.600 14.800 174.400 ;
        RECT 14.000 171.600 14.800 172.400 ;
        RECT 14.100 162.400 14.700 171.600 ;
        RECT 15.600 166.200 16.400 177.800 ;
        RECT 17.200 175.600 18.000 176.400 ;
        RECT 18.800 166.200 19.600 177.800 ;
        RECT 20.400 164.200 21.200 177.800 ;
        RECT 22.000 164.200 22.800 177.800 ;
        RECT 23.600 164.200 24.400 177.800 ;
        RECT 25.300 172.400 25.900 181.700 ;
        RECT 33.300 176.400 33.900 185.600 ;
        RECT 34.800 184.200 35.600 195.800 ;
        RECT 36.400 184.200 37.200 197.800 ;
        RECT 38.000 184.200 38.800 197.800 ;
        RECT 39.600 184.200 40.400 197.800 ;
        RECT 33.200 175.600 34.000 176.400 ;
        RECT 25.200 171.600 26.000 172.400 ;
        RECT 36.400 170.200 37.200 175.800 ;
        RECT 38.000 175.600 38.800 176.400 ;
        RECT 33.200 167.600 34.000 168.400 ;
        RECT 9.200 161.600 10.000 162.400 ;
        RECT 14.000 161.600 14.800 162.400 ;
        RECT 6.000 149.700 8.300 150.300 ;
        RECT 6.000 149.600 6.800 149.700 ;
        RECT 2.800 145.600 3.600 146.400 ;
        RECT 1.200 130.200 2.000 135.800 ;
        RECT 4.400 126.200 5.200 137.800 ;
        RECT 1.200 106.200 2.000 111.800 ;
        RECT 2.800 111.600 3.600 112.400 ;
        RECT 1.200 103.600 2.000 104.400 ;
        RECT 1.300 98.400 1.900 103.600 ;
        RECT 1.200 97.600 2.000 98.400 ;
        RECT 1.200 91.600 2.000 92.400 ;
        RECT 1.300 90.400 1.900 91.600 ;
        RECT 1.200 89.600 2.000 90.400 ;
        RECT 1.200 66.200 2.000 71.800 ;
        RECT 1.200 50.200 2.000 55.800 ;
        RECT 2.900 30.400 3.500 111.600 ;
        RECT 4.400 104.200 5.200 115.800 ;
        RECT 6.100 112.400 6.700 149.600 ;
        RECT 7.600 137.600 8.400 138.400 ;
        RECT 7.700 132.400 8.300 137.600 ;
        RECT 7.600 131.600 8.400 132.400 ;
        RECT 6.000 111.600 6.800 112.400 ;
        RECT 6.000 109.400 6.800 110.200 ;
        RECT 6.100 104.400 6.700 109.400 ;
        RECT 6.000 103.600 6.800 104.400 ;
        RECT 9.300 102.300 9.900 161.600 ;
        RECT 28.400 157.600 29.200 158.400 ;
        RECT 10.800 151.600 11.600 152.400 ;
        RECT 28.500 150.400 29.100 157.600 ;
        RECT 33.300 152.400 33.900 167.600 ;
        RECT 33.200 151.600 34.000 152.400 ;
        RECT 34.800 151.600 35.600 152.400 ;
        RECT 14.000 149.600 14.800 150.400 ;
        RECT 22.000 149.600 22.800 150.400 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 31.600 149.600 32.400 150.400 ;
        RECT 18.800 147.600 19.600 148.400 ;
        RECT 12.400 131.600 13.200 132.400 ;
        RECT 12.500 110.400 13.100 131.600 ;
        RECT 14.000 126.200 14.800 137.800 ;
        RECT 18.800 123.600 19.600 124.400 ;
        RECT 12.400 109.600 13.200 110.400 ;
        RECT 14.000 104.200 14.800 115.800 ;
        RECT 22.100 112.400 22.700 149.600 ;
        RECT 31.700 148.400 32.300 149.600 ;
        RECT 23.600 147.600 24.400 148.400 ;
        RECT 30.000 147.600 30.800 148.400 ;
        RECT 31.600 147.600 32.400 148.400 ;
        RECT 34.800 147.600 35.600 148.400 ;
        RECT 23.700 134.300 24.300 147.600 ;
        RECT 31.600 145.600 32.400 146.400 ;
        RECT 25.200 143.600 26.000 144.400 ;
        RECT 25.300 136.300 25.900 143.600 ;
        RECT 26.800 137.600 27.600 138.400 ;
        RECT 25.300 135.700 27.500 136.300 ;
        RECT 26.900 134.400 27.500 135.700 ;
        RECT 31.700 134.400 32.300 145.600 ;
        RECT 25.200 134.300 26.000 134.400 ;
        RECT 23.700 133.700 26.000 134.300 ;
        RECT 25.200 133.600 26.000 133.700 ;
        RECT 26.800 133.600 27.600 134.400 ;
        RECT 31.600 133.600 32.400 134.400 ;
        RECT 26.900 132.400 27.500 133.600 ;
        RECT 26.800 131.600 27.600 132.400 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 23.600 129.600 24.400 130.400 ;
        RECT 26.800 129.600 27.600 130.400 ;
        RECT 28.400 123.600 29.200 124.400 ;
        RECT 22.000 111.600 22.800 112.400 ;
        RECT 25.200 111.600 26.000 112.400 ;
        RECT 25.300 110.400 25.900 111.600 ;
        RECT 28.500 110.400 29.100 123.600 ;
        RECT 30.100 118.400 30.700 131.600 ;
        RECT 33.200 130.200 34.000 135.800 ;
        RECT 34.900 134.400 35.500 147.600 ;
        RECT 34.800 133.600 35.600 134.400 ;
        RECT 36.400 126.200 37.200 137.800 ;
        RECT 38.100 136.400 38.700 175.600 ;
        RECT 39.600 166.200 40.400 177.800 ;
        RECT 41.300 176.400 41.900 217.700 ;
        RECT 49.300 216.400 49.900 267.600 ;
        RECT 50.900 266.400 51.500 271.600 ;
        RECT 54.000 269.600 54.800 270.400 ;
        RECT 50.800 265.600 51.600 266.400 ;
        RECT 50.800 263.600 51.600 264.400 ;
        RECT 50.900 254.400 51.500 263.600 ;
        RECT 54.100 260.400 54.700 269.600 ;
        RECT 57.300 268.400 57.900 307.600 ;
        RECT 58.800 303.600 59.600 304.400 ;
        RECT 58.900 272.400 59.500 303.600 ;
        RECT 60.500 294.400 61.100 307.600 ;
        RECT 70.000 304.200 70.800 317.800 ;
        RECT 71.600 304.200 72.400 317.800 ;
        RECT 74.800 317.600 75.600 318.400 ;
        RECT 73.200 304.200 74.000 315.800 ;
        RECT 74.900 308.400 75.500 317.600 ;
        RECT 74.800 307.600 75.600 308.400 ;
        RECT 76.400 304.200 77.200 315.800 ;
        RECT 78.000 305.600 78.800 306.400 ;
        RECT 60.400 293.600 61.200 294.400 ;
        RECT 60.400 291.600 61.200 292.400 ;
        RECT 70.000 284.200 70.800 297.800 ;
        RECT 71.600 284.200 72.400 297.800 ;
        RECT 73.200 286.200 74.000 297.800 ;
        RECT 74.800 293.600 75.600 294.400 ;
        RECT 76.400 286.200 77.200 297.800 ;
        RECT 78.100 296.400 78.700 305.600 ;
        RECT 79.600 304.200 80.400 315.800 ;
        RECT 81.200 304.200 82.000 317.800 ;
        RECT 82.800 304.200 83.600 317.800 ;
        RECT 84.400 304.200 85.200 317.800 ;
        RECT 87.700 310.400 88.300 345.600 ;
        RECT 90.900 340.400 91.500 363.600 ;
        RECT 92.400 357.600 93.200 358.400 ;
        RECT 92.400 349.600 93.200 350.400 ;
        RECT 90.800 339.600 91.600 340.400 ;
        RECT 92.500 338.400 93.100 349.600 ;
        RECT 94.100 342.400 94.700 363.600 ;
        RECT 95.700 356.400 96.300 371.600 ;
        RECT 97.300 364.400 97.900 371.600 ;
        RECT 103.700 370.400 104.300 371.600 ;
        RECT 100.400 369.600 101.200 370.400 ;
        RECT 103.600 369.600 104.400 370.400 ;
        RECT 100.500 368.400 101.100 369.600 ;
        RECT 100.400 367.600 101.200 368.400 ;
        RECT 97.200 363.600 98.000 364.400 ;
        RECT 103.600 363.600 104.400 364.400 ;
        RECT 95.600 355.600 96.400 356.400 ;
        RECT 95.700 348.400 96.300 355.600 ;
        RECT 100.400 351.600 101.200 352.400 ;
        RECT 100.500 350.400 101.100 351.600 ;
        RECT 100.400 349.600 101.200 350.400 ;
        RECT 103.600 349.600 104.400 350.400 ;
        RECT 95.600 347.600 96.400 348.400 ;
        RECT 102.000 347.600 102.800 348.400 ;
        RECT 94.000 341.600 94.800 342.400 ;
        RECT 90.800 337.600 91.600 338.400 ;
        RECT 92.400 337.600 93.200 338.400 ;
        RECT 92.400 333.600 93.200 334.400 ;
        RECT 94.100 332.400 94.700 341.600 ;
        RECT 94.000 331.600 94.800 332.400 ;
        RECT 90.800 323.600 91.600 324.400 ;
        RECT 94.000 323.600 94.800 324.400 ;
        RECT 90.900 312.400 91.500 323.600 ;
        RECT 94.100 318.400 94.700 323.600 ;
        RECT 94.000 317.600 94.800 318.400 ;
        RECT 90.800 311.600 91.600 312.400 ;
        RECT 86.000 309.600 86.800 310.400 ;
        RECT 87.600 309.600 88.400 310.400 ;
        RECT 86.100 306.400 86.700 309.600 ;
        RECT 95.700 308.400 96.300 347.600 ;
        RECT 102.100 344.400 102.700 347.600 ;
        RECT 103.700 344.400 104.300 349.600 ;
        RECT 105.300 348.400 105.900 389.600 ;
        RECT 106.900 358.400 107.500 429.600 ;
        RECT 108.500 428.400 109.100 451.600 ;
        RECT 111.700 446.400 112.300 463.600 ;
        RECT 118.100 456.400 118.700 467.600 ;
        RECT 119.700 462.400 120.300 469.600 ;
        RECT 124.500 468.400 125.100 491.600 ;
        RECT 126.100 470.400 126.700 491.700 ;
        RECT 127.600 491.600 128.400 491.700 ;
        RECT 129.200 486.200 130.000 497.800 ;
        RECT 161.200 495.600 162.000 496.400 ;
        RECT 161.300 494.400 161.900 495.600 ;
        RECT 148.400 493.600 149.200 494.400 ;
        RECT 150.000 493.600 150.800 494.400 ;
        RECT 161.200 493.600 162.000 494.400 ;
        RECT 135.600 491.600 136.400 492.400 ;
        RECT 134.000 483.600 134.800 484.400 ;
        RECT 137.200 483.600 138.000 484.400 ;
        RECT 132.400 471.600 133.200 472.400 ;
        RECT 132.500 470.400 133.100 471.600 ;
        RECT 137.300 470.400 137.900 483.600 ;
        RECT 148.500 482.400 149.100 493.600 ;
        RECT 148.400 481.600 149.200 482.400 ;
        RECT 126.000 469.600 126.800 470.400 ;
        RECT 127.600 469.600 128.400 470.400 ;
        RECT 130.800 469.600 131.600 470.400 ;
        RECT 132.400 469.600 133.200 470.400 ;
        RECT 137.200 469.600 138.000 470.400 ;
        RECT 138.800 469.600 139.600 470.400 ;
        RECT 124.400 467.600 125.200 468.400 ;
        RECT 124.400 465.600 125.200 466.400 ;
        RECT 119.600 461.600 120.400 462.400 ;
        RECT 118.000 455.600 118.800 456.400 ;
        RECT 111.600 445.600 112.400 446.400 ;
        RECT 121.200 446.200 122.000 457.800 ;
        RECT 124.500 454.400 125.100 465.600 ;
        RECT 126.100 454.400 126.700 469.600 ;
        RECT 127.700 464.400 128.300 469.600 ;
        RECT 129.200 467.600 130.000 468.400 ;
        RECT 129.300 466.400 129.900 467.600 ;
        RECT 129.200 465.600 130.000 466.400 ;
        RECT 127.600 463.600 128.400 464.400 ;
        RECT 134.000 463.600 134.800 464.400 ;
        RECT 129.200 461.600 130.000 462.400 ;
        RECT 129.300 456.400 129.900 461.600 ;
        RECT 129.200 455.600 130.000 456.400 ;
        RECT 124.400 453.600 125.200 454.400 ;
        RECT 126.000 453.600 126.800 454.400 ;
        RECT 116.400 444.300 117.200 444.400 ;
        RECT 116.400 443.700 118.700 444.300 ;
        RECT 116.400 443.600 117.200 443.700 ;
        RECT 118.100 430.400 118.700 443.700 ;
        RECT 124.500 438.400 125.100 453.600 ;
        RECT 127.600 451.600 128.400 452.400 ;
        RECT 127.600 445.600 128.400 446.400 ;
        RECT 124.400 437.600 125.200 438.400 ;
        RECT 118.000 429.600 118.800 430.400 ;
        RECT 119.600 429.600 120.400 430.400 ;
        RECT 121.200 429.600 122.000 430.400 ;
        RECT 122.800 429.600 123.600 430.400 ;
        RECT 108.400 427.600 109.200 428.400 ;
        RECT 110.000 406.200 110.800 417.800 ;
        RECT 116.400 413.600 117.200 414.400 ;
        RECT 114.800 409.600 115.600 410.400 ;
        RECT 114.900 406.400 115.500 409.600 ;
        RECT 114.800 405.600 115.600 406.400 ;
        RECT 118.100 394.400 118.700 429.600 ;
        RECT 119.700 422.400 120.300 429.600 ;
        RECT 119.600 421.600 120.400 422.400 ;
        RECT 121.200 409.600 122.000 410.400 ;
        RECT 119.600 403.600 120.400 404.400 ;
        RECT 119.700 394.400 120.300 403.600 ;
        RECT 121.300 398.400 121.900 409.600 ;
        RECT 121.200 397.600 122.000 398.400 ;
        RECT 122.900 396.400 123.500 429.600 ;
        RECT 126.000 427.600 126.800 428.400 ;
        RECT 126.100 414.400 126.700 427.600 ;
        RECT 124.400 413.600 125.200 414.400 ;
        RECT 126.000 413.600 126.800 414.400 ;
        RECT 124.500 412.400 125.100 413.600 ;
        RECT 124.400 411.600 125.200 412.400 ;
        RECT 127.700 410.400 128.300 445.600 ;
        RECT 129.300 438.400 129.900 455.600 ;
        RECT 130.800 446.200 131.600 457.800 ;
        RECT 137.300 456.400 137.900 469.600 ;
        RECT 134.000 450.200 134.800 455.800 ;
        RECT 137.200 455.600 138.000 456.400 ;
        RECT 138.900 452.400 139.500 469.600 ;
        RECT 140.400 463.600 141.200 464.400 ;
        RECT 145.200 464.200 146.000 475.800 ;
        RECT 146.800 463.600 147.600 464.400 ;
        RECT 145.200 453.600 146.000 454.400 ;
        RECT 145.300 452.400 145.900 453.600 ;
        RECT 146.900 452.400 147.500 463.600 ;
        RECT 150.100 462.400 150.700 493.600 ;
        RECT 161.300 492.400 161.900 493.600 ;
        RECT 151.600 491.600 152.400 492.400 ;
        RECT 156.400 491.600 157.200 492.400 ;
        RECT 161.200 491.600 162.000 492.400 ;
        RECT 166.000 491.600 166.800 492.400 ;
        RECT 175.600 491.600 176.400 492.400 ;
        RECT 151.700 490.400 152.300 491.600 ;
        RECT 156.500 490.400 157.100 491.600 ;
        RECT 151.600 489.600 152.400 490.400 ;
        RECT 154.800 489.600 155.600 490.400 ;
        RECT 156.400 489.600 157.200 490.400 ;
        RECT 164.400 489.600 165.200 490.400 ;
        RECT 154.900 488.400 155.500 489.600 ;
        RECT 154.800 487.600 155.600 488.400 ;
        RECT 167.600 487.600 168.400 488.400 ;
        RECT 167.700 484.400 168.300 487.600 ;
        RECT 175.700 486.400 176.300 491.600 ;
        RECT 175.600 485.600 176.400 486.400 ;
        RECT 159.600 483.600 160.400 484.400 ;
        RECT 167.600 483.600 168.400 484.400 ;
        RECT 177.200 484.200 178.000 497.800 ;
        RECT 178.800 484.200 179.600 497.800 ;
        RECT 180.400 484.200 181.200 497.800 ;
        RECT 182.000 486.200 182.800 497.800 ;
        RECT 183.600 495.600 184.400 496.400 ;
        RECT 153.200 469.400 154.000 470.200 ;
        RECT 150.000 461.600 150.800 462.400 ;
        RECT 153.300 458.400 153.900 469.400 ;
        RECT 154.800 464.200 155.600 475.800 ;
        RECT 156.400 467.600 157.200 468.400 ;
        RECT 156.500 464.400 157.100 467.600 ;
        RECT 158.000 466.200 158.800 471.800 ;
        RECT 159.700 468.400 160.300 483.600 ;
        RECT 167.700 474.400 168.300 483.600 ;
        RECT 164.400 473.600 165.200 474.400 ;
        RECT 167.600 473.600 168.400 474.400 ;
        RECT 172.400 471.600 173.200 472.400 ;
        RECT 180.400 471.600 181.200 472.400 ;
        RECT 162.800 469.600 163.600 470.400 ;
        RECT 167.600 469.600 168.400 470.400 ;
        RECT 169.200 469.600 170.000 470.400 ;
        RECT 159.600 467.600 160.400 468.400 ;
        RECT 164.400 467.600 165.200 468.400 ;
        RECT 164.500 466.400 165.100 467.600 ;
        RECT 164.400 465.600 165.200 466.400 ;
        RECT 156.400 463.600 157.200 464.400 ;
        RECT 162.800 463.600 163.600 464.400 ;
        RECT 153.200 457.600 154.000 458.400 ;
        RECT 162.900 454.400 163.500 463.600 ;
        RECT 164.500 456.400 165.100 465.600 ;
        RECT 164.400 455.600 165.200 456.400 ;
        RECT 148.400 453.600 149.200 454.400 ;
        RECT 162.800 453.600 163.600 454.400 ;
        RECT 164.400 453.600 165.200 454.400 ;
        RECT 138.800 451.600 139.600 452.400 ;
        RECT 140.400 452.300 141.200 452.400 ;
        RECT 140.400 451.700 142.700 452.300 ;
        RECT 140.400 451.600 141.200 451.700 ;
        RECT 135.600 443.600 136.400 444.400 ;
        RECT 129.200 437.600 130.000 438.400 ;
        RECT 132.400 429.600 133.200 430.400 ;
        RECT 134.000 429.600 134.800 430.400 ;
        RECT 130.800 415.600 131.600 416.400 ;
        RECT 129.200 411.600 130.000 412.400 ;
        RECT 127.600 409.600 128.400 410.400 ;
        RECT 127.600 407.600 128.400 408.400 ;
        RECT 122.800 395.600 123.600 396.400 ;
        RECT 126.000 395.600 126.800 396.400 ;
        RECT 108.400 393.600 109.200 394.400 ;
        RECT 113.200 393.600 114.000 394.400 ;
        RECT 118.000 393.600 118.800 394.400 ;
        RECT 119.600 393.600 120.400 394.400 ;
        RECT 108.500 392.400 109.100 393.600 ;
        RECT 108.400 391.600 109.200 392.400 ;
        RECT 108.400 389.600 109.200 390.400 ;
        RECT 111.600 383.600 112.400 384.400 ;
        RECT 108.400 371.600 109.200 372.400 ;
        RECT 108.500 370.400 109.100 371.600 ;
        RECT 111.700 370.400 112.300 383.600 ;
        RECT 113.300 370.400 113.900 393.600 ;
        RECT 121.200 391.600 122.000 392.400 ;
        RECT 121.300 390.400 121.900 391.600 ;
        RECT 118.000 389.600 118.800 390.400 ;
        RECT 121.200 389.600 122.000 390.400 ;
        RECT 114.800 385.600 115.600 386.400 ;
        RECT 114.900 382.400 115.500 385.600 ;
        RECT 116.400 383.600 117.200 384.400 ;
        RECT 114.800 381.600 115.600 382.400 ;
        RECT 114.900 372.400 115.500 381.600 ;
        RECT 114.800 371.600 115.600 372.400 ;
        RECT 108.400 369.600 109.200 370.400 ;
        RECT 111.600 369.600 112.400 370.400 ;
        RECT 113.200 369.600 114.000 370.400 ;
        RECT 108.500 366.400 109.100 369.600 ;
        RECT 118.100 368.400 118.700 389.600 ;
        RECT 119.600 387.600 120.400 388.400 ;
        RECT 119.600 371.600 120.400 372.400 ;
        RECT 119.700 370.400 120.300 371.600 ;
        RECT 119.600 369.600 120.400 370.400 ;
        RECT 114.800 367.600 115.600 368.400 ;
        RECT 116.400 367.600 117.200 368.400 ;
        RECT 118.000 367.600 118.800 368.400 ;
        RECT 114.900 366.400 115.500 367.600 ;
        RECT 108.400 365.600 109.200 366.400 ;
        RECT 114.800 365.600 115.600 366.400 ;
        RECT 106.800 357.600 107.600 358.400 ;
        RECT 106.800 353.600 107.600 354.400 ;
        RECT 106.900 352.400 107.500 353.600 ;
        RECT 106.800 351.600 107.600 352.400 ;
        RECT 105.200 347.600 106.000 348.400 ;
        RECT 97.200 343.600 98.000 344.400 ;
        RECT 102.000 343.600 102.800 344.400 ;
        RECT 103.600 343.600 104.400 344.400 ;
        RECT 108.500 336.400 109.100 365.600 ;
        RECT 121.300 358.400 121.900 389.600 ;
        RECT 122.900 374.400 123.500 395.600 ;
        RECT 124.400 393.600 125.200 394.400 ;
        RECT 124.500 392.400 125.100 393.600 ;
        RECT 126.100 392.400 126.700 395.600 ;
        RECT 124.400 391.600 125.200 392.400 ;
        RECT 126.000 391.600 126.800 392.400 ;
        RECT 127.700 390.400 128.300 407.600 ;
        RECT 129.200 403.600 130.000 404.400 ;
        RECT 129.300 396.400 129.900 403.600 ;
        RECT 129.200 395.600 130.000 396.400 ;
        RECT 129.200 391.600 130.000 392.400 ;
        RECT 129.300 390.400 129.900 391.600 ;
        RECT 127.600 389.600 128.400 390.400 ;
        RECT 129.200 389.600 130.000 390.400 ;
        RECT 127.600 387.600 128.400 388.400 ;
        RECT 127.700 384.400 128.300 387.600 ;
        RECT 129.300 386.400 129.900 389.600 ;
        RECT 130.900 388.400 131.500 415.600 ;
        RECT 132.500 404.400 133.100 429.600 ;
        RECT 134.000 421.600 134.800 422.400 ;
        RECT 134.100 412.400 134.700 421.600 ;
        RECT 135.700 416.400 136.300 443.600 ;
        RECT 137.200 439.600 138.000 440.400 ;
        RECT 137.300 438.400 137.900 439.600 ;
        RECT 137.200 437.600 138.000 438.400 ;
        RECT 138.900 436.400 139.500 451.600 ;
        RECT 142.100 450.400 142.700 451.700 ;
        RECT 145.200 451.600 146.000 452.400 ;
        RECT 146.800 451.600 147.600 452.400 ;
        RECT 142.000 449.600 142.800 450.400 ;
        RECT 138.800 435.600 139.600 436.400 ;
        RECT 135.600 415.600 136.400 416.400 ;
        RECT 137.200 415.600 138.000 416.400 ;
        RECT 137.300 414.400 137.900 415.600 ;
        RECT 137.200 413.600 138.000 414.400 ;
        RECT 134.000 411.600 134.800 412.400 ;
        RECT 135.600 411.600 136.400 412.400 ;
        RECT 132.400 403.600 133.200 404.400 ;
        RECT 132.400 395.600 133.200 396.400 ;
        RECT 135.700 394.400 136.300 411.600 ;
        RECT 137.200 409.600 138.000 410.400 ;
        RECT 134.000 393.600 134.800 394.400 ;
        RECT 135.600 393.600 136.400 394.400 ;
        RECT 134.100 390.400 134.700 393.600 ;
        RECT 135.700 392.400 136.300 393.600 ;
        RECT 135.600 391.600 136.400 392.400 ;
        RECT 134.000 389.600 134.800 390.400 ;
        RECT 135.600 389.600 136.400 390.400 ;
        RECT 130.800 387.600 131.600 388.400 ;
        RECT 129.200 385.600 130.000 386.400 ;
        RECT 126.000 383.600 126.800 384.400 ;
        RECT 127.600 383.600 128.400 384.400 ;
        RECT 129.200 383.600 130.000 384.400 ;
        RECT 126.100 376.300 126.700 383.600 ;
        RECT 129.300 378.400 129.900 383.600 ;
        RECT 135.700 382.400 136.300 389.600 ;
        RECT 135.600 381.600 136.400 382.400 ;
        RECT 129.200 377.600 130.000 378.400 ;
        RECT 137.300 376.400 137.900 409.600 ;
        RECT 138.900 400.400 139.500 435.600 ;
        RECT 140.400 423.600 141.200 424.400 ;
        RECT 140.500 420.400 141.100 423.600 ;
        RECT 140.400 419.600 141.200 420.400 ;
        RECT 140.400 412.300 141.200 412.400 ;
        RECT 142.100 412.300 142.700 449.600 ;
        RECT 145.200 424.200 146.000 435.800 ;
        RECT 146.900 432.400 147.500 451.600 ;
        RECT 148.500 440.400 149.100 453.600 ;
        RECT 164.500 452.400 165.100 453.600 ;
        RECT 167.700 452.400 168.300 469.600 ;
        RECT 172.500 466.400 173.100 471.600 ;
        RECT 177.200 469.600 178.000 470.400 ;
        RECT 178.800 469.600 179.600 470.400 ;
        RECT 177.300 468.400 177.900 469.600 ;
        RECT 177.200 467.600 178.000 468.400 ;
        RECT 180.400 467.600 181.200 468.400 ;
        RECT 183.700 468.300 184.300 495.600 ;
        RECT 185.200 486.200 186.000 497.800 ;
        RECT 186.800 493.600 187.600 494.400 ;
        RECT 186.900 492.400 187.500 493.600 ;
        RECT 186.800 491.600 187.600 492.400 ;
        RECT 188.400 486.200 189.200 497.800 ;
        RECT 190.000 484.200 190.800 497.800 ;
        RECT 191.600 484.200 192.400 497.800 ;
        RECT 201.200 495.600 202.000 496.400 ;
        RECT 201.300 494.400 201.900 495.600 ;
        RECT 201.200 493.600 202.000 494.400 ;
        RECT 204.400 493.600 205.200 494.400 ;
        RECT 198.000 491.600 198.800 492.400 ;
        RECT 214.000 491.600 214.800 492.400 ;
        RECT 206.000 483.600 206.800 484.400 ;
        RECT 215.600 484.200 216.400 497.800 ;
        RECT 217.200 484.200 218.000 497.800 ;
        RECT 218.800 484.200 219.600 497.800 ;
        RECT 220.400 486.200 221.200 497.800 ;
        RECT 222.000 495.600 222.800 496.400 ;
        RECT 223.600 486.200 224.400 497.800 ;
        RECT 225.200 493.600 226.000 494.400 ;
        RECT 226.800 486.200 227.600 497.800 ;
        RECT 228.400 484.200 229.200 497.800 ;
        RECT 230.000 484.200 230.800 497.800 ;
        RECT 239.600 495.600 240.400 496.400 ;
        RECT 239.700 494.400 240.300 495.600 ;
        RECT 239.600 493.600 240.400 494.400 ;
        RECT 249.200 493.600 250.000 494.400 ;
        RECT 252.400 493.600 253.200 494.400 ;
        RECT 236.400 491.600 237.200 492.400 ;
        RECT 194.800 469.600 195.600 470.400 ;
        RECT 182.100 467.700 184.300 468.300 ;
        RECT 180.500 466.400 181.100 467.600 ;
        RECT 172.400 465.600 173.200 466.400 ;
        RECT 174.000 465.600 174.800 466.400 ;
        RECT 180.400 465.600 181.200 466.400 ;
        RECT 182.100 464.400 182.700 467.700 ;
        RECT 185.200 467.600 186.000 468.400 ;
        RECT 183.600 465.600 184.400 466.400 ;
        RECT 170.800 463.600 171.600 464.400 ;
        RECT 175.600 463.600 176.400 464.400 ;
        RECT 182.000 463.600 182.800 464.400 ;
        RECT 170.900 454.400 171.500 463.600 ;
        RECT 175.700 458.400 176.300 463.600 ;
        RECT 172.400 457.600 173.200 458.400 ;
        RECT 175.600 457.600 176.400 458.400 ;
        RECT 169.200 453.600 170.000 454.400 ;
        RECT 170.800 453.600 171.600 454.400 ;
        RECT 150.000 451.600 150.800 452.400 ;
        RECT 154.800 451.600 155.600 452.400 ;
        RECT 156.400 451.600 157.200 452.400 ;
        RECT 161.200 451.600 162.000 452.400 ;
        RECT 162.800 451.600 163.600 452.400 ;
        RECT 164.400 451.600 165.200 452.400 ;
        RECT 167.600 451.600 168.400 452.400 ;
        RECT 153.200 449.600 154.000 450.400 ;
        RECT 148.400 439.600 149.200 440.400 ;
        RECT 151.600 433.600 152.400 434.400 ;
        RECT 146.800 431.600 147.600 432.400 ;
        RECT 145.200 416.300 146.000 416.400 ;
        RECT 146.900 416.300 147.500 431.600 ;
        RECT 151.700 430.400 152.300 433.600 ;
        RECT 153.300 430.400 153.900 449.600 ;
        RECT 154.900 438.400 155.500 451.600 ;
        RECT 156.500 448.400 157.100 451.600 ;
        RECT 161.300 450.400 161.900 451.600 ;
        RECT 161.200 449.600 162.000 450.400 ;
        RECT 156.400 447.600 157.200 448.400 ;
        RECT 154.800 438.300 155.600 438.400 ;
        RECT 154.800 437.700 157.100 438.300 ;
        RECT 154.800 437.600 155.600 437.700 ;
        RECT 151.600 429.600 152.400 430.400 ;
        RECT 153.200 429.600 154.000 430.400 ;
        RECT 153.200 427.600 154.000 428.400 ;
        RECT 154.800 424.200 155.600 435.800 ;
        RECT 154.800 417.600 155.600 418.400 ;
        RECT 154.900 416.400 155.500 417.600 ;
        RECT 145.200 415.700 147.500 416.300 ;
        RECT 145.200 415.600 146.000 415.700 ;
        RECT 154.800 415.600 155.600 416.400 ;
        RECT 151.600 413.600 152.400 414.400 ;
        RECT 140.400 411.700 142.700 412.300 ;
        RECT 140.400 411.600 141.200 411.700 ;
        RECT 150.000 411.600 150.800 412.400 ;
        RECT 138.800 399.600 139.600 400.400 ;
        RECT 140.500 398.400 141.100 411.600 ;
        RECT 148.400 407.600 149.200 408.400 ;
        RECT 150.100 408.300 150.700 411.600 ;
        RECT 151.700 410.400 152.300 413.600 ;
        RECT 154.800 411.600 155.600 412.400 ;
        RECT 154.900 410.400 155.500 411.600 ;
        RECT 151.600 409.600 152.400 410.400 ;
        RECT 154.800 409.600 155.600 410.400 ;
        RECT 150.100 407.700 152.300 408.300 ;
        RECT 143.600 403.600 144.400 404.400 ;
        RECT 150.000 403.600 150.800 404.400 ;
        RECT 140.400 397.600 141.200 398.400 ;
        RECT 138.800 395.600 139.600 396.400 ;
        RECT 138.900 392.400 139.500 395.600 ;
        RECT 143.700 394.400 144.300 403.600 ;
        RECT 143.600 393.600 144.400 394.400 ;
        RECT 138.800 391.600 139.600 392.400 ;
        RECT 142.000 391.600 142.800 392.400 ;
        RECT 143.600 391.600 144.400 392.400 ;
        RECT 145.200 391.600 146.000 392.400 ;
        RECT 140.400 389.600 141.200 390.400 ;
        RECT 124.500 375.700 126.700 376.300 ;
        RECT 124.500 374.400 125.100 375.700 ;
        RECT 134.000 375.600 134.800 376.400 ;
        RECT 135.600 375.600 136.400 376.400 ;
        RECT 137.200 375.600 138.000 376.400 ;
        RECT 122.800 373.600 123.600 374.400 ;
        RECT 124.400 373.600 125.200 374.400 ;
        RECT 126.000 373.600 126.800 374.400 ;
        RECT 126.100 372.400 126.700 373.600 ;
        RECT 122.800 371.600 123.600 372.400 ;
        RECT 126.000 371.600 126.800 372.400 ;
        RECT 132.400 371.600 133.200 372.400 ;
        RECT 122.900 370.400 123.500 371.600 ;
        RECT 122.800 369.600 123.600 370.400 ;
        RECT 122.800 365.600 123.600 366.400 ;
        RECT 116.400 357.600 117.200 358.400 ;
        RECT 121.200 357.600 122.000 358.400 ;
        RECT 114.800 353.600 115.600 354.400 ;
        RECT 114.800 350.300 115.600 350.400 ;
        RECT 116.500 350.300 117.100 357.600 ;
        RECT 119.600 353.600 120.400 354.400 ;
        RECT 118.000 351.600 118.800 352.400 ;
        RECT 118.100 350.400 118.700 351.600 ;
        RECT 119.700 350.400 120.300 353.600 ;
        RECT 126.100 352.400 126.700 371.600 ;
        RECT 127.600 361.600 128.400 362.400 ;
        RECT 126.000 351.600 126.800 352.400 ;
        RECT 126.100 350.400 126.700 351.600 ;
        RECT 127.700 350.400 128.300 361.600 ;
        RECT 132.500 356.400 133.100 371.600 ;
        RECT 134.000 367.600 134.800 368.400 ;
        RECT 135.700 368.300 136.300 375.600 ;
        RECT 138.800 373.600 139.600 374.400 ;
        RECT 140.500 372.400 141.100 389.600 ;
        RECT 142.100 374.400 142.700 391.600 ;
        RECT 143.700 390.400 144.300 391.600 ;
        RECT 143.600 389.600 144.400 390.400 ;
        RECT 145.300 388.400 145.900 391.600 ;
        RECT 148.400 389.600 149.200 390.400 ;
        RECT 143.600 387.600 144.400 388.400 ;
        RECT 145.200 387.600 146.000 388.400 ;
        RECT 148.400 387.600 149.200 388.400 ;
        RECT 143.700 386.400 144.300 387.600 ;
        RECT 150.100 386.400 150.700 403.600 ;
        RECT 143.600 385.600 144.400 386.400 ;
        RECT 150.000 385.600 150.800 386.400 ;
        RECT 151.700 382.400 152.300 407.700 ;
        RECT 154.800 407.600 155.600 408.400 ;
        RECT 153.200 389.600 154.000 390.400 ;
        RECT 151.600 381.600 152.400 382.400 ;
        RECT 145.200 379.600 146.000 380.400 ;
        RECT 150.000 379.600 150.800 380.400 ;
        RECT 145.300 376.400 145.900 379.600 ;
        RECT 150.100 378.400 150.700 379.600 ;
        RECT 148.400 377.600 149.200 378.400 ;
        RECT 150.000 377.600 150.800 378.400 ;
        RECT 148.500 376.400 149.100 377.600 ;
        RECT 145.200 375.600 146.000 376.400 ;
        RECT 148.400 375.600 149.200 376.400 ;
        RECT 142.000 373.600 142.800 374.400 ;
        RECT 137.200 371.600 138.000 372.400 ;
        RECT 140.400 371.600 141.200 372.400 ;
        RECT 137.300 370.400 137.900 371.600 ;
        RECT 137.200 369.600 138.000 370.400 ;
        RECT 135.700 367.700 137.900 368.300 ;
        RECT 132.400 355.600 133.200 356.400 ;
        RECT 130.800 351.600 131.600 352.400 ;
        RECT 114.800 349.700 117.100 350.300 ;
        RECT 114.800 349.600 115.600 349.700 ;
        RECT 118.000 349.600 118.800 350.400 ;
        RECT 119.600 349.600 120.400 350.400 ;
        RECT 121.200 349.600 122.000 350.400 ;
        RECT 126.000 349.600 126.800 350.400 ;
        RECT 127.600 349.600 128.400 350.400 ;
        RECT 113.200 347.600 114.000 348.400 ;
        RECT 113.300 346.400 113.900 347.600 ;
        RECT 113.200 345.600 114.000 346.400 ;
        RECT 111.600 343.600 112.400 344.400 ;
        RECT 98.800 335.600 99.600 336.400 ;
        RECT 103.600 335.600 104.400 336.400 ;
        RECT 108.400 335.600 109.200 336.400 ;
        RECT 98.900 332.400 99.500 335.600 ;
        RECT 98.800 331.600 99.600 332.400 ;
        RECT 103.700 330.400 104.300 335.600 ;
        RECT 108.400 331.600 109.200 332.400 ;
        RECT 97.200 329.600 98.000 330.400 ;
        RECT 103.600 329.600 104.400 330.400 ;
        RECT 97.300 328.400 97.900 329.600 ;
        RECT 97.200 327.600 98.000 328.400 ;
        RECT 102.000 327.600 102.800 328.400 ;
        RECT 97.200 321.600 98.000 322.400 ;
        RECT 97.300 318.400 97.900 321.600 ;
        RECT 102.100 318.400 102.700 327.600 ;
        RECT 103.600 323.600 104.400 324.400 ;
        RECT 97.200 317.600 98.000 318.400 ;
        RECT 102.000 317.600 102.800 318.400 ;
        RECT 103.700 314.400 104.300 323.600 ;
        RECT 103.600 313.600 104.400 314.400 ;
        RECT 100.400 311.600 101.200 312.400 ;
        RECT 102.000 309.600 102.800 310.400 ;
        RECT 95.600 307.600 96.400 308.400 ;
        RECT 86.000 305.600 86.800 306.400 ;
        RECT 98.800 305.600 99.600 306.400 ;
        RECT 78.000 295.600 78.800 296.400 ;
        RECT 78.100 286.400 78.700 295.600 ;
        RECT 78.000 285.600 78.800 286.400 ;
        RECT 79.600 286.200 80.400 297.800 ;
        RECT 81.200 284.200 82.000 297.800 ;
        RECT 82.800 284.200 83.600 297.800 ;
        RECT 84.400 284.200 85.200 297.800 ;
        RECT 86.100 292.400 86.700 305.600 ;
        RECT 95.600 293.600 96.400 294.400 ;
        RECT 97.200 293.600 98.000 294.400 ;
        RECT 86.000 291.600 86.800 292.400 ;
        RECT 97.300 290.400 97.900 293.600 ;
        RECT 94.000 289.600 94.800 290.400 ;
        RECT 97.200 289.600 98.000 290.400 ;
        RECT 68.400 277.600 69.200 278.400 ;
        RECT 58.800 271.600 59.600 272.400 ;
        RECT 65.200 271.600 66.000 272.400 ;
        RECT 76.400 269.600 77.200 270.400 ;
        RECT 55.600 267.600 56.400 268.400 ;
        RECT 57.200 267.600 58.000 268.400 ;
        RECT 60.400 267.600 61.200 268.400 ;
        RECT 57.200 265.600 58.000 266.400 ;
        RECT 54.000 259.600 54.800 260.400 ;
        RECT 50.800 253.600 51.600 254.400 ;
        RECT 57.300 250.400 57.900 265.600 ;
        RECT 65.200 263.600 66.000 264.400 ;
        RECT 66.800 263.600 67.600 264.400 ;
        RECT 65.300 260.400 65.900 263.600 ;
        RECT 65.200 259.600 66.000 260.400 ;
        RECT 58.800 251.600 59.600 252.400 ;
        RECT 50.800 249.600 51.600 250.400 ;
        RECT 57.200 249.600 58.000 250.400 ;
        RECT 60.400 244.200 61.200 257.800 ;
        RECT 62.000 244.200 62.800 257.800 ;
        RECT 63.600 244.200 64.400 257.800 ;
        RECT 65.200 246.200 66.000 257.800 ;
        RECT 66.900 256.400 67.500 263.600 ;
        RECT 70.000 259.600 70.800 260.400 ;
        RECT 66.800 255.600 67.600 256.400 ;
        RECT 68.400 246.200 69.200 257.800 ;
        RECT 70.100 254.400 70.700 259.600 ;
        RECT 70.000 253.600 70.800 254.400 ;
        RECT 71.600 246.200 72.400 257.800 ;
        RECT 73.200 244.200 74.000 257.800 ;
        RECT 74.800 244.200 75.600 257.800 ;
        RECT 76.500 252.400 77.100 269.600 ;
        RECT 78.000 264.200 78.800 277.800 ;
        RECT 79.600 264.200 80.400 277.800 ;
        RECT 81.200 264.200 82.000 277.800 ;
        RECT 82.800 264.200 83.600 275.800 ;
        RECT 84.400 265.600 85.200 266.400 ;
        RECT 84.500 264.400 85.100 265.600 ;
        RECT 84.400 263.600 85.200 264.400 ;
        RECT 86.000 264.200 86.800 275.800 ;
        RECT 87.600 269.600 88.400 270.400 ;
        RECT 87.700 268.400 88.300 269.600 ;
        RECT 87.600 267.600 88.400 268.400 ;
        RECT 89.200 264.200 90.000 275.800 ;
        RECT 90.800 264.200 91.600 277.800 ;
        RECT 92.400 264.200 93.200 277.800 ;
        RECT 97.200 269.600 98.000 270.400 ;
        RECT 89.200 259.600 90.000 260.400 ;
        RECT 89.300 258.400 89.900 259.600 ;
        RECT 97.300 258.400 97.900 269.600 ;
        RECT 98.900 260.400 99.500 305.600 ;
        RECT 108.500 294.400 109.100 331.600 ;
        RECT 110.000 330.200 110.800 335.800 ;
        RECT 111.700 332.400 112.300 343.600 ;
        RECT 121.300 338.400 121.900 349.600 ;
        RECT 129.200 345.600 130.000 346.400 ;
        RECT 122.800 343.600 123.600 344.400 ;
        RECT 130.900 338.400 131.500 351.600 ;
        RECT 132.400 349.600 133.200 350.400 ;
        RECT 132.400 345.600 133.200 346.400 ;
        RECT 111.600 331.600 112.400 332.400 ;
        RECT 113.200 326.200 114.000 337.800 ;
        RECT 121.200 337.600 122.000 338.400 ;
        RECT 118.000 333.600 118.800 334.400 ;
        RECT 114.800 331.600 115.600 332.600 ;
        RECT 118.100 330.400 118.700 333.600 ;
        RECT 118.000 329.600 118.800 330.400 ;
        RECT 113.200 309.600 114.000 310.400 ;
        RECT 110.000 307.600 110.800 308.400 ;
        RECT 110.100 298.400 110.700 307.600 ;
        RECT 113.300 306.400 113.900 309.600 ;
        RECT 113.200 305.600 114.000 306.400 ;
        RECT 110.000 297.600 110.800 298.400 ;
        RECT 111.600 297.600 112.400 298.400 ;
        RECT 111.700 294.400 112.300 297.600 ;
        RECT 106.800 293.600 107.600 294.400 ;
        RECT 108.400 293.600 109.200 294.400 ;
        RECT 111.600 293.600 112.400 294.400 ;
        RECT 102.000 291.600 102.800 292.400 ;
        RECT 105.200 291.600 106.000 292.400 ;
        RECT 100.400 289.600 101.200 290.400 ;
        RECT 100.500 274.400 101.100 289.600 ;
        RECT 102.100 278.400 102.700 291.600 ;
        RECT 106.900 290.400 107.500 293.600 ;
        RECT 108.500 290.400 109.100 293.600 ;
        RECT 106.800 289.600 107.600 290.400 ;
        RECT 108.400 289.600 109.200 290.400 ;
        RECT 105.200 287.600 106.000 288.400 ;
        RECT 105.300 278.400 105.900 287.600 ;
        RECT 102.000 277.600 102.800 278.400 ;
        RECT 105.200 277.600 106.000 278.400 ;
        RECT 100.400 273.600 101.200 274.400 ;
        RECT 108.400 271.600 109.200 272.400 ;
        RECT 111.600 269.600 112.400 270.400 ;
        RECT 111.700 268.400 112.300 269.600 ;
        RECT 111.600 267.600 112.400 268.400 ;
        RECT 103.600 265.600 104.400 266.400 ;
        RECT 106.800 265.600 107.600 266.400 ;
        RECT 108.400 265.600 109.200 266.400 ;
        RECT 103.700 260.400 104.300 265.600 ;
        RECT 106.900 262.400 107.500 265.600 ;
        RECT 118.100 264.400 118.700 329.600 ;
        RECT 122.800 326.200 123.600 337.800 ;
        RECT 127.600 337.600 128.400 338.400 ;
        RECT 130.800 337.600 131.600 338.400 ;
        RECT 132.500 330.400 133.100 345.600 ;
        RECT 134.100 334.400 134.700 367.600 ;
        RECT 135.600 355.600 136.400 356.400 ;
        RECT 135.700 350.400 136.300 355.600 ;
        RECT 135.600 349.600 136.400 350.400 ;
        RECT 137.300 348.400 137.900 367.700 ;
        RECT 145.200 367.600 146.000 368.400 ;
        RECT 143.600 363.600 144.400 364.400 ;
        RECT 138.800 351.600 139.600 352.400 ;
        RECT 142.000 349.600 142.800 350.400 ;
        RECT 142.100 348.400 142.700 349.600 ;
        RECT 143.700 348.400 144.300 363.600 ;
        RECT 145.300 348.400 145.900 367.600 ;
        RECT 150.000 357.600 150.800 358.400 ;
        RECT 150.100 352.400 150.700 357.600 ;
        RECT 151.700 352.400 152.300 381.600 ;
        RECT 150.000 351.600 150.800 352.400 ;
        RECT 151.600 351.600 152.400 352.400 ;
        RECT 146.800 349.600 147.600 350.400 ;
        RECT 137.200 347.600 138.000 348.400 ;
        RECT 140.400 347.600 141.200 348.400 ;
        RECT 142.000 347.600 142.800 348.400 ;
        RECT 143.600 347.600 144.400 348.400 ;
        RECT 145.200 347.600 146.000 348.400 ;
        RECT 135.600 343.600 136.400 344.400 ;
        RECT 135.700 338.400 136.300 343.600 ;
        RECT 135.600 337.600 136.400 338.400 ;
        RECT 134.000 333.600 134.800 334.400 ;
        RECT 132.400 329.600 133.200 330.400 ;
        RECT 134.100 324.400 134.700 333.600 ;
        RECT 134.000 323.600 134.800 324.400 ;
        RECT 119.600 304.200 120.400 317.800 ;
        RECT 121.200 304.200 122.000 317.800 ;
        RECT 122.800 304.200 123.600 315.800 ;
        RECT 124.400 307.600 125.200 308.400 ;
        RECT 126.000 304.200 126.800 315.800 ;
        RECT 127.600 305.600 128.400 306.400 ;
        RECT 127.700 302.400 128.300 305.600 ;
        RECT 129.200 304.200 130.000 315.800 ;
        RECT 130.800 304.200 131.600 317.800 ;
        RECT 132.400 304.200 133.200 317.800 ;
        RECT 134.000 304.200 134.800 317.800 ;
        RECT 137.300 314.400 137.900 347.600 ;
        RECT 140.500 346.400 141.100 347.600 ;
        RECT 140.400 345.600 141.200 346.400 ;
        RECT 142.100 344.400 142.700 347.600 ;
        RECT 142.000 343.600 142.800 344.400 ;
        RECT 146.900 342.400 147.500 349.600 ;
        RECT 150.000 343.600 150.800 344.400 ;
        RECT 146.800 341.600 147.600 342.400 ;
        RECT 150.100 338.400 150.700 343.600 ;
        RECT 150.000 337.600 150.800 338.400 ;
        RECT 140.400 335.600 141.200 336.400 ;
        RECT 142.000 335.600 142.800 336.400 ;
        RECT 140.500 332.400 141.100 335.600 ;
        RECT 142.100 334.400 142.700 335.600 ;
        RECT 143.400 335.000 144.200 335.800 ;
        RECT 145.200 335.000 149.400 335.600 ;
        RECT 150.000 335.000 150.800 335.800 ;
        RECT 142.000 333.600 142.800 334.400 ;
        RECT 140.400 331.600 141.200 332.400 ;
        RECT 137.200 313.600 138.000 314.400 ;
        RECT 140.500 310.400 141.100 331.600 ;
        RECT 143.400 330.200 144.000 335.000 ;
        RECT 145.200 334.800 146.000 335.000 ;
        RECT 148.600 334.800 149.400 335.000 ;
        RECT 150.200 334.200 150.800 335.000 ;
        RECT 146.000 333.600 150.800 334.200 ;
        RECT 146.000 333.400 146.800 333.600 ;
        RECT 150.200 330.200 150.800 333.600 ;
        RECT 151.700 332.400 152.300 351.600 ;
        RECT 153.300 348.400 153.900 389.600 ;
        RECT 154.900 388.400 155.500 407.600 ;
        RECT 156.500 390.400 157.100 437.700 ;
        RECT 161.300 436.400 161.900 449.600 ;
        RECT 169.300 440.400 169.900 453.600 ;
        RECT 170.800 451.600 171.600 452.400 ;
        RECT 169.200 440.300 170.000 440.400 ;
        RECT 169.200 439.700 171.500 440.300 ;
        RECT 169.200 439.600 170.000 439.700 ;
        RECT 161.200 435.600 162.000 436.400 ;
        RECT 169.200 433.600 170.000 434.400 ;
        RECT 158.000 426.200 158.800 431.800 ;
        RECT 159.600 431.600 160.400 432.400 ;
        RECT 166.000 431.600 166.800 432.400 ;
        RECT 169.200 431.600 170.000 432.400 ;
        RECT 159.600 429.600 160.400 430.400 ;
        RECT 162.800 429.600 163.600 430.400 ;
        RECT 164.400 428.300 165.200 428.400 ;
        RECT 162.900 427.700 165.200 428.300 ;
        RECT 159.600 423.600 160.400 424.400 ;
        RECT 158.000 391.600 158.800 392.400 ;
        RECT 158.100 390.400 158.700 391.600 ;
        RECT 156.400 389.600 157.200 390.400 ;
        RECT 158.000 389.600 158.800 390.400 ;
        RECT 154.800 387.600 155.600 388.400 ;
        RECT 158.100 380.400 158.700 389.600 ;
        RECT 158.000 379.600 158.800 380.400 ;
        RECT 154.800 366.200 155.600 377.800 ;
        RECT 156.400 353.600 157.200 354.400 ;
        RECT 154.800 351.600 155.600 352.400 ;
        RECT 156.500 350.400 157.100 353.600 ;
        RECT 159.700 352.400 160.300 423.600 ;
        RECT 162.900 414.400 163.500 427.700 ;
        RECT 164.400 427.600 165.200 427.700 ;
        RECT 166.100 414.400 166.700 431.600 ;
        RECT 169.300 430.400 169.900 431.600 ;
        RECT 169.200 429.600 170.000 430.400 ;
        RECT 170.900 428.400 171.500 439.700 ;
        RECT 172.500 430.400 173.100 457.600 ;
        RECT 174.000 451.600 174.800 452.400 ;
        RECT 174.000 449.600 174.800 450.400 ;
        RECT 175.600 450.200 176.400 455.800 ;
        RECT 178.800 446.200 179.600 457.800 ;
        RECT 182.100 454.400 182.700 463.600 ;
        RECT 185.300 454.400 185.900 467.600 ;
        RECT 182.000 453.600 182.800 454.400 ;
        RECT 185.200 453.600 186.000 454.400 ;
        RECT 180.400 451.600 181.200 452.600 ;
        RECT 185.200 449.600 186.000 450.400 ;
        RECT 182.000 447.600 182.800 448.400 ;
        RECT 178.800 435.600 179.600 436.400 ;
        RECT 177.200 431.600 178.000 432.400 ;
        RECT 178.900 430.400 179.500 435.600 ;
        RECT 182.100 432.400 182.700 447.600 ;
        RECT 185.300 438.400 185.900 449.600 ;
        RECT 188.400 446.200 189.200 457.800 ;
        RECT 194.900 456.400 195.500 469.600 ;
        RECT 196.400 464.200 197.200 477.800 ;
        RECT 198.000 464.200 198.800 477.800 ;
        RECT 199.600 464.200 200.400 477.800 ;
        RECT 201.200 464.200 202.000 475.800 ;
        RECT 202.800 465.600 203.600 466.400 ;
        RECT 198.000 461.600 198.800 462.400 ;
        RECT 194.800 455.600 195.600 456.400 ;
        RECT 198.100 452.400 198.700 461.600 ;
        RECT 202.900 458.400 203.500 465.600 ;
        RECT 204.400 464.200 205.200 475.800 ;
        RECT 206.000 467.600 206.800 468.400 ;
        RECT 206.100 458.400 206.700 467.600 ;
        RECT 207.600 464.200 208.400 475.800 ;
        RECT 209.200 464.200 210.000 477.800 ;
        RECT 210.800 464.200 211.600 477.800 ;
        RECT 221.800 471.800 222.600 472.600 ;
        RECT 228.400 471.800 229.200 472.600 ;
        RECT 215.600 469.600 216.400 470.400 ;
        RECT 220.400 467.600 221.200 468.400 ;
        RECT 220.500 462.400 221.100 467.600 ;
        RECT 221.800 467.000 222.400 471.800 ;
        RECT 224.400 468.400 225.200 468.600 ;
        RECT 228.600 468.400 229.200 471.800 ;
        RECT 231.600 469.600 232.400 470.400 ;
        RECT 241.200 469.600 242.000 470.400 ;
        RECT 231.700 468.400 232.300 469.600 ;
        RECT 224.400 467.800 229.200 468.400 ;
        RECT 223.600 467.000 224.400 467.200 ;
        RECT 227.000 467.000 227.800 467.200 ;
        RECT 228.600 467.000 229.200 467.800 ;
        RECT 230.000 467.600 230.800 468.400 ;
        RECT 231.600 467.600 232.400 468.400 ;
        RECT 221.800 466.200 222.600 467.000 ;
        RECT 223.600 466.400 227.800 467.000 ;
        RECT 228.400 466.200 229.200 467.000 ;
        RECT 242.800 464.200 243.600 477.800 ;
        RECT 244.400 464.200 245.200 477.800 ;
        RECT 246.000 464.200 246.800 477.800 ;
        RECT 247.600 464.200 248.400 475.800 ;
        RECT 249.300 466.400 249.900 493.600 ;
        RECT 252.500 482.400 253.100 493.600 ;
        RECT 262.000 491.600 262.800 492.400 ;
        RECT 266.800 484.200 267.600 497.800 ;
        RECT 268.400 484.200 269.200 497.800 ;
        RECT 270.000 486.200 270.800 497.800 ;
        RECT 271.600 493.600 272.400 494.400 ;
        RECT 271.700 484.300 272.300 493.600 ;
        RECT 273.200 486.200 274.000 497.800 ;
        RECT 274.800 495.600 275.600 496.400 ;
        RECT 274.900 494.400 275.500 495.600 ;
        RECT 274.800 493.600 275.600 494.400 ;
        RECT 276.400 486.200 277.200 497.800 ;
        RECT 271.700 483.700 273.900 484.300 ;
        RECT 278.000 484.200 278.800 497.800 ;
        RECT 279.600 484.200 280.400 497.800 ;
        RECT 281.200 484.200 282.000 497.800 ;
        RECT 292.400 493.600 293.200 494.400 ;
        RECT 303.600 493.600 304.400 494.400 ;
        RECT 290.800 491.600 291.600 492.400 ;
        RECT 252.400 481.600 253.200 482.400 ;
        RECT 273.300 478.400 273.900 483.700 ;
        RECT 281.200 481.600 282.000 482.400 ;
        RECT 249.200 465.600 250.000 466.400 ;
        RECT 250.800 464.200 251.600 475.800 ;
        RECT 252.400 467.600 253.200 468.400 ;
        RECT 254.000 464.200 254.800 475.800 ;
        RECT 255.600 464.200 256.400 477.800 ;
        RECT 257.200 464.200 258.000 477.800 ;
        RECT 273.200 477.600 274.000 478.400 ;
        RECT 276.400 471.600 277.200 472.400 ;
        RECT 260.400 469.600 261.200 470.400 ;
        RECT 273.200 469.600 274.000 470.400 ;
        RECT 276.400 469.600 277.200 470.400 ;
        RECT 220.400 461.600 221.200 462.400 ;
        RECT 202.800 457.600 203.600 458.400 ;
        RECT 206.000 457.600 206.800 458.400 ;
        RECT 201.200 455.000 202.000 455.800 ;
        RECT 202.600 455.000 206.800 455.600 ;
        RECT 207.800 455.000 208.600 455.800 ;
        RECT 199.600 453.600 200.400 454.400 ;
        RECT 201.200 454.200 201.800 455.000 ;
        RECT 202.600 454.800 203.400 455.000 ;
        RECT 206.000 454.800 206.800 455.000 ;
        RECT 201.200 453.600 206.000 454.200 ;
        RECT 196.400 451.600 197.200 452.400 ;
        RECT 198.000 451.600 198.800 452.400 ;
        RECT 190.000 447.600 190.800 448.400 ;
        RECT 193.200 447.600 194.000 448.400 ;
        RECT 185.200 437.600 186.000 438.400 ;
        RECT 182.000 431.600 182.800 432.400 ;
        RECT 172.400 429.600 173.200 430.400 ;
        RECT 174.000 429.600 174.800 430.400 ;
        RECT 178.800 429.600 179.600 430.400 ;
        RECT 180.400 429.600 181.200 430.400 ;
        RECT 170.800 427.600 171.600 428.400 ;
        RECT 167.600 419.600 168.400 420.400 ;
        RECT 162.800 413.600 163.600 414.400 ;
        RECT 166.000 413.600 166.800 414.400 ;
        RECT 164.400 411.600 165.200 412.400 ;
        RECT 167.700 410.400 168.300 419.600 ;
        RECT 169.200 415.600 170.000 416.400 ;
        RECT 169.300 412.400 169.900 415.600 ;
        RECT 170.800 413.600 171.600 414.400 ;
        RECT 170.900 412.400 171.500 413.600 ;
        RECT 169.200 411.600 170.000 412.400 ;
        RECT 170.800 411.600 171.600 412.400 ;
        RECT 167.600 409.600 168.400 410.400 ;
        RECT 162.800 389.600 163.600 390.400 ;
        RECT 162.900 382.400 163.500 389.600 ;
        RECT 167.700 388.400 168.300 409.600 ;
        RECT 172.500 406.400 173.100 429.600 ;
        RECT 174.100 420.400 174.700 429.600 ;
        RECT 178.800 427.600 179.600 428.400 ;
        RECT 174.000 419.600 174.800 420.400 ;
        RECT 178.900 414.400 179.500 427.600 ;
        RECT 180.500 426.400 181.100 429.600 ;
        RECT 180.400 425.600 181.200 426.400 ;
        RECT 178.800 414.300 179.600 414.400 ;
        RECT 177.300 413.700 179.600 414.300 ;
        RECT 174.000 409.600 174.800 410.400 ;
        RECT 172.400 405.600 173.200 406.400 ;
        RECT 177.300 396.400 177.900 413.700 ;
        RECT 178.800 413.600 179.600 413.700 ;
        RECT 180.500 412.400 181.100 425.600 ;
        RECT 182.100 418.400 182.700 431.600 ;
        RECT 190.100 430.400 190.700 447.600 ;
        RECT 198.100 440.400 198.700 451.600 ;
        RECT 201.200 450.200 201.800 453.600 ;
        RECT 205.200 453.400 206.000 453.600 ;
        RECT 208.000 450.200 208.600 455.000 ;
        RECT 209.200 453.600 210.000 454.400 ;
        RECT 209.300 452.400 209.900 453.600 ;
        RECT 209.200 451.600 210.000 452.400 ;
        RECT 214.000 451.600 214.800 452.400 ;
        RECT 218.800 451.600 219.600 452.400 ;
        RECT 201.200 449.400 202.000 450.200 ;
        RECT 207.800 449.400 208.600 450.200 ;
        RECT 215.600 449.600 216.400 450.400 ;
        RECT 214.000 447.600 214.800 448.400 ;
        RECT 210.800 443.600 211.600 444.400 ;
        RECT 198.000 439.600 198.800 440.400 ;
        RECT 185.200 429.600 186.000 430.400 ;
        RECT 188.400 429.600 189.200 430.400 ;
        RECT 190.000 429.600 190.800 430.400 ;
        RECT 185.300 426.400 185.900 429.600 ;
        RECT 186.800 427.600 187.600 428.400 ;
        RECT 188.500 426.400 189.100 429.600 ;
        RECT 191.600 427.600 192.400 428.400 ;
        RECT 185.200 425.600 186.000 426.400 ;
        RECT 188.400 425.600 189.200 426.400 ;
        RECT 193.200 425.600 194.000 426.400 ;
        RECT 185.200 423.600 186.000 424.400 ;
        RECT 185.300 418.400 185.900 423.600 ;
        RECT 193.300 418.400 193.900 425.600 ;
        RECT 194.800 423.600 195.600 424.400 ;
        RECT 199.600 424.200 200.400 435.800 ;
        RECT 201.200 429.600 202.000 430.400 ;
        RECT 206.000 429.600 206.800 430.400 ;
        RECT 206.100 424.400 206.700 429.600 ;
        RECT 206.000 423.600 206.800 424.400 ;
        RECT 209.200 424.200 210.000 435.800 ;
        RECT 210.900 430.400 211.500 443.600 ;
        RECT 210.800 429.600 211.600 430.400 ;
        RECT 212.400 426.200 213.200 431.800 ;
        RECT 214.100 426.400 214.700 447.600 ;
        RECT 215.700 428.400 216.300 449.600 ;
        RECT 218.900 438.400 219.500 451.600 ;
        RECT 218.800 437.600 219.600 438.400 ;
        RECT 217.200 431.600 218.000 432.400 ;
        RECT 217.300 430.400 217.900 431.600 ;
        RECT 217.200 429.600 218.000 430.400 ;
        RECT 220.500 428.400 221.100 461.600 ;
        RECT 222.000 449.600 222.800 450.400 ;
        RECT 222.100 448.400 222.700 449.600 ;
        RECT 222.000 447.600 222.800 448.400 ;
        RECT 226.800 447.600 227.600 448.400 ;
        RECT 215.600 427.600 216.400 428.400 ;
        RECT 220.400 427.600 221.200 428.400 ;
        RECT 214.000 425.600 214.800 426.400 ;
        RECT 217.200 425.600 218.000 426.400 ;
        RECT 220.400 426.300 221.200 426.400 ;
        RECT 222.100 426.300 222.700 447.600 ;
        RECT 225.200 443.600 226.000 444.400 ;
        RECT 238.000 444.200 238.800 457.800 ;
        RECT 239.600 444.200 240.400 457.800 ;
        RECT 241.200 444.200 242.000 457.800 ;
        RECT 242.800 446.200 243.600 457.800 ;
        RECT 244.400 457.600 245.200 458.400 ;
        RECT 244.500 456.400 245.100 457.600 ;
        RECT 244.400 455.600 245.200 456.400 ;
        RECT 225.300 434.400 225.900 443.600 ;
        RECT 231.600 437.600 232.400 438.400 ;
        RECT 225.200 433.600 226.000 434.400 ;
        RECT 228.400 431.600 229.200 432.400 ;
        RECT 225.200 429.600 226.000 430.400 ;
        RECT 226.800 430.300 227.600 430.400 ;
        RECT 226.800 429.700 229.100 430.300 ;
        RECT 226.800 429.600 227.600 429.700 ;
        RECT 225.300 428.400 225.900 429.600 ;
        RECT 225.200 427.600 226.000 428.400 ;
        RECT 220.400 425.700 222.700 426.300 ;
        RECT 220.400 425.600 221.200 425.700 ;
        RECT 215.600 423.600 216.400 424.400 ;
        RECT 182.000 417.600 182.800 418.400 ;
        RECT 185.200 417.600 186.000 418.400 ;
        RECT 193.200 417.600 194.000 418.400 ;
        RECT 194.900 414.400 195.500 423.600 ;
        RECT 209.200 421.600 210.000 422.400 ;
        RECT 183.600 413.600 184.400 414.400 ;
        RECT 190.000 413.600 190.800 414.400 ;
        RECT 194.800 413.600 195.600 414.400 ;
        RECT 178.800 411.600 179.600 412.400 ;
        RECT 180.400 411.600 181.200 412.400 ;
        RECT 178.900 410.300 179.500 411.600 ;
        RECT 183.700 410.400 184.300 413.600 ;
        RECT 188.400 411.600 189.200 412.400 ;
        RECT 188.500 410.400 189.100 411.600 ;
        RECT 178.900 409.700 181.100 410.300 ;
        RECT 178.800 399.600 179.600 400.400 ;
        RECT 177.200 395.600 178.000 396.400 ;
        RECT 172.400 391.600 173.200 392.400 ;
        RECT 175.600 391.600 176.400 392.400 ;
        RECT 175.700 390.400 176.300 391.600 ;
        RECT 175.600 389.600 176.400 390.400 ;
        RECT 177.300 388.400 177.900 395.600 ;
        RECT 178.900 390.400 179.500 399.600 ;
        RECT 180.500 390.400 181.100 409.700 ;
        RECT 183.600 409.600 184.400 410.400 ;
        RECT 188.400 409.600 189.200 410.400 ;
        RECT 188.400 393.600 189.200 394.400 ;
        RECT 186.800 391.600 187.600 392.400 ;
        RECT 178.800 389.600 179.600 390.400 ;
        RECT 180.400 389.600 181.200 390.400 ;
        RECT 185.200 390.300 186.000 390.400 ;
        RECT 186.900 390.300 187.500 391.600 ;
        RECT 188.500 390.400 189.100 393.600 ;
        RECT 185.200 389.700 187.500 390.300 ;
        RECT 185.200 389.600 186.000 389.700 ;
        RECT 188.400 389.600 189.200 390.400 ;
        RECT 166.000 387.600 166.800 388.400 ;
        RECT 167.600 387.600 168.400 388.400 ;
        RECT 177.200 387.600 178.000 388.400 ;
        RECT 166.100 384.400 166.700 387.600 ;
        RECT 166.000 383.600 166.800 384.400 ;
        RECT 170.800 383.600 171.600 384.400 ;
        RECT 162.800 381.600 163.600 382.400 ;
        RECT 166.000 381.600 166.800 382.400 ;
        RECT 162.800 373.600 163.600 374.400 ;
        RECT 161.200 371.600 162.000 372.400 ;
        RECT 162.900 370.400 163.500 373.600 ;
        RECT 162.800 369.600 163.600 370.400 ;
        RECT 164.400 366.200 165.200 377.800 ;
        RECT 166.100 362.400 166.700 381.600 ;
        RECT 169.200 379.600 170.000 380.400 ;
        RECT 167.600 370.200 168.400 375.800 ;
        RECT 169.300 372.400 169.900 379.600 ;
        RECT 170.900 372.400 171.500 383.600 ;
        RECT 180.500 382.400 181.100 389.600 ;
        RECT 180.400 381.600 181.200 382.400 ;
        RECT 185.300 378.400 185.900 389.600 ;
        RECT 186.800 387.600 187.600 388.400 ;
        RECT 188.400 387.600 189.200 388.400 ;
        RECT 186.900 386.400 187.500 387.600 ;
        RECT 186.800 385.600 187.600 386.400 ;
        RECT 190.100 384.400 190.700 413.600 ;
        RECT 201.200 411.600 202.000 412.400 ;
        RECT 193.200 403.600 194.000 404.400 ;
        RECT 201.300 402.400 201.900 411.600 ;
        RECT 202.800 404.200 203.600 417.800 ;
        RECT 204.400 404.200 205.200 417.800 ;
        RECT 206.000 404.200 206.800 417.800 ;
        RECT 207.600 406.200 208.400 417.800 ;
        RECT 209.300 416.400 209.900 421.600 ;
        RECT 215.700 420.400 216.300 423.600 ;
        RECT 212.400 419.600 213.200 420.400 ;
        RECT 215.600 419.600 216.400 420.400 ;
        RECT 209.200 415.600 210.000 416.400 ;
        RECT 201.200 401.600 202.000 402.400 ;
        RECT 204.400 401.600 205.200 402.400 ;
        RECT 201.200 393.600 202.000 394.400 ;
        RECT 201.300 392.400 201.900 393.600 ;
        RECT 193.200 391.600 194.000 392.400 ;
        RECT 199.600 391.600 200.400 392.400 ;
        RECT 201.200 391.600 202.000 392.400 ;
        RECT 199.700 390.400 200.300 391.600 ;
        RECT 194.800 389.600 195.600 390.400 ;
        RECT 196.400 389.600 197.200 390.400 ;
        RECT 199.600 389.600 200.400 390.400 ;
        RECT 194.800 387.600 195.600 388.400 ;
        RECT 194.900 384.400 195.500 387.600 ;
        RECT 196.500 386.400 197.100 389.600 ;
        RECT 199.600 387.600 200.400 388.400 ;
        RECT 196.400 385.600 197.200 386.400 ;
        RECT 190.000 383.600 190.800 384.400 ;
        RECT 194.800 383.600 195.600 384.400 ;
        RECT 185.200 377.600 186.000 378.400 ;
        RECT 186.800 377.600 187.600 378.400 ;
        RECT 177.200 375.600 178.000 376.400 ;
        RECT 174.000 373.600 174.800 374.400 ;
        RECT 175.600 373.600 176.400 374.400 ;
        RECT 178.800 373.600 179.600 374.400 ;
        RECT 174.100 372.400 174.700 373.600 ;
        RECT 175.700 372.400 176.300 373.600 ;
        RECT 169.200 371.600 170.000 372.400 ;
        RECT 170.800 371.600 171.600 372.400 ;
        RECT 174.000 371.600 174.800 372.400 ;
        RECT 175.600 371.600 176.400 372.400 ;
        RECT 183.600 371.600 184.400 372.400 ;
        RECT 166.000 361.600 166.800 362.400 ;
        RECT 162.800 353.600 163.600 354.400 ;
        RECT 158.000 351.600 158.800 352.400 ;
        RECT 159.600 351.600 160.400 352.400 ;
        RECT 156.400 349.600 157.200 350.400 ;
        RECT 161.200 349.600 162.000 350.400 ;
        RECT 161.300 348.400 161.900 349.600 ;
        RECT 162.900 348.400 163.500 353.600 ;
        RECT 164.400 351.600 165.200 352.400 ;
        RECT 166.100 350.400 166.700 361.600 ;
        RECT 169.200 355.600 170.000 356.400 ;
        RECT 166.000 349.600 166.800 350.400 ;
        RECT 167.600 349.600 168.400 350.400 ;
        RECT 169.300 348.400 169.900 355.600 ;
        RECT 175.700 350.400 176.300 371.600 ;
        RECT 186.900 370.400 187.500 377.600 ;
        RECT 186.800 369.600 187.600 370.400 ;
        RECT 175.600 349.600 176.400 350.400 ;
        RECT 153.200 347.600 154.000 348.400 ;
        RECT 156.400 347.600 157.200 348.400 ;
        RECT 159.600 347.600 160.400 348.400 ;
        RECT 161.200 347.600 162.000 348.400 ;
        RECT 162.800 347.600 163.600 348.400 ;
        RECT 169.200 347.600 170.000 348.400 ;
        RECT 156.500 334.400 157.100 347.600 ;
        RECT 159.700 342.400 160.300 347.600 ;
        RECT 162.800 345.600 163.600 346.400 ;
        RECT 158.000 341.600 158.800 342.400 ;
        RECT 159.600 341.600 160.400 342.400 ;
        RECT 158.100 338.400 158.700 341.600 ;
        RECT 158.000 337.600 158.800 338.400 ;
        RECT 153.200 333.600 154.000 334.400 ;
        RECT 156.400 333.600 157.200 334.400 ;
        RECT 159.600 333.600 160.400 334.400 ;
        RECT 161.200 333.600 162.000 334.400 ;
        RECT 159.700 332.400 160.300 333.600 ;
        RECT 162.900 332.400 163.500 345.600 ;
        RECT 178.800 344.200 179.600 357.800 ;
        RECT 180.400 344.200 181.200 357.800 ;
        RECT 182.000 344.200 182.800 355.800 ;
        RECT 183.600 347.600 184.400 348.400 ;
        RECT 183.700 344.400 184.300 347.600 ;
        RECT 183.600 343.600 184.400 344.400 ;
        RECT 185.200 344.200 186.000 355.800 ;
        RECT 186.900 346.400 187.500 369.600 ;
        RECT 188.400 364.200 189.200 377.800 ;
        RECT 190.000 364.200 190.800 377.800 ;
        RECT 191.600 366.200 192.400 377.800 ;
        RECT 193.200 375.600 194.000 376.400 ;
        RECT 193.300 374.400 193.900 375.600 ;
        RECT 193.200 373.600 194.000 374.400 ;
        RECT 194.800 366.200 195.600 377.800 ;
        RECT 196.400 377.600 197.200 378.400 ;
        RECT 196.500 376.400 197.100 377.600 ;
        RECT 196.400 375.600 197.200 376.400 ;
        RECT 198.000 366.200 198.800 377.800 ;
        RECT 199.600 364.200 200.400 377.800 ;
        RECT 201.200 364.200 202.000 377.800 ;
        RECT 202.800 364.200 203.600 377.800 ;
        RECT 204.500 372.400 205.100 401.600 ;
        RECT 206.000 384.200 206.800 395.800 ;
        RECT 209.300 390.400 209.900 415.600 ;
        RECT 210.800 406.200 211.600 417.800 ;
        RECT 212.500 414.400 213.100 419.600 ;
        RECT 212.400 413.600 213.200 414.400 ;
        RECT 214.000 406.200 214.800 417.800 ;
        RECT 215.600 404.200 216.400 417.800 ;
        RECT 217.200 404.200 218.000 417.800 ;
        RECT 220.500 414.400 221.100 425.600 ;
        RECT 223.600 423.600 224.400 424.400 ;
        RECT 220.400 413.600 221.200 414.400 ;
        RECT 223.700 412.400 224.300 423.600 ;
        RECT 228.500 418.400 229.100 429.700 ;
        RECT 231.700 428.400 232.300 437.600 ;
        RECT 234.800 431.600 235.600 432.400 ;
        RECT 234.900 430.400 235.500 431.600 ;
        RECT 234.800 429.600 235.600 430.400 ;
        RECT 231.600 427.600 232.400 428.400 ;
        RECT 228.400 417.600 229.200 418.400 ;
        RECT 226.800 413.600 227.600 414.400 ;
        RECT 223.600 411.600 224.400 412.400 ;
        RECT 231.700 410.400 232.300 427.600 ;
        RECT 244.500 426.400 245.100 455.600 ;
        RECT 246.000 446.200 246.800 457.800 ;
        RECT 247.600 453.600 248.400 454.400 ;
        RECT 247.700 444.300 248.300 453.600 ;
        RECT 249.200 446.200 250.000 457.800 ;
        RECT 247.700 443.700 249.900 444.300 ;
        RECT 250.800 444.200 251.600 457.800 ;
        RECT 252.400 444.200 253.200 457.800 ;
        RECT 260.500 452.400 261.100 469.600 ;
        RECT 281.300 468.400 281.900 481.600 ;
        RECT 271.600 467.600 272.400 468.400 ;
        RECT 281.200 467.600 282.000 468.400 ;
        RECT 271.700 452.400 272.300 467.600 ;
        RECT 279.600 465.600 280.400 466.400 ;
        RECT 281.300 460.400 281.900 467.600 ;
        RECT 281.200 459.600 282.000 460.400 ;
        RECT 257.200 451.600 258.000 452.400 ;
        RECT 260.400 451.600 261.200 452.400 ;
        RECT 271.600 451.600 272.400 452.400 ;
        RECT 247.600 433.600 248.400 434.400 ;
        RECT 246.000 427.600 246.800 428.400 ;
        RECT 234.800 425.600 235.600 426.400 ;
        RECT 238.000 425.600 238.800 426.400 ;
        RECT 241.200 425.600 242.000 426.400 ;
        RECT 244.400 425.600 245.200 426.400 ;
        RECT 234.900 414.400 235.500 425.600 ;
        RECT 236.400 423.600 237.200 424.400 ;
        RECT 236.500 416.400 237.100 423.600 ;
        RECT 236.400 415.600 237.200 416.400 ;
        RECT 238.100 414.400 238.700 425.600 ;
        RECT 244.500 422.400 245.100 425.600 ;
        RECT 244.400 421.600 245.200 422.400 ;
        RECT 234.800 413.600 235.600 414.400 ;
        RECT 236.400 413.600 237.200 414.400 ;
        RECT 238.000 413.600 238.800 414.400 ;
        RECT 231.600 409.600 232.400 410.400 ;
        RECT 209.200 389.600 210.000 390.400 ;
        RECT 210.800 389.600 211.600 390.400 ;
        RECT 210.900 388.400 211.500 389.600 ;
        RECT 210.800 387.600 211.600 388.400 ;
        RECT 215.600 384.200 216.400 395.800 ;
        RECT 226.800 393.600 227.600 394.400 ;
        RECT 218.800 386.200 219.600 391.800 ;
        RECT 220.400 391.600 221.200 392.400 ;
        RECT 222.200 391.800 223.000 392.600 ;
        RECT 228.400 391.800 229.200 392.600 ;
        RECT 231.700 392.300 232.300 409.600 ;
        RECT 233.200 393.600 234.000 394.400 ;
        RECT 220.500 388.400 221.100 391.600 ;
        RECT 220.400 387.600 221.200 388.400 ;
        RECT 222.200 387.000 222.800 391.800 ;
        RECT 223.400 389.800 224.200 390.600 ;
        RECT 223.600 388.400 224.200 389.800 ;
        RECT 228.600 388.400 229.200 391.800 ;
        RECT 230.100 391.700 232.300 392.300 ;
        RECT 230.100 388.400 230.700 391.700 ;
        RECT 233.300 390.400 233.900 393.600 ;
        RECT 234.900 392.400 235.500 413.600 ;
        RECT 234.800 391.600 235.600 392.400 ;
        RECT 231.600 389.600 232.400 390.400 ;
        RECT 233.200 389.600 234.000 390.400 ;
        RECT 223.600 387.800 229.200 388.400 ;
        RECT 223.600 387.000 224.400 387.200 ;
        RECT 227.000 387.000 227.800 387.200 ;
        RECT 228.600 387.000 229.200 387.800 ;
        RECT 230.000 387.600 230.800 388.400 ;
        RECT 222.200 386.400 227.800 387.000 ;
        RECT 222.200 386.200 223.000 386.400 ;
        RECT 228.400 386.200 229.200 387.000 ;
        RECT 217.200 383.600 218.000 384.400 ;
        RECT 206.000 375.600 206.800 376.400 ;
        RECT 204.400 371.600 205.200 372.400 ;
        RECT 204.500 370.400 205.100 371.600 ;
        RECT 204.400 369.600 205.200 370.400 ;
        RECT 186.800 345.600 187.600 346.400 ;
        RECT 186.900 340.300 187.500 345.600 ;
        RECT 188.400 344.200 189.200 355.800 ;
        RECT 190.000 344.200 190.800 357.800 ;
        RECT 191.600 344.200 192.400 357.800 ;
        RECT 193.200 344.200 194.000 357.800 ;
        RECT 204.400 355.600 205.200 356.400 ;
        RECT 188.400 341.600 189.200 342.400 ;
        RECT 185.300 339.700 187.500 340.300 ;
        RECT 167.600 337.600 168.400 338.400 ;
        RECT 167.700 336.400 168.300 337.600 ;
        RECT 167.600 335.600 168.400 336.400 ;
        RECT 151.600 331.600 152.400 332.400 ;
        RECT 159.600 331.600 160.400 332.400 ;
        RECT 162.800 331.600 163.600 332.400 ;
        RECT 166.000 331.600 166.800 332.400 ;
        RECT 167.700 330.400 168.300 335.600 ;
        RECT 143.400 329.400 144.200 330.200 ;
        RECT 150.000 329.400 150.800 330.200 ;
        RECT 159.600 329.600 160.400 330.400 ;
        RECT 167.600 329.600 168.400 330.400 ;
        RECT 154.800 327.600 155.600 328.400 ;
        RECT 145.200 323.600 146.000 324.400 ;
        RECT 145.300 318.400 145.900 323.600 ;
        RECT 154.900 318.400 155.500 327.600 ;
        RECT 159.700 318.400 160.300 329.600 ;
        RECT 162.800 323.600 163.600 324.400 ;
        RECT 178.800 324.200 179.600 337.800 ;
        RECT 180.400 324.200 181.200 337.800 ;
        RECT 182.000 324.200 182.800 337.800 ;
        RECT 183.600 326.200 184.400 337.800 ;
        RECT 185.300 336.400 185.900 339.700 ;
        RECT 185.200 335.600 186.000 336.400 ;
        RECT 186.800 326.200 187.600 337.800 ;
        RECT 188.500 334.400 189.100 341.600 ;
        RECT 204.500 338.400 205.100 355.600 ;
        RECT 206.100 348.400 206.700 375.600 ;
        RECT 214.000 373.600 214.800 374.400 ;
        RECT 212.400 363.600 213.200 364.400 ;
        RECT 212.500 360.400 213.100 363.600 ;
        RECT 212.400 359.600 213.200 360.400 ;
        RECT 207.600 351.800 208.400 352.600 ;
        RECT 213.800 351.800 214.600 352.600 ;
        RECT 217.300 352.400 217.900 383.600 ;
        RECT 228.400 381.600 229.200 382.400 ;
        RECT 220.400 373.600 221.200 374.400 ;
        RECT 220.400 371.600 221.200 372.400 ;
        RECT 222.000 371.600 222.800 372.400 ;
        RECT 226.800 371.600 227.600 372.400 ;
        RECT 220.500 366.400 221.100 371.600 ;
        RECT 220.400 365.600 221.200 366.400 ;
        RECT 207.600 348.400 208.200 351.800 ;
        RECT 212.600 349.800 213.400 350.600 ;
        RECT 212.600 348.400 213.200 349.800 ;
        RECT 206.000 347.600 206.800 348.400 ;
        RECT 207.600 347.800 213.200 348.400 ;
        RECT 207.600 347.000 208.200 347.800 ;
        RECT 209.000 347.000 209.800 347.200 ;
        RECT 212.400 347.000 213.200 347.200 ;
        RECT 214.000 347.000 214.600 351.800 ;
        RECT 217.200 351.600 218.000 352.400 ;
        RECT 220.500 350.400 221.100 365.600 ;
        RECT 222.100 352.400 222.700 371.600 ;
        RECT 222.000 351.600 222.800 352.400 ;
        RECT 220.400 350.300 221.200 350.400 ;
        RECT 223.600 350.300 224.400 350.400 ;
        RECT 220.400 349.700 224.400 350.300 ;
        RECT 220.400 349.600 221.200 349.700 ;
        RECT 223.600 349.600 224.400 349.700 ;
        RECT 207.600 346.200 208.400 347.000 ;
        RECT 209.000 346.400 214.600 347.000 ;
        RECT 223.700 346.400 224.300 349.600 ;
        RECT 225.200 347.600 226.000 348.400 ;
        RECT 213.800 346.200 214.600 346.400 ;
        RECT 220.400 345.600 221.200 346.400 ;
        RECT 223.600 346.300 224.400 346.400 ;
        RECT 223.600 345.700 225.900 346.300 ;
        RECT 223.600 345.600 224.400 345.700 ;
        RECT 209.200 343.600 210.000 344.400 ;
        RECT 206.000 339.600 206.800 340.400 ;
        RECT 188.400 333.600 189.200 334.400 ;
        RECT 190.000 326.200 190.800 337.800 ;
        RECT 191.600 324.200 192.400 337.800 ;
        RECT 193.200 324.200 194.000 337.800 ;
        RECT 204.400 337.600 205.200 338.400 ;
        RECT 198.000 331.600 198.800 332.400 ;
        RECT 198.100 330.400 198.700 331.600 ;
        RECT 198.000 329.600 198.800 330.400 ;
        RECT 145.200 317.600 146.000 318.400 ;
        RECT 154.800 317.600 155.600 318.400 ;
        RECT 156.400 317.600 157.200 318.400 ;
        RECT 159.600 317.600 160.400 318.400 ;
        RECT 146.800 311.600 147.600 312.400 ;
        RECT 153.200 311.600 154.000 312.400 ;
        RECT 135.600 309.600 136.400 310.400 ;
        RECT 140.400 309.600 141.200 310.400 ;
        RECT 150.000 309.600 150.800 310.400 ;
        RECT 135.700 306.400 136.300 309.600 ;
        RECT 156.500 308.400 157.100 317.600 ;
        RECT 161.200 309.600 162.000 310.400 ;
        RECT 151.600 307.600 152.400 308.400 ;
        RECT 154.800 307.600 155.600 308.400 ;
        RECT 156.400 307.600 157.200 308.400 ;
        RECT 135.600 305.600 136.400 306.400 ;
        RECT 146.800 303.600 147.600 304.400 ;
        RECT 127.600 301.600 128.400 302.400 ;
        RECT 134.000 301.600 134.800 302.400 ;
        RECT 119.600 285.600 120.400 286.400 ;
        RECT 119.700 278.400 120.300 285.600 ;
        RECT 126.000 284.200 126.800 297.800 ;
        RECT 127.600 284.200 128.400 297.800 ;
        RECT 129.200 286.200 130.000 297.800 ;
        RECT 130.800 293.600 131.600 294.400 ;
        RECT 132.400 286.200 133.200 297.800 ;
        RECT 134.100 296.400 134.700 301.600 ;
        RECT 146.900 298.400 147.500 303.600 ;
        RECT 134.000 295.600 134.800 296.400 ;
        RECT 134.100 286.400 134.700 295.600 ;
        RECT 134.000 285.600 134.800 286.400 ;
        RECT 135.600 286.200 136.400 297.800 ;
        RECT 132.400 283.600 133.200 284.400 ;
        RECT 137.200 284.200 138.000 297.800 ;
        RECT 138.800 284.200 139.600 297.800 ;
        RECT 140.400 284.200 141.200 297.800 ;
        RECT 146.800 297.600 147.600 298.400 ;
        RECT 142.000 295.600 142.800 296.400 ;
        RECT 142.100 292.400 142.700 295.600 ;
        RECT 142.000 291.600 142.800 292.400 ;
        RECT 151.700 290.400 152.300 307.600 ;
        RECT 153.200 293.600 154.000 294.400 ;
        RECT 151.600 289.600 152.400 290.400 ;
        RECT 153.200 290.300 154.000 290.400 ;
        RECT 154.900 290.300 155.500 307.600 ;
        RECT 158.000 305.600 158.800 306.400 ;
        RECT 153.200 289.700 155.500 290.300 ;
        RECT 153.200 289.600 154.000 289.700 ;
        RECT 150.000 287.600 150.800 288.400 ;
        RECT 153.200 285.600 154.000 286.400 ;
        RECT 132.500 278.400 133.100 283.600 ;
        RECT 119.600 277.600 120.400 278.400 ;
        RECT 132.400 277.600 133.200 278.400 ;
        RECT 137.200 273.600 138.000 274.400 ;
        RECT 137.300 272.400 137.900 273.600 ;
        RECT 137.200 271.600 138.000 272.400 ;
        RECT 130.800 267.600 131.600 268.400 ;
        RECT 118.000 263.600 118.800 264.400 ;
        RECT 129.200 263.600 130.000 264.400 ;
        RECT 106.800 261.600 107.600 262.400 ;
        RECT 98.800 259.600 99.600 260.400 ;
        RECT 103.600 259.600 104.400 260.400 ;
        RECT 124.400 259.600 125.200 260.400 ;
        RECT 89.200 257.600 90.000 258.400 ;
        RECT 97.200 257.600 98.000 258.400 ;
        RECT 82.800 253.600 83.600 254.400 ;
        RECT 76.400 251.600 77.200 252.400 ;
        RECT 78.000 251.600 78.800 252.400 ;
        RECT 76.400 245.600 77.200 246.400 ;
        RECT 65.200 231.600 66.000 232.400 ;
        RECT 65.300 230.400 65.900 231.600 ;
        RECT 76.500 230.400 77.100 245.600 ;
        RECT 78.100 232.400 78.700 251.600 ;
        RECT 82.900 238.400 83.500 253.600 ;
        RECT 84.400 243.600 85.200 244.400 ;
        RECT 98.800 244.200 99.600 257.800 ;
        RECT 100.400 244.200 101.200 257.800 ;
        RECT 102.000 244.200 102.800 257.800 ;
        RECT 103.600 246.200 104.400 257.800 ;
        RECT 105.200 255.600 106.000 256.400 ;
        RECT 106.800 246.200 107.600 257.800 ;
        RECT 108.400 253.600 109.200 254.400 ;
        RECT 110.000 246.200 110.800 257.800 ;
        RECT 111.600 244.200 112.400 257.800 ;
        RECT 113.200 244.200 114.000 257.800 ;
        RECT 119.600 255.600 120.400 256.400 ;
        RECT 118.000 251.600 118.800 252.400 ;
        RECT 82.800 237.600 83.600 238.400 ;
        RECT 78.000 231.600 78.800 232.400 ;
        RECT 78.100 230.400 78.700 231.600 ;
        RECT 84.500 230.400 85.100 243.600 ;
        RECT 52.400 229.600 53.200 230.400 ;
        RECT 58.800 229.600 59.600 230.400 ;
        RECT 63.600 229.600 64.400 230.400 ;
        RECT 65.200 229.600 66.000 230.400 ;
        RECT 70.000 229.600 70.800 230.400 ;
        RECT 76.400 229.600 77.200 230.400 ;
        RECT 78.000 229.600 78.800 230.400 ;
        RECT 79.600 229.600 80.400 230.400 ;
        RECT 84.400 229.600 85.200 230.400 ;
        RECT 90.800 229.600 91.600 230.400 ;
        RECT 52.500 224.400 53.100 229.600 ;
        RECT 57.200 227.600 58.000 228.400 ;
        RECT 62.000 225.600 62.800 226.400 ;
        RECT 52.400 223.600 53.200 224.400 ;
        RECT 62.100 218.400 62.700 225.600 ;
        RECT 62.000 217.600 62.800 218.400 ;
        RECT 49.200 215.600 50.000 216.400 ;
        RECT 58.800 215.600 59.600 216.400 ;
        RECT 58.900 214.400 59.500 215.600 ;
        RECT 58.800 213.600 59.600 214.400 ;
        RECT 42.800 203.600 43.600 204.400 ;
        RECT 47.600 203.600 48.400 204.400 ;
        RECT 62.000 203.600 62.800 204.400 ;
        RECT 47.700 186.400 48.300 203.600 ;
        RECT 49.200 195.600 50.000 196.400 ;
        RECT 57.200 193.600 58.000 194.400 ;
        RECT 50.800 191.600 51.600 192.400 ;
        RECT 50.900 190.400 51.500 191.600 ;
        RECT 50.800 189.600 51.600 190.400 ;
        RECT 55.600 189.600 56.400 190.400 ;
        RECT 55.700 188.400 56.300 189.600 ;
        RECT 55.600 187.600 56.400 188.400 ;
        RECT 47.600 185.600 48.400 186.400 ;
        RECT 41.200 175.600 42.000 176.400 ;
        RECT 41.200 171.800 42.000 172.600 ;
        RECT 41.300 164.300 41.900 171.800 ;
        RECT 49.200 166.200 50.000 177.800 ;
        RECT 52.400 177.600 53.200 178.400 ;
        RECT 39.700 163.700 41.900 164.300 ;
        RECT 39.700 158.400 40.300 163.700 ;
        RECT 41.200 161.600 42.000 162.400 ;
        RECT 39.600 157.600 40.400 158.400 ;
        RECT 41.300 152.400 41.900 161.600 ;
        RECT 44.400 155.600 45.200 156.400 ;
        RECT 41.200 151.600 42.000 152.400 ;
        RECT 41.300 150.400 41.900 151.600 ;
        RECT 39.600 149.600 40.400 150.400 ;
        RECT 41.200 149.600 42.000 150.400 ;
        RECT 39.700 148.400 40.300 149.600 ;
        RECT 39.600 147.600 40.400 148.400 ;
        RECT 41.200 147.600 42.000 148.400 ;
        RECT 42.800 147.600 43.600 148.400 ;
        RECT 41.300 146.400 41.900 147.600 ;
        RECT 41.200 145.600 42.000 146.400 ;
        RECT 38.000 135.600 38.800 136.400 ;
        RECT 38.100 132.400 38.700 135.600 ;
        RECT 38.000 131.600 38.800 132.400 ;
        RECT 39.600 131.600 40.400 132.400 ;
        RECT 38.000 127.600 38.800 128.400 ;
        RECT 30.000 117.600 30.800 118.400 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 36.500 110.400 37.100 111.600 ;
        RECT 15.600 109.600 16.400 110.400 ;
        RECT 25.200 109.600 26.000 110.400 ;
        RECT 26.800 109.600 27.600 110.400 ;
        RECT 28.400 109.600 29.200 110.400 ;
        RECT 33.200 109.600 34.000 110.400 ;
        RECT 34.800 109.600 35.600 110.400 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 7.700 101.700 9.900 102.300 ;
        RECT 6.000 93.600 6.800 94.400 ;
        RECT 4.400 64.200 5.200 75.800 ;
        RECT 6.100 68.400 6.700 93.600 ;
        RECT 6.000 67.600 6.800 68.400 ;
        RECT 6.000 65.600 6.800 66.400 ;
        RECT 4.400 46.200 5.200 57.800 ;
        RECT 6.100 56.400 6.700 65.600 ;
        RECT 6.000 55.600 6.800 56.400 ;
        RECT 7.700 30.400 8.300 101.700 ;
        RECT 9.200 93.600 10.000 94.400 ;
        RECT 9.300 92.400 9.900 93.600 ;
        RECT 15.700 92.400 16.300 109.600 ;
        RECT 25.300 108.400 25.900 109.600 ;
        RECT 25.200 107.600 26.000 108.400 ;
        RECT 18.800 103.600 19.600 104.400 ;
        RECT 22.000 103.600 22.800 104.400 ;
        RECT 9.200 91.600 10.000 92.400 ;
        RECT 14.000 91.600 14.800 92.400 ;
        RECT 15.600 91.600 16.400 92.400 ;
        RECT 17.200 91.600 18.000 92.400 ;
        RECT 14.100 90.400 14.700 91.600 ;
        RECT 14.000 89.600 14.800 90.400 ;
        RECT 17.200 90.300 18.000 90.400 ;
        RECT 18.900 90.300 19.500 103.600 ;
        RECT 22.100 96.400 22.700 103.600 ;
        RECT 31.600 99.600 32.400 100.400 ;
        RECT 26.800 97.600 27.600 98.400 ;
        RECT 22.000 95.600 22.800 96.400 ;
        RECT 22.100 94.400 22.700 95.600 ;
        RECT 22.000 93.600 22.800 94.400 ;
        RECT 23.600 93.600 24.400 94.400 ;
        RECT 20.400 91.600 21.200 92.400 ;
        RECT 17.200 89.700 19.500 90.300 ;
        RECT 17.200 89.600 18.000 89.700 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 9.300 66.400 9.900 69.600 ;
        RECT 9.200 65.600 10.000 66.400 ;
        RECT 14.000 64.200 14.800 75.800 ;
        RECT 18.800 73.600 19.600 74.400 ;
        RECT 18.900 72.400 19.500 73.600 ;
        RECT 18.800 71.600 19.600 72.400 ;
        RECT 20.500 70.400 21.100 91.600 ;
        RECT 20.400 69.600 21.200 70.400 ;
        RECT 20.400 68.300 21.200 68.400 ;
        RECT 22.100 68.300 22.700 93.600 ;
        RECT 26.900 92.400 27.500 97.600 ;
        RECT 30.000 93.600 30.800 94.400 ;
        RECT 31.700 92.400 32.300 99.600 ;
        RECT 26.800 91.600 27.600 92.400 ;
        RECT 31.600 91.600 32.400 92.400 ;
        RECT 23.600 89.600 24.400 90.400 ;
        RECT 23.700 88.400 24.300 89.600 ;
        RECT 23.600 87.600 24.400 88.400 ;
        RECT 26.800 85.600 27.600 86.400 ;
        RECT 25.200 71.600 26.000 72.400 ;
        RECT 33.300 70.400 33.900 109.600 ;
        RECT 34.900 106.400 35.500 109.600 ;
        RECT 34.800 105.600 35.600 106.400 ;
        RECT 34.900 98.400 35.500 105.600 ;
        RECT 38.100 98.400 38.700 127.600 ;
        RECT 42.800 109.600 43.600 110.400 ;
        RECT 42.900 108.400 43.500 109.600 ;
        RECT 41.200 107.600 42.000 108.400 ;
        RECT 42.800 107.600 43.600 108.400 ;
        RECT 34.800 97.600 35.600 98.400 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 36.400 95.600 37.200 96.400 ;
        RECT 36.500 94.400 37.100 95.600 ;
        RECT 36.400 93.600 37.200 94.400 ;
        RECT 41.300 92.400 41.900 107.600 ;
        RECT 42.900 102.400 43.500 107.600 ;
        RECT 42.800 101.600 43.600 102.400 ;
        RECT 42.800 97.600 43.600 98.400 ;
        RECT 42.900 94.400 43.500 97.600 ;
        RECT 42.800 93.600 43.600 94.400 ;
        RECT 38.000 91.600 38.800 92.400 ;
        RECT 41.200 91.600 42.000 92.400 ;
        RECT 34.800 90.300 35.600 90.400 ;
        RECT 34.800 89.700 37.100 90.300 ;
        RECT 34.800 89.600 35.600 89.700 ;
        RECT 34.800 71.600 35.600 72.400 ;
        RECT 34.900 70.400 35.500 71.600 ;
        RECT 30.000 69.600 30.800 70.400 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 34.800 69.600 35.600 70.400 ;
        RECT 20.400 67.700 22.700 68.300 ;
        RECT 20.400 67.600 21.200 67.700 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 36.500 68.300 37.100 89.700 ;
        RECT 41.200 89.600 42.000 90.400 ;
        RECT 39.600 87.600 40.400 88.400 ;
        RECT 38.000 83.600 38.800 84.400 ;
        RECT 38.100 72.400 38.700 83.600 ;
        RECT 38.000 71.600 38.800 72.400 ;
        RECT 38.000 69.600 38.800 70.400 ;
        RECT 34.900 67.700 37.100 68.300 ;
        RECT 20.500 64.400 21.100 67.600 ;
        RECT 26.800 65.600 27.600 66.400 ;
        RECT 20.400 63.600 21.200 64.400 ;
        RECT 9.200 53.600 10.000 54.400 ;
        RECT 9.300 52.400 9.900 53.600 ;
        RECT 9.200 51.600 10.000 52.400 ;
        RECT 12.400 51.600 13.200 52.400 ;
        RECT 12.500 44.400 13.100 51.600 ;
        RECT 14.000 46.200 14.800 57.800 ;
        RECT 18.800 57.600 19.600 58.400 ;
        RECT 18.900 50.400 19.500 57.600 ;
        RECT 20.500 54.400 21.100 63.600 ;
        RECT 22.000 55.600 22.800 56.400 ;
        RECT 30.000 55.600 30.800 56.400 ;
        RECT 20.400 53.600 21.200 54.400 ;
        RECT 22.100 52.400 22.700 55.600 ;
        RECT 26.800 53.600 27.600 54.400 ;
        RECT 30.100 52.400 30.700 55.600 ;
        RECT 31.700 54.400 32.300 67.600 ;
        RECT 34.900 58.400 35.500 67.700 ;
        RECT 39.700 58.400 40.300 87.600 ;
        RECT 41.300 84.400 41.900 89.600 ;
        RECT 41.200 83.600 42.000 84.400 ;
        RECT 42.800 71.600 43.600 72.400 ;
        RECT 42.800 70.300 43.600 70.400 ;
        RECT 44.500 70.300 45.100 155.600 ;
        RECT 52.500 152.400 53.100 177.600 ;
        RECT 55.700 170.400 56.300 187.600 ;
        RECT 57.300 178.400 57.900 193.600 ;
        RECT 60.400 187.600 61.200 188.400 ;
        RECT 62.100 186.400 62.700 203.600 ;
        RECT 63.700 198.400 64.300 229.600 ;
        RECT 70.100 228.400 70.700 229.600 ;
        RECT 70.000 227.600 70.800 228.400 ;
        RECT 74.800 227.600 75.600 228.400 ;
        RECT 66.800 225.600 67.600 226.400 ;
        RECT 70.000 223.600 70.800 224.400 ;
        RECT 73.200 223.600 74.000 224.400 ;
        RECT 70.100 212.400 70.700 223.600 ;
        RECT 73.300 220.400 73.900 223.600 ;
        RECT 73.200 219.600 74.000 220.400 ;
        RECT 81.200 219.600 82.000 220.400 ;
        RECT 70.000 211.600 70.800 212.400 ;
        RECT 68.400 203.600 69.200 204.400 ;
        RECT 71.600 204.200 72.400 217.800 ;
        RECT 73.200 204.200 74.000 217.800 ;
        RECT 74.800 204.200 75.600 217.800 ;
        RECT 76.400 206.200 77.200 217.800 ;
        RECT 78.000 217.600 78.800 218.400 ;
        RECT 78.100 216.400 78.700 217.600 ;
        RECT 78.000 215.600 78.800 216.400 ;
        RECT 79.600 206.200 80.400 217.800 ;
        RECT 81.300 214.400 81.900 219.600 ;
        RECT 81.200 213.600 82.000 214.400 ;
        RECT 82.800 206.200 83.600 217.800 ;
        RECT 84.400 204.200 85.200 217.800 ;
        RECT 86.000 204.200 86.800 217.800 ;
        RECT 87.600 217.600 88.400 218.400 ;
        RECT 63.600 197.600 64.400 198.400 ;
        RECT 68.500 194.400 69.100 203.600 ;
        RECT 68.400 193.600 69.200 194.400 ;
        RECT 79.600 193.600 80.400 194.400 ;
        RECT 79.700 192.400 80.300 193.600 ;
        RECT 71.600 191.600 72.400 192.400 ;
        RECT 73.200 191.600 74.000 192.400 ;
        RECT 76.400 191.600 77.200 192.400 ;
        RECT 79.600 191.600 80.400 192.400 ;
        RECT 82.800 191.600 83.600 192.400 ;
        RECT 73.300 190.400 73.900 191.600 ;
        RECT 76.500 190.400 77.100 191.600 ;
        RECT 82.900 190.400 83.500 191.600 ;
        RECT 63.600 189.600 64.400 190.400 ;
        RECT 70.000 189.600 70.800 190.400 ;
        RECT 73.200 189.600 74.000 190.400 ;
        RECT 76.400 189.600 77.200 190.400 ;
        RECT 82.800 189.600 83.600 190.400 ;
        RECT 58.800 185.600 59.600 186.400 ;
        RECT 62.000 185.600 62.800 186.400 ;
        RECT 58.900 182.400 59.500 185.600 ;
        RECT 63.700 184.400 64.300 189.600 ;
        RECT 65.200 187.600 66.000 188.400 ;
        RECT 78.000 187.600 78.800 188.400 ;
        RECT 84.400 187.600 85.200 188.400 ;
        RECT 63.600 183.600 64.400 184.400 ;
        RECT 58.800 182.300 59.600 182.400 ;
        RECT 58.800 181.700 61.100 182.300 ;
        RECT 58.800 181.600 59.600 181.700 ;
        RECT 57.200 177.600 58.000 178.400 ;
        RECT 60.500 174.400 61.100 181.700 ;
        RECT 63.700 176.400 64.300 183.600 ;
        RECT 63.600 175.600 64.400 176.400 ;
        RECT 65.300 174.400 65.900 187.600 ;
        RECT 70.000 185.600 70.800 186.400 ;
        RECT 86.000 186.200 86.800 191.800 ;
        RECT 87.700 188.400 88.300 217.600 ;
        RECT 90.900 212.400 91.500 229.600 ;
        RECT 95.600 224.200 96.400 237.800 ;
        RECT 97.200 224.200 98.000 237.800 ;
        RECT 98.800 224.200 99.600 235.800 ;
        RECT 100.400 231.600 101.200 232.400 ;
        RECT 100.500 228.400 101.100 231.600 ;
        RECT 100.400 227.600 101.200 228.400 ;
        RECT 102.000 224.200 102.800 235.800 ;
        RECT 103.600 225.600 104.400 226.400 ;
        RECT 103.700 224.400 104.300 225.600 ;
        RECT 103.600 223.600 104.400 224.400 ;
        RECT 105.200 224.200 106.000 235.800 ;
        RECT 106.800 224.200 107.600 237.800 ;
        RECT 108.400 224.200 109.200 237.800 ;
        RECT 110.000 224.200 110.800 237.800 ;
        RECT 118.100 230.400 118.700 251.600 ;
        RECT 119.700 238.400 120.300 255.600 ;
        RECT 119.600 237.600 120.400 238.400 ;
        RECT 111.600 229.600 112.400 230.400 ;
        RECT 118.000 229.600 118.800 230.400 ;
        RECT 119.600 225.600 120.400 226.400 ;
        RECT 119.700 218.400 120.300 225.600 ;
        RECT 119.600 217.600 120.400 218.400 ;
        RECT 108.400 215.600 109.200 216.400 ;
        RECT 108.500 214.400 109.100 215.600 ;
        RECT 124.500 214.400 125.100 259.600 ;
        RECT 129.300 258.400 129.900 263.600 ;
        RECT 130.900 260.400 131.500 267.600 ;
        RECT 134.000 265.600 134.800 266.400 ;
        RECT 130.800 259.600 131.600 260.400 ;
        RECT 129.200 257.600 130.000 258.400 ;
        RECT 127.600 229.600 128.400 230.400 ;
        RECT 127.700 228.400 128.300 229.600 ;
        RECT 127.600 227.600 128.400 228.400 ;
        RECT 134.100 226.400 134.700 265.600 ;
        RECT 146.800 264.200 147.600 277.800 ;
        RECT 148.400 264.200 149.200 277.800 ;
        RECT 150.000 264.200 150.800 277.800 ;
        RECT 151.600 264.200 152.400 275.800 ;
        RECT 153.300 266.400 153.900 285.600 ;
        RECT 154.900 280.400 155.500 289.700 ;
        RECT 156.400 287.600 157.200 288.400 ;
        RECT 154.800 279.600 155.600 280.400 ;
        RECT 156.500 276.400 157.100 287.600 ;
        RECT 158.100 278.400 158.700 305.600 ;
        RECT 161.300 292.400 161.900 309.600 ;
        RECT 162.900 308.400 163.500 323.600 ;
        RECT 169.200 315.600 170.000 316.400 ;
        RECT 166.000 309.600 166.800 310.400 ;
        RECT 177.200 309.600 178.000 310.400 ;
        RECT 162.800 307.600 163.600 308.400 ;
        RECT 177.300 306.400 177.900 309.600 ;
        RECT 162.800 305.600 163.600 306.400 ;
        RECT 170.800 305.600 171.600 306.400 ;
        RECT 177.200 305.600 178.000 306.400 ;
        RECT 162.900 304.400 163.500 305.600 ;
        RECT 162.800 303.600 163.600 304.400 ;
        RECT 162.900 302.300 163.500 303.600 ;
        RECT 162.900 301.700 165.100 302.300 ;
        RECT 162.800 299.600 163.600 300.400 ;
        RECT 162.900 294.400 163.500 299.600 ;
        RECT 162.800 293.600 163.600 294.400 ;
        RECT 161.200 291.600 162.000 292.400 ;
        RECT 161.300 284.400 161.900 291.600 ;
        RECT 161.200 283.600 162.000 284.400 ;
        RECT 158.000 277.600 158.800 278.400 ;
        RECT 153.200 265.600 154.000 266.400 ;
        RECT 154.800 264.200 155.600 275.800 ;
        RECT 156.400 275.600 157.200 276.400 ;
        RECT 156.400 267.600 157.200 268.400 ;
        RECT 158.000 264.200 158.800 275.800 ;
        RECT 159.600 264.200 160.400 277.800 ;
        RECT 161.200 264.200 162.000 277.800 ;
        RECT 164.500 270.400 165.100 301.700 ;
        RECT 170.900 296.400 171.500 305.600 ;
        RECT 177.200 303.600 178.000 304.400 ;
        RECT 178.800 304.200 179.600 317.800 ;
        RECT 180.400 304.200 181.200 317.800 ;
        RECT 182.000 304.200 182.800 317.800 ;
        RECT 183.600 304.200 184.400 315.800 ;
        RECT 185.200 305.600 186.000 306.400 ;
        RECT 186.800 304.200 187.600 315.800 ;
        RECT 188.400 307.600 189.200 308.400 ;
        RECT 190.000 304.200 190.800 315.800 ;
        RECT 191.600 304.200 192.400 317.800 ;
        RECT 193.200 304.200 194.000 317.800 ;
        RECT 198.100 310.400 198.700 329.600 ;
        RECT 206.100 312.400 206.700 339.600 ;
        RECT 220.500 334.400 221.100 345.600 ;
        RECT 222.000 339.600 222.800 340.400 ;
        RECT 217.200 333.600 218.000 334.400 ;
        RECT 220.400 333.600 221.200 334.400 ;
        RECT 209.200 331.600 210.000 332.400 ;
        RECT 206.000 311.600 206.800 312.400 ;
        RECT 209.300 310.400 209.900 331.600 ;
        RECT 212.400 329.600 213.200 330.400 ;
        RECT 215.600 329.600 216.400 330.400 ;
        RECT 215.700 328.400 216.300 329.600 ;
        RECT 215.600 327.600 216.400 328.400 ;
        RECT 215.600 325.600 216.400 326.400 ;
        RECT 210.800 315.600 211.600 316.400 ;
        RECT 210.900 314.400 211.500 315.600 ;
        RECT 210.800 313.600 211.600 314.400 ;
        RECT 215.700 310.400 216.300 325.600 ;
        RECT 220.500 318.400 221.100 333.600 ;
        RECT 220.400 317.600 221.200 318.400 ;
        RECT 222.100 310.400 222.700 339.600 ;
        RECT 223.600 335.600 224.400 336.400 ;
        RECT 225.300 332.400 225.900 345.700 ;
        RECT 226.900 340.400 227.500 371.600 ;
        RECT 228.500 358.400 229.100 381.600 ;
        RECT 230.100 376.400 230.700 387.600 ;
        RECT 231.700 384.400 232.300 389.600 ;
        RECT 236.500 384.400 237.100 413.600 ;
        RECT 238.100 412.400 238.700 413.600 ;
        RECT 238.000 411.600 238.800 412.400 ;
        RECT 244.400 411.600 245.200 412.400 ;
        RECT 241.200 409.600 242.000 410.400 ;
        RECT 238.000 391.600 238.800 392.400 ;
        RECT 238.100 390.400 238.700 391.600 ;
        RECT 241.300 390.400 241.900 409.600 ;
        RECT 246.100 398.400 246.700 427.600 ;
        RECT 247.700 414.400 248.300 433.600 ;
        RECT 249.300 418.400 249.900 443.700 ;
        RECT 250.800 424.200 251.600 437.800 ;
        RECT 252.400 424.200 253.200 437.800 ;
        RECT 254.000 424.200 254.800 437.800 ;
        RECT 255.600 424.200 256.400 435.800 ;
        RECT 257.200 425.600 258.000 426.400 ;
        RECT 258.800 424.200 259.600 435.800 ;
        RECT 260.500 430.400 261.100 451.600 ;
        RECT 274.800 444.200 275.600 457.800 ;
        RECT 276.400 444.200 277.200 457.800 ;
        RECT 278.000 446.200 278.800 457.800 ;
        RECT 279.600 453.600 280.400 454.400 ;
        RECT 279.600 451.600 280.400 452.400 ;
        RECT 260.400 429.600 261.200 430.400 ;
        RECT 260.400 427.600 261.200 428.400 ;
        RECT 262.000 424.200 262.800 435.800 ;
        RECT 263.600 424.200 264.400 437.800 ;
        RECT 265.200 424.200 266.000 437.800 ;
        RECT 279.700 434.400 280.300 451.600 ;
        RECT 281.200 446.200 282.000 457.800 ;
        RECT 282.800 455.600 283.600 456.400 ;
        RECT 284.400 446.200 285.200 457.800 ;
        RECT 281.200 443.600 282.000 444.400 ;
        RECT 286.000 444.200 286.800 457.800 ;
        RECT 287.600 444.200 288.400 457.800 ;
        RECT 289.200 444.200 290.000 457.800 ;
        RECT 290.900 452.400 291.500 491.600 ;
        RECT 292.500 478.400 293.100 493.600 ;
        RECT 294.000 491.600 294.800 492.400 ;
        RECT 302.000 491.600 302.800 492.400 ;
        RECT 292.400 477.600 293.200 478.400 ;
        RECT 294.100 466.400 294.700 491.600 ;
        RECT 303.700 478.400 304.300 493.600 ;
        RECT 306.800 484.200 307.600 497.800 ;
        RECT 308.400 484.200 309.200 497.800 ;
        RECT 310.000 486.200 310.800 497.800 ;
        RECT 311.600 493.600 312.400 494.400 ;
        RECT 303.600 477.600 304.400 478.400 ;
        RECT 311.700 470.400 312.300 493.600 ;
        RECT 313.200 486.200 314.000 497.800 ;
        RECT 314.800 495.600 315.600 496.400 ;
        RECT 316.400 486.200 317.200 497.800 ;
        RECT 318.000 484.200 318.800 497.800 ;
        RECT 319.600 484.200 320.400 497.800 ;
        RECT 321.200 484.200 322.000 497.800 ;
        RECT 335.400 495.000 336.200 495.800 ;
        RECT 337.200 495.000 341.400 495.600 ;
        RECT 342.000 495.000 342.800 495.800 ;
        RECT 334.000 493.600 334.800 494.400 ;
        RECT 322.800 491.600 323.600 492.400 ;
        RECT 335.400 490.200 336.000 495.000 ;
        RECT 337.200 494.800 338.000 495.000 ;
        RECT 340.600 494.800 341.400 495.000 ;
        RECT 342.200 494.200 342.800 495.000 ;
        RECT 338.000 493.600 342.800 494.200 ;
        RECT 345.200 493.600 346.000 494.400 ;
        RECT 338.000 493.400 338.800 493.600 ;
        RECT 342.200 490.200 342.800 493.600 ;
        RECT 345.300 492.400 345.900 493.600 ;
        RECT 345.200 491.600 346.000 492.400 ;
        RECT 354.800 491.600 355.600 492.400 ;
        RECT 335.400 489.400 336.200 490.200 ;
        RECT 342.000 489.400 342.800 490.200 ;
        RECT 330.800 483.600 331.600 484.400 ;
        RECT 334.000 483.600 334.800 484.400 ;
        RECT 346.800 483.600 347.600 484.400 ;
        RECT 356.400 484.200 357.200 497.800 ;
        RECT 358.000 484.200 358.800 497.800 ;
        RECT 359.600 484.200 360.400 497.800 ;
        RECT 361.200 486.200 362.000 497.800 ;
        RECT 362.800 495.600 363.600 496.400 ;
        RECT 362.900 492.400 363.500 495.600 ;
        RECT 362.800 491.600 363.600 492.400 ;
        RECT 364.400 486.200 365.200 497.800 ;
        RECT 366.000 493.600 366.800 494.400 ;
        RECT 367.600 486.200 368.400 497.800 ;
        RECT 369.200 484.200 370.000 497.800 ;
        RECT 370.800 484.200 371.600 497.800 ;
        RECT 386.800 495.600 387.600 496.400 ;
        RECT 396.400 484.200 397.200 497.800 ;
        RECT 398.000 484.200 398.800 497.800 ;
        RECT 399.600 484.200 400.400 497.800 ;
        RECT 401.200 486.200 402.000 497.800 ;
        RECT 402.800 495.600 403.600 496.400 ;
        RECT 402.900 492.400 403.500 495.600 ;
        RECT 402.800 491.600 403.600 492.400 ;
        RECT 401.200 483.600 402.000 484.400 ;
        RECT 332.400 481.600 333.200 482.400 ;
        RECT 326.000 473.600 326.800 474.400 ;
        RECT 316.400 471.600 317.200 472.400 ;
        RECT 319.600 471.600 320.400 472.400 ;
        RECT 326.100 470.400 326.700 473.600 ;
        RECT 330.800 471.600 331.600 472.400 ;
        RECT 298.800 469.600 299.600 470.400 ;
        RECT 300.400 469.600 301.200 470.400 ;
        RECT 310.000 469.600 310.800 470.400 ;
        RECT 311.600 469.600 312.400 470.400 ;
        RECT 316.400 469.600 317.200 470.400 ;
        RECT 326.000 469.600 326.800 470.400 ;
        RECT 327.600 469.600 328.400 470.400 ;
        RECT 298.900 466.400 299.500 469.600 ;
        RECT 294.000 465.600 294.800 466.400 ;
        RECT 295.600 465.600 296.400 466.400 ;
        RECT 298.800 465.600 299.600 466.400 ;
        RECT 292.400 463.600 293.200 464.400 ;
        RECT 292.500 456.400 293.100 463.600 ;
        RECT 292.400 455.600 293.200 456.400 ;
        RECT 290.800 451.600 291.600 452.400 ;
        RECT 281.300 438.400 281.900 443.600 ;
        RECT 281.200 437.600 282.000 438.400 ;
        RECT 279.600 433.600 280.400 434.400 ;
        RECT 270.000 429.600 270.800 430.400 ;
        RECT 249.200 417.600 250.000 418.400 ;
        RECT 257.200 415.600 258.000 416.400 ;
        RECT 247.600 413.600 248.400 414.400 ;
        RECT 257.300 412.400 257.900 415.600 ;
        RECT 258.800 413.600 259.600 414.400 ;
        RECT 257.200 411.600 258.000 412.400 ;
        RECT 247.600 409.600 248.400 410.400 ;
        RECT 252.400 409.600 253.200 410.400 ;
        RECT 268.400 409.600 269.200 410.400 ;
        RECT 246.000 397.600 246.800 398.400 ;
        RECT 242.800 393.600 243.600 394.400 ;
        RECT 250.800 393.600 251.600 394.400 ;
        RECT 242.900 390.400 243.500 393.600 ;
        RECT 250.900 390.400 251.500 393.600 ;
        RECT 238.000 389.600 238.800 390.400 ;
        RECT 241.200 389.600 242.000 390.400 ;
        RECT 242.800 389.600 243.600 390.400 ;
        RECT 247.600 389.600 248.400 390.400 ;
        RECT 250.800 389.600 251.600 390.400 ;
        RECT 239.600 387.600 240.400 388.400 ;
        RECT 231.600 383.600 232.400 384.400 ;
        RECT 236.400 383.600 237.200 384.400 ;
        RECT 241.300 382.400 241.900 389.600 ;
        RECT 247.700 388.400 248.300 389.600 ;
        RECT 247.600 387.600 248.400 388.400 ;
        RECT 241.200 381.600 242.000 382.400 ;
        RECT 250.900 380.400 251.500 389.600 ;
        RECT 252.500 386.400 253.100 409.600 ;
        RECT 268.500 406.400 269.100 409.600 ;
        RECT 254.000 405.600 254.800 406.400 ;
        RECT 268.400 406.300 269.200 406.400 ;
        RECT 270.100 406.300 270.700 429.600 ;
        RECT 279.700 420.400 280.300 433.600 ;
        RECT 282.800 427.600 283.600 428.400 ;
        RECT 281.200 425.600 282.000 426.400 ;
        RECT 281.300 420.400 281.900 425.600 ;
        RECT 286.000 423.600 286.800 424.400 ;
        RECT 286.100 420.400 286.700 423.600 ;
        RECT 279.600 419.600 280.400 420.400 ;
        RECT 281.200 419.600 282.000 420.400 ;
        RECT 286.000 419.600 286.800 420.400 ;
        RECT 268.400 405.700 270.700 406.300 ;
        RECT 268.400 405.600 269.200 405.700 ;
        RECT 254.100 398.400 254.700 405.600 ;
        RECT 273.200 404.200 274.000 417.800 ;
        RECT 274.800 404.200 275.600 417.800 ;
        RECT 276.400 406.200 277.200 417.800 ;
        RECT 278.000 415.600 278.800 416.400 ;
        RECT 278.100 414.400 278.700 415.600 ;
        RECT 278.000 413.600 278.800 414.400 ;
        RECT 279.600 406.200 280.400 417.800 ;
        RECT 281.300 416.400 281.900 419.600 ;
        RECT 281.200 415.600 282.000 416.400 ;
        RECT 282.800 406.200 283.600 417.800 ;
        RECT 284.400 404.200 285.200 417.800 ;
        RECT 286.000 404.200 286.800 417.800 ;
        RECT 287.600 404.200 288.400 417.800 ;
        RECT 290.900 402.400 291.500 451.600 ;
        RECT 295.700 430.400 296.300 465.600 ;
        RECT 300.500 456.400 301.100 469.600 ;
        RECT 310.100 468.400 310.700 469.600 ;
        RECT 305.200 467.600 306.000 468.400 ;
        RECT 310.000 467.600 310.800 468.400 ;
        RECT 305.300 456.400 305.900 467.600 ;
        RECT 306.800 465.600 307.600 466.400 ;
        RECT 310.000 465.600 310.800 466.400 ;
        RECT 314.800 465.600 315.600 466.400 ;
        RECT 300.400 455.600 301.200 456.400 ;
        RECT 305.200 455.600 306.000 456.400 ;
        RECT 300.400 453.600 301.200 454.400 ;
        RECT 300.400 449.600 301.200 450.400 ;
        RECT 298.800 443.600 299.600 444.400 ;
        RECT 298.900 432.400 299.500 443.600 ;
        RECT 300.500 438.400 301.100 449.600 ;
        RECT 306.900 446.400 307.500 465.600 ;
        RECT 308.400 455.600 309.200 456.400 ;
        RECT 308.400 453.600 309.200 454.400 ;
        RECT 306.800 445.600 307.600 446.400 ;
        RECT 308.500 438.400 309.100 453.600 ;
        RECT 300.400 437.600 301.200 438.400 ;
        RECT 308.400 437.600 309.200 438.400 ;
        RECT 298.800 431.600 299.600 432.400 ;
        RECT 303.600 431.600 304.400 432.400 ;
        RECT 305.200 432.300 306.000 432.400 ;
        RECT 305.200 431.700 307.500 432.300 ;
        RECT 305.200 431.600 306.000 431.700 ;
        RECT 295.600 429.600 296.400 430.400 ;
        RECT 300.400 429.600 301.200 430.400 ;
        RECT 297.200 427.600 298.000 428.400 ;
        RECT 298.800 427.600 299.600 428.400 ;
        RECT 298.900 426.400 299.500 427.600 ;
        RECT 292.400 425.600 293.200 426.400 ;
        RECT 298.800 425.600 299.600 426.400 ;
        RECT 284.400 401.600 285.200 402.400 ;
        RECT 290.800 401.600 291.600 402.400 ;
        RECT 274.800 399.600 275.600 400.400 ;
        RECT 274.900 398.400 275.500 399.600 ;
        RECT 254.000 397.600 254.800 398.400 ;
        RECT 274.800 397.600 275.600 398.400 ;
        RECT 278.000 397.600 278.800 398.400 ;
        RECT 271.600 395.600 272.400 396.400 ;
        RECT 258.800 393.600 259.600 394.400 ;
        RECT 271.700 390.400 272.300 395.600 ;
        RECT 278.100 390.400 278.700 397.600 ;
        RECT 284.500 390.400 285.100 401.600 ;
        RECT 271.600 389.600 272.400 390.400 ;
        RECT 276.400 389.600 277.200 390.400 ;
        RECT 278.000 389.600 278.800 390.400 ;
        RECT 284.400 389.600 285.200 390.400 ;
        RECT 252.400 385.600 253.200 386.400 ;
        RECT 254.000 383.600 254.800 384.400 ;
        RECT 250.800 379.600 251.600 380.400 ;
        RECT 254.100 378.400 254.700 383.600 ;
        RECT 230.000 375.600 230.800 376.400 ;
        RECT 234.800 375.600 235.600 376.400 ;
        RECT 230.000 373.600 230.800 374.400 ;
        RECT 236.400 373.600 237.200 374.400 ;
        RECT 241.200 371.600 242.000 372.400 ;
        RECT 241.300 370.400 241.900 371.600 ;
        RECT 233.200 369.600 234.000 370.400 ;
        RECT 241.200 369.600 242.000 370.400 ;
        RECT 233.300 368.400 233.900 369.600 ;
        RECT 233.200 367.600 234.000 368.400 ;
        RECT 230.000 363.600 230.800 364.400 ;
        RECT 239.600 363.600 240.400 364.400 ;
        RECT 228.400 357.600 229.200 358.400 ;
        RECT 228.500 354.400 229.100 357.600 ;
        RECT 228.400 353.600 229.200 354.400 ;
        RECT 228.400 351.600 229.200 352.400 ;
        RECT 226.800 339.600 227.600 340.400 ;
        RECT 226.800 337.600 227.600 338.400 ;
        RECT 228.500 336.400 229.100 351.600 ;
        RECT 230.100 348.400 230.700 363.600 ;
        RECT 236.400 353.600 237.200 354.400 ;
        RECT 239.700 352.400 240.300 363.600 ;
        RECT 239.600 351.600 240.400 352.400 ;
        RECT 231.600 349.600 232.400 350.400 ;
        RECT 230.000 347.600 230.800 348.400 ;
        RECT 238.000 347.600 238.800 348.400 ;
        RECT 230.100 336.400 230.700 347.600 ;
        RECT 228.400 335.600 229.200 336.400 ;
        RECT 230.000 335.600 230.800 336.400 ;
        RECT 228.500 334.400 229.100 335.600 ;
        RECT 228.400 333.600 229.200 334.400 ;
        RECT 239.700 334.300 240.300 351.600 ;
        RECT 241.300 350.400 241.900 369.600 ;
        RECT 246.000 364.200 246.800 377.800 ;
        RECT 247.600 364.200 248.400 377.800 ;
        RECT 249.200 366.200 250.000 377.800 ;
        RECT 250.800 375.600 251.600 376.400 ;
        RECT 250.900 374.400 251.500 375.600 ;
        RECT 250.800 373.600 251.600 374.400 ;
        RECT 252.400 366.200 253.200 377.800 ;
        RECT 254.000 377.600 254.800 378.400 ;
        RECT 254.100 376.400 254.700 377.600 ;
        RECT 254.000 375.600 254.800 376.400 ;
        RECT 241.200 349.600 242.000 350.400 ;
        RECT 244.400 349.600 245.200 350.400 ;
        RECT 249.200 344.200 250.000 357.800 ;
        RECT 250.800 344.200 251.600 357.800 ;
        RECT 252.400 344.200 253.200 355.800 ;
        RECT 254.100 350.400 254.700 375.600 ;
        RECT 255.600 366.200 256.400 377.800 ;
        RECT 257.200 364.200 258.000 377.800 ;
        RECT 258.800 364.200 259.600 377.800 ;
        RECT 260.400 364.200 261.200 377.800 ;
        RECT 282.800 375.600 283.600 376.400 ;
        RECT 282.900 374.400 283.500 375.600 ;
        RECT 284.500 374.400 285.100 389.600 ;
        RECT 287.600 384.200 288.400 397.800 ;
        RECT 289.200 384.200 290.000 397.800 ;
        RECT 290.800 384.200 291.600 395.800 ;
        RECT 292.500 388.400 293.100 425.600 ;
        RECT 303.700 416.400 304.300 431.600 ;
        RECT 305.200 429.600 306.000 430.400 ;
        RECT 303.600 415.600 304.400 416.400 ;
        RECT 300.400 409.600 301.200 410.400 ;
        RECT 303.600 409.600 304.400 410.400 ;
        RECT 297.200 403.600 298.000 404.400 ;
        RECT 300.500 400.400 301.100 409.600 ;
        RECT 300.400 399.600 301.200 400.400 ;
        RECT 292.400 387.600 293.200 388.400 ;
        RECT 292.400 383.600 293.200 384.400 ;
        RECT 294.000 384.200 294.800 395.800 ;
        RECT 295.600 385.600 296.400 386.400 ;
        RECT 295.700 384.400 296.300 385.600 ;
        RECT 295.600 383.600 296.400 384.400 ;
        RECT 297.200 384.200 298.000 395.800 ;
        RECT 298.800 384.200 299.600 397.800 ;
        RECT 300.400 384.200 301.200 397.800 ;
        RECT 302.000 384.200 302.800 397.800 ;
        RECT 305.300 394.400 305.900 429.600 ;
        RECT 306.900 426.400 307.500 431.700 ;
        RECT 308.400 429.600 309.200 430.400 ;
        RECT 306.800 425.600 307.600 426.400 ;
        RECT 308.500 424.400 309.100 429.600 ;
        RECT 308.400 423.600 309.200 424.400 ;
        RECT 310.100 418.400 310.700 465.600 ;
        RECT 314.900 454.400 315.500 465.600 ;
        RECT 316.500 458.400 317.100 469.600 ;
        RECT 327.700 468.400 328.300 469.600 ;
        RECT 332.500 468.400 333.100 481.600 ;
        RECT 319.600 467.600 320.400 468.400 ;
        RECT 324.400 467.600 325.200 468.400 ;
        RECT 327.600 467.600 328.400 468.400 ;
        RECT 332.400 467.600 333.200 468.400 ;
        RECT 319.700 462.400 320.300 467.600 ;
        RECT 321.200 465.600 322.000 466.400 ;
        RECT 319.600 461.600 320.400 462.400 ;
        RECT 316.400 457.600 317.200 458.400 ;
        RECT 318.000 455.600 318.800 456.400 ;
        RECT 311.600 453.600 312.400 454.400 ;
        RECT 314.800 453.600 315.600 454.400 ;
        RECT 314.800 451.600 315.600 452.400 ;
        RECT 314.900 448.400 315.500 451.600 ;
        RECT 314.800 447.600 315.600 448.400 ;
        RECT 318.100 442.400 318.700 455.600 ;
        RECT 319.600 453.600 320.400 454.400 ;
        RECT 322.800 451.600 323.600 452.400 ;
        RECT 322.800 449.600 323.600 450.400 ;
        RECT 321.200 447.600 322.000 448.400 ;
        RECT 318.000 441.600 318.800 442.400 ;
        RECT 322.900 436.400 323.500 449.600 ;
        RECT 322.800 435.600 323.600 436.400 ;
        RECT 319.600 433.600 320.400 434.400 ;
        RECT 319.700 430.400 320.300 433.600 ;
        RECT 313.200 429.600 314.000 430.400 ;
        RECT 318.000 429.600 318.800 430.400 ;
        RECT 319.600 429.600 320.400 430.400 ;
        RECT 313.200 427.600 314.000 428.400 ;
        RECT 313.300 426.400 313.900 427.600 ;
        RECT 313.200 425.600 314.000 426.400 ;
        RECT 314.800 425.600 315.600 426.400 ;
        RECT 310.000 417.600 310.800 418.400 ;
        RECT 306.800 415.600 307.600 416.400 ;
        RECT 305.200 393.600 306.000 394.400 ;
        RECT 303.600 389.600 304.400 390.400 ;
        RECT 303.600 383.600 304.400 384.400 ;
        RECT 290.800 381.600 291.600 382.400 ;
        RECT 287.600 375.600 288.400 376.400 ;
        RECT 290.900 374.400 291.500 381.600 ;
        RECT 271.600 373.600 272.400 374.400 ;
        RECT 282.800 373.600 283.600 374.400 ;
        RECT 284.400 373.600 285.200 374.400 ;
        RECT 290.800 373.600 291.600 374.400 ;
        RECT 281.200 371.600 282.000 372.400 ;
        RECT 284.400 371.600 285.200 372.400 ;
        RECT 278.000 367.600 278.800 368.400 ;
        RECT 278.100 362.400 278.700 367.600 ;
        RECT 281.300 366.400 281.900 371.600 ;
        RECT 281.200 365.600 282.000 366.400 ;
        RECT 278.000 361.600 278.800 362.400 ;
        RECT 254.000 349.600 254.800 350.400 ;
        RECT 254.000 347.600 254.800 348.400 ;
        RECT 255.600 344.200 256.400 355.800 ;
        RECT 257.200 349.600 258.000 350.400 ;
        RECT 257.300 346.400 257.900 349.600 ;
        RECT 257.200 345.600 258.000 346.400 ;
        RECT 258.800 344.200 259.600 355.800 ;
        RECT 260.400 344.200 261.200 357.800 ;
        RECT 262.000 344.200 262.800 357.800 ;
        RECT 263.600 344.200 264.400 357.800 ;
        RECT 290.900 356.400 291.500 373.600 ;
        RECT 292.500 358.400 293.100 383.600 ;
        RECT 298.800 375.600 299.600 376.400 ;
        RECT 294.000 373.600 294.800 374.400 ;
        RECT 292.400 357.600 293.200 358.400 ;
        RECT 281.200 355.600 282.000 356.400 ;
        RECT 290.800 355.600 291.600 356.400 ;
        RECT 273.200 353.600 274.000 354.400 ;
        RECT 281.300 348.400 281.900 355.600 ;
        RECT 281.200 347.600 282.000 348.400 ;
        RECT 238.100 333.700 240.300 334.300 ;
        RECT 225.200 331.600 226.000 332.400 ;
        RECT 234.800 331.600 235.600 332.400 ;
        RECT 225.300 326.400 225.900 331.600 ;
        RECT 225.200 325.600 226.000 326.400 ;
        RECT 225.300 320.400 225.900 325.600 ;
        RECT 225.200 319.600 226.000 320.400 ;
        RECT 234.900 318.400 235.500 331.600 ;
        RECT 234.800 317.600 235.600 318.400 ;
        RECT 230.000 313.600 230.800 314.400 ;
        RECT 198.000 309.600 198.800 310.400 ;
        RECT 209.200 309.600 210.000 310.400 ;
        RECT 215.600 309.600 216.400 310.400 ;
        RECT 222.000 309.600 222.800 310.400 ;
        RECT 202.800 307.600 203.600 308.400 ;
        RECT 206.000 307.600 206.800 308.400 ;
        RECT 170.800 295.600 171.600 296.400 ;
        RECT 170.900 292.400 171.500 295.600 ;
        RECT 170.800 291.600 171.600 292.400 ;
        RECT 172.400 284.200 173.200 297.800 ;
        RECT 174.000 284.200 174.800 297.800 ;
        RECT 175.600 286.200 176.400 297.800 ;
        RECT 177.300 294.400 177.900 303.600 ;
        RECT 180.400 301.600 181.200 302.400 ;
        RECT 177.200 293.600 178.000 294.400 ;
        RECT 178.800 286.200 179.600 297.800 ;
        RECT 180.500 296.400 181.100 301.600 ;
        RECT 199.600 299.600 200.400 300.400 ;
        RECT 180.400 295.600 181.200 296.400 ;
        RECT 180.400 293.600 181.200 294.400 ;
        RECT 180.500 290.400 181.100 293.600 ;
        RECT 180.400 289.600 181.200 290.400 ;
        RECT 178.800 283.600 179.600 284.400 ;
        RECT 170.800 279.600 171.600 280.400 ;
        RECT 170.900 272.400 171.500 279.600 ;
        RECT 170.800 271.600 171.600 272.400 ;
        RECT 174.000 271.600 174.800 272.400 ;
        RECT 178.900 270.400 179.500 283.600 ;
        RECT 164.400 269.600 165.200 270.400 ;
        RECT 178.800 269.600 179.600 270.400 ;
        RECT 180.500 268.400 181.100 289.600 ;
        RECT 182.000 286.200 182.800 297.800 ;
        RECT 183.600 284.200 184.400 297.800 ;
        RECT 185.200 284.200 186.000 297.800 ;
        RECT 186.800 284.200 187.600 297.800 ;
        RECT 190.000 297.600 190.800 298.400 ;
        RECT 185.200 279.600 186.000 280.400 ;
        RECT 170.800 267.600 171.600 268.400 ;
        RECT 180.400 268.300 181.200 268.400 ;
        RECT 180.400 267.700 182.700 268.300 ;
        RECT 180.400 267.600 181.200 267.700 ;
        RECT 142.000 259.600 142.800 260.400 ;
        RECT 142.100 254.400 142.700 259.600 ;
        RECT 182.100 256.400 182.700 267.700 ;
        RECT 183.600 263.600 184.400 264.400 ;
        RECT 183.700 260.400 184.300 263.600 ;
        RECT 183.600 259.600 184.400 260.400 ;
        RECT 156.400 255.600 157.200 256.400 ;
        RECT 169.200 255.600 170.000 256.400 ;
        RECT 182.000 255.600 182.800 256.400 ;
        RECT 169.300 254.400 169.900 255.600 ;
        RECT 140.400 253.600 141.200 254.400 ;
        RECT 142.000 253.600 142.800 254.400 ;
        RECT 159.600 253.600 160.400 254.400 ;
        RECT 169.200 253.600 170.000 254.400 ;
        RECT 183.600 253.600 184.400 254.400 ;
        RECT 137.200 241.600 138.000 242.400 ;
        RECT 137.300 230.400 137.900 241.600 ;
        RECT 140.500 238.400 141.100 253.600 ;
        RECT 156.400 249.600 157.200 250.400 ;
        RECT 153.200 243.600 154.000 244.400 ;
        RECT 153.300 240.400 153.900 243.600 ;
        RECT 156.500 240.400 157.100 249.600 ;
        RECT 153.200 239.600 154.000 240.400 ;
        RECT 156.400 239.600 157.200 240.400 ;
        RECT 140.400 237.600 141.200 238.400 ;
        RECT 137.200 229.600 138.000 230.400 ;
        RECT 148.400 229.600 149.200 230.400 ;
        RECT 135.600 227.600 136.400 228.400 ;
        RECT 130.800 225.600 131.600 226.400 ;
        RECT 134.000 225.600 134.800 226.400 ;
        RECT 134.000 223.600 134.800 224.400 ;
        RECT 134.100 220.400 134.700 223.600 ;
        RECT 135.700 222.400 136.300 227.600 ;
        RECT 135.600 221.600 136.400 222.400 ;
        RECT 134.000 219.600 134.800 220.400 ;
        RECT 138.800 219.600 139.600 220.400 ;
        RECT 95.600 213.600 96.400 214.400 ;
        RECT 108.400 213.600 109.200 214.400 ;
        RECT 124.400 213.600 125.200 214.400 ;
        RECT 90.800 211.600 91.600 212.400 ;
        RECT 118.000 207.600 118.800 208.400 ;
        RECT 106.800 203.600 107.600 204.400 ;
        RECT 87.600 187.600 88.400 188.400 ;
        RECT 73.200 183.600 74.000 184.400 ;
        RECT 79.600 183.600 80.400 184.400 ;
        RECT 89.200 184.200 90.000 195.800 ;
        RECT 90.800 189.400 91.600 190.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 92.500 186.400 93.100 187.600 ;
        RECT 92.400 185.600 93.200 186.400 ;
        RECT 70.000 175.600 70.800 176.400 ;
        RECT 58.800 173.600 59.600 174.400 ;
        RECT 60.400 173.600 61.200 174.400 ;
        RECT 65.200 173.600 66.000 174.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 70.100 172.400 70.700 175.600 ;
        RECT 62.000 171.600 62.800 172.400 ;
        RECT 70.000 171.600 70.800 172.400 ;
        RECT 62.100 170.400 62.700 171.600 ;
        RECT 55.600 169.600 56.400 170.400 ;
        RECT 62.000 169.600 62.800 170.400 ;
        RECT 65.200 169.600 66.000 170.400 ;
        RECT 55.600 167.600 56.400 168.400 ;
        RECT 54.000 163.600 54.800 164.400 ;
        RECT 54.100 162.400 54.700 163.600 ;
        RECT 54.000 161.600 54.800 162.400 ;
        RECT 73.300 156.400 73.900 183.600 ;
        RECT 79.700 178.400 80.300 183.600 ;
        RECT 79.600 177.600 80.400 178.400 ;
        RECT 74.800 175.600 75.600 176.400 ;
        RECT 74.900 170.400 75.500 175.600 ;
        RECT 79.600 171.600 80.400 172.400 ;
        RECT 74.800 169.600 75.600 170.400 ;
        RECT 84.400 164.200 85.200 177.800 ;
        RECT 86.000 164.200 86.800 177.800 ;
        RECT 87.600 166.200 88.400 177.800 ;
        RECT 89.200 173.600 90.000 174.400 ;
        RECT 90.800 166.200 91.600 177.800 ;
        RECT 92.500 176.400 93.100 185.600 ;
        RECT 98.800 184.200 99.600 195.800 ;
        RECT 105.200 195.600 106.000 196.400 ;
        RECT 105.300 194.400 105.900 195.600 ;
        RECT 105.200 193.600 106.000 194.400 ;
        RECT 103.600 183.600 104.400 184.400 ;
        RECT 92.400 175.600 93.200 176.400 ;
        RECT 94.000 166.200 94.800 177.800 ;
        RECT 90.800 163.600 91.600 164.400 ;
        RECT 95.600 164.200 96.400 177.800 ;
        RECT 97.200 164.200 98.000 177.800 ;
        RECT 98.800 164.200 99.600 177.800 ;
        RECT 87.600 161.600 88.400 162.400 ;
        RECT 73.200 155.600 74.000 156.400 ;
        RECT 79.600 155.600 80.400 156.400 ;
        RECT 49.200 151.600 50.000 152.400 ;
        RECT 52.400 151.600 53.200 152.400 ;
        RECT 58.800 151.600 59.600 152.400 ;
        RECT 68.400 151.600 69.200 152.400 ;
        RECT 49.300 150.400 49.900 151.600 ;
        RECT 52.500 150.400 53.100 151.600 ;
        RECT 58.900 150.400 59.500 151.600 ;
        RECT 79.700 150.400 80.300 155.600 ;
        RECT 86.000 151.600 86.800 152.400 ;
        RECT 49.200 149.600 50.000 150.400 ;
        RECT 50.800 149.600 51.600 150.400 ;
        RECT 52.400 149.600 53.200 150.400 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 58.800 149.600 59.600 150.400 ;
        RECT 60.400 149.600 61.200 150.400 ;
        RECT 63.600 149.600 64.400 150.400 ;
        RECT 66.800 149.600 67.600 150.400 ;
        RECT 71.600 149.600 72.400 150.400 ;
        RECT 79.600 149.600 80.400 150.400 ;
        RECT 82.800 149.600 83.600 150.400 ;
        RECT 49.300 138.400 49.900 149.600 ;
        RECT 50.900 140.400 51.500 149.600 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 52.400 141.600 53.200 142.400 ;
        RECT 50.800 139.600 51.600 140.400 ;
        RECT 46.000 126.200 46.800 137.800 ;
        RECT 49.200 137.600 50.000 138.400 ;
        RECT 50.800 137.600 51.600 138.400 ;
        RECT 50.900 130.400 51.500 137.600 ;
        RECT 52.500 134.400 53.100 141.600 ;
        RECT 54.100 134.400 54.700 143.600 ;
        RECT 60.500 136.400 61.100 149.600 ;
        RECT 66.900 148.400 67.500 149.600 ;
        RECT 62.000 147.600 62.800 148.400 ;
        RECT 66.800 147.600 67.600 148.400 ;
        RECT 62.100 146.400 62.700 147.600 ;
        RECT 62.000 145.600 62.800 146.400 ;
        RECT 60.400 135.600 61.200 136.400 ;
        RECT 52.400 133.600 53.200 134.400 ;
        RECT 54.000 133.600 54.800 134.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 50.800 129.600 51.600 130.400 ;
        RECT 47.600 127.600 48.400 128.400 ;
        RECT 46.000 119.600 46.800 120.400 ;
        RECT 46.100 118.400 46.700 119.600 ;
        RECT 46.000 117.600 46.800 118.400 ;
        RECT 47.700 108.400 48.300 127.600 ;
        RECT 52.500 120.400 53.100 133.600 ;
        RECT 54.100 132.400 54.700 133.600 ;
        RECT 58.900 132.400 59.500 133.600 ;
        RECT 54.000 131.600 54.800 132.400 ;
        RECT 58.800 131.600 59.600 132.400 ;
        RECT 57.200 129.600 58.000 130.400 ;
        RECT 52.400 119.600 53.200 120.400 ;
        RECT 47.600 107.600 48.400 108.400 ;
        RECT 49.200 106.200 50.000 111.800 ;
        RECT 50.800 107.600 51.600 108.400 ;
        RECT 46.000 103.600 46.800 104.400 ;
        RECT 52.400 104.200 53.200 115.800 ;
        RECT 55.600 111.600 56.400 112.400 ;
        RECT 55.700 110.400 56.300 111.600 ;
        RECT 60.500 110.400 61.100 135.600 ;
        RECT 62.100 134.300 62.700 145.600 ;
        RECT 71.700 144.400 72.300 149.600 ;
        RECT 73.200 147.600 74.000 148.400 ;
        RECT 74.800 147.600 75.600 148.400 ;
        RECT 71.600 143.600 72.400 144.400 ;
        RECT 73.300 142.400 73.900 147.600 ;
        RECT 74.900 146.400 75.500 147.600 ;
        RECT 74.800 145.600 75.600 146.400 ;
        RECT 73.200 141.600 74.000 142.400 ;
        RECT 68.400 139.600 69.200 140.400 ;
        RECT 66.800 137.600 67.600 138.400 ;
        RECT 63.600 134.300 64.400 134.400 ;
        RECT 62.100 133.700 64.400 134.300 ;
        RECT 63.600 133.600 64.400 133.700 ;
        RECT 66.900 132.400 67.500 137.600 ;
        RECT 66.800 131.600 67.600 132.400 ;
        RECT 55.600 109.600 56.400 110.400 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 62.000 104.200 62.800 115.800 ;
        RECT 66.800 113.600 67.600 114.400 ;
        RECT 68.500 110.400 69.100 139.600 ;
        RECT 71.600 137.600 72.400 138.400 ;
        RECT 71.700 132.400 72.300 137.600 ;
        RECT 74.900 134.400 75.500 145.600 ;
        RECT 76.400 135.600 77.200 136.400 ;
        RECT 74.800 133.600 75.600 134.400 ;
        RECT 71.600 131.600 72.400 132.400 ;
        RECT 73.200 131.600 74.000 132.400 ;
        RECT 74.800 131.600 75.600 132.400 ;
        RECT 71.700 130.400 72.300 131.600 ;
        RECT 71.600 129.600 72.400 130.400 ;
        RECT 73.300 128.300 73.900 131.600 ;
        RECT 71.700 127.700 73.900 128.300 ;
        RECT 71.700 110.400 72.300 127.700 ;
        RECT 74.900 126.300 75.500 131.600 ;
        RECT 76.500 130.400 77.100 135.600 ;
        RECT 76.400 129.600 77.200 130.400 ;
        RECT 73.300 125.700 75.500 126.300 ;
        RECT 73.300 118.400 73.900 125.700 ;
        RECT 76.400 123.600 77.200 124.400 ;
        RECT 73.200 117.600 74.000 118.400 ;
        RECT 76.500 112.400 77.100 123.600 ;
        RECT 78.000 113.600 78.800 114.400 ;
        RECT 76.400 111.600 77.200 112.400 ;
        RECT 78.100 110.400 78.700 113.600 ;
        RECT 66.800 109.600 67.600 110.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 70.000 109.600 70.800 110.400 ;
        RECT 71.600 109.600 72.400 110.400 ;
        RECT 78.000 109.600 78.800 110.400 ;
        RECT 46.100 98.400 46.700 103.600 ;
        RECT 46.000 97.600 46.800 98.400 ;
        RECT 52.400 97.600 53.200 98.400 ;
        RECT 58.800 97.600 59.600 98.400 ;
        RECT 47.600 95.600 48.400 96.400 ;
        RECT 47.700 90.400 48.300 95.600 ;
        RECT 52.500 92.400 53.100 97.600 ;
        RECT 65.200 95.600 66.000 96.400 ;
        RECT 54.000 93.600 54.800 94.400 ;
        RECT 63.600 93.600 64.400 94.400 ;
        RECT 52.400 91.600 53.200 92.400 ;
        RECT 54.000 91.600 54.800 92.400 ;
        RECT 57.200 91.600 58.000 92.400 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 52.400 87.600 53.200 88.400 ;
        RECT 50.800 85.600 51.600 86.400 ;
        RECT 46.000 71.600 46.800 72.400 ;
        RECT 50.900 70.400 51.500 85.600 ;
        RECT 42.800 69.700 45.100 70.300 ;
        RECT 42.800 69.600 43.600 69.700 ;
        RECT 34.800 57.600 35.600 58.400 ;
        RECT 39.600 57.600 40.400 58.400 ;
        RECT 41.200 55.600 42.000 56.400 ;
        RECT 41.300 54.400 41.900 55.600 ;
        RECT 44.500 54.400 45.100 69.700 ;
        RECT 50.800 69.600 51.600 70.400 ;
        RECT 47.600 67.600 48.400 68.400 ;
        RECT 52.400 63.600 53.200 64.400 ;
        RECT 50.800 59.600 51.600 60.400 ;
        RECT 49.200 57.600 50.000 58.400 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 36.400 53.600 37.200 54.400 ;
        RECT 38.000 53.600 38.800 54.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 44.400 53.600 45.200 54.400 ;
        RECT 22.000 51.600 22.800 52.400 ;
        RECT 30.000 51.600 30.800 52.400 ;
        RECT 18.800 49.600 19.600 50.400 ;
        RECT 25.200 49.600 26.000 50.400 ;
        RECT 33.200 47.600 34.000 48.400 ;
        RECT 12.400 43.600 13.200 44.400 ;
        RECT 17.200 43.600 18.000 44.400 ;
        RECT 2.800 29.600 3.600 30.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 1.200 16.300 2.000 16.400 ;
        RECT 2.900 16.300 3.500 29.600 ;
        RECT 1.200 15.700 3.500 16.300 ;
        RECT 1.200 15.600 2.000 15.700 ;
        RECT 2.800 13.600 3.600 14.400 ;
        RECT 7.700 12.400 8.300 29.600 ;
        RECT 9.200 24.200 10.000 37.800 ;
        RECT 10.800 24.200 11.600 37.800 ;
        RECT 12.400 24.200 13.200 35.800 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 15.600 24.200 16.400 35.800 ;
        RECT 17.300 26.400 17.900 43.600 ;
        RECT 33.300 38.400 33.900 47.600 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 12.400 4.200 13.200 17.800 ;
        RECT 14.000 4.200 14.800 17.800 ;
        RECT 15.600 6.200 16.400 17.800 ;
        RECT 17.300 16.400 17.900 25.600 ;
        RECT 18.800 24.200 19.600 35.800 ;
        RECT 20.400 24.200 21.200 37.800 ;
        RECT 22.000 24.200 22.800 37.800 ;
        RECT 23.600 24.200 24.400 37.800 ;
        RECT 33.200 37.600 34.000 38.400 ;
        RECT 33.300 32.400 33.900 37.600 ;
        RECT 33.200 31.600 34.000 32.400 ;
        RECT 38.100 26.400 38.700 53.600 ;
        RECT 44.500 52.400 45.100 53.600 ;
        RECT 49.300 52.400 49.900 57.600 ;
        RECT 50.900 52.400 51.500 59.600 ;
        RECT 52.500 54.400 53.100 63.600 ;
        RECT 54.100 56.400 54.700 91.600 ;
        RECT 57.300 86.400 57.900 91.600 ;
        RECT 57.200 85.600 58.000 86.400 ;
        RECT 58.800 85.600 59.600 86.400 ;
        RECT 55.600 83.600 56.400 84.400 ;
        RECT 55.700 70.400 56.300 83.600 ;
        RECT 58.900 70.400 59.500 85.600 ;
        RECT 55.600 69.600 56.400 70.400 ;
        RECT 58.800 69.600 59.600 70.400 ;
        RECT 60.400 69.600 61.200 70.400 ;
        RECT 57.200 61.600 58.000 62.400 ;
        RECT 54.000 55.600 54.800 56.400 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 44.400 51.600 45.200 52.400 ;
        RECT 49.200 51.600 50.000 52.400 ;
        RECT 50.800 51.600 51.600 52.400 ;
        RECT 49.300 50.400 49.900 51.600 ;
        RECT 49.200 49.600 50.000 50.400 ;
        RECT 50.800 49.600 51.600 50.400 ;
        RECT 41.200 47.600 42.000 48.400 ;
        RECT 41.300 34.400 41.900 47.600 ;
        RECT 41.200 33.600 42.000 34.400 ;
        RECT 49.200 33.600 50.000 34.400 ;
        RECT 46.000 31.600 46.800 32.400 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 46.000 27.600 46.800 28.400 ;
        RECT 38.000 25.600 38.800 26.400 ;
        RECT 17.200 15.600 18.000 16.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 20.400 15.600 21.200 16.400 ;
        RECT 22.000 6.200 22.800 17.800 ;
        RECT 23.600 4.200 24.400 17.800 ;
        RECT 25.200 4.200 26.000 17.800 ;
        RECT 26.800 4.200 27.600 17.800 ;
        RECT 38.100 16.400 38.700 25.600 ;
        RECT 46.100 18.400 46.700 27.600 ;
        RECT 49.300 18.400 49.900 33.600 ;
        RECT 50.900 30.400 51.500 49.600 ;
        RECT 50.800 29.600 51.600 30.400 ;
        RECT 46.000 17.600 46.800 18.400 ;
        RECT 49.200 17.600 50.000 18.400 ;
        RECT 38.000 15.600 38.800 16.400 ;
        RECT 50.900 14.400 51.500 29.600 ;
        RECT 52.500 28.400 53.100 53.600 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 57.300 50.400 57.900 61.600 ;
        RECT 58.900 60.400 59.500 69.600 ;
        RECT 63.700 68.400 64.300 93.600 ;
        RECT 65.300 92.400 65.900 95.600 ;
        RECT 65.200 91.600 66.000 92.400 ;
        RECT 66.900 70.400 67.500 109.600 ;
        RECT 68.500 92.400 69.100 109.600 ;
        RECT 70.100 108.400 70.700 109.600 ;
        RECT 70.000 107.600 70.800 108.400 ;
        RECT 78.100 106.400 78.700 109.600 ;
        RECT 79.700 106.400 80.300 149.600 ;
        RECT 81.200 147.600 82.000 148.400 ;
        RECT 81.300 142.400 81.900 147.600 ;
        RECT 82.900 144.400 83.500 149.600 ;
        RECT 82.800 144.300 83.600 144.400 ;
        RECT 82.800 143.700 85.100 144.300 ;
        RECT 82.800 143.600 83.600 143.700 ;
        RECT 81.200 141.600 82.000 142.400 ;
        RECT 84.500 132.400 85.100 143.700 ;
        RECT 86.000 141.600 86.800 142.400 ;
        RECT 86.100 134.400 86.700 141.600 ;
        RECT 87.700 136.400 88.300 161.600 ;
        RECT 90.900 158.400 91.500 163.600 ;
        RECT 90.800 157.600 91.600 158.400 ;
        RECT 94.000 153.600 94.800 154.400 ;
        RECT 90.800 149.600 91.600 150.400 ;
        RECT 90.900 148.400 91.500 149.600 ;
        RECT 90.800 147.600 91.600 148.400 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 92.500 146.400 93.100 147.600 ;
        RECT 92.400 145.600 93.200 146.400 ;
        RECT 98.800 144.200 99.600 155.800 ;
        RECT 103.700 152.400 104.300 183.600 ;
        RECT 103.600 151.600 104.400 152.400 ;
        RECT 105.200 149.600 106.000 150.400 ;
        RECT 106.900 148.400 107.500 203.600 ;
        RECT 118.100 190.400 118.700 207.600 ;
        RECT 129.200 204.200 130.000 217.800 ;
        RECT 130.800 204.200 131.600 217.800 ;
        RECT 132.400 204.200 133.200 217.800 ;
        RECT 134.000 206.200 134.800 217.800 ;
        RECT 135.600 215.600 136.400 216.400 ;
        RECT 137.200 206.200 138.000 217.800 ;
        RECT 138.900 214.400 139.500 219.600 ;
        RECT 138.800 213.600 139.600 214.400 ;
        RECT 140.400 206.200 141.200 217.800 ;
        RECT 142.000 204.200 142.800 217.800 ;
        RECT 143.600 204.200 144.400 217.800 ;
        RECT 148.500 212.400 149.100 229.600 ;
        RECT 150.000 224.200 150.800 237.800 ;
        RECT 151.600 224.200 152.400 237.800 ;
        RECT 153.200 224.200 154.000 237.800 ;
        RECT 154.800 224.200 155.600 235.800 ;
        RECT 156.500 226.400 157.100 239.600 ;
        RECT 156.400 225.600 157.200 226.400 ;
        RECT 156.500 224.400 157.100 225.600 ;
        RECT 156.400 223.600 157.200 224.400 ;
        RECT 158.000 224.200 158.800 235.800 ;
        RECT 159.700 232.400 160.300 253.600 ;
        RECT 166.000 251.600 166.800 252.400 ;
        RECT 167.600 251.600 168.400 252.400 ;
        RECT 178.800 251.600 179.600 252.400 ;
        RECT 180.400 251.600 181.200 252.400 ;
        RECT 166.100 250.300 166.700 251.600 ;
        RECT 166.100 249.700 168.300 250.300 ;
        RECT 167.700 242.400 168.300 249.700 ;
        RECT 175.600 243.600 176.400 244.400 ;
        RECT 167.600 241.600 168.400 242.400 ;
        RECT 167.700 238.400 168.300 241.600 ;
        RECT 159.600 231.600 160.400 232.400 ;
        RECT 159.600 227.600 160.400 228.400 ;
        RECT 161.200 224.200 162.000 235.800 ;
        RECT 162.800 224.200 163.600 237.800 ;
        RECT 164.400 224.200 165.200 237.800 ;
        RECT 167.600 237.600 168.400 238.400 ;
        RECT 167.600 233.600 168.400 234.400 ;
        RECT 167.700 230.400 168.300 233.600 ;
        RECT 167.600 229.600 168.400 230.400 ;
        RECT 175.700 228.400 176.300 243.600 ;
        RECT 175.600 227.600 176.400 228.400 ;
        RECT 174.000 225.600 174.800 226.400 ;
        RECT 174.000 223.600 174.800 224.400 ;
        RECT 154.800 217.600 155.600 218.400 ;
        RECT 156.500 216.400 157.100 223.600 ;
        RECT 158.000 221.600 158.800 222.400 ;
        RECT 150.000 215.600 150.800 216.400 ;
        RECT 156.400 215.600 157.200 216.400 ;
        RECT 148.400 211.600 149.200 212.400 ;
        RECT 118.000 189.600 118.800 190.400 ;
        RECT 108.400 187.600 109.200 188.400 ;
        RECT 119.600 187.600 120.400 188.400 ;
        RECT 114.800 183.600 115.600 184.400 ;
        RECT 108.400 169.600 109.200 170.400 ;
        RECT 111.600 165.600 112.400 166.400 ;
        RECT 114.900 164.400 115.500 183.600 ;
        RECT 118.000 177.600 118.800 178.400 ;
        RECT 118.100 176.400 118.700 177.600 ;
        RECT 118.000 175.600 118.800 176.400 ;
        RECT 119.700 172.400 120.300 187.600 ;
        RECT 121.200 186.200 122.000 191.800 ;
        RECT 122.800 187.600 123.600 188.400 ;
        RECT 122.900 186.400 123.500 187.600 ;
        RECT 122.800 185.600 123.600 186.400 ;
        RECT 124.400 184.200 125.200 195.800 ;
        RECT 130.800 189.600 131.600 190.400 ;
        RECT 130.900 178.400 131.500 189.600 ;
        RECT 134.000 184.200 134.800 195.800 ;
        RECT 140.400 191.600 141.200 192.400 ;
        RECT 142.000 187.600 142.800 188.400 ;
        RECT 142.100 186.400 142.700 187.600 ;
        RECT 142.000 185.600 142.800 186.400 ;
        RECT 143.600 186.200 144.400 191.800 ;
        RECT 138.800 183.600 139.600 184.400 ;
        RECT 146.800 184.200 147.600 195.800 ;
        RECT 150.100 190.400 150.700 215.600 ;
        RECT 150.000 189.600 150.800 190.400 ;
        RECT 153.200 189.600 154.000 190.400 ;
        RECT 150.100 188.400 150.700 189.600 ;
        RECT 150.000 187.600 150.800 188.400 ;
        RECT 130.800 177.600 131.600 178.400 ;
        RECT 134.000 175.600 134.800 176.400 ;
        RECT 122.800 173.600 123.600 174.400 ;
        RECT 122.900 172.400 123.500 173.600 ;
        RECT 134.100 172.400 134.700 175.600 ;
        RECT 135.600 173.600 136.400 174.400 ;
        RECT 137.200 173.600 138.000 174.400 ;
        RECT 119.600 171.600 120.400 172.400 ;
        RECT 122.800 171.600 123.600 172.400 ;
        RECT 124.400 171.600 125.200 172.400 ;
        RECT 134.000 171.600 134.800 172.400 ;
        RECT 124.500 170.400 125.100 171.600 ;
        RECT 118.000 169.600 118.800 170.400 ;
        RECT 124.400 170.300 125.200 170.400 ;
        RECT 122.900 169.700 125.200 170.300 ;
        RECT 121.200 167.600 122.000 168.400 ;
        RECT 114.800 163.600 115.600 164.400 ;
        RECT 122.900 158.400 123.500 169.700 ;
        RECT 124.400 169.600 125.200 169.700 ;
        RECT 130.800 169.600 131.600 170.400 ;
        RECT 135.700 170.300 136.300 173.600 ;
        RECT 137.300 172.400 137.900 173.600 ;
        RECT 138.900 172.400 139.500 183.600 ;
        RECT 140.400 175.600 141.200 176.400 ;
        RECT 150.000 175.600 150.800 176.400 ;
        RECT 137.200 171.600 138.000 172.400 ;
        RECT 138.800 171.600 139.600 172.400 ;
        RECT 143.600 171.600 144.400 172.400 ;
        RECT 146.800 171.600 147.600 172.400 ;
        RECT 135.700 169.700 137.900 170.300 ;
        RECT 124.400 163.600 125.200 164.400 ;
        RECT 127.600 163.600 128.400 164.400 ;
        RECT 122.800 157.600 123.600 158.400 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 100.400 145.600 101.200 146.400 ;
        RECT 87.600 135.600 88.400 136.400 ;
        RECT 86.000 133.600 86.800 134.400 ;
        RECT 90.800 133.600 91.600 134.400 ;
        RECT 84.400 131.600 85.200 132.400 ;
        RECT 92.400 131.600 93.200 132.400 ;
        RECT 97.200 131.600 98.000 132.400 ;
        RECT 98.800 131.600 99.600 132.400 ;
        RECT 81.200 129.600 82.000 130.400 ;
        RECT 81.300 114.400 81.900 129.600 ;
        RECT 95.600 123.600 96.400 124.400 ;
        RECT 81.200 113.600 82.000 114.400 ;
        RECT 70.000 105.600 70.800 106.400 ;
        RECT 78.000 105.600 78.800 106.400 ;
        RECT 79.600 105.600 80.400 106.400 ;
        RECT 81.200 106.200 82.000 111.800 ;
        RECT 70.100 92.400 70.700 105.600 ;
        RECT 79.600 103.600 80.400 104.400 ;
        RECT 84.400 104.200 85.200 115.800 ;
        RECT 87.600 111.600 88.400 112.400 ;
        RECT 87.700 110.400 88.300 111.600 ;
        RECT 87.600 109.600 88.400 110.400 ;
        RECT 87.600 107.600 88.400 108.400 ;
        RECT 79.700 100.400 80.300 103.600 ;
        RECT 79.600 99.600 80.400 100.400 ;
        RECT 71.600 97.600 72.400 98.400 ;
        RECT 71.700 96.400 72.300 97.600 ;
        RECT 71.600 95.600 72.400 96.400 ;
        RECT 68.400 91.600 69.200 92.400 ;
        RECT 70.000 91.600 70.800 92.400 ;
        RECT 76.400 86.200 77.200 97.800 ;
        RECT 82.800 91.600 83.600 92.400 ;
        RECT 82.900 88.400 83.500 91.600 ;
        RECT 82.800 87.600 83.600 88.400 ;
        RECT 86.000 86.200 86.800 97.800 ;
        RECT 87.700 94.400 88.300 107.600 ;
        RECT 94.000 104.200 94.800 115.800 ;
        RECT 95.700 110.400 96.300 123.600 ;
        RECT 97.300 118.300 97.900 131.600 ;
        RECT 100.500 130.400 101.100 145.600 ;
        RECT 108.400 144.200 109.200 155.800 ;
        RECT 111.600 146.200 112.400 151.800 ;
        RECT 119.600 151.600 120.400 152.400 ;
        RECT 119.700 150.400 120.300 151.600 ;
        RECT 118.000 149.600 118.800 150.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 118.100 146.400 118.700 149.600 ;
        RECT 118.000 145.600 118.800 146.400 ;
        RECT 105.200 141.600 106.000 142.400 ;
        RECT 102.000 131.600 102.800 132.400 ;
        RECT 100.400 129.600 101.200 130.400 ;
        RECT 102.100 124.400 102.700 131.600 ;
        RECT 103.600 127.600 104.400 128.400 ;
        RECT 102.000 123.600 102.800 124.400 ;
        RECT 98.800 118.300 99.600 118.400 ;
        RECT 97.300 117.700 99.600 118.300 ;
        RECT 98.800 117.600 99.600 117.700 ;
        RECT 98.800 115.600 99.600 116.400 ;
        RECT 95.600 109.600 96.400 110.400 ;
        RECT 98.900 102.400 99.500 115.600 ;
        RECT 102.000 111.600 102.800 112.400 ;
        RECT 102.000 109.600 102.800 110.400 ;
        RECT 100.400 107.600 101.200 108.400 ;
        RECT 100.500 102.400 101.100 107.600 ;
        RECT 102.000 105.600 102.800 106.400 ;
        RECT 94.000 101.600 94.800 102.400 ;
        RECT 98.800 101.600 99.600 102.400 ;
        RECT 100.400 101.600 101.200 102.400 ;
        RECT 87.600 93.600 88.400 94.400 ;
        RECT 86.000 83.600 86.800 84.400 ;
        RECT 86.100 78.400 86.700 83.600 ;
        RECT 87.700 82.400 88.300 93.600 ;
        RECT 89.200 90.200 90.000 95.800 ;
        RECT 90.800 95.600 91.600 96.400 ;
        RECT 94.100 92.400 94.700 101.600 ;
        RECT 97.200 93.600 98.000 94.400 ;
        RECT 92.400 91.600 93.200 92.400 ;
        RECT 94.000 91.600 94.800 92.400 ;
        RECT 97.300 88.400 97.900 93.600 ;
        RECT 102.100 92.400 102.700 105.600 ;
        RECT 103.700 92.400 104.300 127.600 ;
        RECT 105.300 112.400 105.900 141.600 ;
        RECT 108.400 135.600 109.200 136.400 ;
        RECT 108.500 134.400 109.100 135.600 ;
        RECT 108.400 133.600 109.200 134.400 ;
        RECT 111.600 133.600 112.400 134.400 ;
        RECT 118.000 134.300 118.800 134.400 ;
        RECT 119.700 134.300 120.300 149.600 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 121.300 146.400 121.900 147.600 ;
        RECT 121.200 145.600 122.000 146.400 ;
        RECT 118.000 133.700 120.300 134.300 ;
        RECT 118.000 133.600 118.800 133.700 ;
        RECT 110.000 132.300 110.800 132.400 ;
        RECT 108.500 131.700 110.800 132.300 ;
        RECT 106.800 117.600 107.600 118.400 ;
        RECT 106.900 112.400 107.500 117.600 ;
        RECT 105.200 111.600 106.000 112.400 ;
        RECT 106.800 111.600 107.600 112.400 ;
        RECT 106.900 110.400 107.500 111.600 ;
        RECT 106.800 109.600 107.600 110.400 ;
        RECT 108.500 98.300 109.100 131.700 ;
        RECT 110.000 131.600 110.800 131.700 ;
        RECT 121.200 129.600 122.000 130.400 ;
        RECT 118.000 117.600 118.800 118.400 ;
        RECT 111.600 111.600 112.400 112.400 ;
        RECT 114.800 111.600 115.600 112.400 ;
        RECT 111.700 108.400 112.300 111.600 ;
        RECT 114.900 110.400 115.500 111.600 ;
        RECT 118.100 110.400 118.700 117.600 ;
        RECT 121.300 114.400 121.900 129.600 ;
        RECT 122.900 118.400 123.500 157.600 ;
        RECT 124.500 150.400 125.100 163.600 ;
        RECT 127.700 154.400 128.300 163.600 ;
        RECT 127.600 153.600 128.400 154.400 ;
        RECT 127.700 150.400 128.300 153.600 ;
        RECT 130.900 150.400 131.500 169.600 ;
        RECT 137.300 158.400 137.900 169.700 ;
        RECT 138.900 158.400 139.500 171.600 ;
        RECT 143.700 164.400 144.300 171.600 ;
        RECT 153.300 170.400 153.900 189.600 ;
        RECT 156.400 184.200 157.200 195.800 ;
        RECT 154.800 179.600 155.600 180.400 ;
        RECT 154.900 172.400 155.500 179.600 ;
        RECT 158.100 176.400 158.700 221.600 ;
        RECT 164.400 204.200 165.200 217.800 ;
        RECT 166.000 204.200 166.800 217.800 ;
        RECT 167.600 204.200 168.400 217.800 ;
        RECT 169.200 206.200 170.000 217.800 ;
        RECT 170.800 215.600 171.600 216.400 ;
        RECT 162.800 186.200 163.600 191.800 ;
        RECT 164.400 189.600 165.200 190.400 ;
        RECT 164.500 188.400 165.100 189.600 ;
        RECT 164.400 187.600 165.200 188.400 ;
        RECT 161.200 183.600 162.000 184.400 ;
        RECT 161.300 176.400 161.900 183.600 ;
        RECT 158.000 175.600 158.800 176.400 ;
        RECT 161.200 175.600 162.000 176.400 ;
        RECT 158.100 174.400 158.700 175.600 ;
        RECT 158.000 173.600 158.800 174.400 ;
        RECT 162.800 173.600 163.600 174.400 ;
        RECT 154.800 171.600 155.600 172.400 ;
        RECT 156.400 171.600 157.200 172.400 ;
        RECT 148.400 169.600 149.200 170.400 ;
        RECT 151.600 169.600 152.400 170.400 ;
        RECT 153.200 169.600 154.000 170.400 ;
        RECT 151.700 168.400 152.300 169.600 ;
        RECT 151.600 167.600 152.400 168.400 ;
        RECT 154.800 167.600 155.600 168.400 ;
        RECT 143.600 163.600 144.400 164.400 ;
        RECT 150.000 163.600 150.800 164.400 ;
        RECT 142.000 159.600 142.800 160.400 ;
        RECT 132.400 157.600 133.200 158.400 ;
        RECT 137.200 157.600 138.000 158.400 ;
        RECT 138.800 157.600 139.600 158.400 ;
        RECT 132.500 152.400 133.100 157.600 ;
        RECT 134.000 155.600 134.800 156.400 ;
        RECT 132.400 151.600 133.200 152.400 ;
        RECT 124.400 149.600 125.200 150.400 ;
        RECT 127.600 149.600 128.400 150.400 ;
        RECT 130.800 149.600 131.600 150.400 ;
        RECT 127.600 147.600 128.400 148.400 ;
        RECT 127.700 142.400 128.300 147.600 ;
        RECT 129.200 145.600 130.000 146.400 ;
        RECT 127.600 141.600 128.400 142.400 ;
        RECT 126.000 131.600 126.800 132.400 ;
        RECT 124.400 127.600 125.200 128.400 ;
        RECT 122.800 117.600 123.600 118.400 ;
        RECT 124.500 114.400 125.100 127.600 ;
        RECT 126.000 123.600 126.800 124.400 ;
        RECT 126.100 118.400 126.700 123.600 ;
        RECT 126.000 117.600 126.800 118.400 ;
        RECT 121.200 113.600 122.000 114.400 ;
        RECT 124.400 113.600 125.200 114.400 ;
        RECT 121.200 111.600 122.000 112.400 ;
        RECT 127.600 111.600 128.400 112.400 ;
        RECT 114.800 109.600 115.600 110.400 ;
        RECT 118.000 109.600 118.800 110.400 ;
        RECT 124.400 109.600 125.200 110.400 ;
        RECT 124.500 108.400 125.100 109.600 ;
        RECT 111.600 107.600 112.400 108.400 ;
        RECT 122.800 107.600 123.600 108.400 ;
        RECT 124.400 107.600 125.200 108.400 ;
        RECT 127.600 107.600 128.400 108.400 ;
        RECT 121.200 101.600 122.000 102.400 ;
        RECT 121.300 98.400 121.900 101.600 ;
        RECT 110.000 98.300 110.800 98.400 ;
        RECT 108.500 97.700 110.800 98.300 ;
        RECT 110.000 97.600 110.800 97.700 ;
        RECT 121.200 97.600 122.000 98.400 ;
        RECT 110.100 92.400 110.700 97.600 ;
        RECT 118.000 95.600 118.800 96.400 ;
        RECT 111.600 93.600 112.400 94.400 ;
        RECT 102.000 91.600 102.800 92.400 ;
        RECT 103.600 91.600 104.400 92.400 ;
        RECT 110.000 91.600 110.800 92.400 ;
        RECT 100.400 89.600 101.200 90.400 ;
        RECT 103.700 88.400 104.300 91.600 ;
        RECT 111.700 90.400 112.300 93.600 ;
        RECT 118.100 92.400 118.700 95.600 ;
        RECT 118.000 91.600 118.800 92.400 ;
        RECT 122.900 90.400 123.500 107.600 ;
        RECT 126.000 103.600 126.800 104.400 ;
        RECT 126.100 92.400 126.700 103.600 ;
        RECT 127.700 100.400 128.300 107.600 ;
        RECT 127.600 99.600 128.400 100.400 ;
        RECT 126.000 91.600 126.800 92.400 ;
        RECT 111.600 89.600 112.400 90.400 ;
        RECT 122.800 89.600 123.600 90.400 ;
        RECT 92.400 87.600 93.200 88.400 ;
        RECT 97.200 87.600 98.000 88.400 ;
        RECT 103.600 87.600 104.400 88.400 ;
        RECT 90.800 83.600 91.600 84.400 ;
        RECT 87.600 81.600 88.400 82.400 ;
        RECT 86.000 77.600 86.800 78.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 66.800 69.600 67.600 70.400 ;
        RECT 63.600 67.600 64.400 68.400 ;
        RECT 62.000 63.600 62.800 64.400 ;
        RECT 58.800 59.600 59.600 60.400 ;
        RECT 62.100 52.400 62.700 63.600 ;
        RECT 63.700 54.400 64.300 67.600 ;
        RECT 65.300 62.400 65.900 69.600 ;
        RECT 66.900 64.400 67.500 69.600 ;
        RECT 68.400 66.200 69.200 71.800 ;
        RECT 70.000 67.600 70.800 68.400 ;
        RECT 66.800 63.600 67.600 64.400 ;
        RECT 65.200 61.600 66.000 62.400 ;
        RECT 63.600 53.600 64.400 54.400 ;
        RECT 60.400 51.600 61.200 52.400 ;
        RECT 62.000 51.600 62.800 52.400 ;
        RECT 57.200 49.600 58.000 50.400 ;
        RECT 65.200 50.200 66.000 55.800 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 66.900 38.400 67.500 53.600 ;
        RECT 68.400 46.200 69.200 57.800 ;
        RECT 70.100 56.400 70.700 67.600 ;
        RECT 71.600 64.200 72.400 75.800 ;
        RECT 73.200 71.600 74.000 72.400 ;
        RECT 73.300 70.200 73.900 71.600 ;
        RECT 73.200 69.400 74.000 70.200 ;
        RECT 81.200 64.200 82.000 75.800 ;
        RECT 86.000 75.600 86.800 76.400 ;
        RECT 82.800 61.600 83.600 62.400 ;
        RECT 82.900 58.400 83.500 61.600 ;
        RECT 86.100 58.400 86.700 75.600 ;
        RECT 90.900 68.400 91.500 83.600 ;
        RECT 90.800 67.600 91.600 68.400 ;
        RECT 87.600 65.600 88.400 66.400 ;
        RECT 87.700 62.400 88.300 65.600 ;
        RECT 89.200 63.600 90.000 64.400 ;
        RECT 89.300 62.400 89.900 63.600 ;
        RECT 87.600 61.600 88.400 62.400 ;
        RECT 89.200 61.600 90.000 62.400 ;
        RECT 70.000 55.600 70.800 56.400 ;
        RECT 70.000 51.600 70.800 52.600 ;
        RECT 78.000 46.200 78.800 57.800 ;
        RECT 82.800 57.600 83.600 58.400 ;
        RECT 84.400 57.600 85.200 58.400 ;
        RECT 86.000 57.600 86.800 58.400 ;
        RECT 84.500 54.400 85.100 57.600 ;
        RECT 92.500 54.400 93.100 87.600 ;
        RECT 129.300 86.400 129.900 145.600 ;
        RECT 130.800 136.300 131.600 136.400 ;
        RECT 132.500 136.300 133.100 151.600 ;
        RECT 134.100 150.400 134.700 155.600 ;
        RECT 142.100 150.400 142.700 159.600 ;
        RECT 134.000 149.600 134.800 150.400 ;
        RECT 140.400 149.600 141.200 150.400 ;
        RECT 142.000 149.600 142.800 150.400 ;
        RECT 146.800 149.600 147.600 150.400 ;
        RECT 148.400 149.600 149.200 150.400 ;
        RECT 138.800 147.600 139.600 148.400 ;
        RECT 138.800 137.600 139.600 138.400 ;
        RECT 138.900 136.400 139.500 137.600 ;
        RECT 130.800 135.700 133.100 136.300 ;
        RECT 130.800 135.600 131.600 135.700 ;
        RECT 138.800 135.600 139.600 136.400 ;
        RECT 134.000 131.600 134.800 132.400 ;
        RECT 132.400 129.600 133.200 130.400 ;
        RECT 132.500 126.400 133.100 129.600 ;
        RECT 134.100 126.400 134.700 131.600 ;
        RECT 135.600 127.600 136.400 128.400 ;
        RECT 132.400 125.600 133.200 126.400 ;
        RECT 134.000 125.600 134.800 126.400 ;
        RECT 134.000 123.600 134.800 124.400 ;
        RECT 134.100 112.400 134.700 123.600 ;
        RECT 134.000 111.600 134.800 112.400 ;
        RECT 130.800 109.600 131.600 110.400 ;
        RECT 130.900 98.400 131.500 109.600 ;
        RECT 134.000 105.600 134.800 106.400 ;
        RECT 130.800 97.600 131.600 98.400 ;
        RECT 134.000 93.600 134.800 94.400 ;
        RECT 135.700 92.400 136.300 127.600 ;
        RECT 137.200 109.600 138.000 110.400 ;
        RECT 138.800 109.600 139.600 110.400 ;
        RECT 137.300 104.400 137.900 109.600 ;
        RECT 140.500 108.300 141.100 149.600 ;
        RECT 146.900 148.400 147.500 149.600 ;
        RECT 146.800 147.600 147.600 148.400 ;
        RECT 148.500 146.400 149.100 149.600 ;
        RECT 150.100 148.400 150.700 163.600 ;
        RECT 154.900 160.400 155.500 167.600 ;
        RECT 154.800 159.600 155.600 160.400 ;
        RECT 161.200 159.600 162.000 160.400 ;
        RECT 159.600 153.600 160.400 154.400 ;
        RECT 156.400 151.600 157.200 152.400 ;
        RECT 151.600 149.600 152.400 150.400 ;
        RECT 154.800 149.600 155.600 150.400 ;
        RECT 154.900 148.400 155.500 149.600 ;
        RECT 150.000 147.600 150.800 148.400 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 156.500 146.400 157.100 151.600 ;
        RECT 159.700 150.400 160.300 153.600 ;
        RECT 159.600 149.600 160.400 150.400 ;
        RECT 158.000 147.600 158.800 148.400 ;
        RECT 148.400 145.600 149.200 146.400 ;
        RECT 156.400 145.600 157.200 146.400 ;
        RECT 151.600 143.600 152.400 144.400 ;
        RECT 151.700 132.400 152.300 143.600 ;
        RECT 153.200 141.600 154.000 142.400 ;
        RECT 153.300 134.400 153.900 141.600 ;
        RECT 154.800 135.600 155.600 136.400 ;
        RECT 154.900 134.400 155.500 135.600 ;
        RECT 153.200 133.600 154.000 134.400 ;
        RECT 154.800 133.600 155.600 134.400 ;
        RECT 143.600 131.600 144.400 132.400 ;
        RECT 148.400 131.600 149.200 132.400 ;
        RECT 150.000 131.600 150.800 132.400 ;
        RECT 151.600 131.600 152.400 132.400 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 142.000 123.600 142.800 124.400 ;
        RECT 142.100 110.400 142.700 123.600 ;
        RECT 143.700 120.400 144.300 131.600 ;
        RECT 146.800 129.600 147.600 130.400 ;
        RECT 148.400 129.600 149.200 130.400 ;
        RECT 146.900 128.400 147.500 129.600 ;
        RECT 146.800 127.600 147.600 128.400 ;
        RECT 148.500 124.400 149.100 129.600 ;
        RECT 148.400 123.600 149.200 124.400 ;
        RECT 143.600 119.600 144.400 120.400 ;
        RECT 150.100 112.400 150.700 131.600 ;
        RECT 158.100 130.400 158.700 147.600 ;
        RECT 159.700 144.400 160.300 149.600 ;
        RECT 161.300 148.400 161.900 159.600 ;
        RECT 162.900 156.400 163.500 173.600 ;
        RECT 162.800 155.600 163.600 156.400 ;
        RECT 161.200 147.600 162.000 148.400 ;
        RECT 159.600 143.600 160.400 144.400 ;
        RECT 161.300 142.400 161.900 147.600 ;
        RECT 162.800 146.200 163.600 151.800 ;
        RECT 164.500 148.400 165.100 187.600 ;
        RECT 166.000 184.200 166.800 195.800 ;
        RECT 169.200 189.600 170.000 190.400 ;
        RECT 169.300 182.400 169.900 189.600 ;
        RECT 170.900 186.400 171.500 215.600 ;
        RECT 172.400 206.200 173.200 217.800 ;
        RECT 174.100 214.400 174.700 223.600 ;
        RECT 178.900 222.300 179.500 251.600 ;
        RECT 180.500 240.400 181.100 251.600 ;
        RECT 185.300 242.300 185.900 279.600 ;
        RECT 190.100 278.400 190.700 297.600 ;
        RECT 199.700 294.400 200.300 299.600 ;
        RECT 202.900 294.400 203.500 307.600 ;
        RECT 215.700 304.400 216.300 309.600 ;
        RECT 217.200 307.600 218.000 308.400 ;
        RECT 226.800 307.600 227.600 308.400 ;
        RECT 204.400 303.600 205.200 304.400 ;
        RECT 215.600 303.600 216.400 304.400 ;
        RECT 217.300 300.400 217.900 307.600 ;
        RECT 226.900 304.400 227.500 307.600 ;
        RECT 218.800 303.600 219.600 304.400 ;
        RECT 226.800 303.600 227.600 304.400 ;
        RECT 217.200 299.600 218.000 300.400 ;
        RECT 199.600 293.600 200.400 294.400 ;
        RECT 202.800 293.600 203.600 294.400 ;
        RECT 201.200 291.600 202.000 292.400 ;
        RECT 196.400 289.600 197.200 290.400 ;
        RECT 201.300 284.400 201.900 291.600 ;
        RECT 204.400 289.600 205.200 290.400 ;
        RECT 201.200 283.600 202.000 284.400 ;
        RECT 204.500 282.400 205.100 289.600 ;
        RECT 214.000 284.200 214.800 297.800 ;
        RECT 215.600 284.200 216.400 297.800 ;
        RECT 217.200 286.200 218.000 297.800 ;
        RECT 218.900 296.400 219.500 303.600 ;
        RECT 222.000 301.600 222.800 302.400 ;
        RECT 218.800 295.600 219.600 296.400 ;
        RECT 218.800 293.600 219.600 294.400 ;
        RECT 218.800 291.600 219.600 292.400 ;
        RECT 218.900 290.400 219.500 291.600 ;
        RECT 218.800 289.600 219.600 290.400 ;
        RECT 220.400 286.200 221.200 297.800 ;
        RECT 222.100 296.400 222.700 301.600 ;
        RECT 222.000 295.600 222.800 296.400 ;
        RECT 223.600 286.200 224.400 297.800 ;
        RECT 223.600 283.600 224.400 284.400 ;
        RECT 225.200 284.200 226.000 297.800 ;
        RECT 226.800 284.200 227.600 297.800 ;
        RECT 228.400 284.200 229.200 297.800 ;
        RECT 204.400 281.600 205.200 282.400 ;
        RECT 223.700 278.400 224.300 283.600 ;
        RECT 230.100 278.400 230.700 313.600 ;
        RECT 238.100 312.400 238.700 333.700 ;
        RECT 239.600 331.600 240.400 332.400 ;
        RECT 241.200 324.200 242.000 337.800 ;
        RECT 242.800 324.200 243.600 337.800 ;
        RECT 244.400 324.200 245.200 337.800 ;
        RECT 246.000 326.200 246.800 337.800 ;
        RECT 247.600 335.600 248.400 336.400 ;
        RECT 247.700 320.400 248.300 335.600 ;
        RECT 249.200 326.200 250.000 337.800 ;
        RECT 250.800 333.600 251.600 334.400 ;
        RECT 252.400 326.200 253.200 337.800 ;
        RECT 254.000 324.200 254.800 337.800 ;
        RECT 255.600 324.200 256.400 337.800 ;
        RECT 257.200 329.600 258.000 330.400 ;
        RECT 244.400 319.600 245.200 320.400 ;
        RECT 247.600 319.600 248.400 320.400 ;
        RECT 238.000 311.600 238.800 312.400 ;
        RECT 244.500 310.400 245.100 319.600 ;
        RECT 242.800 309.600 243.600 310.400 ;
        RECT 244.400 309.600 245.200 310.400 ;
        RECT 241.200 307.600 242.000 308.400 ;
        RECT 242.800 307.600 243.600 308.400 ;
        RECT 246.000 307.600 246.800 308.400 ;
        RECT 241.300 306.400 241.900 307.600 ;
        RECT 241.200 305.600 242.000 306.400 ;
        RECT 242.900 304.400 243.500 307.600 ;
        RECT 246.100 306.400 246.700 307.600 ;
        RECT 246.000 305.600 246.800 306.400 ;
        RECT 231.600 303.600 232.400 304.400 ;
        RECT 242.800 303.600 243.600 304.400 ;
        RECT 190.000 277.600 190.800 278.400 ;
        RECT 190.100 270.400 190.700 277.600 ;
        RECT 190.000 269.600 190.800 270.400 ;
        RECT 199.600 264.200 200.400 277.800 ;
        RECT 201.200 264.200 202.000 277.800 ;
        RECT 202.800 264.200 203.600 277.800 ;
        RECT 204.400 264.200 205.200 275.800 ;
        RECT 206.000 265.600 206.800 266.400 ;
        RECT 207.600 264.200 208.400 275.800 ;
        RECT 209.200 267.600 210.000 268.400 ;
        RECT 209.300 258.400 209.900 267.600 ;
        RECT 210.800 264.200 211.600 275.800 ;
        RECT 212.400 264.200 213.200 277.800 ;
        RECT 214.000 264.200 214.800 277.800 ;
        RECT 223.600 277.600 224.400 278.400 ;
        RECT 230.000 277.600 230.800 278.400 ;
        RECT 231.700 270.400 232.300 303.600 ;
        RECT 247.700 302.400 248.300 319.600 ;
        RECT 252.400 313.600 253.200 314.400 ;
        RECT 257.300 310.400 257.900 329.600 ;
        RECT 278.000 324.200 278.800 337.800 ;
        RECT 279.600 324.200 280.400 337.800 ;
        RECT 281.200 326.200 282.000 337.800 ;
        RECT 282.800 333.600 283.600 334.400 ;
        RECT 284.400 326.200 285.200 337.800 ;
        RECT 286.000 335.600 286.800 336.400 ;
        RECT 282.800 321.600 283.600 322.400 ;
        RECT 270.000 319.600 270.800 320.400 ;
        RECT 257.200 309.600 258.000 310.400 ;
        RECT 262.000 304.200 262.800 317.800 ;
        RECT 263.600 304.200 264.400 317.800 ;
        RECT 265.200 304.200 266.000 315.800 ;
        RECT 266.800 309.600 267.600 310.400 ;
        RECT 266.900 308.400 267.500 309.600 ;
        RECT 266.800 307.600 267.600 308.400 ;
        RECT 268.400 304.200 269.200 315.800 ;
        RECT 270.100 306.400 270.700 319.600 ;
        RECT 270.000 305.600 270.800 306.400 ;
        RECT 270.100 302.400 270.700 305.600 ;
        RECT 271.600 304.200 272.400 315.800 ;
        RECT 273.200 304.200 274.000 317.800 ;
        RECT 274.800 304.200 275.600 317.800 ;
        RECT 276.400 304.200 277.200 317.800 ;
        RECT 247.600 301.600 248.400 302.400 ;
        RECT 270.000 301.600 270.800 302.400 ;
        RECT 274.800 301.600 275.600 302.400 ;
        RECT 247.600 297.600 248.400 298.400 ;
        RECT 241.200 293.600 242.000 294.400 ;
        RECT 244.400 293.600 245.200 294.400 ;
        RECT 247.700 290.400 248.300 297.600 ;
        RECT 250.800 295.600 251.600 296.400 ;
        RECT 238.000 289.600 238.800 290.400 ;
        RECT 247.600 289.600 248.400 290.400 ;
        RECT 252.400 289.600 253.200 290.400 ;
        RECT 233.200 273.600 234.000 274.400 ;
        RECT 218.800 269.600 219.600 270.400 ;
        RECT 223.600 269.600 224.400 270.400 ;
        RECT 231.600 269.600 232.400 270.400 ;
        RECT 186.800 257.600 187.600 258.400 ;
        RECT 186.900 252.400 187.500 257.600 ;
        RECT 186.800 251.600 187.600 252.400 ;
        RECT 193.200 244.200 194.000 257.800 ;
        RECT 194.800 244.200 195.600 257.800 ;
        RECT 196.400 246.200 197.200 257.800 ;
        RECT 198.000 253.600 198.800 254.400 ;
        RECT 199.600 246.200 200.400 257.800 ;
        RECT 201.200 255.600 202.000 256.400 ;
        RECT 201.300 250.400 201.900 255.600 ;
        RECT 201.200 249.600 202.000 250.400 ;
        RECT 202.800 246.200 203.600 257.800 ;
        RECT 204.400 244.200 205.200 257.800 ;
        RECT 206.000 244.200 206.800 257.800 ;
        RECT 207.600 244.200 208.400 257.800 ;
        RECT 209.200 257.600 210.000 258.400 ;
        RECT 217.200 257.600 218.000 258.400 ;
        RECT 218.900 252.400 219.500 269.600 ;
        RECT 220.400 261.600 221.200 262.400 ;
        RECT 220.500 256.400 221.100 261.600 ;
        RECT 223.700 258.400 224.300 269.600 ;
        RECT 228.400 265.600 229.200 266.400 ;
        RECT 225.200 261.600 226.000 262.400 ;
        RECT 225.300 258.400 225.900 261.600 ;
        RECT 228.500 258.400 229.100 265.600 ;
        RECT 230.000 263.600 230.800 264.400 ;
        RECT 230.100 262.400 230.700 263.600 ;
        RECT 230.000 261.600 230.800 262.400 ;
        RECT 223.600 257.600 224.400 258.400 ;
        RECT 225.200 257.600 226.000 258.400 ;
        RECT 228.400 257.600 229.200 258.400 ;
        RECT 220.400 255.600 221.200 256.400 ;
        RECT 226.800 253.600 227.600 254.400 ;
        RECT 209.200 251.600 210.000 252.400 ;
        RECT 218.800 251.600 219.600 252.400 ;
        RECT 222.000 243.600 222.800 244.400 ;
        RECT 183.700 241.700 185.900 242.300 ;
        RECT 180.400 239.600 181.200 240.400 ;
        RECT 183.700 230.400 184.300 241.700 ;
        RECT 185.200 239.600 186.000 240.400 ;
        RECT 185.300 230.400 185.900 239.600 ;
        RECT 183.600 229.600 184.400 230.400 ;
        RECT 185.200 229.600 186.000 230.400 ;
        RECT 180.400 223.600 181.200 224.400 ;
        RECT 178.900 221.700 181.100 222.300 ;
        RECT 174.000 213.600 174.800 214.400 ;
        RECT 175.600 206.200 176.400 217.800 ;
        RECT 177.200 204.200 178.000 217.800 ;
        RECT 178.800 204.200 179.600 217.800 ;
        RECT 180.500 196.400 181.100 221.700 ;
        RECT 183.700 216.400 184.300 229.600 ;
        RECT 188.400 223.600 189.200 224.400 ;
        RECT 198.000 224.200 198.800 237.800 ;
        RECT 199.600 224.200 200.400 237.800 ;
        RECT 201.200 224.200 202.000 237.800 ;
        RECT 202.800 224.200 203.600 235.800 ;
        RECT 204.400 225.600 205.200 226.400 ;
        RECT 188.500 222.400 189.100 223.600 ;
        RECT 188.400 221.600 189.200 222.400 ;
        RECT 183.600 215.600 184.400 216.400 ;
        RECT 183.600 213.600 184.400 214.400 ;
        RECT 190.000 213.600 190.800 214.400 ;
        RECT 183.700 212.400 184.300 213.600 ;
        RECT 190.100 212.400 190.700 213.600 ;
        RECT 183.600 211.600 184.400 212.400 ;
        RECT 190.000 211.600 190.800 212.400 ;
        RECT 196.400 204.200 197.200 217.800 ;
        RECT 198.000 204.200 198.800 217.800 ;
        RECT 199.600 206.200 200.400 217.800 ;
        RECT 201.200 213.600 202.000 214.400 ;
        RECT 202.800 206.200 203.600 217.800 ;
        RECT 204.500 216.400 205.100 225.600 ;
        RECT 206.000 224.200 206.800 235.800 ;
        RECT 207.600 229.600 208.400 230.400 ;
        RECT 207.700 228.400 208.300 229.600 ;
        RECT 207.600 227.600 208.400 228.400 ;
        RECT 209.200 224.200 210.000 235.800 ;
        RECT 210.800 224.200 211.600 237.800 ;
        RECT 212.400 224.200 213.200 237.800 ;
        RECT 217.200 235.600 218.000 236.400 ;
        RECT 217.300 230.400 217.900 235.600 ;
        RECT 222.100 230.400 222.700 243.600 ;
        RECT 226.900 238.400 227.500 253.600 ;
        RECT 233.300 252.400 233.900 273.600 ;
        RECT 238.100 270.400 238.700 289.600 ;
        RECT 242.800 285.600 243.600 286.400 ;
        RECT 242.900 284.400 243.500 285.600 ;
        RECT 242.800 283.600 243.600 284.400 ;
        RECT 242.900 280.400 243.500 283.600 ;
        RECT 242.800 279.600 243.600 280.400 ;
        RECT 247.700 278.400 248.300 289.600 ;
        RECT 266.800 284.200 267.600 297.800 ;
        RECT 268.400 284.200 269.200 297.800 ;
        RECT 270.000 286.200 270.800 297.800 ;
        RECT 271.600 293.600 272.400 294.400 ;
        RECT 273.200 286.200 274.000 297.800 ;
        RECT 274.900 296.400 275.500 301.600 ;
        RECT 274.800 295.600 275.600 296.400 ;
        RECT 274.900 278.400 275.500 295.600 ;
        RECT 276.400 286.200 277.200 297.800 ;
        RECT 278.000 284.200 278.800 297.800 ;
        RECT 279.600 284.200 280.400 297.800 ;
        RECT 281.200 284.200 282.000 297.800 ;
        RECT 282.900 292.400 283.500 321.600 ;
        RECT 286.100 320.400 286.700 335.600 ;
        RECT 287.600 326.200 288.400 337.800 ;
        RECT 289.200 324.200 290.000 337.800 ;
        RECT 290.800 324.200 291.600 337.800 ;
        RECT 292.400 324.200 293.200 337.800 ;
        RECT 294.100 332.400 294.700 373.600 ;
        RECT 297.200 351.600 298.000 352.400 ;
        RECT 298.900 348.400 299.500 375.600 ;
        RECT 300.400 365.600 301.200 366.400 ;
        RECT 297.200 347.600 298.000 348.400 ;
        RECT 298.800 347.600 299.600 348.400 ;
        RECT 297.300 346.400 297.900 347.600 ;
        RECT 297.200 345.600 298.000 346.400 ;
        RECT 294.000 331.600 294.800 332.400 ;
        RECT 294.100 322.400 294.700 331.600 ;
        RECT 298.900 324.400 299.500 347.600 ;
        RECT 298.800 323.600 299.600 324.400 ;
        RECT 290.800 321.600 291.600 322.400 ;
        RECT 294.000 321.600 294.800 322.400 ;
        RECT 286.000 319.600 286.800 320.400 ;
        RECT 290.900 318.400 291.500 321.600 ;
        RECT 290.800 317.600 291.600 318.400 ;
        RECT 295.600 317.600 296.400 318.400 ;
        RECT 300.500 316.400 301.100 365.600 ;
        RECT 302.000 363.600 302.800 364.400 ;
        RECT 303.700 352.400 304.300 383.600 ;
        RECT 305.300 376.400 305.900 393.600 ;
        RECT 306.900 376.400 307.500 415.600 ;
        RECT 308.400 413.600 309.200 414.400 ;
        RECT 308.500 384.400 309.100 413.600 ;
        RECT 311.600 409.600 312.400 410.400 ;
        RECT 311.700 408.400 312.300 409.600 ;
        RECT 311.600 407.600 312.400 408.400 ;
        RECT 313.300 406.400 313.900 425.600 ;
        RECT 313.200 405.600 314.000 406.400 ;
        RECT 314.900 396.400 315.500 425.600 ;
        RECT 316.400 415.600 317.200 416.400 ;
        RECT 318.100 400.400 318.700 429.600 ;
        RECT 324.500 428.400 325.100 467.600 ;
        RECT 330.800 463.600 331.600 464.400 ;
        RECT 330.900 458.400 331.500 463.600 ;
        RECT 330.800 457.600 331.600 458.400 ;
        RECT 330.800 453.600 331.600 454.400 ;
        RECT 332.400 453.600 333.200 454.400 ;
        RECT 332.500 452.400 333.100 453.600 ;
        RECT 327.600 451.600 328.400 452.400 ;
        RECT 329.200 451.600 330.000 452.400 ;
        RECT 332.400 451.600 333.200 452.400 ;
        RECT 326.000 449.600 326.800 450.400 ;
        RECT 326.100 446.400 326.700 449.600 ;
        RECT 327.700 448.400 328.300 451.600 ;
        RECT 327.600 447.600 328.400 448.400 ;
        RECT 326.000 445.600 326.800 446.400 ;
        RECT 329.300 444.400 329.900 451.600 ;
        RECT 332.400 450.300 333.200 450.400 ;
        RECT 330.900 449.700 333.200 450.300 ;
        RECT 329.200 443.600 330.000 444.400 ;
        RECT 330.900 438.400 331.500 449.700 ;
        RECT 332.400 449.600 333.200 449.700 ;
        RECT 330.800 437.600 331.600 438.400 ;
        RECT 330.800 435.600 331.600 436.400 ;
        RECT 327.600 433.600 328.400 434.400 ;
        RECT 327.700 432.400 328.300 433.600 ;
        RECT 327.600 431.600 328.400 432.400 ;
        RECT 324.400 427.600 325.200 428.400 ;
        RECT 319.600 425.600 320.400 426.400 ;
        RECT 321.200 425.600 322.000 426.400 ;
        RECT 319.700 418.400 320.300 425.600 ;
        RECT 322.800 423.600 323.600 424.400 ;
        RECT 321.200 421.600 322.000 422.400 ;
        RECT 319.600 417.600 320.400 418.400 ;
        RECT 321.300 416.400 321.900 421.600 ;
        RECT 322.900 418.400 323.500 423.600 ;
        RECT 322.800 417.600 323.600 418.400 ;
        RECT 321.200 415.600 322.000 416.400 ;
        RECT 322.800 409.600 323.600 410.400 ;
        RECT 322.900 408.400 323.500 409.600 ;
        RECT 322.800 407.600 323.600 408.400 ;
        RECT 318.000 399.600 318.800 400.400 ;
        RECT 321.200 399.600 322.000 400.400 ;
        RECT 318.000 397.600 318.800 398.400 ;
        RECT 314.800 395.600 315.600 396.400 ;
        RECT 313.200 391.600 314.000 392.400 ;
        RECT 314.800 391.600 315.600 392.400 ;
        RECT 313.300 388.400 313.900 391.600 ;
        RECT 314.900 390.400 315.500 391.600 ;
        RECT 314.800 389.600 315.600 390.400 ;
        RECT 318.100 388.400 318.700 397.600 ;
        RECT 319.600 395.600 320.400 396.400 ;
        RECT 319.700 388.400 320.300 395.600 ;
        RECT 321.300 390.400 321.900 399.600 ;
        RECT 324.500 392.400 325.100 427.600 ;
        RECT 326.000 425.600 326.800 426.400 ;
        RECT 326.100 414.400 326.700 425.600 ;
        RECT 327.700 416.300 328.300 431.600 ;
        RECT 329.200 427.600 330.000 428.400 ;
        RECT 329.300 426.400 329.900 427.600 ;
        RECT 329.200 425.600 330.000 426.400 ;
        RECT 330.900 418.400 331.500 435.600 ;
        RECT 332.400 431.600 333.200 432.400 ;
        RECT 332.400 427.600 333.200 428.400 ;
        RECT 330.800 417.600 331.600 418.400 ;
        RECT 329.200 416.300 330.000 416.400 ;
        RECT 332.500 416.300 333.100 427.600 ;
        RECT 334.100 416.400 334.700 483.600 ;
        RECT 346.900 482.400 347.500 483.600 ;
        RECT 346.800 481.600 347.600 482.400 ;
        RECT 359.600 481.600 360.400 482.400 ;
        RECT 343.700 473.700 349.100 474.300 ;
        RECT 335.600 471.600 336.400 472.400 ;
        RECT 335.700 470.400 336.300 471.600 ;
        RECT 343.700 470.400 344.300 473.700 ;
        RECT 346.800 471.600 347.600 472.400 ;
        RECT 346.900 470.400 347.500 471.600 ;
        RECT 348.500 470.400 349.100 473.700 ;
        RECT 353.200 471.600 354.000 472.400 ;
        RECT 358.000 471.600 358.800 472.400 ;
        RECT 353.300 470.400 353.900 471.600 ;
        RECT 335.600 469.600 336.400 470.400 ;
        RECT 338.800 469.600 339.600 470.400 ;
        RECT 343.600 469.600 344.400 470.400 ;
        RECT 346.800 469.600 347.600 470.400 ;
        RECT 348.400 469.600 349.200 470.400 ;
        RECT 353.200 469.600 354.000 470.400 ;
        RECT 335.700 468.400 336.300 469.600 ;
        RECT 335.600 467.600 336.400 468.400 ;
        RECT 338.900 464.400 339.500 469.600 ;
        RECT 346.900 468.400 347.500 469.600 ;
        RECT 343.600 467.600 344.400 468.400 ;
        RECT 346.800 467.600 347.600 468.400 ;
        RECT 346.900 466.400 347.500 467.600 ;
        RECT 340.400 465.600 341.200 466.400 ;
        RECT 346.800 465.600 347.600 466.400 ;
        RECT 353.200 465.600 354.000 466.400 ;
        RECT 335.600 463.600 336.400 464.400 ;
        RECT 338.800 463.600 339.600 464.400 ;
        RECT 335.700 456.400 336.300 463.600 ;
        RECT 340.500 458.400 341.100 465.600 ;
        RECT 343.600 463.600 344.400 464.400 ;
        RECT 350.000 463.600 350.800 464.400 ;
        RECT 340.400 457.600 341.200 458.400 ;
        RECT 335.600 455.600 336.400 456.400 ;
        RECT 338.800 455.600 339.600 456.400 ;
        RECT 338.900 454.400 339.500 455.600 ;
        RECT 343.700 454.400 344.300 463.600 ;
        RECT 350.100 462.400 350.700 463.600 ;
        RECT 350.000 461.600 350.800 462.400 ;
        RECT 350.100 460.400 350.700 461.600 ;
        RECT 350.000 459.600 350.800 460.400 ;
        RECT 348.400 457.600 349.200 458.400 ;
        RECT 345.200 455.600 346.000 456.400 ;
        RECT 338.800 453.600 339.600 454.400 ;
        RECT 343.600 453.600 344.400 454.400 ;
        RECT 335.600 451.600 336.400 452.400 ;
        RECT 342.000 451.600 342.800 452.400 ;
        RECT 335.700 444.400 336.300 451.600 ;
        RECT 342.100 444.400 342.700 451.600 ;
        RECT 335.600 443.600 336.400 444.400 ;
        RECT 342.000 443.600 342.800 444.400 ;
        RECT 340.400 441.600 341.200 442.400 ;
        RECT 340.500 432.300 341.100 441.600 ;
        RECT 342.000 437.600 342.800 438.400 ;
        RECT 342.100 434.400 342.700 437.600 ;
        RECT 342.000 433.600 342.800 434.400 ;
        RECT 340.500 431.700 342.700 432.300 ;
        RECT 337.200 430.300 338.000 430.400 ;
        RECT 335.700 429.700 338.000 430.300 ;
        RECT 335.700 426.400 336.300 429.700 ;
        RECT 337.200 429.600 338.000 429.700 ;
        RECT 340.400 429.600 341.200 430.400 ;
        RECT 337.200 427.600 338.000 428.400 ;
        RECT 337.300 426.400 337.900 427.600 ;
        RECT 335.600 425.600 336.400 426.400 ;
        RECT 337.200 425.600 338.000 426.400 ;
        RECT 340.400 421.600 341.200 422.400 ;
        RECT 340.500 418.400 341.100 421.600 ;
        RECT 340.400 417.600 341.200 418.400 ;
        RECT 327.700 415.700 330.000 416.300 ;
        RECT 329.200 415.600 330.000 415.700 ;
        RECT 330.900 415.700 333.100 416.300 ;
        RECT 326.000 413.600 326.800 414.400 ;
        RECT 327.600 413.600 328.400 414.400 ;
        RECT 326.100 412.400 326.700 413.600 ;
        RECT 327.700 412.400 328.300 413.600 ;
        RECT 326.000 411.600 326.800 412.400 ;
        RECT 327.600 411.600 328.400 412.400 ;
        RECT 326.000 393.600 326.800 394.400 ;
        RECT 326.100 392.400 326.700 393.600 ;
        RECT 324.400 391.600 325.200 392.400 ;
        RECT 326.000 391.600 326.800 392.400 ;
        RECT 321.200 389.600 322.000 390.400 ;
        RECT 313.200 387.600 314.000 388.400 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 319.600 387.600 320.400 388.400 ;
        RECT 308.400 383.600 309.200 384.400 ;
        RECT 311.600 383.600 312.400 384.400 ;
        RECT 313.200 383.600 314.000 384.400 ;
        RECT 314.800 383.600 315.600 384.400 ;
        RECT 313.300 378.400 313.900 383.600 ;
        RECT 313.200 377.600 314.000 378.400 ;
        RECT 305.200 375.600 306.000 376.400 ;
        RECT 306.800 375.600 307.600 376.400 ;
        RECT 310.000 375.600 310.800 376.400 ;
        RECT 308.400 374.300 309.200 374.400 ;
        RECT 306.900 373.700 309.200 374.300 ;
        RECT 306.900 358.400 307.500 373.700 ;
        RECT 308.400 373.600 309.200 373.700 ;
        RECT 310.100 372.400 310.700 375.600 ;
        RECT 314.900 374.300 315.500 383.600 ;
        RECT 319.700 380.400 320.300 387.600 ;
        RECT 319.600 379.600 320.400 380.400 ;
        RECT 321.300 376.400 321.900 389.600 ;
        RECT 329.200 387.600 330.000 388.400 ;
        RECT 324.400 385.600 325.200 386.400 ;
        RECT 324.400 379.600 325.200 380.400 ;
        RECT 324.500 376.400 325.100 379.600 ;
        RECT 316.400 375.600 317.200 376.400 ;
        RECT 321.200 375.600 322.000 376.400 ;
        RECT 324.400 375.600 325.200 376.400 ;
        RECT 326.000 375.600 326.800 376.400 ;
        RECT 313.300 373.700 315.500 374.300 ;
        RECT 308.400 371.600 309.200 372.400 ;
        RECT 310.000 371.600 310.800 372.400 ;
        RECT 306.800 357.600 307.600 358.400 ;
        RECT 302.000 351.600 302.800 352.400 ;
        RECT 303.600 351.600 304.400 352.400 ;
        RECT 305.200 351.600 306.000 352.400 ;
        RECT 303.700 348.400 304.300 351.600 ;
        RECT 303.600 347.600 304.400 348.400 ;
        RECT 302.000 343.600 302.800 344.400 ;
        RECT 302.100 330.300 302.700 343.600 ;
        RECT 303.600 333.600 304.400 334.400 ;
        RECT 303.600 330.300 304.400 330.400 ;
        RECT 302.100 329.700 304.400 330.300 ;
        RECT 303.600 329.600 304.400 329.700 ;
        RECT 302.000 323.600 302.800 324.400 ;
        RECT 297.200 315.600 298.000 316.400 ;
        RECT 300.400 315.600 301.200 316.400 ;
        RECT 286.000 313.600 286.800 314.400 ;
        RECT 295.600 313.600 296.400 314.400 ;
        RECT 294.000 311.600 294.800 312.400 ;
        RECT 290.800 305.600 291.600 306.400 ;
        RECT 290.900 298.400 291.500 305.600 ;
        RECT 294.100 298.400 294.700 311.600 ;
        RECT 290.800 297.600 291.600 298.400 ;
        RECT 294.000 297.600 294.800 298.400 ;
        RECT 295.700 292.400 296.300 313.600 ;
        RECT 297.300 308.400 297.900 315.600 ;
        RECT 298.800 313.600 299.600 314.400 ;
        RECT 298.900 308.400 299.500 313.600 ;
        RECT 300.400 311.600 301.200 312.400 ;
        RECT 300.400 309.600 301.200 310.400 ;
        RECT 297.200 307.600 298.000 308.400 ;
        RECT 298.800 307.600 299.600 308.400 ;
        RECT 297.200 295.600 298.000 296.400 ;
        RECT 282.800 291.600 283.600 292.400 ;
        RECT 295.600 291.600 296.400 292.400 ;
        RECT 289.200 289.600 290.000 290.400 ;
        RECT 278.000 281.600 278.800 282.400 ;
        RECT 238.000 269.600 238.800 270.400 ;
        RECT 239.600 264.200 240.400 277.800 ;
        RECT 241.200 264.200 242.000 277.800 ;
        RECT 242.800 264.200 243.600 277.800 ;
        RECT 247.600 277.600 248.400 278.400 ;
        RECT 244.400 264.200 245.200 275.800 ;
        RECT 246.000 265.600 246.800 266.400 ;
        RECT 246.100 260.400 246.700 265.600 ;
        RECT 247.600 264.200 248.400 275.800 ;
        RECT 249.200 267.600 250.000 268.400 ;
        RECT 249.300 266.400 249.900 267.600 ;
        RECT 249.200 265.600 250.000 266.400 ;
        RECT 250.800 264.200 251.600 275.800 ;
        RECT 252.400 264.200 253.200 277.800 ;
        RECT 254.000 264.200 254.800 277.800 ;
        RECT 274.800 277.600 275.600 278.400 ;
        RECT 276.400 273.600 277.200 274.400 ;
        RECT 274.800 271.600 275.600 272.400 ;
        RECT 278.100 270.400 278.700 281.600 ;
        RECT 282.800 279.600 283.600 280.400 ;
        RECT 281.200 271.600 282.000 272.400 ;
        RECT 258.800 269.600 259.600 270.400 ;
        RECT 260.400 269.600 261.200 270.400 ;
        RECT 268.400 269.600 269.200 270.400 ;
        RECT 271.600 269.600 272.400 270.400 ;
        RECT 278.000 269.600 278.800 270.400 ;
        RECT 258.800 261.600 259.600 262.400 ;
        RECT 241.200 259.600 242.000 260.400 ;
        RECT 246.000 259.600 246.800 260.400 ;
        RECT 233.200 251.600 234.000 252.400 ;
        RECT 234.800 244.200 235.600 257.800 ;
        RECT 236.400 244.200 237.200 257.800 ;
        RECT 238.000 244.200 238.800 257.800 ;
        RECT 239.600 246.200 240.400 257.800 ;
        RECT 241.300 256.400 241.900 259.600 ;
        RECT 241.200 255.600 242.000 256.400 ;
        RECT 230.000 239.600 230.800 240.400 ;
        RECT 226.800 237.600 227.600 238.400 ;
        RECT 230.100 230.400 230.700 239.600 ;
        RECT 239.600 235.600 240.400 236.400 ;
        RECT 231.600 231.600 232.400 232.400 ;
        RECT 236.400 231.600 237.200 232.400 ;
        RECT 217.200 229.600 218.000 230.400 ;
        RECT 222.000 229.600 222.800 230.400 ;
        RECT 228.400 229.600 229.200 230.400 ;
        RECT 230.000 229.600 230.800 230.400 ;
        RECT 228.500 228.400 229.100 229.600 ;
        RECT 228.400 227.600 229.200 228.400 ;
        RECT 231.700 218.400 232.300 231.600 ;
        RECT 233.200 229.600 234.000 230.400 ;
        RECT 234.800 229.600 235.600 230.400 ;
        RECT 233.200 227.600 234.000 228.400 ;
        RECT 204.400 215.600 205.200 216.400 ;
        RECT 206.000 206.200 206.800 217.800 ;
        RECT 207.600 204.200 208.400 217.800 ;
        RECT 209.200 204.200 210.000 217.800 ;
        RECT 210.800 204.200 211.600 217.800 ;
        RECT 231.600 217.600 232.400 218.400 ;
        RECT 215.600 215.600 216.400 216.400 ;
        RECT 212.400 211.600 213.200 212.400 ;
        RECT 212.500 202.300 213.100 211.600 ;
        RECT 210.900 201.700 213.100 202.300 ;
        RECT 170.800 185.600 171.600 186.400 ;
        RECT 175.600 184.200 176.400 195.800 ;
        RECT 180.400 195.600 181.200 196.400 ;
        RECT 180.400 183.600 181.200 184.400 ;
        RECT 183.600 183.600 184.400 184.400 ;
        RECT 193.200 184.200 194.000 197.800 ;
        RECT 194.800 184.200 195.600 197.800 ;
        RECT 196.400 184.200 197.200 197.800 ;
        RECT 198.000 184.200 198.800 195.800 ;
        RECT 199.600 185.600 200.400 186.400 ;
        RECT 201.200 184.200 202.000 195.800 ;
        RECT 202.800 187.600 203.600 188.400 ;
        RECT 202.900 186.400 203.500 187.600 ;
        RECT 202.800 185.600 203.600 186.400 ;
        RECT 204.400 184.200 205.200 195.800 ;
        RECT 206.000 184.200 206.800 197.800 ;
        RECT 207.600 184.200 208.400 197.800 ;
        RECT 209.200 197.600 210.000 198.400 ;
        RECT 169.200 181.600 170.000 182.400 ;
        RECT 166.000 175.600 166.800 176.400 ;
        RECT 169.200 175.600 170.000 176.400 ;
        RECT 166.100 174.400 166.700 175.600 ;
        RECT 166.000 173.600 166.800 174.400 ;
        RECT 166.100 160.400 166.700 173.600 ;
        RECT 169.300 172.400 169.900 175.600 ;
        RECT 177.200 173.600 178.000 174.400 ;
        RECT 167.600 171.600 168.400 172.400 ;
        RECT 169.200 171.600 170.000 172.400 ;
        RECT 174.000 171.600 174.800 172.400 ;
        RECT 174.100 168.400 174.700 171.600 ;
        RECT 174.000 167.600 174.800 168.400 ;
        RECT 166.000 159.600 166.800 160.400 ;
        RECT 164.400 147.600 165.200 148.400 ;
        RECT 162.800 143.600 163.600 144.400 ;
        RECT 166.000 144.200 166.800 155.800 ;
        RECT 170.800 155.600 171.600 156.400 ;
        RECT 167.600 149.400 168.400 150.400 ;
        RECT 161.200 141.600 162.000 142.400 ;
        RECT 159.600 137.600 160.400 138.400 ;
        RECT 162.900 136.400 163.500 143.600 ;
        RECT 167.600 141.600 168.400 142.400 ;
        RECT 167.700 138.400 168.300 141.600 ;
        RECT 167.600 137.600 168.400 138.400 ;
        RECT 162.800 135.600 163.600 136.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 162.800 131.600 163.600 132.400 ;
        RECT 158.000 129.600 158.800 130.400 ;
        RECT 159.600 129.600 160.400 130.400 ;
        RECT 148.400 111.600 149.200 112.400 ;
        RECT 150.000 111.600 150.800 112.400 ;
        RECT 142.000 109.600 142.800 110.400 ;
        RECT 143.600 109.600 144.400 110.400 ;
        RECT 146.800 109.600 147.600 110.400 ;
        RECT 140.500 107.700 142.700 108.300 ;
        RECT 137.200 103.600 138.000 104.400 ;
        RECT 137.200 95.600 138.000 96.400 ;
        RECT 130.800 91.600 131.600 92.400 ;
        RECT 132.400 91.600 133.200 92.400 ;
        RECT 134.000 91.600 134.800 92.400 ;
        RECT 135.600 91.600 136.400 92.400 ;
        RECT 130.900 88.400 131.500 91.600 ;
        RECT 130.800 87.600 131.600 88.400 ;
        RECT 132.500 86.400 133.100 91.600 ;
        RECT 134.100 90.400 134.700 91.600 ;
        RECT 134.000 89.600 134.800 90.400 ;
        RECT 129.200 85.600 130.000 86.400 ;
        RECT 132.400 85.600 133.200 86.400 ;
        RECT 110.000 83.600 110.800 84.400 ;
        RECT 127.600 83.600 128.400 84.400 ;
        RECT 129.200 83.600 130.000 84.400 ;
        RECT 97.200 81.600 98.000 82.400 ;
        RECT 94.000 71.600 94.800 72.400 ;
        RECT 95.600 66.200 96.400 71.800 ;
        RECT 97.300 68.400 97.900 81.600 ;
        RECT 127.700 80.400 128.300 83.600 ;
        RECT 127.600 79.600 128.400 80.400 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 94.000 63.600 94.800 64.400 ;
        RECT 94.100 58.400 94.700 63.600 ;
        RECT 94.000 57.600 94.800 58.400 ;
        RECT 94.000 55.600 94.800 56.400 ;
        RECT 84.400 53.600 85.200 54.400 ;
        RECT 92.400 53.600 93.200 54.400 ;
        RECT 87.600 49.600 88.400 50.400 ;
        RECT 89.200 49.600 90.000 50.400 ;
        RECT 79.600 45.600 80.400 46.400 ;
        RECT 66.800 37.600 67.600 38.400 ;
        RECT 57.200 33.600 58.000 34.400 ;
        RECT 57.300 32.400 57.900 33.600 ;
        RECT 57.200 31.600 58.000 32.400 ;
        RECT 58.800 31.600 59.600 32.400 ;
        RECT 63.600 31.600 64.400 32.400 ;
        RECT 58.900 30.400 59.500 31.600 ;
        RECT 58.800 29.600 59.600 30.400 ;
        RECT 60.400 29.600 61.200 30.400 ;
        RECT 79.700 28.400 80.300 45.600 ;
        RECT 52.400 27.600 53.200 28.400 ;
        RECT 58.800 27.600 59.600 28.400 ;
        RECT 65.200 27.600 66.000 28.400 ;
        RECT 79.600 27.600 80.400 28.400 ;
        RECT 63.600 23.600 64.400 24.400 ;
        RECT 63.700 20.400 64.300 23.600 ;
        RECT 63.600 19.600 64.400 20.400 ;
        RECT 44.400 13.600 45.200 14.400 ;
        RECT 50.800 13.600 51.600 14.400 ;
        RECT 44.500 12.400 45.100 13.600 ;
        RECT 28.400 11.600 29.200 12.400 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 57.200 11.600 58.000 12.400 ;
        RECT 58.800 4.200 59.600 17.800 ;
        RECT 60.400 4.200 61.200 17.800 ;
        RECT 62.000 4.200 62.800 17.800 ;
        RECT 63.600 6.200 64.400 17.800 ;
        RECT 65.300 16.400 65.900 27.600 ;
        RECT 68.400 19.600 69.200 20.400 ;
        RECT 65.200 15.600 66.000 16.400 ;
        RECT 66.800 6.200 67.600 17.800 ;
        RECT 68.500 14.400 69.100 19.600 ;
        RECT 68.400 13.600 69.200 14.400 ;
        RECT 70.000 6.200 70.800 17.800 ;
        RECT 71.600 4.200 72.400 17.800 ;
        RECT 73.200 4.200 74.000 17.800 ;
        RECT 89.300 14.400 89.900 49.600 ;
        RECT 90.800 43.600 91.600 44.400 ;
        RECT 90.800 41.600 91.600 42.400 ;
        RECT 90.900 38.400 91.500 41.600 ;
        RECT 90.800 37.600 91.600 38.400 ;
        RECT 92.500 28.400 93.100 53.600 ;
        RECT 94.100 52.400 94.700 55.600 ;
        RECT 94.000 51.600 94.800 52.400 ;
        RECT 95.600 51.600 96.400 52.400 ;
        RECT 94.100 50.400 94.700 51.600 ;
        RECT 94.000 49.600 94.800 50.400 ;
        RECT 94.000 43.600 94.800 44.400 ;
        RECT 94.100 32.400 94.700 43.600 ;
        RECT 97.300 42.400 97.900 67.600 ;
        RECT 98.800 64.200 99.600 75.800 ;
        RECT 102.000 69.600 102.800 70.400 ;
        RECT 106.800 67.600 107.600 68.400 ;
        RECT 106.900 58.400 107.500 67.600 ;
        RECT 108.400 64.200 109.200 75.800 ;
        RECT 119.600 71.600 120.400 72.400 ;
        RECT 130.800 71.600 131.600 72.400 ;
        RECT 132.400 71.600 133.200 72.400 ;
        RECT 114.800 69.600 115.600 70.400 ;
        RECT 113.200 65.600 114.000 66.400 ;
        RECT 113.300 64.400 113.900 65.600 ;
        RECT 119.700 64.400 120.300 71.600 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 127.600 69.600 128.400 70.400 ;
        RECT 122.900 68.400 123.500 69.600 ;
        RECT 122.800 67.600 123.600 68.400 ;
        RECT 124.400 67.600 125.200 68.400 ;
        RECT 126.000 67.600 126.800 68.400 ;
        RECT 111.600 63.600 112.400 64.400 ;
        RECT 113.200 63.600 114.000 64.400 ;
        RECT 119.600 63.600 120.400 64.400 ;
        RECT 122.800 63.600 123.600 64.400 ;
        RECT 110.000 59.600 110.800 60.400 ;
        RECT 106.800 57.600 107.600 58.400 ;
        RECT 110.100 52.400 110.700 59.600 ;
        RECT 111.700 52.400 112.300 63.600 ;
        RECT 113.300 60.400 113.900 63.600 ;
        RECT 113.200 59.600 114.000 60.400 ;
        RECT 113.300 56.400 113.900 59.600 ;
        RECT 122.900 58.400 123.500 63.600 ;
        RECT 122.800 57.600 123.600 58.400 ;
        RECT 113.200 55.600 114.000 56.400 ;
        RECT 122.800 55.600 123.600 56.400 ;
        RECT 118.000 53.600 118.800 54.400 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 105.200 51.600 106.000 52.400 ;
        RECT 110.000 51.600 110.800 52.400 ;
        RECT 111.600 51.600 112.400 52.400 ;
        RECT 118.000 51.600 118.800 52.400 ;
        RECT 119.600 51.600 120.400 52.400 ;
        RECT 98.800 43.600 99.600 44.400 ;
        RECT 97.200 41.600 98.000 42.400 ;
        RECT 94.000 31.600 94.800 32.400 ;
        RECT 98.900 30.400 99.500 43.600 ;
        RECT 100.500 38.400 101.100 51.600 ;
        RECT 118.100 42.400 118.700 51.600 ;
        RECT 118.000 41.600 118.800 42.400 ;
        RECT 100.400 37.600 101.200 38.400 ;
        RECT 100.500 32.400 101.100 37.600 ;
        RECT 103.600 35.600 104.400 36.400 ;
        RECT 106.800 35.600 107.600 36.400 ;
        RECT 103.600 33.600 104.400 34.400 ;
        RECT 100.400 31.600 101.200 32.400 ;
        RECT 103.700 30.400 104.300 33.600 ;
        RECT 106.900 32.400 107.500 35.600 ;
        RECT 119.700 34.400 120.300 51.600 ;
        RECT 122.900 50.400 123.500 55.600 ;
        RECT 124.500 54.400 125.100 67.600 ;
        RECT 126.100 62.400 126.700 67.600 ;
        RECT 126.000 61.600 126.800 62.400 ;
        RECT 130.900 58.400 131.500 71.600 ;
        RECT 132.500 68.400 133.100 71.600 ;
        RECT 132.400 67.600 133.200 68.400 ;
        RECT 132.400 65.600 133.200 66.400 ;
        RECT 130.800 57.600 131.600 58.400 ;
        RECT 126.000 55.600 126.800 56.400 ;
        RECT 124.400 53.600 125.200 54.400 ;
        RECT 122.800 49.600 123.600 50.400 ;
        RECT 124.500 50.300 125.100 53.600 ;
        RECT 126.100 52.400 126.700 55.600 ;
        RECT 130.800 53.600 131.600 54.400 ;
        RECT 126.000 51.600 126.800 52.400 ;
        RECT 127.600 51.600 128.400 52.400 ;
        RECT 132.400 52.300 133.200 52.400 ;
        RECT 134.100 52.300 134.700 89.600 ;
        RECT 137.300 70.400 137.900 95.600 ;
        RECT 138.800 89.600 139.600 90.400 ;
        RECT 138.900 88.400 139.500 89.600 ;
        RECT 138.800 87.600 139.600 88.400 ;
        RECT 138.900 84.400 139.500 87.600 ;
        RECT 138.800 83.600 139.600 84.400 ;
        RECT 142.100 78.400 142.700 107.700 ;
        RECT 143.700 104.400 144.300 109.600 ;
        RECT 145.200 107.600 146.000 108.400 ;
        RECT 143.600 103.600 144.400 104.400 ;
        RECT 145.300 102.400 145.900 107.600 ;
        RECT 145.200 101.600 146.000 102.400 ;
        RECT 145.300 94.400 145.900 101.600 ;
        RECT 148.500 98.400 149.100 111.600 ;
        RECT 150.000 109.600 150.800 110.400 ;
        RECT 151.600 106.200 152.400 111.800 ;
        RECT 153.200 107.600 154.000 108.400 ;
        RECT 154.800 104.200 155.600 115.800 ;
        RECT 156.400 109.400 157.200 110.400 ;
        RECT 148.400 97.600 149.200 98.400 ;
        RECT 150.000 95.600 150.800 96.400 ;
        RECT 143.600 93.600 144.400 94.400 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 146.800 93.600 147.600 94.400 ;
        RECT 143.700 92.400 144.300 93.600 ;
        RECT 146.900 92.400 147.500 93.600 ;
        RECT 143.600 91.600 144.400 92.400 ;
        RECT 145.200 92.300 146.000 92.400 ;
        RECT 146.800 92.300 147.600 92.400 ;
        RECT 145.200 91.700 147.600 92.300 ;
        RECT 145.200 91.600 146.000 91.700 ;
        RECT 146.800 91.600 147.600 91.700 ;
        RECT 143.600 89.600 144.400 90.400 ;
        RECT 143.600 81.600 144.400 82.400 ;
        RECT 142.000 77.600 142.800 78.400 ;
        RECT 140.400 75.600 141.200 76.400 ;
        RECT 140.500 72.400 141.100 75.600 ;
        RECT 142.000 73.600 142.800 74.400 ;
        RECT 142.100 72.400 142.700 73.600 ;
        RECT 140.400 71.600 141.200 72.400 ;
        RECT 142.000 71.600 142.800 72.400 ;
        RECT 143.700 70.400 144.300 81.600 ;
        RECT 145.300 74.400 145.900 91.600 ;
        RECT 148.400 87.600 149.200 88.400 ;
        RECT 150.100 82.400 150.700 95.600 ;
        RECT 151.600 90.200 152.400 95.800 ;
        RECT 154.800 86.200 155.600 97.800 ;
        RECT 156.400 91.800 157.200 92.600 ;
        RECT 156.500 90.400 157.100 91.800 ;
        RECT 156.400 89.600 157.200 90.400 ;
        RECT 150.000 81.600 150.800 82.400 ;
        RECT 154.800 79.600 155.600 80.400 ;
        RECT 145.200 73.600 146.000 74.400 ;
        RECT 146.800 71.600 147.600 72.400 ;
        RECT 153.200 71.600 154.000 72.400 ;
        RECT 137.200 69.600 138.000 70.400 ;
        RECT 140.400 69.600 141.200 70.400 ;
        RECT 143.600 69.600 144.400 70.400 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 143.700 68.400 144.300 69.600 ;
        RECT 143.600 67.600 144.400 68.400 ;
        RECT 148.400 67.600 149.200 68.400 ;
        RECT 148.500 58.400 149.100 67.600 ;
        RECT 150.100 58.400 150.700 69.600 ;
        RECT 154.900 68.400 155.500 79.600 ;
        RECT 156.400 73.600 157.200 74.400 ;
        RECT 156.500 70.400 157.100 73.600 ;
        RECT 156.400 69.600 157.200 70.400 ;
        RECT 154.800 67.600 155.600 68.400 ;
        RECT 153.200 65.600 154.000 66.400 ;
        RECT 148.400 57.600 149.200 58.400 ;
        RECT 150.000 57.600 150.800 58.400 ;
        RECT 140.400 55.600 141.200 56.400 ;
        RECT 146.800 55.600 147.600 56.400 ;
        RECT 132.400 51.700 134.700 52.300 ;
        RECT 132.400 51.600 133.200 51.700 ;
        RECT 124.500 49.700 126.700 50.300 ;
        RECT 119.600 33.600 120.400 34.400 ;
        RECT 106.800 31.600 107.600 32.400 ;
        RECT 110.000 31.600 110.800 32.400 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 98.800 29.600 99.600 30.400 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 110.000 29.600 110.800 30.400 ;
        RECT 92.400 27.600 93.200 28.400 ;
        RECT 97.300 26.400 97.900 29.600 ;
        RECT 98.800 27.600 99.600 28.400 ;
        RECT 105.200 27.600 106.000 28.400 ;
        RECT 111.600 27.600 112.400 28.400 ;
        RECT 111.700 26.400 112.300 27.600 ;
        RECT 97.200 25.600 98.000 26.400 ;
        RECT 111.600 25.600 112.400 26.400 ;
        RECT 118.000 26.200 118.800 31.800 ;
        RECT 90.800 23.600 91.600 24.400 ;
        RECT 94.000 23.600 94.800 24.400 ;
        RECT 121.200 24.200 122.000 35.800 ;
        RECT 122.800 31.600 123.600 32.400 ;
        RECT 122.900 30.200 123.500 31.600 ;
        RECT 122.800 29.400 123.600 30.200 ;
        RECT 124.400 27.600 125.200 28.400 ;
        RECT 90.900 16.400 91.500 23.600 ;
        RECT 94.100 20.400 94.700 23.600 ;
        RECT 94.000 19.600 94.800 20.400 ;
        RECT 103.600 19.600 104.400 20.400 ;
        RECT 90.800 15.600 91.600 16.400 ;
        RECT 84.200 13.600 85.200 14.400 ;
        RECT 89.200 13.600 90.000 14.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 92.400 11.600 93.200 12.400 ;
        RECT 94.000 4.200 94.800 17.800 ;
        RECT 95.600 4.200 96.400 17.800 ;
        RECT 97.200 4.200 98.000 17.800 ;
        RECT 98.800 6.200 99.600 17.800 ;
        RECT 100.400 15.600 101.200 16.400 ;
        RECT 102.000 6.200 102.800 17.800 ;
        RECT 103.700 14.400 104.300 19.600 ;
        RECT 103.600 13.600 104.400 14.400 ;
        RECT 105.200 6.200 106.000 17.800 ;
        RECT 106.800 4.200 107.600 17.800 ;
        RECT 108.400 4.200 109.200 17.800 ;
        RECT 124.500 16.400 125.100 27.600 ;
        RECT 126.100 26.400 126.700 49.700 ;
        RECT 126.000 25.600 126.800 26.400 ;
        RECT 111.600 11.600 112.400 12.400 ;
        RECT 111.700 10.400 112.300 11.600 ;
        RECT 111.600 9.600 112.400 10.400 ;
        RECT 122.800 10.200 123.600 15.800 ;
        RECT 124.400 15.600 125.200 16.400 ;
        RECT 124.500 14.400 125.100 15.600 ;
        RECT 124.400 13.600 125.200 14.400 ;
        RECT 126.000 6.200 126.800 17.800 ;
        RECT 127.700 12.600 128.300 51.600 ;
        RECT 129.200 49.600 130.000 50.400 ;
        RECT 129.300 48.400 129.900 49.600 ;
        RECT 129.200 47.600 130.000 48.400 ;
        RECT 132.400 47.600 133.200 48.400 ;
        RECT 130.800 24.200 131.600 35.800 ;
        RECT 134.100 30.400 134.700 51.700 ;
        RECT 137.200 51.600 138.000 52.400 ;
        RECT 138.800 51.600 139.600 52.400 ;
        RECT 143.600 51.600 144.400 52.400 ;
        RECT 137.300 50.400 137.900 51.600 ;
        RECT 135.600 49.600 136.400 50.400 ;
        RECT 137.200 49.600 138.000 50.400 ;
        RECT 135.700 48.400 136.300 49.600 ;
        RECT 143.700 48.400 144.300 51.600 ;
        RECT 145.200 49.600 146.000 50.400 ;
        RECT 135.600 47.600 136.400 48.400 ;
        RECT 140.400 47.600 141.200 48.400 ;
        RECT 143.600 47.600 144.400 48.400 ;
        RECT 135.600 37.600 136.400 38.400 ;
        RECT 134.000 29.600 134.800 30.400 ;
        RECT 137.200 29.600 138.000 30.400 ;
        RECT 137.200 27.600 138.000 28.400 ;
        RECT 140.500 18.400 141.100 47.600 ;
        RECT 145.300 38.400 145.900 49.600 ;
        RECT 146.900 38.400 147.500 55.600 ;
        RECT 158.100 52.400 158.700 129.600 ;
        RECT 159.700 128.400 160.300 129.600 ;
        RECT 159.600 127.600 160.400 128.400 ;
        RECT 159.700 72.400 160.300 127.600 ;
        RECT 162.900 116.400 163.500 131.600 ;
        RECT 169.200 123.600 170.000 124.400 ;
        RECT 169.300 118.400 169.900 123.600 ;
        RECT 167.600 117.600 168.400 118.400 ;
        RECT 169.200 117.600 170.000 118.400 ;
        RECT 162.800 115.600 163.600 116.400 ;
        RECT 164.400 104.200 165.200 115.800 ;
        RECT 162.800 91.600 163.600 92.400 ;
        RECT 164.400 86.200 165.200 97.800 ;
        RECT 162.800 79.600 163.600 80.400 ;
        RECT 162.900 78.400 163.500 79.600 ;
        RECT 162.800 77.600 163.600 78.400 ;
        RECT 159.600 71.600 160.400 72.400 ;
        RECT 166.000 71.600 166.800 72.400 ;
        RECT 167.700 70.400 168.300 117.600 ;
        RECT 169.200 83.600 170.000 84.400 ;
        RECT 169.200 73.600 170.000 74.400 ;
        RECT 170.900 70.400 171.500 155.600 ;
        RECT 174.100 150.400 174.700 167.600 ;
        RECT 177.300 164.400 177.900 173.600 ;
        RECT 180.500 170.400 181.100 183.600 ;
        RECT 188.400 181.600 189.200 182.400 ;
        RECT 206.000 181.600 206.800 182.400 ;
        RECT 188.500 178.400 189.100 181.600 ;
        RECT 188.400 177.600 189.200 178.400 ;
        RECT 206.100 176.400 206.700 181.600 ;
        RECT 209.300 176.400 209.900 197.600 ;
        RECT 210.900 192.400 211.500 201.700 ;
        RECT 210.800 191.600 211.600 192.400 ;
        RECT 210.900 190.400 211.500 191.600 ;
        RECT 210.800 189.600 211.600 190.400 ;
        RECT 214.000 189.600 214.800 190.400 ;
        RECT 212.400 185.600 213.200 186.400 ;
        RECT 212.500 178.400 213.100 185.600 ;
        RECT 212.400 177.600 213.200 178.400 ;
        RECT 198.000 175.600 198.800 176.400 ;
        RECT 206.000 175.600 206.800 176.400 ;
        RECT 209.200 175.600 210.000 176.400 ;
        RECT 183.600 173.600 184.400 174.400 ;
        RECT 194.800 173.600 195.600 174.400 ;
        RECT 178.800 169.600 179.600 170.400 ;
        RECT 180.400 169.600 181.200 170.400 ;
        RECT 182.000 169.600 182.800 170.400 ;
        RECT 182.100 168.400 182.700 169.600 ;
        RECT 182.000 167.600 182.800 168.400 ;
        RECT 183.700 164.400 184.300 173.600 ;
        RECT 185.200 171.600 186.000 172.400 ;
        RECT 188.400 171.600 189.200 172.400 ;
        RECT 194.800 171.600 195.600 172.400 ;
        RECT 186.800 169.600 187.600 170.400 ;
        RECT 177.200 163.600 178.000 164.400 ;
        RECT 183.600 163.600 184.400 164.400 ;
        RECT 174.000 149.600 174.800 150.400 ;
        RECT 175.600 144.200 176.400 155.800 ;
        RECT 182.000 153.600 182.800 154.400 ;
        RECT 182.100 146.400 182.700 153.600 ;
        RECT 186.900 150.400 187.500 169.600 ;
        RECT 188.500 158.400 189.100 171.600 ;
        RECT 190.000 169.600 190.800 170.400 ;
        RECT 188.400 157.600 189.200 158.400 ;
        RECT 193.200 155.600 194.000 156.400 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 186.800 149.600 187.600 150.400 ;
        RECT 191.600 149.600 192.400 150.400 ;
        RECT 185.300 148.400 185.900 149.600 ;
        RECT 185.200 147.600 186.000 148.400 ;
        RECT 182.000 145.600 182.800 146.400 ;
        RECT 183.600 143.600 184.400 144.400 ;
        RECT 175.600 139.600 176.400 140.400 ;
        RECT 172.400 133.600 173.200 134.400 ;
        RECT 172.500 130.400 173.100 133.600 ;
        RECT 174.000 131.600 174.800 132.400 ;
        RECT 172.400 129.600 173.200 130.400 ;
        RECT 172.400 127.600 173.200 128.400 ;
        RECT 172.500 108.400 173.100 127.600 ;
        RECT 174.100 126.400 174.700 131.600 ;
        RECT 175.700 130.400 176.300 139.600 ;
        RECT 183.700 134.400 184.300 143.600 ;
        RECT 186.900 140.400 187.500 149.600 ;
        RECT 186.800 139.600 187.600 140.400 ;
        RECT 186.800 135.600 187.600 136.400 ;
        RECT 186.900 134.400 187.500 135.600 ;
        RECT 193.300 134.400 193.900 155.600 ;
        RECT 194.900 154.400 195.500 171.600 ;
        RECT 198.100 170.400 198.700 175.600 ;
        RECT 214.100 174.400 214.700 189.600 ;
        RECT 204.400 173.600 205.200 174.400 ;
        RECT 209.200 173.600 210.000 174.400 ;
        RECT 214.000 173.600 214.800 174.400 ;
        RECT 198.000 169.600 198.800 170.400 ;
        RECT 202.800 167.600 203.600 168.400 ;
        RECT 196.400 163.600 197.200 164.400 ;
        RECT 196.500 156.400 197.100 163.600 ;
        RECT 196.400 155.600 197.200 156.400 ;
        RECT 194.800 153.600 195.600 154.400 ;
        RECT 201.200 151.600 202.000 152.400 ;
        RECT 201.300 150.400 201.900 151.600 ;
        RECT 194.800 149.600 195.600 150.400 ;
        RECT 196.400 149.600 197.200 150.400 ;
        RECT 201.200 149.600 202.000 150.400 ;
        RECT 194.900 142.400 195.500 149.600 ;
        RECT 194.800 141.600 195.600 142.400 ;
        RECT 196.500 136.400 197.100 149.600 ;
        RECT 204.500 148.400 205.100 173.600 ;
        RECT 209.300 172.400 209.900 173.600 ;
        RECT 215.700 172.400 216.300 215.600 ;
        RECT 226.800 213.600 227.600 214.400 ;
        RECT 231.600 213.600 232.400 214.400 ;
        RECT 233.300 212.400 233.900 227.600 ;
        RECT 234.900 224.400 235.500 229.600 ;
        RECT 236.500 228.400 237.100 231.600 ;
        RECT 239.700 230.400 240.300 235.600 ;
        RECT 239.600 229.600 240.400 230.400 ;
        RECT 236.400 227.600 237.200 228.400 ;
        RECT 234.800 223.600 235.600 224.400 ;
        RECT 234.800 221.600 235.600 222.400 ;
        RECT 234.900 214.400 235.500 221.600 ;
        RECT 236.500 220.400 237.100 227.600 ;
        RECT 241.300 226.400 241.900 255.600 ;
        RECT 242.800 246.200 243.600 257.800 ;
        RECT 244.400 253.600 245.200 254.400 ;
        RECT 244.400 251.600 245.200 252.400 ;
        RECT 244.500 244.300 245.100 251.600 ;
        RECT 246.000 246.200 246.800 257.800 ;
        RECT 242.900 243.700 245.100 244.300 ;
        RECT 247.600 244.200 248.400 257.800 ;
        RECT 249.200 244.200 250.000 257.800 ;
        RECT 258.900 256.400 259.500 261.600 ;
        RECT 258.800 255.600 259.600 256.400 ;
        RECT 242.900 234.400 243.500 243.700 ;
        RECT 260.500 240.300 261.100 269.600 ;
        RECT 268.500 268.400 269.100 269.600 ;
        RECT 271.700 268.400 272.300 269.600 ;
        RECT 268.400 267.600 269.200 268.400 ;
        RECT 271.600 267.600 272.400 268.400 ;
        RECT 270.000 265.600 270.800 266.400 ;
        RECT 270.100 254.400 270.700 265.600 ;
        RECT 274.800 257.600 275.600 258.400 ;
        RECT 270.000 253.600 270.800 254.400 ;
        RECT 268.400 251.600 269.200 252.400 ;
        RECT 268.500 244.400 269.100 251.600 ;
        RECT 271.600 249.600 272.400 250.400 ;
        RECT 268.400 243.600 269.200 244.400 ;
        RECT 271.700 240.400 272.300 249.600 ;
        RECT 260.500 239.700 262.700 240.300 ;
        RECT 242.800 233.600 243.600 234.400 ;
        RECT 242.900 228.300 243.500 233.600 ;
        RECT 242.900 227.700 245.100 228.300 ;
        RECT 241.200 225.600 242.000 226.400 ;
        RECT 242.800 223.600 243.600 224.400 ;
        RECT 236.400 219.600 237.200 220.400 ;
        RECT 239.600 219.600 240.400 220.400 ;
        RECT 236.400 217.600 237.200 218.400 ;
        RECT 239.700 216.400 240.300 219.600 ;
        RECT 239.600 215.600 240.400 216.400 ;
        RECT 234.800 213.600 235.600 214.400 ;
        RECT 238.000 213.600 238.800 214.400 ;
        RECT 242.900 212.400 243.500 223.600 ;
        RECT 244.500 214.400 245.100 227.700 ;
        RECT 246.000 224.200 246.800 237.800 ;
        RECT 247.600 224.200 248.400 237.800 ;
        RECT 249.200 224.200 250.000 235.800 ;
        RECT 250.800 227.600 251.600 228.400 ;
        RECT 250.900 218.400 251.500 227.600 ;
        RECT 252.400 224.200 253.200 235.800 ;
        RECT 254.000 225.600 254.800 226.400 ;
        RECT 250.800 217.600 251.600 218.400 ;
        RECT 244.400 213.600 245.200 214.400 ;
        RECT 226.800 212.300 227.600 212.400 ;
        RECT 225.300 211.700 227.600 212.300 ;
        RECT 220.400 204.300 221.200 204.400 ;
        RECT 218.900 203.700 221.200 204.300 ;
        RECT 217.200 189.600 218.000 190.400 ;
        RECT 217.200 179.600 218.000 180.400 ;
        RECT 217.300 178.400 217.900 179.600 ;
        RECT 217.200 177.600 218.000 178.400 ;
        RECT 218.900 176.400 219.500 203.700 ;
        RECT 220.400 203.600 221.200 203.700 ;
        RECT 225.300 190.400 225.900 211.700 ;
        RECT 226.800 211.600 227.600 211.700 ;
        RECT 233.200 211.600 234.000 212.400 ;
        RECT 242.800 211.600 243.600 212.400 ;
        RECT 249.200 211.600 250.000 212.400 ;
        RECT 238.000 209.600 238.800 210.400 ;
        RECT 254.100 208.400 254.700 225.600 ;
        RECT 255.600 224.200 256.400 235.800 ;
        RECT 257.200 224.200 258.000 237.800 ;
        RECT 258.800 224.200 259.600 237.800 ;
        RECT 260.400 224.200 261.200 237.800 ;
        RECT 262.100 230.400 262.700 239.700 ;
        RECT 271.600 239.600 272.400 240.400 ;
        RECT 262.000 229.600 262.800 230.400 ;
        RECT 270.000 229.600 271.000 230.400 ;
        RECT 282.900 226.400 283.500 279.600 ;
        RECT 289.300 278.400 289.900 289.600 ;
        RECT 297.300 288.400 297.900 295.600 ;
        RECT 300.400 292.300 301.200 292.400 ;
        RECT 302.100 292.300 302.700 323.600 ;
        RECT 303.600 312.300 304.400 312.400 ;
        RECT 305.300 312.300 305.900 351.600 ;
        RECT 306.800 350.300 307.600 350.400 ;
        RECT 308.500 350.300 309.100 371.600 ;
        RECT 313.300 370.400 313.900 373.700 ;
        RECT 316.400 373.600 317.200 374.400 ;
        RECT 319.600 373.600 320.400 374.400 ;
        RECT 324.400 373.600 325.200 374.400 ;
        RECT 314.800 371.600 315.600 372.400 ;
        RECT 313.200 369.600 314.000 370.400 ;
        RECT 314.900 368.300 315.500 371.600 ;
        RECT 316.500 368.400 317.100 373.600 ;
        RECT 326.000 371.600 326.800 372.400 ;
        RECT 329.200 371.600 330.000 372.400 ;
        RECT 319.600 369.600 320.400 370.400 ;
        RECT 313.300 367.700 315.500 368.300 ;
        RECT 310.000 359.600 310.800 360.400 ;
        RECT 306.800 349.700 309.100 350.300 ;
        RECT 306.800 349.600 307.600 349.700 ;
        RECT 306.900 332.400 307.500 349.600 ;
        RECT 308.400 347.600 309.200 348.400 ;
        RECT 308.500 346.400 309.100 347.600 ;
        RECT 308.400 345.600 309.200 346.400 ;
        RECT 308.400 339.600 309.200 340.400 ;
        RECT 308.500 332.400 309.100 339.600 ;
        RECT 306.800 331.600 307.600 332.400 ;
        RECT 308.400 331.600 309.200 332.400 ;
        RECT 308.400 329.600 309.200 330.400 ;
        RECT 303.600 311.700 305.900 312.300 ;
        RECT 303.600 311.600 304.400 311.700 ;
        RECT 303.600 309.600 304.400 310.400 ;
        RECT 306.800 309.600 307.600 310.400 ;
        RECT 306.900 306.400 307.500 309.600 ;
        RECT 308.500 308.400 309.100 329.600 ;
        RECT 308.400 307.600 309.200 308.400 ;
        RECT 306.800 305.600 307.600 306.400 ;
        RECT 308.500 302.400 309.100 307.600 ;
        RECT 308.400 301.600 309.200 302.400 ;
        RECT 306.800 295.600 307.600 296.400 ;
        RECT 300.400 291.700 302.700 292.300 ;
        RECT 300.400 291.600 301.200 291.700 ;
        RECT 297.200 287.600 298.000 288.400 ;
        RECT 295.600 283.600 296.400 284.400 ;
        RECT 289.200 277.600 290.000 278.400 ;
        RECT 284.400 272.300 285.200 272.400 ;
        RECT 284.400 271.700 286.700 272.300 ;
        RECT 284.400 271.600 285.200 271.700 ;
        RECT 286.100 270.400 286.700 271.700 ;
        RECT 292.400 271.600 293.200 272.400 ;
        RECT 284.400 269.600 285.200 270.400 ;
        RECT 286.000 269.600 286.800 270.400 ;
        RECT 284.500 262.400 285.100 269.600 ;
        RECT 286.000 267.600 286.800 268.400 ;
        RECT 287.600 267.600 288.400 268.400 ;
        RECT 287.700 264.400 288.300 267.600 ;
        RECT 287.600 263.600 288.400 264.400 ;
        RECT 284.400 261.600 285.200 262.400 ;
        RECT 295.700 260.400 296.300 283.600 ;
        RECT 297.300 274.400 297.900 287.600 ;
        RECT 300.500 280.400 301.100 291.600 ;
        RECT 306.900 288.400 307.500 295.600 ;
        RECT 308.400 292.300 309.200 292.400 ;
        RECT 310.100 292.300 310.700 359.600 ;
        RECT 313.300 358.400 313.900 367.700 ;
        RECT 316.400 367.600 317.200 368.400 ;
        RECT 313.200 357.600 314.000 358.400 ;
        RECT 314.800 357.600 315.600 358.400 ;
        RECT 311.600 355.600 312.400 356.400 ;
        RECT 311.700 354.400 312.300 355.600 ;
        RECT 311.600 353.600 312.400 354.400 ;
        RECT 314.900 352.400 315.500 357.600 ;
        RECT 316.400 353.600 317.200 354.400 ;
        RECT 314.800 351.600 315.600 352.400 ;
        RECT 316.500 350.400 317.100 353.600 ;
        RECT 313.200 349.600 314.000 350.400 ;
        RECT 316.400 349.600 317.200 350.400 ;
        RECT 319.700 348.400 320.300 369.600 ;
        RECT 327.600 365.600 328.400 366.400 ;
        RECT 326.000 361.600 326.800 362.400 ;
        RECT 321.200 351.600 322.000 352.400 ;
        RECT 322.800 351.600 323.600 352.400 ;
        RECT 321.300 350.400 321.900 351.600 ;
        RECT 322.900 350.400 323.500 351.600 ;
        RECT 321.200 349.600 322.000 350.400 ;
        RECT 322.800 349.600 323.600 350.400 ;
        RECT 324.400 349.600 325.200 350.400 ;
        RECT 326.100 348.400 326.700 361.600 ;
        RECT 311.600 347.600 312.400 348.400 ;
        RECT 313.200 347.600 314.000 348.400 ;
        RECT 318.000 347.600 318.800 348.400 ;
        RECT 319.600 347.600 320.400 348.400 ;
        RECT 321.200 347.600 322.000 348.400 ;
        RECT 324.400 347.600 325.200 348.400 ;
        RECT 326.000 347.600 326.800 348.400 ;
        RECT 311.700 330.400 312.300 347.600 ;
        RECT 311.600 329.600 312.400 330.400 ;
        RECT 311.700 314.400 312.300 329.600 ;
        RECT 313.300 318.400 313.900 347.600 ;
        RECT 318.100 342.400 318.700 347.600 ;
        RECT 319.600 345.600 320.400 346.400 ;
        RECT 318.000 341.600 318.800 342.400 ;
        RECT 319.700 338.400 320.300 345.600 ;
        RECT 322.800 343.600 323.600 344.400 ;
        RECT 318.000 337.600 318.800 338.400 ;
        RECT 319.600 337.600 320.400 338.400 ;
        RECT 316.400 335.600 317.200 336.400 ;
        RECT 316.500 334.400 317.100 335.600 ;
        RECT 316.400 333.600 317.200 334.400 ;
        RECT 314.800 331.600 315.600 332.400 ;
        RECT 318.100 330.400 318.700 337.600 ;
        RECT 319.600 333.600 320.400 334.400 ;
        RECT 321.200 333.600 322.000 334.400 ;
        RECT 318.000 329.600 318.800 330.400 ;
        RECT 313.200 317.600 314.000 318.400 ;
        RECT 314.800 315.600 315.600 316.400 ;
        RECT 314.900 314.400 315.500 315.600 ;
        RECT 311.600 313.600 312.400 314.400 ;
        RECT 314.800 313.600 315.600 314.400 ;
        RECT 318.000 313.600 318.800 314.400 ;
        RECT 318.100 312.400 318.700 313.600 ;
        RECT 319.700 312.400 320.300 333.600 ;
        RECT 321.300 328.400 321.900 333.600 ;
        RECT 322.900 332.400 323.500 343.600 ;
        RECT 324.500 334.400 325.100 347.600 ;
        RECT 326.100 340.400 326.700 347.600 ;
        RECT 326.000 339.600 326.800 340.400 ;
        RECT 327.700 338.300 328.300 365.600 ;
        RECT 330.900 358.400 331.500 415.700 ;
        RECT 334.000 415.600 334.800 416.400 ;
        RECT 332.400 413.600 333.200 414.400 ;
        RECT 332.500 410.400 333.100 413.600 ;
        RECT 334.000 411.600 334.800 412.400 ;
        RECT 340.400 411.600 341.200 412.400 ;
        RECT 332.400 409.600 333.200 410.400 ;
        RECT 334.100 406.400 334.700 411.600 ;
        RECT 335.600 409.600 336.400 410.400 ;
        RECT 338.800 409.600 339.600 410.400 ;
        RECT 337.200 407.600 338.000 408.400 ;
        RECT 334.000 405.600 334.800 406.400 ;
        RECT 334.000 399.600 334.800 400.400 ;
        RECT 334.100 398.400 334.700 399.600 ;
        RECT 334.000 397.600 334.800 398.400 ;
        RECT 334.000 393.600 334.800 394.400 ;
        RECT 334.100 390.400 334.700 393.600 ;
        RECT 337.200 392.300 338.000 392.400 ;
        RECT 338.900 392.300 339.500 409.600 ;
        RECT 340.500 406.400 341.100 411.600 ;
        RECT 340.400 405.600 341.200 406.400 ;
        RECT 340.400 399.600 341.200 400.400 ;
        RECT 337.200 391.700 339.500 392.300 ;
        RECT 337.200 391.600 338.000 391.700 ;
        RECT 340.500 390.400 341.100 399.600 ;
        RECT 334.000 389.600 334.800 390.400 ;
        RECT 340.400 389.600 341.200 390.400 ;
        RECT 335.600 387.600 336.400 388.400 ;
        RECT 335.700 386.400 336.300 387.600 ;
        RECT 335.600 385.600 336.400 386.400 ;
        RECT 337.200 383.600 338.000 384.400 ;
        RECT 337.300 382.400 337.900 383.600 ;
        RECT 342.100 382.400 342.700 431.700 ;
        RECT 343.700 428.400 344.300 453.600 ;
        RECT 345.300 452.400 345.900 455.600 ;
        RECT 346.800 453.600 347.600 454.400 ;
        RECT 348.500 452.400 349.100 457.600 ;
        RECT 351.600 455.600 352.400 456.400 ;
        RECT 350.000 453.600 350.800 454.400 ;
        RECT 345.200 451.600 346.000 452.400 ;
        RECT 348.400 451.600 349.200 452.400 ;
        RECT 345.300 436.400 345.900 451.600 ;
        RECT 350.100 450.300 350.700 453.600 ;
        RECT 351.700 452.400 352.300 455.600 ;
        RECT 351.600 451.600 352.400 452.400 ;
        RECT 350.100 449.700 352.300 450.300 ;
        RECT 350.000 441.600 350.800 442.400 ;
        RECT 345.200 435.600 346.000 436.400 ;
        RECT 348.400 435.600 349.200 436.400 ;
        RECT 345.200 431.600 346.000 432.400 ;
        RECT 345.300 430.400 345.900 431.600 ;
        RECT 348.500 430.400 349.100 435.600 ;
        RECT 345.200 429.600 346.000 430.400 ;
        RECT 348.400 429.600 349.200 430.400 ;
        RECT 348.500 428.400 349.100 429.600 ;
        RECT 350.100 428.400 350.700 441.600 ;
        RECT 351.700 438.400 352.300 449.700 ;
        RECT 351.600 437.600 352.400 438.400 ;
        RECT 343.600 427.600 344.400 428.400 ;
        RECT 346.800 427.600 347.600 428.400 ;
        RECT 348.400 427.600 349.200 428.400 ;
        RECT 350.000 427.600 350.800 428.400 ;
        RECT 353.300 428.300 353.900 465.600 ;
        RECT 358.100 464.400 358.700 471.600 ;
        RECT 359.700 468.400 360.300 481.600 ;
        RECT 377.200 473.600 378.000 474.400 ;
        RECT 366.000 471.600 366.800 472.400 ;
        RECT 372.400 471.600 373.200 472.400 ;
        RECT 375.600 471.600 376.400 472.400 ;
        RECT 369.200 469.600 370.000 470.400 ;
        RECT 359.600 467.600 360.400 468.400 ;
        RECT 361.200 467.600 362.000 468.400 ;
        RECT 354.800 463.600 355.600 464.400 ;
        RECT 358.000 463.600 358.800 464.400 ;
        RECT 354.900 454.400 355.500 463.600 ;
        RECT 356.400 455.600 357.200 456.400 ;
        RECT 354.800 453.600 355.600 454.400 ;
        RECT 358.100 452.400 358.700 463.600 ;
        RECT 359.700 462.400 360.300 467.600 ;
        RECT 359.600 461.600 360.400 462.400 ;
        RECT 361.300 456.400 361.900 467.600 ;
        RECT 364.400 463.600 365.200 464.400 ;
        RECT 361.200 455.600 362.000 456.400 ;
        RECT 356.400 451.600 357.200 452.400 ;
        RECT 358.000 451.600 358.800 452.400 ;
        RECT 354.800 441.600 355.600 442.400 ;
        RECT 354.900 428.400 355.500 441.600 ;
        RECT 356.500 432.400 357.100 451.600 ;
        RECT 359.600 443.600 360.400 444.400 ;
        RECT 356.400 431.600 357.200 432.400 ;
        RECT 359.700 432.300 360.300 443.600 ;
        RECT 361.300 434.300 361.900 455.600 ;
        RECT 364.500 448.400 365.100 463.600 ;
        RECT 366.000 453.600 366.800 454.400 ;
        RECT 366.100 452.400 366.700 453.600 ;
        RECT 366.000 451.600 366.800 452.400 ;
        RECT 367.600 449.600 368.400 450.400 ;
        RECT 364.400 447.600 365.200 448.400 ;
        RECT 362.800 445.600 363.600 446.400 ;
        RECT 366.000 443.600 366.800 444.400 ;
        RECT 362.800 439.600 363.600 440.400 ;
        RECT 362.900 438.400 363.500 439.600 ;
        RECT 366.100 438.400 366.700 443.600 ;
        RECT 369.300 442.400 369.900 469.600 ;
        RECT 370.800 467.600 371.600 468.400 ;
        RECT 370.900 466.400 371.500 467.600 ;
        RECT 370.800 465.600 371.600 466.400 ;
        RECT 370.800 459.600 371.600 460.400 ;
        RECT 370.900 448.400 371.500 459.600 ;
        RECT 377.300 458.400 377.900 473.600 ;
        RECT 385.200 464.200 386.000 477.800 ;
        RECT 386.800 464.200 387.600 477.800 ;
        RECT 388.400 464.200 389.200 475.800 ;
        RECT 390.000 467.600 390.800 468.400 ;
        RECT 391.600 464.200 392.400 475.800 ;
        RECT 393.200 465.600 394.000 466.400 ;
        RECT 393.300 462.400 393.900 465.600 ;
        RECT 394.800 464.200 395.600 475.800 ;
        RECT 396.400 464.200 397.200 477.800 ;
        RECT 398.000 464.200 398.800 477.800 ;
        RECT 399.600 464.200 400.400 477.800 ;
        RECT 401.300 470.400 401.900 483.600 ;
        RECT 401.200 469.600 402.000 470.400 ;
        RECT 386.800 461.600 387.600 462.400 ;
        RECT 393.200 461.600 394.000 462.400 ;
        RECT 377.200 457.600 378.000 458.400 ;
        RECT 375.600 455.600 376.400 456.400 ;
        RECT 378.800 453.600 379.600 454.400 ;
        RECT 382.000 453.600 382.800 454.400 ;
        RECT 378.900 452.400 379.500 453.600 ;
        RECT 372.400 451.600 373.200 452.400 ;
        RECT 374.000 451.600 374.800 452.400 ;
        RECT 378.800 451.600 379.600 452.400 ;
        RECT 382.000 451.600 382.800 452.400 ;
        RECT 374.100 450.400 374.700 451.600 ;
        RECT 374.000 449.600 374.800 450.400 ;
        RECT 377.200 449.600 378.000 450.400 ;
        RECT 380.400 449.600 381.200 450.400 ;
        RECT 370.800 447.600 371.600 448.400 ;
        RECT 369.200 441.600 370.000 442.400 ;
        RECT 369.300 438.400 369.900 441.600 ;
        RECT 362.800 437.600 363.600 438.400 ;
        RECT 366.000 437.600 366.800 438.400 ;
        RECT 369.200 437.600 370.000 438.400 ;
        RECT 366.000 435.600 366.800 436.400 ;
        RECT 361.300 433.700 363.500 434.300 ;
        RECT 359.700 431.700 361.900 432.300 ;
        RECT 356.500 430.400 357.100 431.600 ;
        RECT 356.400 429.600 357.200 430.400 ;
        RECT 359.600 429.600 360.400 430.400 ;
        RECT 359.700 428.400 360.300 429.600 ;
        RECT 361.300 428.400 361.900 431.700 ;
        RECT 351.700 427.700 353.900 428.300 ;
        RECT 343.700 426.400 344.300 427.600 ;
        RECT 346.900 426.400 347.500 427.600 ;
        RECT 343.600 425.600 344.400 426.400 ;
        RECT 346.800 425.600 347.600 426.400 ;
        RECT 348.400 423.600 349.200 424.400 ;
        RECT 345.200 421.600 346.000 422.400 ;
        RECT 346.800 421.600 347.600 422.400 ;
        RECT 343.600 419.600 344.400 420.400 ;
        RECT 343.700 412.400 344.300 419.600 ;
        RECT 343.600 411.600 344.400 412.400 ;
        RECT 343.700 408.400 344.300 411.600 ;
        RECT 343.600 407.600 344.400 408.400 ;
        RECT 345.300 394.400 345.900 421.600 ;
        RECT 346.900 416.400 347.500 421.600 ;
        RECT 348.500 418.400 349.100 423.600 ;
        RECT 350.000 419.600 350.800 420.400 ;
        RECT 348.400 417.600 349.200 418.400 ;
        RECT 346.800 415.600 347.600 416.400 ;
        RECT 348.400 415.600 349.200 416.400 ;
        RECT 346.800 413.600 347.600 414.400 ;
        RECT 346.900 402.400 347.500 413.600 ;
        RECT 346.800 401.600 347.600 402.400 ;
        RECT 343.600 393.600 344.400 394.400 ;
        RECT 345.200 393.600 346.000 394.400 ;
        RECT 343.600 391.600 344.400 392.400 ;
        RECT 343.700 388.400 344.300 391.600 ;
        RECT 348.500 390.400 349.100 415.600 ;
        RECT 350.100 414.400 350.700 419.600 ;
        RECT 351.700 416.300 352.300 427.700 ;
        RECT 354.800 427.600 355.600 428.400 ;
        RECT 358.000 427.600 358.800 428.400 ;
        RECT 359.600 427.600 360.400 428.400 ;
        RECT 361.200 427.600 362.000 428.400 ;
        RECT 353.200 425.600 354.000 426.400 ;
        RECT 354.800 425.600 355.600 426.400 ;
        RECT 353.300 420.400 353.900 425.600 ;
        RECT 353.200 419.600 354.000 420.400 ;
        RECT 353.200 416.300 354.000 416.400 ;
        RECT 351.700 415.700 354.000 416.300 ;
        RECT 353.200 415.600 354.000 415.700 ;
        RECT 350.000 413.600 350.800 414.400 ;
        RECT 351.600 411.600 352.400 412.400 ;
        RECT 353.200 411.600 354.000 412.400 ;
        RECT 351.700 410.400 352.300 411.600 ;
        RECT 351.600 409.600 352.400 410.400 ;
        RECT 351.600 407.600 352.400 408.400 ;
        RECT 350.000 401.600 350.800 402.400 ;
        RECT 350.100 396.400 350.700 401.600 ;
        RECT 350.000 395.600 350.800 396.400 ;
        RECT 348.400 389.600 349.200 390.400 ;
        RECT 343.600 387.600 344.400 388.400 ;
        RECT 346.800 387.600 347.600 388.400 ;
        RECT 343.600 385.600 344.400 386.400 ;
        RECT 337.200 381.600 338.000 382.400 ;
        RECT 342.000 381.600 342.800 382.400 ;
        RECT 346.900 378.400 347.500 387.600 ;
        RECT 332.400 377.600 333.200 378.400 ;
        RECT 338.800 377.600 339.600 378.400 ;
        RECT 346.800 378.300 347.600 378.400 ;
        RECT 345.300 377.700 347.600 378.300 ;
        RECT 334.000 373.600 334.800 374.400 ;
        RECT 334.100 362.400 334.700 373.600 ;
        RECT 338.900 372.400 339.500 377.600 ;
        RECT 342.000 375.600 342.800 376.400 ;
        RECT 335.600 371.600 336.400 372.400 ;
        RECT 338.800 371.600 339.600 372.400 ;
        RECT 334.000 361.600 334.800 362.400 ;
        RECT 335.700 360.400 336.300 371.600 ;
        RECT 337.200 369.600 338.000 370.400 ;
        RECT 343.600 369.600 344.400 370.400 ;
        RECT 340.400 367.600 341.200 368.400 ;
        RECT 343.700 366.400 344.300 369.600 ;
        RECT 345.300 368.400 345.900 377.700 ;
        RECT 346.800 377.600 347.600 377.700 ;
        RECT 346.800 371.600 347.600 372.400 ;
        RECT 348.500 368.400 349.100 389.600 ;
        RECT 350.100 388.400 350.700 395.600 ;
        RECT 351.700 390.400 352.300 407.600 ;
        RECT 354.900 402.300 355.500 425.600 ;
        RECT 356.400 423.600 357.200 424.400 ;
        RECT 356.500 412.400 357.100 423.600 ;
        RECT 358.100 420.300 358.700 427.600 ;
        RECT 361.200 425.600 362.000 426.400 ;
        RECT 358.100 419.700 360.300 420.300 ;
        RECT 358.000 417.600 358.800 418.400 ;
        RECT 358.100 414.400 358.700 417.600 ;
        RECT 358.000 413.600 358.800 414.400 ;
        RECT 356.400 411.600 357.200 412.400 ;
        RECT 359.700 410.300 360.300 419.700 ;
        RECT 361.300 416.400 361.900 425.600 ;
        RECT 362.900 418.400 363.500 433.700 ;
        RECT 364.400 433.600 365.200 434.400 ;
        RECT 366.100 430.400 366.700 435.600 ;
        RECT 370.900 434.400 371.500 447.600 ;
        RECT 372.400 446.300 373.200 446.400 ;
        RECT 372.400 445.700 374.700 446.300 ;
        RECT 372.400 445.600 373.200 445.700 ;
        RECT 372.400 443.600 373.200 444.400 ;
        RECT 372.500 438.400 373.100 443.600 ;
        RECT 372.400 437.600 373.200 438.400 ;
        RECT 374.100 434.400 374.700 445.700 ;
        RECT 370.800 433.600 371.600 434.400 ;
        RECT 374.000 433.600 374.800 434.400 ;
        RECT 377.300 432.400 377.900 449.600 ;
        RECT 382.100 448.400 382.700 451.600 ;
        RECT 386.900 450.400 387.500 461.600 ;
        RECT 390.000 459.600 390.800 460.400 ;
        RECT 393.200 459.600 394.000 460.400 ;
        RECT 388.400 451.600 389.200 452.400 ;
        RECT 386.800 449.600 387.600 450.400 ;
        RECT 382.000 447.600 382.800 448.400 ;
        RECT 383.600 447.600 384.400 448.400 ;
        RECT 378.800 443.600 379.600 444.400 ;
        RECT 367.600 431.600 368.400 432.400 ;
        RECT 374.000 431.600 374.800 432.400 ;
        RECT 377.200 431.600 378.000 432.400 ;
        RECT 366.000 429.600 366.800 430.400 ;
        RECT 367.600 429.600 368.400 430.400 ;
        RECT 366.100 424.400 366.700 429.600 ;
        RECT 366.000 423.600 366.800 424.400 ;
        RECT 362.800 417.600 363.600 418.400 ;
        RECT 361.200 415.600 362.000 416.400 ;
        RECT 362.800 413.600 363.600 414.400 ;
        RECT 358.100 409.700 360.300 410.300 ;
        RECT 358.100 402.400 358.700 409.700 ;
        RECT 361.200 409.600 362.000 410.400 ;
        RECT 359.600 407.600 360.400 408.400 ;
        RECT 361.300 402.400 361.900 409.600 ;
        RECT 362.900 406.300 363.500 413.600 ;
        RECT 366.000 411.600 366.800 412.400 ;
        RECT 366.100 408.400 366.700 411.600 ;
        RECT 364.400 407.600 365.200 408.400 ;
        RECT 366.000 407.600 366.800 408.400 ;
        RECT 362.900 405.700 365.100 406.300 ;
        RECT 362.800 403.600 363.600 404.400 ;
        RECT 354.900 401.700 357.100 402.300 ;
        RECT 354.800 399.600 355.600 400.400 ;
        RECT 351.600 389.600 352.400 390.400 ;
        RECT 350.000 387.600 350.800 388.400 ;
        RECT 351.600 383.600 352.400 384.400 ;
        RECT 351.700 382.400 352.300 383.600 ;
        RECT 351.600 381.600 352.400 382.400 ;
        RECT 353.200 375.600 354.000 376.400 ;
        RECT 353.300 372.400 353.900 375.600 ;
        RECT 353.200 371.600 354.000 372.400 ;
        RECT 354.900 370.400 355.500 399.600 ;
        RECT 356.500 388.400 357.100 401.700 ;
        RECT 358.000 401.600 358.800 402.400 ;
        RECT 361.200 401.600 362.000 402.400 ;
        RECT 358.000 395.600 358.800 396.400 ;
        RECT 361.200 395.600 362.000 396.400 ;
        RECT 358.100 390.400 358.700 395.600 ;
        RECT 361.300 394.300 361.900 395.600 ;
        RECT 362.900 394.300 363.500 403.600 ;
        RECT 361.300 393.700 363.500 394.300 ;
        RECT 361.300 390.400 361.900 393.700 ;
        RECT 362.800 391.600 363.600 392.400 ;
        RECT 358.000 389.600 358.800 390.400 ;
        RECT 361.200 389.600 362.000 390.400 ;
        RECT 356.400 387.600 357.200 388.400 ;
        RECT 356.500 376.400 357.100 387.600 ;
        RECT 359.600 385.600 360.400 386.400 ;
        RECT 358.000 379.600 358.800 380.400 ;
        RECT 356.400 375.600 357.200 376.400 ;
        RECT 358.100 372.300 358.700 379.600 ;
        RECT 361.300 376.400 361.900 389.600 ;
        RECT 362.800 385.600 363.600 386.400 ;
        RECT 362.900 382.400 363.500 385.600 ;
        RECT 362.800 381.600 363.600 382.400 ;
        RECT 362.800 379.600 363.600 380.400 ;
        RECT 362.900 378.400 363.500 379.600 ;
        RECT 362.800 377.600 363.600 378.400 ;
        RECT 361.200 375.600 362.000 376.400 ;
        RECT 361.200 373.600 362.000 374.400 ;
        RECT 361.300 372.400 361.900 373.600 ;
        RECT 356.500 371.700 358.700 372.300 ;
        RECT 350.000 369.600 350.800 370.400 ;
        RECT 354.800 369.600 355.600 370.400 ;
        RECT 356.500 368.400 357.100 371.700 ;
        RECT 359.600 371.600 360.400 372.400 ;
        RECT 361.200 371.600 362.000 372.400 ;
        RECT 358.000 369.600 358.800 370.400 ;
        RECT 345.200 367.600 346.000 368.400 ;
        RECT 348.400 367.600 349.200 368.400 ;
        RECT 356.400 367.600 357.200 368.400 ;
        RECT 359.700 368.300 360.300 371.600 ;
        RECT 358.100 367.700 360.300 368.300 ;
        RECT 343.600 365.600 344.400 366.400 ;
        RECT 348.400 365.600 349.200 366.400 ;
        RECT 332.400 359.600 333.200 360.400 ;
        RECT 335.600 359.600 336.400 360.400 ;
        RECT 342.000 359.600 342.800 360.400 ;
        RECT 329.200 357.600 330.000 358.400 ;
        RECT 330.800 357.600 331.600 358.400 ;
        RECT 332.500 354.400 333.100 359.600 ;
        RECT 342.100 358.400 342.700 359.600 ;
        RECT 358.100 358.400 358.700 367.700 ;
        RECT 342.000 357.600 342.800 358.400 ;
        RECT 358.000 357.600 358.800 358.400 ;
        RECT 343.600 355.600 344.400 356.400 ;
        RECT 348.400 355.600 349.200 356.400 ;
        RECT 356.400 355.600 357.200 356.400 ;
        RECT 343.700 354.400 344.300 355.600 ;
        RECT 356.500 354.400 357.100 355.600 ;
        RECT 332.400 353.600 333.200 354.400 ;
        RECT 337.200 354.300 338.000 354.400 ;
        RECT 337.200 353.700 341.100 354.300 ;
        RECT 337.200 353.600 338.000 353.700 ;
        RECT 332.500 350.400 333.100 353.600 ;
        RECT 340.500 352.400 341.100 353.700 ;
        RECT 343.600 353.600 344.400 354.400 ;
        RECT 356.400 353.600 357.200 354.400 ;
        RECT 338.800 351.600 339.600 352.400 ;
        RECT 340.400 351.600 341.200 352.400 ;
        RECT 359.600 351.600 360.400 352.400 ;
        RECT 361.200 352.300 362.000 352.400 ;
        RECT 364.500 352.300 365.100 405.700 ;
        RECT 366.000 403.600 366.800 404.400 ;
        RECT 366.100 392.400 366.700 403.600 ;
        RECT 366.000 391.600 366.800 392.400 ;
        RECT 367.700 380.400 368.300 429.600 ;
        RECT 370.800 425.600 371.600 426.400 ;
        RECT 370.900 424.400 371.500 425.600 ;
        RECT 370.800 423.600 371.600 424.400 ;
        RECT 370.800 419.600 371.600 420.400 ;
        RECT 370.900 412.400 371.500 419.600 ;
        RECT 370.800 411.600 371.600 412.400 ;
        RECT 372.400 411.600 373.200 412.400 ;
        RECT 369.200 409.600 370.000 410.400 ;
        RECT 372.500 410.300 373.100 411.600 ;
        RECT 370.900 409.700 373.100 410.300 ;
        RECT 370.900 408.400 371.500 409.700 ;
        RECT 369.200 407.600 370.000 408.400 ;
        RECT 370.800 407.600 371.600 408.400 ;
        RECT 372.400 407.600 373.200 408.400 ;
        RECT 369.300 406.300 369.900 407.600 ;
        RECT 370.800 406.300 371.600 406.400 ;
        RECT 369.300 405.700 371.600 406.300 ;
        RECT 370.800 405.600 371.600 405.700 ;
        RECT 374.100 404.400 374.700 431.600 ;
        RECT 375.600 429.600 376.400 430.400 ;
        RECT 375.700 428.400 376.300 429.600 ;
        RECT 375.600 427.600 376.400 428.400 ;
        RECT 377.300 422.300 377.900 431.600 ;
        RECT 378.900 426.400 379.500 443.600 ;
        RECT 383.700 440.400 384.300 447.600 ;
        RECT 383.600 439.600 384.400 440.400 ;
        RECT 382.000 435.600 382.800 436.400 ;
        RECT 380.400 431.600 381.200 432.400 ;
        RECT 378.800 425.600 379.600 426.400 ;
        RECT 378.800 423.600 379.600 424.400 ;
        RECT 375.700 421.700 377.900 422.300 ;
        RECT 375.700 412.400 376.300 421.700 ;
        RECT 378.900 420.300 379.500 423.600 ;
        RECT 377.300 419.700 379.500 420.300 ;
        RECT 377.300 416.400 377.900 419.700 ;
        RECT 378.800 417.600 379.600 418.400 ;
        RECT 377.200 415.600 378.000 416.400 ;
        RECT 378.900 412.400 379.500 417.600 ;
        RECT 375.600 411.600 376.400 412.400 ;
        RECT 378.800 411.600 379.600 412.400 ;
        RECT 380.500 410.400 381.100 431.600 ;
        RECT 382.100 430.400 382.700 435.600 ;
        RECT 386.900 432.400 387.500 449.600 ;
        RECT 390.100 448.400 390.700 459.600 ;
        RECT 388.400 447.600 389.200 448.400 ;
        RECT 390.000 447.600 390.800 448.400 ;
        RECT 388.500 446.400 389.100 447.600 ;
        RECT 388.400 445.600 389.200 446.400 ;
        RECT 390.000 443.600 390.800 444.400 ;
        RECT 390.100 434.400 390.700 443.600 ;
        RECT 390.000 433.600 390.800 434.400 ;
        RECT 383.600 431.600 384.400 432.400 ;
        RECT 386.800 431.600 387.600 432.400 ;
        RECT 388.400 431.600 389.200 432.400 ;
        RECT 382.000 429.600 382.800 430.400 ;
        RECT 383.700 428.400 384.300 431.600 ;
        RECT 388.500 430.400 389.100 431.600 ;
        RECT 390.100 430.400 390.700 433.600 ;
        RECT 393.300 430.400 393.900 459.600 ;
        RECT 398.000 453.600 398.800 454.400 ;
        RECT 394.800 443.600 395.600 444.400 ;
        RECT 398.100 438.400 398.700 453.600 ;
        RECT 399.600 445.600 400.400 446.400 ;
        RECT 398.000 437.600 398.800 438.400 ;
        RECT 399.700 432.400 400.300 445.600 ;
        RECT 401.300 442.400 401.900 469.600 ;
        RECT 402.900 456.400 403.500 491.600 ;
        RECT 404.400 486.200 405.200 497.800 ;
        RECT 406.000 493.600 406.800 494.400 ;
        RECT 406.000 491.600 406.800 492.400 ;
        RECT 406.100 484.400 406.700 491.600 ;
        RECT 407.600 486.200 408.400 497.800 ;
        RECT 406.000 483.600 406.800 484.400 ;
        RECT 409.200 484.200 410.000 497.800 ;
        RECT 410.800 484.200 411.600 497.800 ;
        RECT 430.000 495.600 430.800 496.400 ;
        RECT 433.200 493.600 434.000 494.400 ;
        RECT 439.600 493.600 440.400 494.400 ;
        RECT 422.000 491.600 422.800 492.400 ;
        RECT 422.100 478.400 422.700 491.600 ;
        RECT 433.300 478.400 433.900 493.600 ;
        RECT 436.400 491.600 437.200 492.400 ;
        RECT 442.800 489.600 443.600 490.400 ;
        RECT 409.200 477.600 410.000 478.400 ;
        RECT 422.000 477.600 422.800 478.400 ;
        RECT 426.800 477.600 427.600 478.400 ;
        RECT 433.200 477.600 434.000 478.400 ;
        RECT 426.900 472.400 427.500 477.600 ;
        RECT 442.900 474.400 443.500 489.600 ;
        RECT 455.600 484.200 456.400 497.800 ;
        RECT 457.200 484.200 458.000 497.800 ;
        RECT 458.800 484.200 459.600 497.800 ;
        RECT 460.400 486.200 461.200 497.800 ;
        RECT 462.000 495.600 462.800 496.400 ;
        RECT 463.600 486.200 464.400 497.800 ;
        RECT 465.200 493.600 466.000 494.400 ;
        RECT 466.800 486.200 467.600 497.800 ;
        RECT 468.400 484.200 469.200 497.800 ;
        RECT 470.000 484.200 470.800 497.800 ;
        RECT 476.400 493.600 477.200 494.400 ;
        RECT 471.600 491.600 472.400 492.400 ;
        RECT 442.800 473.600 443.600 474.400 ;
        RECT 420.400 471.600 421.200 472.400 ;
        RECT 426.800 471.600 427.600 472.400 ;
        RECT 428.400 471.600 429.200 472.400 ;
        RECT 430.000 471.600 430.800 472.400 ;
        RECT 420.400 469.600 421.200 470.400 ;
        RECT 423.600 469.600 424.400 470.400 ;
        RECT 426.900 468.400 427.500 471.600 ;
        RECT 430.100 470.400 430.700 471.600 ;
        RECT 430.000 469.600 430.800 470.400 ;
        RECT 434.800 469.600 435.600 470.400 ;
        RECT 445.800 469.600 446.800 470.400 ;
        RECT 454.000 469.600 454.800 470.400 ;
        RECT 430.100 468.400 430.700 469.600 ;
        RECT 415.600 467.600 416.400 468.400 ;
        RECT 426.800 467.600 427.600 468.400 ;
        RECT 430.000 467.600 430.800 468.400 ;
        RECT 423.600 465.600 424.400 466.400 ;
        RECT 402.800 455.600 403.600 456.400 ;
        RECT 404.400 444.200 405.200 457.800 ;
        RECT 406.000 444.200 406.800 457.800 ;
        RECT 407.600 444.200 408.400 457.800 ;
        RECT 409.200 446.200 410.000 457.800 ;
        RECT 410.800 455.600 411.600 456.400 ;
        RECT 412.400 446.200 413.200 457.800 ;
        RECT 414.000 453.600 414.800 454.400 ;
        RECT 415.600 446.200 416.400 457.800 ;
        RECT 417.200 444.200 418.000 457.800 ;
        RECT 418.800 444.200 419.600 457.800 ;
        RECT 423.700 452.400 424.300 465.600 ;
        RECT 423.600 451.600 424.400 452.400 ;
        RECT 401.200 441.600 402.000 442.400 ;
        RECT 407.600 441.600 408.400 442.400 ;
        RECT 406.000 435.600 406.800 436.400 ;
        RECT 399.600 431.600 400.400 432.400 ;
        RECT 388.400 429.600 389.200 430.400 ;
        RECT 390.000 429.600 390.800 430.400 ;
        RECT 393.200 429.600 394.000 430.400 ;
        RECT 383.600 427.600 384.400 428.400 ;
        RECT 391.600 427.600 392.400 428.400 ;
        RECT 385.200 423.600 386.000 424.400 ;
        RECT 383.600 421.600 384.400 422.400 ;
        RECT 383.700 418.400 384.300 421.600 ;
        RECT 385.300 420.400 385.900 423.600 ;
        RECT 385.200 419.600 386.000 420.400 ;
        RECT 383.600 417.600 384.400 418.400 ;
        RECT 383.700 414.400 384.300 417.600 ;
        RECT 383.600 413.600 384.400 414.400 ;
        RECT 385.300 412.400 385.900 419.600 ;
        RECT 390.000 415.600 390.800 416.400 ;
        RECT 390.100 414.400 390.700 415.600 ;
        RECT 393.300 414.400 393.900 429.600 ;
        RECT 394.800 427.600 395.600 428.400 ;
        RECT 396.400 427.600 397.200 428.400 ;
        RECT 394.900 426.400 395.500 427.600 ;
        RECT 394.800 425.600 395.600 426.400 ;
        RECT 399.600 417.600 400.400 418.400 ;
        RECT 399.700 416.400 400.300 417.600 ;
        RECT 394.800 415.600 395.600 416.400 ;
        RECT 399.600 415.600 400.400 416.400 ;
        RECT 401.200 415.600 402.000 416.400 ;
        RECT 386.800 413.600 387.600 414.400 ;
        RECT 390.000 413.600 390.800 414.400 ;
        RECT 393.200 413.600 394.000 414.400 ;
        RECT 394.900 412.400 395.500 415.600 ;
        RECT 402.800 413.600 403.600 414.400 ;
        RECT 402.900 412.400 403.500 413.600 ;
        RECT 406.100 412.400 406.700 435.600 ;
        RECT 407.700 430.400 408.300 441.600 ;
        RECT 426.900 440.400 427.500 467.600 ;
        RECT 434.900 464.400 435.500 469.600 ;
        RECT 436.400 467.600 437.200 468.400 ;
        RECT 438.000 467.600 438.800 468.400 ;
        RECT 431.600 463.600 432.400 464.400 ;
        RECT 434.800 463.600 435.600 464.400 ;
        RECT 431.700 454.400 432.300 463.600 ;
        RECT 434.900 460.400 435.500 463.600 ;
        RECT 434.800 459.600 435.600 460.400 ;
        RECT 436.500 458.400 437.100 467.600 ;
        RECT 436.400 457.600 437.200 458.400 ;
        RECT 431.600 453.600 432.400 454.400 ;
        RECT 436.400 449.600 437.200 450.400 ;
        RECT 436.500 446.400 437.100 449.600 ;
        RECT 436.400 445.600 437.200 446.400 ;
        RECT 438.100 442.400 438.700 467.600 ;
        RECT 454.100 466.400 454.700 469.600 ;
        RECT 454.000 465.600 454.800 466.400 ;
        RECT 442.800 463.600 443.600 464.400 ;
        RECT 455.600 464.200 456.400 477.800 ;
        RECT 457.200 464.200 458.000 477.800 ;
        RECT 458.800 464.200 459.600 477.800 ;
        RECT 460.400 464.200 461.200 475.800 ;
        RECT 462.000 465.600 462.800 466.400 ;
        RECT 442.900 454.400 443.500 463.600 ;
        RECT 462.100 462.400 462.700 465.600 ;
        RECT 463.600 464.200 464.400 475.800 ;
        RECT 465.200 467.600 466.000 468.400 ;
        RECT 466.800 464.200 467.600 475.800 ;
        RECT 468.400 464.200 469.200 477.800 ;
        RECT 470.000 464.200 470.800 477.800 ;
        RECT 471.700 470.400 472.300 491.600 ;
        RECT 471.600 469.600 472.400 470.400 ;
        RECT 474.800 469.600 475.600 470.400 ;
        RECT 474.900 466.400 475.500 469.600 ;
        RECT 474.800 465.600 475.600 466.400 ;
        RECT 454.000 461.600 454.800 462.400 ;
        RECT 462.000 461.600 462.800 462.400 ;
        RECT 442.800 453.600 443.600 454.400 ;
        RECT 446.000 444.200 446.800 457.800 ;
        RECT 447.600 444.200 448.400 457.800 ;
        RECT 449.200 446.200 450.000 457.800 ;
        RECT 450.800 455.600 451.600 456.400 ;
        RECT 450.900 454.400 451.500 455.600 ;
        RECT 450.800 453.600 451.600 454.400 ;
        RECT 450.800 451.600 451.600 452.400 ;
        RECT 438.000 441.600 438.800 442.400 ;
        RECT 446.000 441.600 446.800 442.400 ;
        RECT 426.800 439.600 427.600 440.400 ;
        RECT 438.000 439.600 438.800 440.400 ;
        RECT 438.100 438.400 438.700 439.600 ;
        RECT 446.100 438.400 446.700 441.600 ;
        RECT 407.600 429.600 408.400 430.400 ;
        RECT 414.000 424.200 414.800 437.800 ;
        RECT 415.600 424.200 416.400 437.800 ;
        RECT 417.200 424.200 418.000 435.800 ;
        RECT 418.800 427.600 419.600 428.400 ;
        RECT 418.900 422.300 419.500 427.600 ;
        RECT 420.400 424.200 421.200 435.800 ;
        RECT 422.000 425.600 422.800 426.400 ;
        RECT 417.300 421.700 419.500 422.300 ;
        RECT 417.300 418.400 417.900 421.700 ;
        RECT 417.200 417.600 418.000 418.400 ;
        RECT 422.100 416.400 422.700 425.600 ;
        RECT 423.600 424.200 424.400 435.800 ;
        RECT 425.200 424.200 426.000 437.800 ;
        RECT 426.800 424.200 427.600 437.800 ;
        RECT 428.400 424.200 429.200 437.800 ;
        RECT 438.000 437.600 438.800 438.400 ;
        RECT 446.000 437.600 446.800 438.400 ;
        RECT 449.200 431.600 450.000 432.400 ;
        RECT 449.300 430.400 449.900 431.600 ;
        RECT 450.900 430.400 451.500 451.600 ;
        RECT 452.400 446.200 453.200 457.800 ;
        RECT 454.100 456.400 454.700 461.600 ;
        RECT 476.500 458.400 477.100 493.600 ;
        RECT 486.000 491.600 486.800 492.400 ;
        RECT 492.200 491.600 493.200 492.400 ;
        RECT 500.400 491.600 501.200 492.400 ;
        RECT 481.200 483.600 482.000 484.400 ;
        RECT 482.800 483.600 483.600 484.400 ;
        RECT 454.000 455.600 454.800 456.400 ;
        RECT 454.100 444.300 454.700 455.600 ;
        RECT 455.600 446.200 456.400 457.800 ;
        RECT 452.500 443.700 454.700 444.300 ;
        RECT 457.200 444.200 458.000 457.800 ;
        RECT 458.800 444.200 459.600 457.800 ;
        RECT 460.400 444.200 461.200 457.800 ;
        RECT 476.400 457.600 477.200 458.400 ;
        RECT 481.300 456.400 481.900 483.600 ;
        RECT 478.000 455.600 478.800 456.400 ;
        RECT 479.600 455.600 480.400 456.400 ;
        RECT 481.200 455.600 482.000 456.400 ;
        RECT 473.200 453.600 474.000 454.400 ;
        RECT 479.700 452.400 480.300 455.600 ;
        RECT 481.200 454.300 482.000 454.400 ;
        RECT 482.900 454.300 483.500 483.600 ;
        RECT 500.500 482.400 501.100 491.600 ;
        RECT 502.000 484.200 502.800 497.800 ;
        RECT 503.600 484.200 504.400 497.800 ;
        RECT 505.200 484.200 506.000 497.800 ;
        RECT 506.800 486.200 507.600 497.800 ;
        RECT 508.400 495.600 509.200 496.400 ;
        RECT 500.400 481.600 501.200 482.400 ;
        RECT 503.600 481.600 504.400 482.400 ;
        RECT 484.400 469.600 485.200 470.400 ;
        RECT 484.500 466.400 485.100 469.600 ;
        RECT 484.400 465.600 485.200 466.400 ;
        RECT 487.600 464.200 488.400 477.800 ;
        RECT 489.200 464.200 490.000 477.800 ;
        RECT 490.800 464.200 491.600 475.800 ;
        RECT 492.400 467.600 493.200 468.400 ;
        RECT 492.400 465.600 493.200 466.400 ;
        RECT 492.500 458.400 493.100 465.600 ;
        RECT 494.000 464.200 494.800 475.800 ;
        RECT 495.600 465.600 496.400 466.400 ;
        RECT 497.200 464.200 498.000 475.800 ;
        RECT 498.800 464.200 499.600 477.800 ;
        RECT 500.400 464.200 501.200 477.800 ;
        RECT 502.000 464.200 502.800 477.800 ;
        RECT 492.400 457.600 493.200 458.400 ;
        RECT 497.200 455.600 498.000 456.400 ;
        RECT 481.200 453.700 483.500 454.300 ;
        RECT 481.200 453.600 482.000 453.700 ;
        RECT 479.600 451.600 480.400 452.400 ;
        RECT 482.800 451.600 483.600 452.400 ;
        RECT 484.400 451.600 485.200 452.400 ;
        RECT 495.600 451.600 496.400 452.400 ;
        RECT 476.400 449.600 477.200 450.400 ;
        RECT 452.500 438.400 453.100 443.700 ;
        RECT 470.000 443.600 470.800 444.400 ;
        RECT 452.400 437.600 453.200 438.400 ;
        RECT 430.000 429.600 430.800 430.400 ;
        RECT 449.200 429.600 450.000 430.400 ;
        RECT 450.800 429.600 451.600 430.400 ;
        RECT 468.400 429.600 469.200 430.400 ;
        RECT 430.100 422.400 430.700 429.600 ;
        RECT 442.800 425.600 443.600 426.400 ;
        RECT 441.200 423.600 442.000 424.400 ;
        RECT 425.200 421.600 426.000 422.400 ;
        RECT 430.000 421.600 430.800 422.400 ;
        RECT 409.200 415.600 410.000 416.400 ;
        RECT 422.000 415.600 422.800 416.400 ;
        RECT 382.000 411.600 382.800 412.400 ;
        RECT 385.200 411.600 386.000 412.400 ;
        RECT 391.600 411.600 392.400 412.400 ;
        RECT 394.800 411.600 395.600 412.400 ;
        RECT 402.800 411.600 403.600 412.400 ;
        RECT 406.000 411.600 406.800 412.400 ;
        RECT 380.400 409.600 381.200 410.400 ;
        RECT 377.200 407.600 378.000 408.400 ;
        RECT 378.800 407.600 379.600 408.400 ;
        RECT 378.900 406.400 379.500 407.600 ;
        RECT 378.800 405.600 379.600 406.400 ;
        RECT 382.000 405.600 382.800 406.400 ;
        RECT 386.800 405.600 387.600 406.400 ;
        RECT 374.000 403.600 374.800 404.400 ;
        RECT 375.600 399.600 376.400 400.400 ;
        RECT 377.200 399.600 378.000 400.400 ;
        RECT 375.700 398.400 376.300 399.600 ;
        RECT 374.000 397.600 374.800 398.400 ;
        RECT 375.600 397.600 376.400 398.400 ;
        RECT 374.100 394.400 374.700 397.600 ;
        RECT 377.300 394.400 377.900 399.600 ;
        RECT 382.100 398.400 382.700 405.600 ;
        RECT 391.700 404.400 392.300 411.600 ;
        RECT 409.300 410.400 409.900 415.600 ;
        RECT 425.300 412.400 425.900 421.600 ;
        RECT 441.300 420.400 441.900 423.600 ;
        RECT 449.300 420.400 449.900 429.600 ;
        RECT 436.400 419.600 437.200 420.400 ;
        RECT 441.200 419.600 442.000 420.400 ;
        RECT 449.200 419.600 450.000 420.400 ;
        RECT 425.200 411.600 426.000 412.400 ;
        RECT 393.200 409.600 394.000 410.400 ;
        RECT 409.200 409.600 410.000 410.400 ;
        RECT 393.300 408.400 393.900 409.600 ;
        RECT 393.200 407.600 394.000 408.400 ;
        RECT 396.400 407.600 397.200 408.400 ;
        RECT 412.400 407.600 413.200 408.400 ;
        RECT 396.500 406.400 397.100 407.600 ;
        RECT 396.400 405.600 397.200 406.400 ;
        RECT 391.600 403.600 392.400 404.400 ;
        RECT 394.800 403.600 395.600 404.400 ;
        RECT 406.000 403.600 406.800 404.400 ;
        RECT 390.000 401.600 390.800 402.400 ;
        RECT 382.000 397.600 382.800 398.400 ;
        RECT 369.200 393.600 370.000 394.400 ;
        RECT 374.000 393.600 374.800 394.400 ;
        RECT 377.200 393.600 378.000 394.400 ;
        RECT 369.300 392.400 369.900 393.600 ;
        RECT 374.100 392.400 374.700 393.600 ;
        RECT 369.200 391.600 370.000 392.400 ;
        RECT 374.000 391.600 374.800 392.400 ;
        RECT 375.600 391.600 376.400 392.400 ;
        RECT 375.700 390.400 376.300 391.600 ;
        RECT 369.200 389.600 370.000 390.400 ;
        RECT 375.600 389.600 376.400 390.400 ;
        RECT 367.600 379.600 368.400 380.400 ;
        RECT 367.600 375.600 368.400 376.400 ;
        RECT 366.000 371.600 366.800 372.400 ;
        RECT 366.100 370.400 366.700 371.600 ;
        RECT 366.000 369.600 366.800 370.400 ;
        RECT 369.300 366.400 369.900 389.600 ;
        RECT 372.400 387.600 373.200 388.400 ;
        RECT 377.300 378.400 377.900 393.600 ;
        RECT 383.600 391.600 384.400 392.400 ;
        RECT 386.800 391.600 387.600 392.400 ;
        RECT 383.700 388.400 384.300 391.600 ;
        RECT 380.400 387.600 381.200 388.400 ;
        RECT 383.600 387.600 384.400 388.400 ;
        RECT 377.200 377.600 378.000 378.400 ;
        RECT 375.600 373.600 376.400 374.400 ;
        RECT 375.700 372.400 376.300 373.600 ;
        RECT 370.800 371.600 371.600 372.400 ;
        RECT 375.600 371.600 376.400 372.400 ;
        RECT 377.200 371.600 378.000 372.400 ;
        RECT 370.900 370.400 371.500 371.600 ;
        RECT 370.800 369.600 371.600 370.400 ;
        RECT 372.400 369.600 373.200 370.400 ;
        RECT 369.200 365.600 370.000 366.400 ;
        RECT 372.500 362.400 373.100 369.600 ;
        RECT 375.600 365.600 376.400 366.400 ;
        RECT 372.400 361.600 373.200 362.400 ;
        RECT 377.300 360.400 377.900 371.600 ;
        RECT 380.500 370.400 381.100 387.600 ;
        RECT 386.900 372.400 387.500 391.600 ;
        RECT 388.400 389.600 389.200 390.400 ;
        RECT 382.000 371.600 382.800 372.400 ;
        RECT 386.800 371.600 387.600 372.400 ;
        RECT 378.800 369.600 379.600 370.400 ;
        RECT 380.400 369.600 381.200 370.400 ;
        RECT 380.400 367.600 381.200 368.400 ;
        RECT 380.500 366.400 381.100 367.600 ;
        RECT 382.100 366.400 382.700 371.600 ;
        RECT 385.200 369.600 386.000 370.400 ;
        RECT 388.400 369.600 389.200 370.400 ;
        RECT 388.500 368.400 389.100 369.600 ;
        RECT 388.400 367.600 389.200 368.400 ;
        RECT 380.400 365.600 381.200 366.400 ;
        RECT 382.000 365.600 382.800 366.400 ;
        RECT 377.200 359.600 378.000 360.400 ;
        RECT 380.400 359.600 381.200 360.400 ;
        RECT 380.500 358.400 381.100 359.600 ;
        RECT 380.400 357.600 381.200 358.400 ;
        RECT 374.000 353.600 374.800 354.400 ;
        RECT 375.600 353.600 376.400 354.400 ;
        RECT 382.000 353.600 382.800 354.400 ;
        RECT 366.000 352.300 366.800 352.400 ;
        RECT 361.200 351.700 363.500 352.300 ;
        RECT 364.500 351.700 366.800 352.300 ;
        RECT 361.200 351.600 362.000 351.700 ;
        RECT 338.900 350.400 339.500 351.600 ;
        RECT 330.800 349.600 331.600 350.400 ;
        RECT 332.400 349.600 333.200 350.400 ;
        RECT 334.000 349.600 334.800 350.400 ;
        RECT 338.800 349.600 339.600 350.400 ;
        RECT 342.000 349.600 342.800 350.400 ;
        RECT 343.600 349.600 344.400 350.400 ;
        RECT 346.800 350.300 347.600 350.400 ;
        RECT 345.300 349.700 347.600 350.300 ;
        RECT 329.200 347.600 330.000 348.400 ;
        RECT 329.300 346.400 329.900 347.600 ;
        RECT 329.200 345.600 330.000 346.400 ;
        RECT 330.900 344.400 331.500 349.600 ;
        RECT 334.100 348.400 334.700 349.600 ;
        RECT 334.000 347.600 334.800 348.400 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 330.800 343.600 331.600 344.400 ;
        RECT 334.100 344.300 334.700 347.600 ;
        RECT 342.100 346.400 342.700 349.600 ;
        RECT 340.400 345.600 341.200 346.400 ;
        RECT 342.000 345.600 342.800 346.400 ;
        RECT 334.100 343.700 336.300 344.300 ;
        RECT 329.200 341.600 330.000 342.400 ;
        RECT 326.100 337.700 328.300 338.300 ;
        RECT 324.400 333.600 325.200 334.400 ;
        RECT 322.800 331.600 323.600 332.400 ;
        RECT 322.800 329.600 323.600 330.400 ;
        RECT 321.200 327.600 322.000 328.400 ;
        RECT 321.200 315.600 322.000 316.400 ;
        RECT 311.600 311.600 312.400 312.400 ;
        RECT 313.200 311.600 314.000 312.400 ;
        RECT 316.400 311.600 317.200 312.400 ;
        RECT 318.000 311.600 318.800 312.400 ;
        RECT 319.600 311.600 320.400 312.400 ;
        RECT 311.600 310.300 312.400 310.400 ;
        RECT 313.300 310.300 313.900 311.600 ;
        RECT 316.500 310.400 317.100 311.600 ;
        RECT 311.600 309.700 313.900 310.300 ;
        RECT 311.600 309.600 312.400 309.700 ;
        RECT 316.400 309.600 317.200 310.400 ;
        RECT 322.900 308.400 323.500 329.600 ;
        RECT 324.400 327.600 325.200 328.400 ;
        RECT 326.100 312.300 326.700 337.700 ;
        RECT 327.600 333.600 328.400 334.400 ;
        RECT 327.700 332.400 328.300 333.600 ;
        RECT 329.300 332.400 329.900 341.600 ;
        RECT 332.400 337.600 333.200 338.400 ;
        RECT 332.400 333.600 333.200 334.400 ;
        RECT 335.700 332.400 336.300 343.700 ;
        RECT 338.800 341.600 339.600 342.400 ;
        RECT 337.200 339.600 338.000 340.400 ;
        RECT 337.300 332.400 337.900 339.600 ;
        RECT 338.900 332.400 339.500 341.600 ;
        RECT 340.500 336.400 341.100 345.600 ;
        RECT 340.400 335.600 341.200 336.400 ;
        RECT 340.500 334.400 341.100 335.600 ;
        RECT 343.700 334.400 344.300 349.600 ;
        RECT 345.300 340.400 345.900 349.700 ;
        RECT 346.800 349.600 347.600 349.700 ;
        RECT 353.200 349.600 354.000 350.400 ;
        RECT 358.000 349.600 358.800 350.400 ;
        RECT 359.700 350.300 360.300 351.600 ;
        RECT 361.200 350.300 362.000 350.400 ;
        RECT 359.700 349.700 362.000 350.300 ;
        RECT 361.200 349.600 362.000 349.700 ;
        RECT 346.800 347.600 347.600 348.400 ;
        RECT 351.600 347.600 352.400 348.400 ;
        RECT 345.200 339.600 346.000 340.400 ;
        RECT 346.900 334.400 347.500 347.600 ;
        RECT 348.400 345.600 349.200 346.400 ;
        RECT 348.500 338.400 349.100 345.600 ;
        RECT 348.400 337.600 349.200 338.400 ;
        RECT 351.700 336.400 352.300 347.600 ;
        RECT 358.100 344.400 358.700 349.600 ;
        RECT 358.000 343.600 358.800 344.400 ;
        RECT 354.800 337.600 355.600 338.400 ;
        RECT 351.600 335.600 352.400 336.400 ;
        RECT 351.700 334.400 352.300 335.600 ;
        RECT 340.400 333.600 341.200 334.400 ;
        RECT 343.600 333.600 344.400 334.400 ;
        RECT 346.800 333.600 347.600 334.400 ;
        RECT 348.400 333.600 349.200 334.400 ;
        RECT 351.600 333.600 352.400 334.400 ;
        RECT 327.600 331.600 328.400 332.400 ;
        RECT 329.200 331.600 330.000 332.400 ;
        RECT 330.800 331.600 331.600 332.400 ;
        RECT 335.600 331.600 336.400 332.400 ;
        RECT 337.200 331.600 338.000 332.400 ;
        RECT 338.800 331.600 339.600 332.400 ;
        RECT 327.600 312.300 328.400 312.400 ;
        RECT 326.100 311.700 328.400 312.300 ;
        RECT 327.600 311.600 328.400 311.700 ;
        RECT 324.400 309.600 325.200 310.400 ;
        RECT 322.800 307.600 323.600 308.400 ;
        RECT 313.200 295.600 314.000 296.400 ;
        RECT 318.000 295.600 318.800 296.400 ;
        RECT 308.400 291.700 310.700 292.300 ;
        RECT 308.400 291.600 309.200 291.700 ;
        RECT 313.300 288.400 313.900 295.600 ;
        RECT 314.800 293.600 315.600 294.400 ;
        RECT 314.900 292.400 315.500 293.600 ;
        RECT 314.800 291.600 315.600 292.400 ;
        RECT 306.800 287.600 307.600 288.400 ;
        RECT 313.200 287.600 314.000 288.400 ;
        RECT 308.400 283.600 309.200 284.400 ;
        RECT 314.800 283.600 315.600 284.400 ;
        RECT 308.500 282.400 309.100 283.600 ;
        RECT 308.400 281.600 309.200 282.400 ;
        RECT 314.900 280.400 315.500 283.600 ;
        RECT 300.400 279.600 301.200 280.400 ;
        RECT 314.800 279.600 315.600 280.400 ;
        RECT 297.200 273.600 298.000 274.400 ;
        RECT 297.200 269.600 298.000 270.400 ;
        RECT 297.300 260.400 297.900 269.600 ;
        RECT 302.000 264.200 302.800 277.800 ;
        RECT 303.600 264.200 304.400 277.800 ;
        RECT 310.000 277.600 310.800 278.400 ;
        RECT 305.200 264.200 306.000 275.800 ;
        RECT 306.800 267.600 307.600 268.400 ;
        RECT 306.900 266.400 307.500 267.600 ;
        RECT 306.800 265.600 307.600 266.400 ;
        RECT 308.400 264.200 309.200 275.800 ;
        RECT 310.100 270.400 310.700 277.600 ;
        RECT 310.000 269.600 310.800 270.400 ;
        RECT 310.100 266.400 310.700 269.600 ;
        RECT 310.000 265.600 310.800 266.400 ;
        RECT 311.600 264.200 312.400 275.800 ;
        RECT 313.200 264.200 314.000 277.800 ;
        RECT 314.800 264.200 315.600 277.800 ;
        RECT 316.400 264.200 317.200 277.800 ;
        RECT 313.200 261.600 314.000 262.400 ;
        RECT 295.600 259.600 296.400 260.400 ;
        RECT 297.200 259.600 298.000 260.400 ;
        RECT 302.000 259.600 302.800 260.400 ;
        RECT 284.400 244.200 285.200 257.800 ;
        RECT 286.000 244.200 286.800 257.800 ;
        RECT 287.600 244.200 288.400 257.800 ;
        RECT 289.200 246.200 290.000 257.800 ;
        RECT 290.800 255.600 291.600 256.400 ;
        RECT 290.900 250.400 291.500 255.600 ;
        RECT 290.800 249.600 291.600 250.400 ;
        RECT 290.800 245.600 291.600 246.400 ;
        RECT 292.400 246.200 293.200 257.800 ;
        RECT 294.000 255.600 294.800 256.400 ;
        RECT 294.100 254.400 294.700 255.600 ;
        RECT 294.000 253.600 294.800 254.400 ;
        RECT 295.600 246.200 296.400 257.800 ;
        RECT 284.400 241.600 285.200 242.400 ;
        RECT 284.500 238.400 285.100 241.600 ;
        RECT 284.400 237.600 285.200 238.400 ;
        RECT 290.900 234.400 291.500 245.600 ;
        RECT 297.200 244.200 298.000 257.800 ;
        RECT 298.800 244.200 299.600 257.800 ;
        RECT 302.100 252.400 302.700 259.600 ;
        RECT 302.000 251.600 302.800 252.400 ;
        RECT 310.000 251.600 310.800 252.400 ;
        RECT 311.600 247.600 312.400 248.400 ;
        RECT 310.000 243.600 310.800 244.400 ;
        RECT 295.600 241.600 296.400 242.400 ;
        RECT 290.800 233.600 291.600 234.400 ;
        RECT 295.700 232.400 296.300 241.600 ;
        RECT 310.100 232.400 310.700 243.600 ;
        RECT 294.000 231.600 294.800 232.400 ;
        RECT 295.600 231.600 296.400 232.400 ;
        RECT 310.000 231.600 310.800 232.400 ;
        RECT 287.600 229.600 288.400 230.400 ;
        RECT 290.800 229.600 291.600 230.400 ;
        RECT 287.700 228.400 288.300 229.600 ;
        RECT 290.900 228.400 291.500 229.600 ;
        RECT 287.600 227.600 288.400 228.400 ;
        RECT 290.800 227.600 291.600 228.400 ;
        RECT 294.100 226.400 294.700 231.600 ;
        RECT 313.300 230.400 313.900 261.600 ;
        RECT 316.400 251.600 317.200 252.400 ;
        RECT 318.100 248.400 318.700 295.600 ;
        RECT 322.900 294.400 323.500 307.600 ;
        RECT 324.500 306.400 325.100 309.600 ;
        RECT 324.400 305.600 325.200 306.400 ;
        RECT 327.700 298.400 328.300 311.600 ;
        RECT 324.400 297.600 325.200 298.400 ;
        RECT 327.600 297.600 328.400 298.400 ;
        RECT 322.800 293.600 323.600 294.400 ;
        RECT 321.200 291.600 322.000 292.400 ;
        RECT 324.500 292.300 325.100 297.600 ;
        RECT 327.600 293.600 328.400 294.400 ;
        RECT 322.900 291.700 325.100 292.300 ;
        RECT 322.900 290.400 323.500 291.700 ;
        RECT 329.300 290.400 329.900 331.600 ;
        RECT 330.900 320.400 331.500 331.600 ;
        RECT 337.300 330.400 337.900 331.600 ;
        RECT 337.200 329.600 338.000 330.400 ;
        RECT 343.700 330.300 344.300 333.600 ;
        RECT 354.900 332.400 355.500 337.600 ;
        RECT 359.600 336.300 360.400 336.400 ;
        RECT 359.600 335.700 361.900 336.300 ;
        RECT 359.600 335.600 360.400 335.700 ;
        RECT 361.300 334.400 361.900 335.700 ;
        RECT 356.400 333.600 357.200 334.400 ;
        RECT 359.600 333.600 360.400 334.400 ;
        RECT 361.200 333.600 362.000 334.400 ;
        RECT 356.500 332.400 357.100 333.600 ;
        RECT 362.900 332.400 363.500 351.700 ;
        RECT 366.000 351.600 366.800 351.700 ;
        RECT 366.100 348.400 366.700 351.600 ;
        RECT 370.800 349.600 371.600 350.400 ;
        RECT 364.400 347.600 365.200 348.400 ;
        RECT 366.000 347.600 366.800 348.400 ;
        RECT 367.600 347.600 368.400 348.400 ;
        RECT 369.200 347.600 370.000 348.400 ;
        RECT 372.400 347.600 373.200 348.400 ;
        RECT 364.500 346.400 365.100 347.600 ;
        RECT 364.400 345.600 365.200 346.400 ;
        RECT 366.000 343.600 366.800 344.400 ;
        RECT 364.400 339.600 365.200 340.400 ;
        RECT 364.500 338.400 365.100 339.600 ;
        RECT 364.400 337.600 365.200 338.400 ;
        RECT 367.700 334.400 368.300 347.600 ;
        RECT 369.300 344.400 369.900 347.600 ;
        RECT 369.200 343.600 370.000 344.400 ;
        RECT 372.500 336.400 373.100 347.600 ;
        RECT 374.100 340.400 374.700 353.600 ;
        RECT 378.800 351.600 379.600 352.400 ;
        RECT 377.200 349.600 378.000 350.400 ;
        RECT 375.600 347.600 376.400 348.400 ;
        RECT 374.000 339.600 374.800 340.400 ;
        RECT 372.400 335.600 373.200 336.400 ;
        RECT 372.500 334.400 373.100 335.600 ;
        RECT 367.600 333.600 368.400 334.400 ;
        RECT 372.400 333.600 373.200 334.400 ;
        RECT 374.100 332.400 374.700 339.600 ;
        RECT 377.300 338.400 377.900 349.600 ;
        RECT 378.900 338.400 379.500 351.600 ;
        RECT 380.400 349.600 381.200 350.400 ;
        RECT 382.000 349.600 382.800 350.400 ;
        RECT 380.500 338.400 381.100 349.600 ;
        RECT 377.200 337.600 378.000 338.400 ;
        RECT 378.800 337.600 379.600 338.400 ;
        RECT 380.400 337.600 381.200 338.400 ;
        RECT 375.600 333.600 376.400 334.400 ;
        RECT 380.400 333.600 381.200 334.400 ;
        RECT 345.200 331.600 346.000 332.400 ;
        RECT 346.800 331.600 347.600 332.400 ;
        RECT 353.200 331.600 354.000 332.400 ;
        RECT 354.800 331.600 355.600 332.400 ;
        RECT 356.400 331.600 357.200 332.400 ;
        RECT 361.200 331.600 362.000 332.400 ;
        RECT 362.800 331.600 363.600 332.400 ;
        RECT 367.600 331.600 368.400 332.400 ;
        RECT 374.000 331.600 374.800 332.400 ;
        RECT 343.700 329.700 345.900 330.300 ;
        RECT 340.400 323.600 341.200 324.400 ;
        RECT 338.800 321.600 339.600 322.400 ;
        RECT 330.800 319.600 331.600 320.400 ;
        RECT 334.000 315.600 334.800 316.400 ;
        RECT 334.100 314.400 334.700 315.600 ;
        RECT 334.000 313.600 334.800 314.400 ;
        RECT 330.800 311.600 331.600 312.400 ;
        RECT 337.200 307.600 338.000 308.400 ;
        RECT 332.400 303.600 333.200 304.400 ;
        RECT 330.800 297.600 331.600 298.400 ;
        RECT 330.800 295.600 331.600 296.400 ;
        RECT 321.200 289.600 322.000 290.400 ;
        RECT 322.800 289.600 323.600 290.400 ;
        RECT 324.400 289.600 325.200 290.400 ;
        RECT 329.200 289.600 330.000 290.400 ;
        RECT 321.300 286.400 321.900 289.600 ;
        RECT 322.800 287.600 323.600 288.400 ;
        RECT 321.200 285.600 322.000 286.400 ;
        RECT 319.600 275.600 320.400 276.400 ;
        RECT 318.000 247.600 318.800 248.400 ;
        RECT 316.400 243.600 317.200 244.400 ;
        RECT 316.500 232.400 317.100 243.600 ;
        RECT 318.000 241.600 318.800 242.400 ;
        RECT 316.400 231.600 317.200 232.400 ;
        RECT 300.400 229.600 301.200 230.400 ;
        RECT 306.800 229.600 307.600 230.400 ;
        RECT 313.200 229.600 314.000 230.400 ;
        RECT 316.400 229.600 317.200 230.400 ;
        RECT 300.400 227.600 301.200 228.400 ;
        RECT 311.600 227.600 312.400 228.400 ;
        RECT 282.800 225.600 283.600 226.400 ;
        RECT 286.000 225.600 286.800 226.400 ;
        RECT 294.000 225.600 294.800 226.400 ;
        RECT 273.200 223.600 274.000 224.400 ;
        RECT 294.000 223.600 294.800 224.400 ;
        RECT 295.600 223.600 296.400 224.400 ;
        RECT 258.800 215.600 259.600 216.400 ;
        RECT 255.600 211.600 256.400 212.400 ;
        RECT 270.000 211.600 270.800 212.400 ;
        RECT 257.200 209.600 258.000 210.400 ;
        RECT 254.000 207.600 254.800 208.400 ;
        RECT 252.400 203.600 253.200 204.400 ;
        RECT 252.500 200.400 253.100 203.600 ;
        RECT 270.100 200.400 270.700 211.600 ;
        RECT 273.200 204.200 274.000 217.800 ;
        RECT 274.800 204.200 275.600 217.800 ;
        RECT 276.400 206.200 277.200 217.800 ;
        RECT 278.000 213.600 278.800 214.400 ;
        RECT 278.100 210.400 278.700 213.600 ;
        RECT 278.000 209.600 278.800 210.400 ;
        RECT 279.600 206.200 280.400 217.800 ;
        RECT 281.200 215.600 282.000 216.400 ;
        RECT 281.300 200.400 281.900 215.600 ;
        RECT 282.800 206.200 283.600 217.800 ;
        RECT 284.400 204.200 285.200 217.800 ;
        RECT 286.000 204.200 286.800 217.800 ;
        RECT 287.600 204.200 288.400 217.800 ;
        RECT 294.100 216.400 294.700 223.600 ;
        RECT 294.000 215.600 294.800 216.400 ;
        RECT 295.700 214.400 296.300 223.600 ;
        RECT 298.800 215.600 299.600 216.400 ;
        RECT 298.900 214.400 299.500 215.600 ;
        RECT 295.600 213.600 296.400 214.400 ;
        RECT 298.800 213.600 299.600 214.400 ;
        RECT 298.800 211.600 299.600 212.400 ;
        RECT 300.500 206.400 301.100 227.600 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 302.100 224.400 302.700 225.600 ;
        RECT 302.000 223.600 302.800 224.400 ;
        RECT 308.400 223.600 309.200 224.400 ;
        RECT 310.000 223.600 310.800 224.400 ;
        RECT 302.000 217.600 302.800 218.400 ;
        RECT 305.200 215.600 306.000 216.400 ;
        RECT 305.300 214.400 305.900 215.600 ;
        RECT 303.600 213.600 304.400 214.400 ;
        RECT 305.200 213.600 306.000 214.400 ;
        RECT 303.700 212.400 304.300 213.600 ;
        RECT 303.600 211.600 304.400 212.400 ;
        RECT 303.600 209.600 304.400 210.400 ;
        RECT 306.800 209.600 307.600 210.400 ;
        RECT 300.400 205.600 301.200 206.400 ;
        RECT 303.600 205.600 304.400 206.400 ;
        RECT 252.400 199.600 253.200 200.400 ;
        RECT 255.600 199.600 256.400 200.400 ;
        RECT 270.000 199.600 270.800 200.400 ;
        RECT 278.000 199.600 278.800 200.400 ;
        RECT 281.200 199.600 282.000 200.400 ;
        RECT 226.800 195.600 227.600 196.400 ;
        RECT 226.900 190.400 227.500 195.600 ;
        RECT 238.000 191.600 238.800 192.400 ;
        RECT 238.100 190.400 238.700 191.600 ;
        RECT 225.200 189.600 226.000 190.400 ;
        RECT 226.800 189.600 227.600 190.400 ;
        RECT 238.000 189.600 238.800 190.400 ;
        RECT 225.300 188.400 225.900 189.600 ;
        RECT 220.400 187.600 221.200 188.400 ;
        RECT 225.200 187.600 226.000 188.400 ;
        RECT 229.800 187.600 230.800 188.400 ;
        RECT 220.500 186.400 221.100 187.600 ;
        RECT 220.400 185.600 221.200 186.400 ;
        RECT 223.600 185.600 224.400 186.400 ;
        RECT 239.600 184.200 240.400 197.800 ;
        RECT 241.200 184.200 242.000 197.800 ;
        RECT 242.800 184.200 243.600 197.800 ;
        RECT 244.400 184.200 245.200 195.800 ;
        RECT 246.000 185.600 246.800 186.400 ;
        RECT 246.100 184.400 246.700 185.600 ;
        RECT 246.000 183.600 246.800 184.400 ;
        RECT 247.600 184.200 248.400 195.800 ;
        RECT 249.200 187.600 250.000 188.400 ;
        RECT 249.300 186.400 249.900 187.600 ;
        RECT 249.200 185.600 250.000 186.400 ;
        RECT 250.800 184.200 251.600 195.800 ;
        RECT 252.400 184.200 253.200 197.800 ;
        RECT 254.000 184.200 254.800 197.800 ;
        RECT 255.700 190.400 256.300 199.600 ;
        RECT 278.100 190.400 278.700 199.600 ;
        RECT 303.700 198.400 304.300 205.600 ;
        RECT 255.600 189.600 256.400 190.400 ;
        RECT 278.000 189.600 278.800 190.400 ;
        RECT 260.400 187.600 261.200 188.400 ;
        RECT 218.800 175.600 219.600 176.400 ;
        RECT 206.000 171.600 206.800 172.400 ;
        RECT 209.200 171.600 210.000 172.400 ;
        RECT 215.600 171.600 216.400 172.400 ;
        RECT 230.000 171.600 230.800 172.400 ;
        RECT 206.100 154.400 206.700 171.600 ;
        RECT 220.400 167.600 221.200 168.400 ;
        RECT 215.600 163.600 216.400 164.400 ;
        RECT 206.000 153.600 206.800 154.400 ;
        RECT 209.200 153.600 210.000 154.400 ;
        RECT 206.100 150.400 206.700 153.600 ;
        RECT 209.300 152.400 209.900 153.600 ;
        RECT 215.700 152.400 216.300 163.600 ;
        RECT 217.200 153.600 218.000 154.400 ;
        RECT 209.200 151.600 210.000 152.400 ;
        RECT 215.600 151.600 216.400 152.400 ;
        RECT 209.300 150.400 209.900 151.600 ;
        RECT 206.000 149.600 206.800 150.400 ;
        RECT 209.200 149.600 210.000 150.400 ;
        RECT 212.400 149.600 213.200 150.400 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 214.100 148.400 214.700 149.600 ;
        RECT 215.700 148.400 216.300 151.600 ;
        RECT 202.800 147.600 203.600 148.400 ;
        RECT 204.400 147.600 205.200 148.400 ;
        RECT 214.000 147.600 214.800 148.400 ;
        RECT 215.600 147.600 216.400 148.400 ;
        RECT 218.800 145.600 219.600 146.400 ;
        RECT 196.400 135.600 197.200 136.400 ;
        RECT 178.800 133.600 179.600 134.400 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 186.800 133.600 187.600 134.400 ;
        RECT 193.200 133.600 194.000 134.400 ;
        RECT 194.800 133.600 195.600 134.400 ;
        RECT 180.400 131.600 181.200 132.400 ;
        RECT 191.600 131.600 192.400 132.400 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 175.600 129.600 176.400 130.400 ;
        RECT 177.200 129.600 178.000 130.400 ;
        RECT 174.000 125.600 174.800 126.400 ;
        RECT 174.100 124.400 174.700 125.600 ;
        RECT 174.000 123.600 174.800 124.400 ;
        RECT 175.600 119.600 176.400 120.400 ;
        RECT 174.000 111.600 174.800 112.400 ;
        RECT 172.400 107.600 173.200 108.400 ;
        RECT 172.500 94.400 173.100 107.600 ;
        RECT 174.100 98.400 174.700 111.600 ;
        RECT 175.700 110.400 176.300 119.600 ;
        RECT 177.200 115.600 178.000 116.400 ;
        RECT 175.600 109.600 176.400 110.400 ;
        RECT 174.000 97.600 174.800 98.400 ;
        RECT 175.700 96.400 176.300 109.600 ;
        RECT 177.300 98.400 177.900 115.600 ;
        RECT 178.800 111.600 179.600 112.400 ;
        RECT 180.500 110.300 181.100 131.600 ;
        RECT 183.600 129.600 184.400 130.400 ;
        RECT 191.600 130.300 192.400 130.400 ;
        RECT 193.300 130.300 193.900 131.600 ;
        RECT 191.600 129.700 193.900 130.300 ;
        RECT 191.600 129.600 192.400 129.700 ;
        RECT 199.600 129.600 200.400 130.400 ;
        RECT 182.000 115.600 182.800 116.400 ;
        RECT 178.900 109.700 181.100 110.300 ;
        RECT 178.900 98.400 179.500 109.700 ;
        RECT 180.400 107.600 181.200 108.400 ;
        RECT 180.500 106.400 181.100 107.600 ;
        RECT 180.400 105.600 181.200 106.400 ;
        RECT 177.200 97.600 178.000 98.400 ;
        RECT 178.800 97.600 179.600 98.400 ;
        RECT 175.600 95.600 176.400 96.400 ;
        RECT 172.400 93.600 173.200 94.400 ;
        RECT 172.500 76.400 173.100 93.600 ;
        RECT 174.000 89.600 174.800 90.400 ;
        RECT 174.100 88.400 174.700 89.600 ;
        RECT 174.000 87.600 174.800 88.400 ;
        RECT 175.700 82.400 176.300 95.600 ;
        RECT 175.600 81.600 176.400 82.400 ;
        RECT 172.400 75.600 173.200 76.400 ;
        RECT 175.600 75.600 176.400 76.400 ;
        RECT 175.700 72.400 176.300 75.600 ;
        RECT 172.400 71.600 173.200 72.400 ;
        RECT 175.600 71.600 176.400 72.400 ;
        RECT 162.800 69.600 163.600 70.400 ;
        RECT 167.600 69.600 168.400 70.400 ;
        RECT 170.800 69.600 171.600 70.400 ;
        RECT 172.500 68.400 173.100 71.600 ;
        RECT 174.000 69.600 174.800 70.400 ;
        RECT 161.200 67.600 162.000 68.400 ;
        RECT 167.600 67.600 168.400 68.400 ;
        RECT 172.400 67.600 173.200 68.400 ;
        RECT 161.300 66.400 161.900 67.600 ;
        RECT 161.200 65.600 162.000 66.400 ;
        RECT 159.600 63.600 160.400 64.400 ;
        RECT 167.700 58.400 168.300 67.600 ;
        RECT 170.800 65.600 171.600 66.400 ;
        RECT 164.400 57.600 165.200 58.400 ;
        RECT 167.600 57.600 168.400 58.400 ;
        RECT 159.600 55.600 160.400 56.400 ;
        RECT 151.600 51.600 152.400 52.400 ;
        RECT 156.400 51.600 157.200 52.400 ;
        RECT 158.000 51.600 158.800 52.400 ;
        RECT 156.500 50.400 157.100 51.600 ;
        RECT 156.400 49.600 157.200 50.400 ;
        RECT 153.200 43.600 154.000 44.400 ;
        RECT 145.200 37.600 146.000 38.400 ;
        RECT 146.800 37.600 147.600 38.400 ;
        RECT 142.000 31.600 142.800 32.400 ;
        RECT 143.600 32.300 144.400 32.400 ;
        RECT 143.600 31.700 145.900 32.300 ;
        RECT 143.600 31.600 144.400 31.700 ;
        RECT 143.600 29.600 144.400 30.400 ;
        RECT 142.000 27.600 142.800 28.400 ;
        RECT 142.100 26.400 142.700 27.600 ;
        RECT 142.000 25.600 142.800 26.400 ;
        RECT 127.600 11.800 128.400 12.600 ;
        RECT 135.600 6.200 136.400 17.800 ;
        RECT 140.400 17.600 141.200 18.400 ;
        RECT 142.100 12.400 142.700 25.600 ;
        RECT 145.300 20.400 145.900 31.700 ;
        RECT 148.400 31.600 149.200 32.400 ;
        RECT 148.500 30.400 149.100 31.600 ;
        RECT 153.300 30.400 153.900 43.600 ;
        RECT 156.500 32.400 157.100 49.600 ;
        RECT 159.700 48.400 160.300 55.600 ;
        RECT 164.500 52.400 165.100 57.600 ;
        RECT 170.900 52.400 171.500 65.600 ;
        RECT 175.700 56.400 176.300 71.600 ;
        RECT 178.900 70.400 179.500 97.600 ;
        RECT 183.700 88.400 184.300 129.600 ;
        RECT 199.700 128.400 200.300 129.600 ;
        RECT 185.200 127.600 186.000 128.400 ;
        RECT 199.600 127.600 200.400 128.400 ;
        RECT 185.300 112.400 185.900 127.600 ;
        RECT 196.400 125.600 197.200 126.400 ;
        RECT 190.000 123.600 190.800 124.400 ;
        RECT 202.800 123.600 203.600 124.400 ;
        RECT 212.400 124.200 213.200 137.800 ;
        RECT 214.000 124.200 214.800 137.800 ;
        RECT 215.600 124.200 216.400 137.800 ;
        RECT 217.200 126.200 218.000 137.800 ;
        RECT 218.900 136.400 219.500 145.600 ;
        RECT 220.500 144.400 221.100 167.600 ;
        RECT 220.400 143.600 221.200 144.400 ;
        RECT 222.000 144.200 222.800 155.800 ;
        RECT 228.400 149.600 229.200 150.400 ;
        RECT 218.800 135.600 219.600 136.400 ;
        RECT 220.400 126.200 221.200 137.800 ;
        RECT 222.000 133.600 222.800 134.400 ;
        RECT 190.100 112.400 190.700 123.600 ;
        RECT 212.400 121.600 213.200 122.400 ;
        RECT 199.600 119.600 200.400 120.400 ;
        RECT 199.700 118.400 200.300 119.600 ;
        RECT 199.600 117.600 200.400 118.400 ;
        RECT 185.200 111.600 186.000 112.400 ;
        RECT 190.000 111.600 190.800 112.400 ;
        RECT 193.200 111.600 194.000 112.400 ;
        RECT 196.400 111.600 197.200 112.400 ;
        RECT 207.600 111.600 208.400 112.400 ;
        RECT 193.200 109.600 194.000 110.400 ;
        RECT 199.600 109.600 200.400 110.400 ;
        RECT 202.800 109.600 203.600 110.400 ;
        RECT 193.300 108.400 193.900 109.600 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 193.200 107.600 194.000 108.400 ;
        RECT 194.800 107.600 195.600 108.400 ;
        RECT 201.200 107.600 202.000 108.400 ;
        RECT 194.900 106.400 195.500 107.600 ;
        RECT 202.900 106.400 203.500 109.600 ;
        RECT 210.800 107.600 211.600 108.400 ;
        RECT 186.800 106.300 187.600 106.400 ;
        RECT 185.300 105.700 187.600 106.300 ;
        RECT 183.600 87.600 184.400 88.400 ;
        RECT 182.000 85.600 182.800 86.400 ;
        RECT 178.800 69.600 179.600 70.400 ;
        RECT 180.400 67.600 181.200 68.400 ;
        RECT 182.100 68.300 182.700 85.600 ;
        RECT 185.300 74.300 185.900 105.700 ;
        RECT 186.800 105.600 187.600 105.700 ;
        RECT 194.800 105.600 195.600 106.400 ;
        RECT 202.800 105.600 203.600 106.400 ;
        RECT 204.400 103.600 205.200 104.400 ;
        RECT 186.800 84.200 187.600 97.800 ;
        RECT 188.400 84.200 189.200 97.800 ;
        RECT 190.000 84.200 190.800 97.800 ;
        RECT 191.600 86.200 192.400 97.800 ;
        RECT 193.200 95.600 194.000 96.400 ;
        RECT 193.300 92.400 193.900 95.600 ;
        RECT 193.200 91.600 194.000 92.400 ;
        RECT 186.800 81.600 187.600 82.400 ;
        RECT 186.900 78.400 187.500 81.600 ;
        RECT 186.800 77.600 187.600 78.400 ;
        RECT 183.700 73.700 185.900 74.300 ;
        RECT 183.700 72.400 184.300 73.700 ;
        RECT 193.300 72.400 193.900 91.600 ;
        RECT 194.800 86.200 195.600 97.800 ;
        RECT 196.400 93.600 197.200 94.400 ;
        RECT 198.000 86.200 198.800 97.800 ;
        RECT 199.600 84.200 200.400 97.800 ;
        RECT 201.200 84.200 202.000 97.800 ;
        RECT 204.500 94.400 205.100 103.600 ;
        RECT 210.900 96.400 211.500 107.600 ;
        RECT 212.500 106.400 213.100 121.600 ;
        RECT 222.100 120.400 222.700 133.600 ;
        RECT 223.600 126.200 224.400 137.800 ;
        RECT 225.200 124.200 226.000 137.800 ;
        RECT 226.800 124.200 227.600 137.800 ;
        RECT 230.100 132.400 230.700 171.600 ;
        RECT 231.600 164.200 232.400 177.800 ;
        RECT 233.200 164.200 234.000 177.800 ;
        RECT 234.800 164.200 235.600 177.800 ;
        RECT 236.400 166.200 237.200 177.800 ;
        RECT 238.000 175.600 238.800 176.400 ;
        RECT 238.100 162.400 238.700 175.600 ;
        RECT 239.600 166.200 240.400 177.800 ;
        RECT 241.200 173.600 242.000 174.400 ;
        RECT 233.200 161.600 234.000 162.400 ;
        RECT 238.000 161.600 238.800 162.400 ;
        RECT 231.600 144.200 232.400 155.800 ;
        RECT 233.300 148.400 233.900 161.600 ;
        RECT 241.300 158.400 241.900 173.600 ;
        RECT 242.800 166.200 243.600 177.800 ;
        RECT 244.400 164.200 245.200 177.800 ;
        RECT 246.000 164.200 246.800 177.800 ;
        RECT 258.800 177.600 259.600 178.400 ;
        RECT 260.500 178.300 261.100 187.600 ;
        RECT 270.000 183.600 270.800 184.400 ;
        RECT 279.600 184.200 280.400 197.800 ;
        RECT 281.200 184.200 282.000 197.800 ;
        RECT 282.800 184.200 283.600 197.800 ;
        RECT 284.400 184.200 285.200 195.800 ;
        RECT 286.000 185.600 286.800 186.400 ;
        RECT 270.100 178.400 270.700 183.600 ;
        RECT 286.100 182.300 286.700 185.600 ;
        RECT 287.600 184.200 288.400 195.800 ;
        RECT 289.200 187.600 290.000 188.400 ;
        RECT 290.800 184.200 291.600 195.800 ;
        RECT 292.400 184.200 293.200 197.800 ;
        RECT 294.000 184.200 294.800 197.800 ;
        RECT 303.600 197.600 304.400 198.400 ;
        RECT 300.400 189.600 301.200 190.400 ;
        RECT 305.200 185.600 306.000 186.400 ;
        RECT 286.100 181.700 288.300 182.300 ;
        RECT 262.000 178.300 262.800 178.400 ;
        RECT 260.500 177.700 262.800 178.300 ;
        RECT 262.000 177.600 262.800 177.700 ;
        RECT 270.000 177.600 270.800 178.400 ;
        RECT 258.900 176.400 259.500 177.600 ;
        RECT 258.800 175.600 259.600 176.400 ;
        RECT 265.200 175.600 266.000 176.400 ;
        RECT 255.600 173.600 256.400 174.400 ;
        RECT 263.600 173.600 264.400 174.400 ;
        RECT 255.700 172.400 256.300 173.600 ;
        RECT 265.300 172.400 265.900 175.600 ;
        RECT 250.800 171.600 251.600 172.400 ;
        RECT 255.600 171.600 256.400 172.400 ;
        RECT 265.200 171.600 266.000 172.400 ;
        RECT 274.800 171.600 275.600 172.400 ;
        RECT 255.600 169.600 256.400 170.400 ;
        RECT 241.200 157.600 242.000 158.400 ;
        RECT 233.200 147.600 234.000 148.400 ;
        RECT 233.300 146.400 233.900 147.600 ;
        RECT 233.200 145.600 234.000 146.400 ;
        RECT 234.800 146.200 235.600 151.800 ;
        RECT 246.000 151.600 246.800 152.400 ;
        RECT 246.100 150.400 246.700 151.600 ;
        RECT 236.400 149.600 237.200 150.400 ;
        RECT 238.000 149.600 238.800 150.400 ;
        RECT 242.800 149.600 243.600 150.400 ;
        RECT 246.000 149.600 246.800 150.400 ;
        RECT 247.600 149.600 248.400 150.400 ;
        RECT 252.400 149.600 253.200 150.400 ;
        RECT 236.500 140.400 237.100 149.600 ;
        RECT 242.900 148.400 243.500 149.600 ;
        RECT 242.800 147.600 243.600 148.400 ;
        RECT 249.200 147.600 250.000 148.400 ;
        RECT 249.300 146.400 249.900 147.600 ;
        RECT 249.200 145.600 250.000 146.400 ;
        RECT 252.500 144.400 253.100 149.600 ;
        RECT 241.200 143.600 242.000 144.400 ;
        RECT 252.400 143.600 253.200 144.400 ;
        RECT 239.600 141.600 240.400 142.400 ;
        RECT 236.400 139.600 237.200 140.400 ;
        RECT 239.700 132.400 240.300 141.600 ;
        RECT 230.000 131.600 230.800 132.400 ;
        RECT 239.600 131.600 240.400 132.400 ;
        RECT 238.000 127.600 238.800 128.400 ;
        RECT 230.000 123.600 230.800 124.400 ;
        RECT 236.400 123.600 237.200 124.400 ;
        RECT 222.000 119.600 222.800 120.400 ;
        RECT 223.600 119.600 224.400 120.400 ;
        RECT 223.700 118.400 224.300 119.600 ;
        RECT 218.800 117.600 219.600 118.400 ;
        RECT 223.600 117.600 224.400 118.400 ;
        RECT 214.000 111.600 214.800 112.400 ;
        RECT 217.200 112.300 218.000 112.400 ;
        RECT 217.200 111.700 219.500 112.300 ;
        RECT 217.200 111.600 218.000 111.700 ;
        RECT 212.400 105.600 213.200 106.400 ;
        RECT 210.800 95.600 211.600 96.400 ;
        RECT 204.400 93.600 205.200 94.400 ;
        RECT 210.800 94.300 211.600 94.400 ;
        RECT 212.500 94.300 213.100 105.600 ;
        RECT 214.100 98.400 214.700 111.600 ;
        RECT 218.900 110.400 219.500 111.700 ;
        RECT 222.000 111.600 222.800 112.400 ;
        RECT 222.100 110.400 222.700 111.600 ;
        RECT 217.200 109.600 218.000 110.400 ;
        RECT 218.800 109.600 219.600 110.400 ;
        RECT 222.000 109.600 222.800 110.400 ;
        RECT 226.800 109.600 227.600 110.400 ;
        RECT 217.200 107.600 218.000 108.400 ;
        RECT 228.400 108.300 229.200 108.400 ;
        RECT 230.100 108.300 230.700 123.600 ;
        RECT 238.100 122.300 238.700 127.600 ;
        RECT 236.500 121.700 238.700 122.300 ;
        RECT 236.500 118.400 237.100 121.700 ;
        RECT 236.400 117.600 237.200 118.400 ;
        RECT 238.000 117.600 238.800 118.400 ;
        RECT 238.100 112.400 238.700 117.600 ;
        RECT 239.700 114.400 240.300 131.600 ;
        RECT 241.300 130.400 241.900 143.600 ;
        RECT 242.800 139.600 243.600 140.400 ;
        RECT 242.900 138.400 243.500 139.600 ;
        RECT 255.700 138.400 256.300 169.600 ;
        RECT 257.400 151.800 258.200 152.600 ;
        RECT 263.600 151.800 264.400 152.600 ;
        RECT 274.900 152.400 275.500 171.600 ;
        RECT 279.600 164.200 280.400 177.800 ;
        RECT 281.200 164.200 282.000 177.800 ;
        RECT 282.800 166.200 283.600 177.800 ;
        RECT 284.400 173.600 285.200 174.400 ;
        RECT 286.000 166.200 286.800 177.800 ;
        RECT 287.700 176.400 288.300 181.700 ;
        RECT 287.600 175.600 288.400 176.400 ;
        RECT 257.400 147.000 258.000 151.800 ;
        RECT 258.600 149.800 259.400 150.600 ;
        RECT 258.800 148.400 259.400 149.800 ;
        RECT 260.400 149.600 261.200 150.400 ;
        RECT 263.800 148.400 264.400 151.800 ;
        RECT 274.800 151.600 275.600 152.400 ;
        RECT 258.800 147.800 264.400 148.400 ;
        RECT 258.800 147.000 259.600 147.200 ;
        RECT 262.200 147.000 263.000 147.200 ;
        RECT 263.800 147.000 264.400 147.800 ;
        RECT 265.200 147.600 266.000 148.400 ;
        RECT 257.400 146.400 263.000 147.000 ;
        RECT 257.400 146.200 258.200 146.400 ;
        RECT 263.600 146.200 264.400 147.000 ;
        RECT 265.300 144.400 265.900 147.600 ;
        RECT 273.200 145.600 274.000 146.400 ;
        RECT 265.200 143.600 266.000 144.400 ;
        RECT 242.800 137.600 243.600 138.400 ;
        RECT 255.600 137.600 256.400 138.400 ;
        RECT 268.400 137.600 269.200 138.400 ;
        RECT 246.000 135.600 246.800 136.400 ;
        RECT 249.200 135.600 250.000 136.400 ;
        RECT 252.400 135.600 253.200 136.400 ;
        RECT 246.100 134.400 246.700 135.600 ;
        RECT 246.000 133.600 246.800 134.400 ;
        RECT 249.300 132.400 249.900 135.600 ;
        RECT 249.200 131.600 250.000 132.400 ;
        RECT 255.600 131.600 256.400 132.400 ;
        RECT 271.600 131.600 272.400 132.400 ;
        RECT 241.200 129.600 242.000 130.400 ;
        RECT 241.300 124.400 241.900 129.600 ;
        RECT 244.400 127.600 245.200 128.400 ;
        RECT 244.500 124.400 245.100 127.600 ;
        RECT 241.200 123.600 242.000 124.400 ;
        RECT 242.800 123.600 243.600 124.400 ;
        RECT 244.400 123.600 245.200 124.400 ;
        RECT 241.200 119.600 242.000 120.400 ;
        RECT 239.600 113.600 240.400 114.400 ;
        RECT 238.000 111.600 238.800 112.400 ;
        RECT 239.600 111.600 240.400 112.400 ;
        RECT 238.100 108.400 238.700 111.600 ;
        RECT 239.700 110.400 240.300 111.600 ;
        RECT 241.300 110.400 241.900 119.600 ;
        RECT 242.900 118.400 243.500 123.600 ;
        RECT 242.800 117.600 243.600 118.400 ;
        RECT 244.500 112.400 245.100 123.600 ;
        RECT 249.300 120.400 249.900 131.600 ;
        RECT 260.400 129.600 261.200 130.400 ;
        RECT 250.800 123.600 251.600 124.400 ;
        RECT 249.200 119.600 250.000 120.400 ;
        RECT 252.400 119.600 253.200 120.400 ;
        RECT 244.400 111.600 245.200 112.400 ;
        RECT 249.200 111.600 250.000 112.400 ;
        RECT 252.500 110.400 253.100 119.600 ;
        RECT 260.500 116.400 261.100 129.600 ;
        RECT 273.300 128.300 273.900 145.600 ;
        RECT 274.900 138.400 275.500 151.600 ;
        RECT 279.600 144.200 280.400 157.800 ;
        RECT 281.200 144.200 282.000 157.800 ;
        RECT 282.800 144.200 283.600 155.800 ;
        RECT 284.400 147.600 285.200 148.400 ;
        RECT 279.600 141.600 280.400 142.400 ;
        RECT 284.500 142.300 285.100 147.600 ;
        RECT 286.000 144.200 286.800 155.800 ;
        RECT 287.700 146.400 288.300 175.600 ;
        RECT 289.200 166.200 290.000 177.800 ;
        RECT 290.800 164.200 291.600 177.800 ;
        RECT 292.400 164.200 293.200 177.800 ;
        RECT 294.000 164.200 294.800 177.800 ;
        RECT 295.600 171.600 296.400 172.400 ;
        RECT 305.200 171.600 306.000 172.400 ;
        RECT 295.700 164.400 296.300 171.600 ;
        RECT 295.600 163.600 296.400 164.400 ;
        RECT 303.600 164.300 304.400 164.400 ;
        RECT 302.100 163.700 304.400 164.300 ;
        RECT 287.600 145.600 288.400 146.400 ;
        RECT 289.200 144.200 290.000 155.800 ;
        RECT 290.800 144.200 291.600 157.800 ;
        RECT 292.400 144.200 293.200 157.800 ;
        RECT 294.000 144.200 294.800 157.800 ;
        RECT 282.900 141.700 285.100 142.300 ;
        RECT 279.700 138.400 280.300 141.600 ;
        RECT 274.800 137.600 275.600 138.400 ;
        RECT 279.600 137.600 280.400 138.400 ;
        RECT 274.800 135.600 275.600 136.400 ;
        RECT 279.600 133.600 280.400 134.400 ;
        RECT 279.700 132.400 280.300 133.600 ;
        RECT 279.600 131.600 280.400 132.400 ;
        RECT 279.600 129.600 280.400 130.400 ;
        RECT 279.700 128.400 280.300 129.600 ;
        RECT 271.700 127.700 273.900 128.300 ;
        RECT 260.400 115.600 261.200 116.400 ;
        RECT 257.200 113.600 258.000 114.400 ;
        RECT 258.800 113.600 259.600 114.400 ;
        RECT 239.600 109.600 240.400 110.400 ;
        RECT 241.200 109.600 242.000 110.400 ;
        RECT 252.400 109.600 253.200 110.400 ;
        RECT 228.400 107.700 230.700 108.300 ;
        RECT 228.400 107.600 229.200 107.700 ;
        RECT 233.200 107.600 234.000 108.400 ;
        RECT 238.000 107.600 238.800 108.400 ;
        RECT 239.600 107.600 240.400 108.400 ;
        RECT 250.800 107.600 251.600 108.400 ;
        RECT 217.300 106.400 217.900 107.600 ;
        RECT 217.200 105.600 218.000 106.400 ;
        RECT 220.400 105.600 221.200 106.400 ;
        RECT 225.200 106.300 226.000 106.400 ;
        RECT 225.200 105.700 227.500 106.300 ;
        RECT 225.200 105.600 226.000 105.700 ;
        RECT 214.000 97.600 214.800 98.400 ;
        RECT 217.200 95.600 218.000 96.400 ;
        RECT 214.000 94.300 214.800 94.400 ;
        RECT 210.800 93.700 214.800 94.300 ;
        RECT 210.800 93.600 211.600 93.700 ;
        RECT 214.000 93.600 214.800 93.700 ;
        RECT 217.300 92.400 217.900 95.600 ;
        RECT 206.000 91.600 206.800 92.400 ;
        RECT 217.200 91.600 218.000 92.400 ;
        RECT 183.600 71.600 184.400 72.400 ;
        RECT 185.200 71.600 186.000 72.400 ;
        RECT 193.200 71.600 194.000 72.400 ;
        RECT 194.800 71.800 195.600 72.600 ;
        RECT 201.400 71.800 202.200 72.600 ;
        RECT 183.700 70.400 184.300 71.600 ;
        RECT 183.600 69.600 184.400 70.400 ;
        RECT 185.300 68.400 185.900 71.600 ;
        RECT 193.200 69.600 194.000 70.400 ;
        RECT 193.300 68.400 193.900 69.600 ;
        RECT 194.800 68.400 195.400 71.800 ;
        RECT 198.800 68.400 199.600 68.600 ;
        RECT 182.100 67.700 184.300 68.300 ;
        RECT 180.500 66.400 181.100 67.600 ;
        RECT 180.400 65.600 181.200 66.400 ;
        RECT 177.200 63.600 178.000 64.400 ;
        RECT 182.000 63.600 182.800 64.400 ;
        RECT 175.600 55.600 176.400 56.400 ;
        RECT 162.800 51.600 163.600 52.400 ;
        RECT 164.400 51.600 165.200 52.400 ;
        RECT 170.800 51.600 171.600 52.400 ;
        RECT 159.600 47.600 160.400 48.400 ;
        RECT 148.400 29.600 149.200 30.400 ;
        RECT 150.000 29.600 150.800 30.400 ;
        RECT 153.200 29.600 154.000 30.400 ;
        RECT 146.800 27.600 147.600 28.400 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 145.200 19.600 146.000 20.400 ;
        RECT 145.300 16.400 145.900 19.600 ;
        RECT 146.900 16.400 147.500 27.600 ;
        RECT 154.800 26.200 155.600 31.800 ;
        RECT 156.400 31.600 157.200 32.400 ;
        RECT 158.000 24.200 158.800 35.800 ;
        RECT 159.600 29.400 160.400 30.400 ;
        RECT 162.900 18.400 163.500 51.600 ;
        RECT 167.600 49.600 168.400 50.400 ;
        RECT 169.200 49.600 170.000 50.400 ;
        RECT 167.700 48.400 168.300 49.600 ;
        RECT 167.600 47.600 168.400 48.400 ;
        RECT 169.300 38.400 169.900 49.600 ;
        RECT 175.700 48.400 176.300 55.600 ;
        RECT 170.800 47.600 171.600 48.400 ;
        RECT 172.400 47.600 173.200 48.400 ;
        RECT 175.600 47.600 176.400 48.400 ;
        RECT 170.900 46.400 171.500 47.600 ;
        RECT 170.800 45.600 171.600 46.400 ;
        RECT 175.600 41.600 176.400 42.400 ;
        RECT 175.700 38.400 176.300 41.600 ;
        RECT 169.200 37.600 170.000 38.400 ;
        RECT 172.400 37.600 173.200 38.400 ;
        RECT 175.600 37.600 176.400 38.400 ;
        RECT 166.000 29.600 166.800 30.400 ;
        RECT 164.400 19.600 165.200 20.400 ;
        RECT 162.800 17.600 163.600 18.400 ;
        RECT 145.200 15.600 146.000 16.400 ;
        RECT 146.800 15.600 147.600 16.400 ;
        RECT 148.200 15.000 149.000 15.800 ;
        RECT 150.000 15.000 154.200 15.600 ;
        RECT 154.800 15.000 155.600 15.800 ;
        RECT 159.600 15.600 160.400 16.400 ;
        RECT 142.000 11.600 142.800 12.400 ;
        RECT 148.200 10.200 148.800 15.000 ;
        RECT 150.000 14.800 150.800 15.000 ;
        RECT 153.400 14.800 154.200 15.000 ;
        RECT 155.000 14.200 155.600 15.000 ;
        RECT 150.800 13.600 155.600 14.200 ;
        RECT 156.400 13.600 157.200 14.400 ;
        RECT 150.800 13.400 151.600 13.600 ;
        RECT 155.000 10.200 155.600 13.600 ;
        RECT 156.500 12.400 157.100 13.600 ;
        RECT 164.500 12.400 165.100 19.600 ;
        RECT 166.100 18.400 166.700 29.600 ;
        RECT 167.600 24.200 168.400 35.800 ;
        RECT 177.300 30.400 177.900 63.600 ;
        RECT 182.100 52.400 182.700 63.600 ;
        RECT 182.000 51.600 182.800 52.400 ;
        RECT 183.700 38.400 184.300 67.700 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 193.200 67.600 194.000 68.400 ;
        RECT 194.800 67.800 199.600 68.400 ;
        RECT 194.800 67.000 195.400 67.800 ;
        RECT 196.200 67.000 197.000 67.200 ;
        RECT 199.600 67.000 200.400 67.200 ;
        RECT 201.600 67.000 202.200 71.800 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 204.400 67.600 205.200 68.400 ;
        RECT 191.600 65.600 192.400 66.400 ;
        RECT 194.800 66.200 195.600 67.000 ;
        RECT 196.200 66.400 200.400 67.000 ;
        RECT 201.400 66.200 202.200 67.000 ;
        RECT 206.100 66.400 206.700 91.600 ;
        RECT 220.500 90.400 221.100 105.600 ;
        RECT 225.200 101.600 226.000 102.400 ;
        RECT 223.600 99.600 224.400 100.400 ;
        RECT 223.700 98.400 224.300 99.600 ;
        RECT 223.600 97.600 224.400 98.400 ;
        RECT 225.300 94.400 225.900 101.600 ;
        RECT 225.200 93.600 226.000 94.400 ;
        RECT 226.900 92.400 227.500 105.700 ;
        RECT 231.600 105.600 232.400 106.400 ;
        RECT 231.700 104.400 232.300 105.600 ;
        RECT 231.600 103.600 232.400 104.400 ;
        RECT 233.300 102.400 233.900 107.600 ;
        RECT 230.000 101.600 230.800 102.400 ;
        RECT 233.200 101.600 234.000 102.400 ;
        RECT 230.100 98.400 230.700 101.600 ;
        RECT 239.700 100.400 240.300 107.600 ;
        RECT 242.800 103.600 243.600 104.400 ;
        RECT 249.200 103.600 250.000 104.400 ;
        RECT 239.600 99.600 240.400 100.400 ;
        RECT 230.000 97.600 230.800 98.400 ;
        RECT 231.600 95.600 232.400 96.400 ;
        RECT 231.700 94.400 232.300 95.600 ;
        RECT 233.200 95.000 234.000 95.800 ;
        RECT 239.400 95.600 240.200 95.800 ;
        RECT 234.600 95.000 240.200 95.600 ;
        RECT 231.600 93.600 232.400 94.400 ;
        RECT 233.200 94.200 233.800 95.000 ;
        RECT 234.600 94.800 235.400 95.000 ;
        RECT 238.000 94.800 238.800 95.000 ;
        RECT 233.200 93.600 238.800 94.200 ;
        RECT 226.800 91.600 227.600 92.400 ;
        RECT 220.400 89.600 221.200 90.400 ;
        RECT 233.200 90.200 233.800 93.600 ;
        RECT 238.200 92.200 238.800 93.600 ;
        RECT 238.200 91.400 239.000 92.200 ;
        RECT 239.600 90.200 240.200 95.000 ;
        RECT 242.900 90.400 243.500 103.600 ;
        RECT 249.300 94.400 249.900 103.600 ;
        RECT 250.900 94.400 251.500 107.600 ;
        RECT 247.600 93.600 248.400 94.400 ;
        RECT 249.200 93.600 250.000 94.400 ;
        RECT 250.800 93.600 251.600 94.400 ;
        RECT 252.500 92.400 253.100 109.600 ;
        RECT 255.600 105.600 256.400 106.400 ;
        RECT 255.700 98.400 256.300 105.600 ;
        RECT 255.600 97.600 256.400 98.400 ;
        RECT 252.400 91.600 253.200 92.400 ;
        RECT 233.200 89.400 234.000 90.200 ;
        RECT 239.400 89.400 240.200 90.200 ;
        RECT 242.800 89.600 243.600 90.400 ;
        RECT 238.000 83.600 238.800 84.400 ;
        RECT 249.200 83.600 250.000 84.400 ;
        RECT 231.600 73.600 232.400 74.400 ;
        RECT 231.700 72.400 232.300 73.600 ;
        RECT 231.600 71.600 232.400 72.400 ;
        RECT 223.600 69.600 224.400 70.400 ;
        RECT 230.000 69.600 230.800 70.400 ;
        RECT 239.600 69.600 240.400 70.400 ;
        RECT 212.400 67.600 213.200 68.400 ;
        RECT 234.800 67.600 235.600 68.400 ;
        RECT 206.000 65.600 206.800 66.400 ;
        RECT 196.400 63.600 197.200 64.400 ;
        RECT 186.800 44.200 187.600 57.800 ;
        RECT 188.400 44.200 189.200 57.800 ;
        RECT 190.000 44.200 190.800 57.800 ;
        RECT 191.600 46.200 192.400 57.800 ;
        RECT 193.200 55.600 194.000 56.400 ;
        RECT 194.800 46.200 195.600 57.800 ;
        RECT 196.500 54.400 197.100 63.600 ;
        RECT 212.500 58.400 213.100 67.600 ;
        RECT 226.800 65.600 227.600 66.400 ;
        RECT 215.600 63.600 216.400 64.400 ;
        RECT 220.400 63.600 221.200 64.400 ;
        RECT 231.600 63.600 232.400 64.400 ;
        RECT 196.400 53.600 197.200 54.400 ;
        RECT 198.000 46.200 198.800 57.800 ;
        RECT 199.600 44.200 200.400 57.800 ;
        RECT 201.200 44.200 202.000 57.800 ;
        RECT 212.400 57.600 213.200 58.400 ;
        RECT 215.700 56.400 216.300 63.600 ;
        RECT 214.000 55.600 214.800 56.400 ;
        RECT 215.600 55.600 216.400 56.400 ;
        RECT 206.000 51.600 206.800 52.400 ;
        RECT 206.100 50.400 206.700 51.600 ;
        RECT 206.000 49.600 206.800 50.400 ;
        RECT 212.400 45.600 213.200 46.400 ;
        RECT 183.600 37.600 184.400 38.400 ;
        RECT 214.100 38.300 214.700 55.600 ;
        RECT 220.500 52.400 221.100 63.600 ;
        RECT 231.700 60.300 232.300 63.600 ;
        RECT 234.900 62.400 235.500 67.600 ;
        RECT 239.700 66.400 240.300 69.600 ;
        RECT 239.600 65.600 240.400 66.400 ;
        RECT 244.400 64.200 245.200 77.800 ;
        RECT 246.000 64.200 246.800 77.800 ;
        RECT 247.600 64.200 248.400 75.800 ;
        RECT 249.300 68.400 249.900 83.600 ;
        RECT 258.900 80.400 259.500 113.600 ;
        RECT 260.500 112.400 261.100 115.600 ;
        RECT 268.400 113.600 269.200 114.400 ;
        RECT 260.400 111.600 261.200 112.400 ;
        RECT 266.800 107.600 267.600 108.400 ;
        RECT 263.600 91.600 264.400 92.400 ;
        RECT 258.800 79.600 259.600 80.400 ;
        RECT 249.200 67.600 250.000 68.400 ;
        RECT 249.200 65.600 250.000 66.400 ;
        RECT 234.800 61.600 235.600 62.400 ;
        RECT 230.100 59.700 232.300 60.300 ;
        RECT 218.800 51.600 219.600 52.400 ;
        RECT 220.400 51.600 221.200 52.400 ;
        RECT 218.900 50.400 219.500 51.600 ;
        RECT 218.800 49.600 219.600 50.400 ;
        RECT 188.200 31.800 189.000 32.600 ;
        RECT 194.800 31.800 195.600 32.600 ;
        RECT 177.200 29.600 178.000 30.400 ;
        RECT 185.200 29.600 186.000 30.400 ;
        RECT 186.800 29.600 187.600 30.400 ;
        RECT 185.300 28.400 185.900 29.600 ;
        RECT 186.900 28.400 187.500 29.600 ;
        RECT 180.400 27.600 181.200 28.400 ;
        RECT 185.200 27.600 186.000 28.400 ;
        RECT 186.800 27.600 187.600 28.400 ;
        RECT 180.500 26.400 181.100 27.600 ;
        RECT 188.200 27.000 188.800 31.800 ;
        RECT 190.800 28.400 191.600 28.600 ;
        RECT 195.000 28.400 195.600 31.800 ;
        RECT 198.000 29.600 198.800 30.400 ;
        RECT 207.600 29.600 208.400 30.400 ;
        RECT 198.100 28.400 198.700 29.600 ;
        RECT 190.800 27.800 195.600 28.400 ;
        RECT 190.000 27.000 190.800 27.200 ;
        RECT 193.400 27.000 194.200 27.200 ;
        RECT 195.000 27.000 195.600 27.800 ;
        RECT 196.400 27.600 197.200 28.400 ;
        RECT 198.000 27.600 198.800 28.400 ;
        RECT 174.000 25.600 174.800 26.400 ;
        RECT 180.400 25.600 181.200 26.400 ;
        RECT 182.000 25.600 182.800 26.400 ;
        RECT 188.200 26.200 189.000 27.000 ;
        RECT 190.000 26.400 194.200 27.000 ;
        RECT 194.800 26.200 195.600 27.000 ;
        RECT 166.000 17.600 166.800 18.400 ;
        RECT 174.100 16.400 174.700 25.600 ;
        RECT 178.800 23.600 179.600 24.400 ;
        RECT 178.900 20.400 179.500 23.600 ;
        RECT 178.800 19.600 179.600 20.400 ;
        RECT 167.600 15.600 168.400 16.400 ;
        RECT 174.000 15.600 174.800 16.400 ;
        RECT 156.400 11.600 157.200 12.400 ;
        RECT 164.400 11.600 165.200 12.400 ;
        RECT 148.200 9.400 149.000 10.200 ;
        RECT 154.800 9.400 155.600 10.200 ;
        RECT 177.200 4.200 178.000 17.800 ;
        RECT 178.800 4.200 179.600 17.800 ;
        RECT 180.400 4.200 181.200 17.800 ;
        RECT 182.000 6.200 182.800 17.800 ;
        RECT 183.600 17.600 184.400 18.400 ;
        RECT 183.700 16.400 184.300 17.600 ;
        RECT 183.600 15.600 184.400 16.400 ;
        RECT 185.200 6.200 186.000 17.800 ;
        RECT 186.800 13.600 187.600 14.400 ;
        RECT 188.400 6.200 189.200 17.800 ;
        RECT 190.000 4.200 190.800 17.800 ;
        RECT 191.600 4.200 192.400 17.800 ;
        RECT 207.700 16.400 208.300 29.600 ;
        RECT 209.200 24.200 210.000 37.800 ;
        RECT 210.800 24.200 211.600 37.800 ;
        RECT 212.400 24.200 213.200 37.800 ;
        RECT 214.100 37.700 216.300 38.300 ;
        RECT 214.000 24.200 214.800 35.800 ;
        RECT 215.700 26.400 216.300 37.700 ;
        RECT 215.600 25.600 216.400 26.400 ;
        RECT 215.700 20.300 216.300 25.600 ;
        RECT 217.200 24.200 218.000 35.800 ;
        RECT 218.900 30.400 219.500 49.600 ;
        RECT 225.200 44.200 226.000 57.800 ;
        RECT 226.800 44.200 227.600 57.800 ;
        RECT 228.400 46.200 229.200 57.800 ;
        RECT 230.100 54.400 230.700 59.700 ;
        RECT 230.000 53.600 230.800 54.400 ;
        RECT 231.600 46.200 232.400 57.800 ;
        RECT 233.200 55.600 234.000 56.400 ;
        RECT 233.300 38.400 233.900 55.600 ;
        RECT 234.800 46.200 235.600 57.800 ;
        RECT 236.400 44.200 237.200 57.800 ;
        RECT 238.000 44.200 238.800 57.800 ;
        RECT 239.600 44.200 240.400 57.800 ;
        RECT 249.300 38.400 249.900 65.600 ;
        RECT 250.800 64.200 251.600 75.800 ;
        RECT 252.400 65.600 253.200 66.400 ;
        RECT 254.000 64.200 254.800 75.800 ;
        RECT 255.600 64.200 256.400 77.800 ;
        RECT 257.200 64.200 258.000 77.800 ;
        RECT 258.800 64.200 259.600 77.800 ;
        RECT 263.700 76.400 264.300 91.600 ;
        RECT 265.200 84.200 266.000 97.800 ;
        RECT 266.800 84.200 267.600 97.800 ;
        RECT 268.400 84.200 269.200 97.800 ;
        RECT 270.000 86.200 270.800 97.800 ;
        RECT 271.700 96.400 272.300 127.700 ;
        RECT 279.600 127.600 280.400 128.400 ;
        RECT 282.900 122.400 283.500 141.700 ;
        RECT 289.200 141.600 290.000 142.400 ;
        RECT 284.400 139.600 285.200 140.400 ;
        RECT 284.500 130.400 285.100 139.600 ;
        RECT 289.300 136.400 289.900 141.600 ;
        RECT 302.100 140.400 302.700 163.700 ;
        RECT 303.600 163.600 304.400 163.700 ;
        RECT 305.300 154.400 305.900 171.600 ;
        RECT 305.200 153.600 306.000 154.400 ;
        RECT 306.800 151.600 307.600 152.400 ;
        RECT 306.900 150.400 307.500 151.600 ;
        RECT 306.800 149.600 307.600 150.400 ;
        RECT 303.600 147.600 304.600 148.400 ;
        RECT 305.200 147.600 306.000 148.400 ;
        RECT 303.600 145.600 304.400 146.400 ;
        RECT 302.000 139.600 302.800 140.400 ;
        RECT 303.700 138.400 304.300 145.600 ;
        RECT 305.300 142.400 305.900 147.600 ;
        RECT 305.200 141.600 306.000 142.400 ;
        RECT 303.600 137.600 304.400 138.400 ;
        RECT 289.200 135.600 290.000 136.400 ;
        RECT 295.600 135.600 296.400 136.400 ;
        RECT 305.200 135.600 306.000 136.400 ;
        RECT 289.300 134.400 289.900 135.600 ;
        RECT 295.700 134.400 296.300 135.600 ;
        RECT 305.300 134.400 305.900 135.600 ;
        RECT 289.200 133.600 290.000 134.400 ;
        RECT 294.000 133.600 294.800 134.400 ;
        RECT 295.600 133.600 296.400 134.400 ;
        RECT 305.200 133.600 306.000 134.400 ;
        RECT 287.600 131.600 288.400 132.400 ;
        RECT 294.100 130.400 294.700 133.600 ;
        RECT 295.600 131.600 296.400 132.400 ;
        RECT 284.400 129.600 285.200 130.400 ;
        RECT 290.800 129.600 291.600 130.400 ;
        RECT 294.000 129.600 294.800 130.400 ;
        RECT 294.000 127.600 294.800 128.400 ;
        RECT 282.800 121.600 283.600 122.400 ;
        RECT 295.700 120.400 296.300 131.600 ;
        RECT 297.200 129.600 298.000 130.400 ;
        RECT 300.400 129.600 301.200 130.400 ;
        RECT 302.000 129.600 302.800 130.400 ;
        RECT 302.100 126.400 302.700 129.600 ;
        RECT 302.000 125.600 302.800 126.400 ;
        RECT 306.900 120.400 307.500 149.600 ;
        RECT 308.500 130.400 309.100 223.600 ;
        RECT 310.100 218.400 310.700 223.600 ;
        RECT 310.000 217.600 310.800 218.400 ;
        RECT 310.000 211.600 310.800 212.400 ;
        RECT 310.000 189.600 310.800 190.400 ;
        RECT 311.700 168.300 312.300 227.600 ;
        RECT 313.200 225.600 314.000 226.400 ;
        RECT 313.300 218.400 313.900 225.600 ;
        RECT 318.100 220.400 318.700 241.600 ;
        RECT 319.700 228.400 320.300 275.600 ;
        RECT 321.200 257.600 322.000 258.400 ;
        RECT 321.300 250.400 321.900 257.600 ;
        RECT 322.900 252.300 323.500 287.600 ;
        RECT 326.000 283.600 326.800 284.400 ;
        RECT 330.900 272.300 331.500 295.600 ;
        RECT 332.500 294.400 333.100 303.600 ;
        RECT 335.600 301.600 336.400 302.400 ;
        RECT 335.700 294.400 336.300 301.600 ;
        RECT 332.400 293.600 333.200 294.400 ;
        RECT 335.600 293.600 336.400 294.400 ;
        RECT 337.300 290.400 337.900 307.600 ;
        RECT 332.400 289.600 333.200 290.400 ;
        RECT 337.200 289.600 338.000 290.400 ;
        RECT 332.500 288.400 333.100 289.600 ;
        RECT 338.900 288.400 339.500 321.600 ;
        RECT 340.500 314.400 341.100 323.600 ;
        RECT 345.300 320.400 345.900 329.700 ;
        RECT 346.900 326.400 347.500 331.600 ;
        RECT 353.300 328.400 353.900 331.600 ;
        RECT 353.200 327.600 354.000 328.400 ;
        RECT 354.900 326.400 355.500 331.600 ;
        RECT 361.300 330.400 361.900 331.600 ;
        RECT 367.700 330.400 368.300 331.600 ;
        RECT 375.700 330.400 376.300 333.600 ;
        RECT 378.800 331.600 379.600 332.400 ;
        RECT 378.900 330.400 379.500 331.600 ;
        RECT 380.500 330.400 381.100 333.600 ;
        RECT 382.100 330.400 382.700 349.600 ;
        RECT 386.800 347.600 387.600 348.400 ;
        RECT 385.200 345.600 386.000 346.400 ;
        RECT 383.600 339.600 384.400 340.400 ;
        RECT 383.700 334.400 384.300 339.600 ;
        RECT 386.900 334.400 387.500 347.600 ;
        RECT 390.100 334.400 390.700 401.600 ;
        RECT 394.900 400.400 395.500 403.600 ;
        RECT 406.100 402.400 406.700 403.600 ;
        RECT 406.000 401.600 406.800 402.400 ;
        RECT 391.600 399.600 392.400 400.400 ;
        RECT 394.800 399.600 395.600 400.400 ;
        RECT 391.700 374.300 392.300 399.600 ;
        RECT 393.200 384.200 394.000 397.800 ;
        RECT 394.800 384.200 395.600 397.800 ;
        RECT 396.400 384.200 397.200 395.800 ;
        RECT 398.000 387.600 398.800 388.400 ;
        RECT 398.100 384.400 398.700 387.600 ;
        RECT 398.000 383.600 398.800 384.400 ;
        RECT 399.600 384.200 400.400 395.800 ;
        RECT 401.200 385.600 402.000 386.400 ;
        RECT 399.600 381.600 400.400 382.400 ;
        RECT 399.700 378.400 400.300 381.600 ;
        RECT 399.600 377.600 400.400 378.400 ;
        RECT 398.000 375.600 398.800 376.400 ;
        RECT 391.700 373.700 393.900 374.300 ;
        RECT 393.300 372.400 393.900 373.700 ;
        RECT 393.200 371.600 394.000 372.400 ;
        RECT 393.300 370.400 393.900 371.600 ;
        RECT 391.600 369.600 392.400 370.400 ;
        RECT 393.200 369.600 394.000 370.400 ;
        RECT 391.700 334.400 392.300 369.600 ;
        RECT 394.800 367.600 395.600 368.400 ;
        RECT 393.200 365.600 394.000 366.400 ;
        RECT 398.100 362.400 398.700 375.600 ;
        RECT 401.300 370.300 401.900 385.600 ;
        RECT 402.800 384.200 403.600 395.800 ;
        RECT 404.400 384.200 405.200 397.800 ;
        RECT 406.000 384.200 406.800 397.800 ;
        RECT 407.600 384.200 408.400 397.800 ;
        RECT 407.600 381.600 408.400 382.400 ;
        RECT 407.700 378.400 408.300 381.600 ;
        RECT 407.600 377.600 408.400 378.400 ;
        RECT 412.500 372.400 413.100 407.600 ;
        RECT 417.200 393.600 418.000 394.400 ;
        RECT 425.300 382.400 425.900 411.600 ;
        RECT 426.800 404.200 427.600 417.800 ;
        RECT 428.400 404.200 429.200 417.800 ;
        RECT 430.000 404.200 430.800 417.800 ;
        RECT 431.600 406.200 432.400 417.800 ;
        RECT 433.200 415.600 434.000 416.400 ;
        RECT 434.800 406.200 435.600 417.800 ;
        RECT 436.500 414.400 437.100 419.600 ;
        RECT 436.400 413.600 437.200 414.400 ;
        RECT 438.000 406.200 438.800 417.800 ;
        RECT 439.600 404.200 440.400 417.800 ;
        RECT 441.200 404.200 442.000 417.800 ;
        RECT 447.600 411.600 448.400 412.400 ;
        RECT 431.600 399.600 432.400 400.400 ;
        RECT 431.700 390.400 432.300 399.600 ;
        RECT 449.300 390.400 449.900 419.600 ;
        RECT 450.900 412.400 451.500 429.600 ;
        RECT 463.600 427.600 464.400 428.400 ;
        RECT 452.400 423.600 453.200 424.400 ;
        RECT 452.500 416.400 453.100 423.600 ;
        RECT 470.100 422.400 470.700 443.600 ;
        RECT 478.000 439.600 478.800 440.400 ;
        RECT 473.200 424.200 474.000 437.800 ;
        RECT 474.800 424.200 475.600 437.800 ;
        RECT 476.400 424.200 477.200 435.800 ;
        RECT 478.100 428.400 478.700 439.600 ;
        RECT 482.900 438.400 483.500 451.600 ;
        RECT 484.500 440.400 485.100 451.600 ;
        RECT 486.000 449.600 486.800 450.400 ;
        RECT 486.100 444.400 486.700 449.600 ;
        RECT 495.700 448.400 496.300 451.600 ;
        RECT 489.200 447.600 490.000 448.400 ;
        RECT 495.600 448.300 496.400 448.400 ;
        RECT 494.100 447.700 496.400 448.300 ;
        RECT 486.000 443.600 486.800 444.400 ;
        RECT 484.400 439.600 485.200 440.400 ;
        RECT 482.800 437.600 483.600 438.400 ;
        RECT 478.000 427.600 478.800 428.400 ;
        RECT 479.600 424.200 480.400 435.800 ;
        RECT 481.200 425.600 482.000 426.400 ;
        RECT 482.800 424.200 483.600 435.800 ;
        RECT 484.400 424.200 485.200 437.800 ;
        RECT 486.000 424.200 486.800 437.800 ;
        RECT 487.600 424.200 488.400 437.800 ;
        RECT 470.000 421.600 470.800 422.400 ;
        RECT 484.400 421.600 485.200 422.400 ;
        RECT 452.400 415.600 453.200 416.400 ;
        RECT 450.800 411.600 451.600 412.400 ;
        RECT 454.000 411.600 454.800 412.400 ;
        RECT 455.600 411.600 456.400 412.400 ;
        RECT 426.800 389.600 427.600 390.400 ;
        RECT 431.600 389.600 432.400 390.400 ;
        RECT 439.600 389.600 440.400 390.400 ;
        RECT 442.800 389.600 443.600 390.400 ;
        RECT 449.200 389.600 450.000 390.400 ;
        RECT 425.200 381.600 426.000 382.400 ;
        RECT 426.900 380.400 427.500 389.600 ;
        RECT 428.400 387.600 429.200 388.400 ;
        RECT 436.400 387.600 437.200 388.400 ;
        RECT 441.200 387.600 442.000 388.400 ;
        RECT 428.500 386.400 429.100 387.600 ;
        RECT 428.400 385.600 429.200 386.400 ;
        RECT 426.800 379.600 427.600 380.400 ;
        RECT 402.800 371.600 403.600 372.400 ;
        RECT 412.400 371.600 413.200 372.400 ;
        RECT 425.200 371.600 426.000 372.400 ;
        RECT 401.300 369.700 403.500 370.300 ;
        RECT 402.900 364.400 403.500 369.700 ;
        RECT 417.200 365.600 418.000 366.400 ;
        RECT 422.000 365.600 422.800 366.400 ;
        RECT 401.200 363.600 402.000 364.400 ;
        RECT 402.800 363.600 403.600 364.400 ;
        RECT 398.000 361.600 398.800 362.400 ;
        RECT 401.300 358.400 401.900 363.600 ;
        RECT 396.400 344.200 397.200 357.800 ;
        RECT 398.000 344.200 398.800 357.800 ;
        RECT 399.600 344.200 400.400 357.800 ;
        RECT 401.200 357.600 402.000 358.400 ;
        RECT 401.200 344.200 402.000 355.800 ;
        RECT 402.900 346.400 403.500 363.600 ;
        RECT 402.800 345.600 403.600 346.400 ;
        RECT 404.400 344.200 405.200 355.800 ;
        RECT 406.000 347.600 406.800 348.400 ;
        RECT 406.000 345.600 406.800 346.400 ;
        RECT 398.000 337.600 398.800 338.400 ;
        RECT 383.600 333.600 384.400 334.400 ;
        RECT 386.800 333.600 387.600 334.400 ;
        RECT 390.000 333.600 390.800 334.400 ;
        RECT 391.600 333.600 392.400 334.400 ;
        RECT 396.400 333.600 397.200 334.400 ;
        RECT 390.100 332.400 390.700 333.600 ;
        RECT 398.100 332.400 398.700 337.600 ;
        RECT 399.600 335.600 400.400 336.400 ;
        RECT 399.700 334.400 400.300 335.600 ;
        RECT 399.600 333.600 400.400 334.400 ;
        RECT 401.200 333.600 402.000 334.400 ;
        RECT 402.800 333.600 403.600 334.400 ;
        RECT 402.900 332.400 403.500 333.600 ;
        RECT 388.400 331.600 389.200 332.400 ;
        RECT 390.000 331.600 390.800 332.400 ;
        RECT 391.600 331.600 392.400 332.400 ;
        RECT 398.000 331.600 398.800 332.400 ;
        RECT 402.800 331.600 403.600 332.400 ;
        RECT 404.400 331.600 405.200 332.400 ;
        RECT 361.200 329.600 362.000 330.400 ;
        RECT 366.000 329.600 366.800 330.400 ;
        RECT 367.600 329.600 368.400 330.400 ;
        RECT 375.600 329.600 376.400 330.400 ;
        RECT 378.800 329.600 379.600 330.400 ;
        RECT 380.400 329.600 381.200 330.400 ;
        RECT 382.000 329.600 382.800 330.400 ;
        RECT 366.100 326.400 366.700 329.600 ;
        RECT 375.700 328.400 376.300 329.600 ;
        RECT 375.600 327.600 376.400 328.400 ;
        RECT 388.500 328.300 389.100 331.600 ;
        RECT 391.700 330.400 392.300 331.600 ;
        RECT 391.600 329.600 392.400 330.400 ;
        RECT 393.200 329.600 394.000 330.400 ;
        RECT 393.300 328.300 393.900 329.600 ;
        RECT 404.500 328.400 405.100 331.600 ;
        RECT 406.100 330.400 406.700 345.600 ;
        RECT 407.600 344.200 408.400 355.800 ;
        RECT 409.200 344.200 410.000 357.800 ;
        RECT 410.800 344.200 411.600 357.800 ;
        RECT 422.100 354.400 422.700 365.600 ;
        RECT 423.600 357.600 424.400 358.400 ;
        RECT 422.000 353.600 422.800 354.400 ;
        RECT 415.600 349.600 416.400 350.400 ;
        RECT 414.000 347.600 414.800 348.400 ;
        RECT 414.100 338.400 414.700 347.600 ;
        RECT 422.100 338.400 422.700 353.600 ;
        RECT 414.000 337.600 414.800 338.400 ;
        RECT 422.000 337.600 422.800 338.400 ;
        RECT 407.600 335.600 408.400 336.400 ;
        RECT 412.400 335.600 413.200 336.400 ;
        RECT 407.700 334.400 408.300 335.600 ;
        RECT 412.500 334.400 413.100 335.600 ;
        RECT 407.600 333.600 408.400 334.400 ;
        RECT 410.800 333.600 411.600 334.400 ;
        RECT 412.400 333.600 413.200 334.400 ;
        RECT 422.000 333.600 422.800 334.400 ;
        RECT 423.700 332.400 424.300 357.600 ;
        RECT 425.300 350.400 425.900 371.600 ;
        RECT 426.800 364.200 427.600 377.800 ;
        RECT 428.400 364.200 429.200 377.800 ;
        RECT 430.000 364.200 430.800 377.800 ;
        RECT 431.600 366.200 432.400 377.800 ;
        RECT 433.200 375.600 434.000 376.400 ;
        RECT 433.300 364.400 433.900 375.600 ;
        RECT 434.800 366.200 435.600 377.800 ;
        RECT 436.400 373.600 437.200 374.400 ;
        RECT 433.200 363.600 434.000 364.400 ;
        RECT 436.500 362.400 437.100 373.600 ;
        RECT 438.000 366.200 438.800 377.800 ;
        RECT 439.600 364.200 440.400 377.800 ;
        RECT 441.200 364.200 442.000 377.800 ;
        RECT 433.200 361.600 434.000 362.400 ;
        RECT 436.400 361.600 437.200 362.400 ;
        RECT 433.300 358.400 433.900 361.600 ;
        RECT 442.900 358.400 443.500 389.600 ;
        RECT 447.600 387.600 448.400 388.400 ;
        RECT 449.200 383.600 450.000 384.400 ;
        RECT 446.000 371.600 446.800 372.400 ;
        RECT 449.300 368.400 449.900 383.600 ;
        RECT 452.400 375.600 453.200 376.400 ;
        RECT 449.200 367.600 450.000 368.400 ;
        RECT 428.400 357.600 429.200 358.400 ;
        RECT 433.200 357.600 434.000 358.400 ;
        RECT 442.800 357.600 443.600 358.400 ;
        RECT 452.500 358.300 453.100 375.600 ;
        RECT 455.700 372.400 456.300 411.600 ;
        RECT 458.800 404.200 459.600 417.800 ;
        RECT 460.400 404.200 461.200 417.800 ;
        RECT 462.000 406.200 462.800 417.800 ;
        RECT 463.600 417.600 464.400 418.400 ;
        RECT 463.700 414.400 464.300 417.600 ;
        RECT 463.600 413.600 464.400 414.400 ;
        RECT 465.200 406.200 466.000 417.800 ;
        RECT 466.800 415.600 467.600 416.400 ;
        RECT 468.400 406.200 469.200 417.800 ;
        RECT 470.000 404.200 470.800 417.800 ;
        RECT 471.600 404.200 472.400 417.800 ;
        RECT 473.200 404.200 474.000 417.800 ;
        RECT 474.800 407.600 475.600 408.400 ;
        RECT 457.200 389.600 458.000 390.400 ;
        RECT 457.300 372.400 457.900 389.600 ;
        RECT 458.800 384.200 459.600 397.800 ;
        RECT 460.400 384.200 461.200 397.800 ;
        RECT 462.000 384.200 462.800 397.800 ;
        RECT 463.600 384.200 464.400 395.800 ;
        RECT 465.200 385.600 466.000 386.400 ;
        RECT 463.600 381.600 464.400 382.400 ;
        RECT 465.300 382.300 465.900 385.600 ;
        RECT 466.800 384.200 467.600 395.800 ;
        RECT 468.400 387.600 469.200 388.400 ;
        RECT 468.500 384.400 469.100 387.600 ;
        RECT 468.400 383.600 469.200 384.400 ;
        RECT 470.000 384.200 470.800 395.800 ;
        RECT 471.600 384.200 472.400 397.800 ;
        RECT 473.200 384.200 474.000 397.800 ;
        RECT 465.300 381.700 467.500 382.300 ;
        RECT 455.600 371.600 456.400 372.400 ;
        RECT 457.200 371.600 458.000 372.400 ;
        RECT 428.500 350.400 429.100 357.600 ;
        RECT 434.800 351.600 435.600 352.400 ;
        RECT 425.200 349.600 426.000 350.400 ;
        RECT 428.400 349.600 429.200 350.400 ;
        RECT 426.800 347.600 427.600 348.400 ;
        RECT 430.000 348.300 430.800 348.400 ;
        RECT 428.500 347.700 430.800 348.300 ;
        RECT 426.900 346.400 427.500 347.600 ;
        RECT 426.800 345.600 427.600 346.400 ;
        RECT 426.800 335.600 427.600 336.400 ;
        RECT 428.500 334.400 429.100 347.700 ;
        RECT 430.000 347.600 430.800 347.700 ;
        RECT 431.600 347.600 432.400 348.400 ;
        RECT 431.700 346.400 432.300 347.600 ;
        RECT 431.600 345.600 432.400 346.400 ;
        RECT 433.200 343.600 434.000 344.400 ;
        RECT 438.000 343.600 438.800 344.400 ;
        RECT 447.600 344.200 448.400 357.800 ;
        RECT 449.200 344.200 450.000 357.800 ;
        RECT 450.800 344.200 451.600 357.800 ;
        RECT 452.500 357.700 454.700 358.300 ;
        RECT 452.400 344.200 453.200 355.800 ;
        RECT 454.100 346.400 454.700 357.700 ;
        RECT 454.000 345.600 454.800 346.400 ;
        RECT 428.400 333.600 429.200 334.400 ;
        RECT 409.200 331.600 410.000 332.400 ;
        RECT 423.600 331.600 424.400 332.400 ;
        RECT 430.000 331.600 430.800 332.400 ;
        RECT 433.300 330.400 433.900 343.600 ;
        RECT 454.100 340.300 454.700 345.600 ;
        RECT 455.600 344.200 456.400 355.800 ;
        RECT 457.300 350.400 457.900 371.600 ;
        RECT 458.800 364.200 459.600 377.800 ;
        RECT 460.400 364.200 461.200 377.800 ;
        RECT 462.000 366.200 462.800 377.800 ;
        RECT 463.700 374.400 464.300 381.600 ;
        RECT 463.600 373.600 464.400 374.400 ;
        RECT 465.200 366.200 466.000 377.800 ;
        RECT 466.900 376.400 467.500 381.700 ;
        RECT 466.800 375.600 467.600 376.400 ;
        RECT 468.400 366.200 469.200 377.800 ;
        RECT 470.000 364.200 470.800 377.800 ;
        RECT 471.600 364.200 472.400 377.800 ;
        RECT 473.200 364.200 474.000 377.800 ;
        RECT 457.200 349.600 458.000 350.400 ;
        RECT 457.200 347.600 458.000 348.400 ;
        RECT 457.300 346.400 457.900 347.600 ;
        RECT 457.200 345.600 458.000 346.400 ;
        RECT 458.800 344.200 459.600 355.800 ;
        RECT 460.400 344.200 461.200 357.800 ;
        RECT 462.000 344.200 462.800 357.800 ;
        RECT 474.900 354.400 475.500 407.600 ;
        RECT 482.800 403.600 483.600 404.400 ;
        RECT 478.000 389.600 478.800 390.400 ;
        RECT 478.100 386.400 478.700 389.600 ;
        RECT 484.500 388.400 485.100 421.600 ;
        RECT 489.300 414.400 489.900 447.600 ;
        RECT 492.400 417.600 493.200 418.400 ;
        RECT 486.000 413.600 486.800 414.400 ;
        RECT 489.200 413.600 490.000 414.400 ;
        RECT 487.600 411.600 488.400 412.400 ;
        RECT 489.200 411.600 490.000 412.400 ;
        RECT 487.600 403.600 488.400 404.400 ;
        RECT 487.700 396.400 488.300 403.600 ;
        RECT 487.600 395.600 488.400 396.400 ;
        RECT 487.700 394.400 488.300 395.600 ;
        RECT 486.000 393.600 486.800 394.400 ;
        RECT 487.600 393.600 488.400 394.400 ;
        RECT 486.100 392.400 486.700 393.600 ;
        RECT 486.000 391.600 486.800 392.400 ;
        RECT 486.000 389.600 486.800 390.400 ;
        RECT 482.800 387.600 483.600 388.400 ;
        RECT 484.400 387.600 485.200 388.400 ;
        RECT 478.000 385.600 478.800 386.400 ;
        RECT 484.400 383.600 485.200 384.400 ;
        RECT 486.100 374.400 486.700 389.600 ;
        RECT 487.600 383.600 488.400 384.400 ;
        RECT 486.000 373.600 486.800 374.400 ;
        RECT 482.800 369.600 483.600 370.400 ;
        RECT 481.200 357.600 482.000 358.400 ;
        RECT 474.800 353.600 475.600 354.400 ;
        RECT 481.300 352.400 481.900 357.600 ;
        RECT 481.200 351.600 482.000 352.400 ;
        RECT 463.600 349.600 464.400 350.400 ;
        RECT 466.800 349.600 467.600 350.400 ;
        RECT 478.000 349.600 478.800 350.400 ;
        RECT 452.500 339.700 454.700 340.300 ;
        RECT 434.800 333.600 435.600 334.400 ;
        RECT 406.000 329.600 406.800 330.400 ;
        RECT 415.600 329.600 416.400 330.400 ;
        RECT 426.800 329.600 427.600 330.400 ;
        RECT 433.200 329.600 434.000 330.400 ;
        RECT 436.400 329.600 437.200 330.400 ;
        RECT 388.500 327.700 393.900 328.300 ;
        RECT 404.400 327.600 405.200 328.400 ;
        RECT 346.800 325.600 347.600 326.400 ;
        RECT 354.800 325.600 355.600 326.400 ;
        RECT 366.000 325.600 366.800 326.400 ;
        RECT 369.200 325.600 370.000 326.400 ;
        RECT 345.200 319.600 346.000 320.400 ;
        RECT 340.400 313.600 341.200 314.400 ;
        RECT 343.600 311.600 344.400 312.400 ;
        RECT 342.000 309.600 342.800 310.400 ;
        RECT 342.100 306.400 342.700 309.600 ;
        RECT 343.700 308.400 344.300 311.600 ;
        RECT 343.600 307.600 344.400 308.400 ;
        RECT 345.300 306.400 345.900 319.600 ;
        RECT 346.900 316.400 347.500 325.600 ;
        RECT 353.200 317.600 354.000 318.400 ;
        RECT 369.200 317.600 370.000 318.400 ;
        RECT 346.800 315.600 347.600 316.400 ;
        RECT 348.400 309.600 349.200 310.400 ;
        RECT 353.300 308.400 353.900 317.600 ;
        RECT 358.000 311.600 358.800 312.400 ;
        RECT 362.800 311.600 363.600 312.400 ;
        RECT 358.100 310.400 358.700 311.600 ;
        RECT 358.000 309.600 358.800 310.400 ;
        RECT 361.200 309.600 362.000 310.400 ;
        RECT 362.800 309.600 363.600 310.400 ;
        RECT 361.300 308.400 361.900 309.600 ;
        RECT 346.800 307.600 347.600 308.400 ;
        RECT 353.200 307.600 354.000 308.400 ;
        RECT 359.600 307.600 360.400 308.400 ;
        RECT 361.200 307.600 362.000 308.400 ;
        RECT 342.000 305.600 342.800 306.400 ;
        RECT 345.200 305.600 346.000 306.400 ;
        RECT 332.400 287.600 333.200 288.400 ;
        RECT 338.800 287.600 339.600 288.400 ;
        RECT 337.200 283.600 338.000 284.400 ;
        RECT 334.000 275.600 334.800 276.400 ;
        RECT 332.400 272.300 333.200 272.400 ;
        RECT 330.900 271.700 333.200 272.300 ;
        RECT 332.400 271.600 333.200 271.700 ;
        RECT 326.000 267.600 327.000 268.400 ;
        RECT 335.600 267.600 336.400 268.400 ;
        RECT 332.400 263.600 333.200 264.400 ;
        RECT 327.600 257.600 328.400 258.400 ;
        RECT 327.700 254.400 328.300 257.600 ;
        RECT 329.200 255.600 330.000 256.400 ;
        RECT 326.000 253.600 326.800 254.400 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 324.400 252.300 325.200 252.400 ;
        RECT 322.900 251.700 325.200 252.300 ;
        RECT 321.200 249.600 322.000 250.400 ;
        RECT 322.900 242.400 323.500 251.700 ;
        RECT 324.400 251.600 325.200 251.700 ;
        RECT 326.000 251.600 326.800 252.400 ;
        RECT 324.400 250.300 325.200 250.400 ;
        RECT 326.100 250.300 326.700 251.600 ;
        RECT 324.400 249.700 326.700 250.300 ;
        RECT 324.400 249.600 325.200 249.700 ;
        RECT 327.700 248.400 328.300 253.600 ;
        RECT 332.500 252.400 333.100 263.600 ;
        RECT 334.000 253.600 334.800 254.400 ;
        RECT 335.600 253.600 336.400 254.400 ;
        RECT 329.200 251.600 330.000 252.400 ;
        RECT 332.400 251.600 333.200 252.400 ;
        RECT 327.600 247.600 328.400 248.400 ;
        RECT 335.700 246.400 336.300 253.600 ;
        RECT 337.300 248.400 337.900 283.600 ;
        RECT 342.100 282.400 342.700 305.600 ;
        RECT 345.200 303.600 346.000 304.400 ;
        RECT 343.600 301.600 344.400 302.400 ;
        RECT 343.700 288.400 344.300 301.600 ;
        RECT 345.300 296.400 345.900 303.600 ;
        RECT 345.200 295.600 346.000 296.400 ;
        RECT 345.200 293.600 346.000 294.400 ;
        RECT 345.300 292.400 345.900 293.600 ;
        RECT 345.200 291.600 346.000 292.400 ;
        RECT 343.600 287.600 344.400 288.400 ;
        RECT 340.400 281.600 341.200 282.400 ;
        RECT 342.000 281.600 342.800 282.400 ;
        RECT 340.500 274.400 341.100 281.600 ;
        RECT 343.600 277.600 344.400 278.400 ;
        RECT 342.000 275.600 342.800 276.400 ;
        RECT 340.400 273.600 341.200 274.400 ;
        RECT 340.400 271.600 341.200 272.400 ;
        RECT 342.100 270.400 342.700 275.600 ;
        RECT 343.700 272.300 344.300 277.600 ;
        RECT 345.300 276.400 345.900 291.600 ;
        RECT 346.900 290.400 347.500 307.600 ;
        RECT 358.000 305.600 358.800 306.400 ;
        RECT 362.900 302.400 363.500 309.600 ;
        RECT 362.800 301.600 363.600 302.400 ;
        RECT 369.200 301.600 370.000 302.400 ;
        RECT 369.300 298.400 369.900 301.600 ;
        RECT 369.200 297.600 370.000 298.400 ;
        RECT 370.800 297.600 371.600 298.400 ;
        RECT 356.400 295.600 357.200 296.400 ;
        RECT 359.600 295.600 360.400 296.400 ;
        RECT 364.400 295.600 365.200 296.400 ;
        RECT 356.500 292.400 357.100 295.600 ;
        RECT 359.700 294.400 360.300 295.600 ;
        RECT 359.600 293.600 360.400 294.400 ;
        RECT 356.400 291.600 357.200 292.400 ;
        RECT 361.200 291.600 362.000 292.400 ;
        RECT 362.800 291.600 363.600 292.400 ;
        RECT 346.800 289.600 347.600 290.400 ;
        RECT 348.400 287.600 349.200 288.400 ;
        RECT 351.600 287.600 352.400 288.400 ;
        RECT 348.500 284.400 349.100 287.600 ;
        RECT 361.300 286.400 361.900 291.600 ;
        RECT 361.200 285.600 362.000 286.400 ;
        RECT 346.800 283.600 347.600 284.400 ;
        RECT 348.400 283.600 349.200 284.400 ;
        RECT 350.000 283.600 350.800 284.400 ;
        RECT 346.900 282.300 347.500 283.600 ;
        RECT 346.900 281.700 349.100 282.300 ;
        RECT 346.800 279.600 347.600 280.400 ;
        RECT 345.200 275.600 346.000 276.400 ;
        RECT 346.900 272.400 347.500 279.600 ;
        RECT 348.500 278.300 349.100 281.700 ;
        RECT 350.100 280.400 350.700 283.600 ;
        RECT 350.000 279.600 350.800 280.400 ;
        RECT 362.900 278.400 363.500 291.600 ;
        RECT 348.500 277.700 350.700 278.300 ;
        RECT 350.100 276.300 350.700 277.700 ;
        RECT 358.000 277.600 358.800 278.400 ;
        RECT 362.800 277.600 363.600 278.400 ;
        RECT 350.100 275.700 352.300 276.300 ;
        RECT 345.200 272.300 346.000 272.400 ;
        RECT 343.700 271.700 346.000 272.300 ;
        RECT 345.200 271.600 346.000 271.700 ;
        RECT 346.800 271.600 347.600 272.400 ;
        RECT 340.400 269.600 341.200 270.400 ;
        RECT 342.000 269.600 342.800 270.400 ;
        RECT 350.000 269.600 350.800 270.400 ;
        RECT 340.500 254.400 341.100 269.600 ;
        RECT 343.600 265.600 344.400 266.400 ;
        RECT 348.400 265.600 349.200 266.400 ;
        RECT 346.800 263.600 347.600 264.400 ;
        RECT 346.900 256.400 347.500 263.600 ;
        RECT 346.800 255.600 347.600 256.400 ;
        RECT 338.800 253.600 339.600 254.400 ;
        RECT 340.400 253.600 341.200 254.400 ;
        RECT 338.900 250.400 339.500 253.600 ;
        RECT 338.800 249.600 339.600 250.400 ;
        RECT 337.200 247.600 338.000 248.400 ;
        RECT 342.000 247.600 342.800 248.400 ;
        RECT 335.600 245.600 336.400 246.400 ;
        RECT 337.200 243.600 338.000 244.400 ;
        RECT 322.800 241.600 323.600 242.400 ;
        RECT 337.300 240.400 337.900 243.600 ;
        RECT 337.200 239.600 338.000 240.400 ;
        RECT 322.800 229.600 323.600 230.400 ;
        RECT 319.600 227.600 320.400 228.400 ;
        RECT 322.900 228.300 323.500 229.600 ;
        RECT 322.900 227.700 325.100 228.300 ;
        RECT 321.200 221.600 322.000 222.400 ;
        RECT 318.000 219.600 318.800 220.400 ;
        RECT 318.100 218.400 318.700 219.600 ;
        RECT 313.200 217.600 314.000 218.400 ;
        RECT 318.000 217.600 318.800 218.400 ;
        RECT 313.300 210.400 313.900 217.600 ;
        RECT 321.300 212.400 321.900 221.600 ;
        RECT 324.500 218.400 325.100 227.700 ;
        RECT 326.000 224.200 326.800 237.800 ;
        RECT 327.600 224.200 328.400 237.800 ;
        RECT 329.200 224.200 330.000 235.800 ;
        RECT 330.800 231.600 331.600 232.400 ;
        RECT 330.900 228.400 331.500 231.600 ;
        RECT 330.800 227.600 331.600 228.400 ;
        RECT 332.400 224.200 333.200 235.800 ;
        RECT 334.000 225.600 334.800 226.400 ;
        RECT 334.100 220.300 334.700 225.600 ;
        RECT 335.600 224.200 336.400 235.800 ;
        RECT 337.200 224.200 338.000 237.800 ;
        RECT 338.800 224.200 339.600 237.800 ;
        RECT 340.400 224.200 341.200 237.800 ;
        RECT 334.100 219.700 336.300 220.300 ;
        RECT 324.400 217.600 325.200 218.400 ;
        RECT 330.800 217.600 331.600 218.400 ;
        RECT 330.900 212.400 331.500 217.600 ;
        RECT 334.000 215.600 334.800 216.400 ;
        RECT 332.400 213.600 333.200 214.400 ;
        RECT 332.500 212.400 333.100 213.600 ;
        RECT 321.200 211.600 322.000 212.400 ;
        RECT 327.600 211.600 328.400 212.400 ;
        RECT 330.800 211.600 331.600 212.400 ;
        RECT 332.400 211.600 333.200 212.400 ;
        RECT 327.700 210.400 328.300 211.600 ;
        RECT 313.200 209.600 314.000 210.400 ;
        RECT 327.600 209.600 328.400 210.400 ;
        RECT 334.000 209.600 334.800 210.400 ;
        RECT 334.100 206.400 334.700 209.600 ;
        RECT 335.700 208.400 336.300 219.700 ;
        RECT 342.100 216.400 342.700 247.600 ;
        RECT 348.500 224.400 349.100 265.600 ;
        RECT 350.100 262.400 350.700 269.600 ;
        RECT 351.700 268.300 352.300 275.700 ;
        RECT 362.800 273.600 363.600 274.400 ;
        RECT 362.900 272.400 363.500 273.600 ;
        RECT 361.200 271.600 362.000 272.400 ;
        RECT 362.800 271.600 363.600 272.400 ;
        RECT 358.000 270.300 358.800 270.400 ;
        RECT 361.200 270.300 362.000 270.400 ;
        RECT 358.000 269.700 362.000 270.300 ;
        RECT 358.000 269.600 358.800 269.700 ;
        RECT 361.200 269.600 362.000 269.700 ;
        RECT 367.600 269.600 368.400 270.400 ;
        RECT 354.800 268.300 355.600 268.400 ;
        RECT 351.700 267.700 355.600 268.300 ;
        RECT 354.800 267.600 355.600 267.700 ;
        RECT 354.800 265.600 355.600 266.400 ;
        RECT 367.700 262.400 368.300 269.600 ;
        RECT 370.900 268.400 371.500 297.600 ;
        RECT 375.700 292.400 376.300 327.600 ;
        RECT 378.800 304.200 379.600 317.800 ;
        RECT 380.400 304.200 381.200 317.800 ;
        RECT 382.000 304.200 382.800 317.800 ;
        RECT 383.600 304.200 384.400 315.800 ;
        RECT 385.200 305.600 386.000 306.400 ;
        RECT 375.600 291.600 376.400 292.400 ;
        RECT 375.600 283.600 376.400 284.400 ;
        RECT 378.800 284.200 379.600 297.800 ;
        RECT 380.400 284.200 381.200 297.800 ;
        RECT 382.000 284.200 382.800 297.800 ;
        RECT 383.600 286.200 384.400 297.800 ;
        RECT 385.300 296.400 385.900 305.600 ;
        RECT 386.800 304.200 387.600 315.800 ;
        RECT 388.400 307.600 389.200 308.400 ;
        RECT 388.500 306.400 389.100 307.600 ;
        RECT 388.400 305.600 389.200 306.400 ;
        RECT 390.000 304.200 390.800 315.800 ;
        RECT 391.600 304.200 392.400 317.800 ;
        RECT 393.200 304.200 394.000 317.800 ;
        RECT 394.800 309.600 395.600 310.400 ;
        RECT 385.200 295.600 386.000 296.400 ;
        RECT 386.800 286.200 387.600 297.800 ;
        RECT 388.400 293.600 389.200 294.400 ;
        RECT 390.000 286.200 390.800 297.800 ;
        RECT 391.600 284.200 392.400 297.800 ;
        RECT 393.200 284.200 394.000 297.800 ;
        RECT 394.900 292.400 395.500 309.600 ;
        RECT 394.800 291.600 395.600 292.400 ;
        RECT 402.800 291.600 403.600 292.400 ;
        RECT 404.400 291.600 405.200 292.400 ;
        RECT 375.700 272.400 376.300 283.600 ;
        RECT 394.900 278.400 395.500 291.600 ;
        RECT 398.000 281.600 398.800 282.400 ;
        RECT 378.800 277.600 379.600 278.400 ;
        RECT 394.800 277.600 395.600 278.400 ;
        RECT 375.600 271.600 376.400 272.400 ;
        RECT 377.200 271.600 378.000 272.400 ;
        RECT 370.800 267.600 371.600 268.400 ;
        RECT 370.800 265.600 371.600 266.400 ;
        RECT 374.000 263.600 374.800 264.400 ;
        RECT 350.000 261.600 350.800 262.400 ;
        RECT 361.300 261.700 365.100 262.300 ;
        RECT 361.300 256.300 361.900 261.700 ;
        RECT 364.500 260.400 365.100 261.700 ;
        RECT 367.600 261.600 368.400 262.400 ;
        RECT 364.400 259.600 365.200 260.400 ;
        RECT 359.700 255.700 361.900 256.300 ;
        RECT 359.700 254.400 360.300 255.700 ;
        RECT 367.700 254.400 368.300 261.600 ;
        RECT 369.200 257.600 370.000 258.400 ;
        RECT 369.300 254.400 369.900 257.600 ;
        RECT 372.400 255.600 373.200 256.400 ;
        RECT 353.200 253.600 354.000 254.400 ;
        RECT 359.600 253.600 360.400 254.400 ;
        RECT 361.200 253.600 362.000 254.400 ;
        RECT 367.600 253.600 368.400 254.400 ;
        RECT 369.200 253.600 370.000 254.400 ;
        RECT 351.600 247.600 352.400 248.400 ;
        RECT 350.000 227.600 350.800 228.400 ;
        RECT 348.400 223.600 349.200 224.400 ;
        RECT 350.100 218.400 350.700 227.600 ;
        RECT 351.700 226.400 352.300 247.600 ;
        RECT 353.300 236.300 353.900 253.600 ;
        RECT 359.600 251.600 360.400 252.400 ;
        RECT 354.800 249.600 355.600 250.400 ;
        RECT 358.000 250.300 358.800 250.400 ;
        RECT 359.700 250.300 360.300 251.600 ;
        RECT 358.000 249.700 360.300 250.300 ;
        RECT 358.000 249.600 358.800 249.700 ;
        RECT 354.900 248.400 355.500 249.600 ;
        RECT 354.800 247.600 355.600 248.400 ;
        RECT 361.300 242.400 361.900 253.600 ;
        RECT 372.500 252.400 373.100 255.600 ;
        RECT 374.100 254.400 374.700 263.600 ;
        RECT 374.000 253.600 374.800 254.400 ;
        RECT 366.000 251.600 366.800 252.400 ;
        RECT 367.600 251.600 368.400 252.400 ;
        RECT 372.400 251.600 373.200 252.400 ;
        RECT 366.100 244.400 366.700 251.600 ;
        RECT 362.800 243.600 363.600 244.400 ;
        RECT 366.000 243.600 366.800 244.400 ;
        RECT 361.200 241.600 362.000 242.400 ;
        RECT 354.800 239.600 355.600 240.400 ;
        RECT 354.900 238.400 355.500 239.600 ;
        RECT 354.800 237.600 355.600 238.400 ;
        RECT 353.300 235.700 355.500 236.300 ;
        RECT 353.200 227.600 354.000 228.400 ;
        RECT 351.600 225.600 352.400 226.400 ;
        RECT 350.000 217.600 350.800 218.400 ;
        RECT 337.200 215.600 338.000 216.400 ;
        RECT 342.000 215.600 342.800 216.400 ;
        RECT 337.300 214.400 337.900 215.600 ;
        RECT 337.200 213.600 338.000 214.400 ;
        RECT 342.000 213.600 342.800 214.400 ;
        RECT 345.200 213.600 346.000 214.400 ;
        RECT 342.100 212.400 342.700 213.600 ;
        RECT 345.300 212.400 345.900 213.600 ;
        RECT 337.200 211.600 338.000 212.400 ;
        RECT 342.000 211.600 342.800 212.400 ;
        RECT 345.200 211.600 346.000 212.400 ;
        RECT 338.800 209.600 339.600 210.400 ;
        RECT 346.800 209.600 347.600 210.400 ;
        RECT 348.400 209.600 349.200 210.400 ;
        RECT 350.000 209.600 350.800 210.400 ;
        RECT 335.600 207.600 336.400 208.400 ;
        RECT 334.000 205.600 334.800 206.400 ;
        RECT 324.400 203.600 325.200 204.400 ;
        RECT 330.800 203.600 331.600 204.400 ;
        RECT 322.800 199.600 323.600 200.400 ;
        RECT 314.800 184.200 315.600 197.800 ;
        RECT 316.400 184.200 317.200 197.800 ;
        RECT 318.000 184.200 318.800 195.800 ;
        RECT 319.600 189.600 320.400 190.400 ;
        RECT 319.700 188.400 320.300 189.600 ;
        RECT 319.600 187.600 320.400 188.400 ;
        RECT 321.200 184.200 322.000 195.800 ;
        RECT 322.900 186.400 323.500 199.600 ;
        RECT 324.500 198.400 325.100 203.600 ;
        RECT 324.400 197.600 325.200 198.400 ;
        RECT 322.800 185.600 323.600 186.400 ;
        RECT 324.400 184.200 325.200 195.800 ;
        RECT 326.000 184.200 326.800 197.800 ;
        RECT 327.600 184.200 328.400 197.800 ;
        RECT 329.200 184.200 330.000 197.800 ;
        RECT 330.900 192.400 331.500 203.600 ;
        RECT 330.800 191.600 331.600 192.400 ;
        RECT 335.700 180.400 336.300 207.600 ;
        RECT 338.900 204.400 339.500 209.600 ;
        RECT 338.800 203.600 339.600 204.400 ;
        RECT 345.200 203.600 346.000 204.400 ;
        RECT 340.400 191.600 341.200 192.400 ;
        RECT 345.300 190.400 345.900 203.600 ;
        RECT 346.900 192.400 347.500 209.600 ;
        RECT 346.800 191.600 347.600 192.400 ;
        RECT 340.400 189.600 341.200 190.400 ;
        RECT 345.200 189.600 346.000 190.400 ;
        RECT 338.800 187.600 339.800 188.400 ;
        RECT 335.600 179.600 336.400 180.400 ;
        RECT 340.400 179.600 341.200 180.400 ;
        RECT 314.800 175.600 315.600 176.400 ;
        RECT 313.200 173.600 314.000 174.400 ;
        RECT 316.400 173.600 317.200 174.400 ;
        RECT 318.000 173.600 318.800 174.400 ;
        RECT 316.500 172.400 317.100 173.600 ;
        RECT 316.400 171.600 317.200 172.400 ;
        RECT 319.600 171.600 320.400 172.400 ;
        RECT 321.200 171.600 322.000 172.400 ;
        RECT 329.200 171.600 330.000 172.400 ;
        RECT 313.200 169.600 314.000 170.400 ;
        RECT 311.700 167.700 313.900 168.300 ;
        RECT 311.600 153.600 312.400 154.400 ;
        RECT 311.600 143.600 312.400 144.400 ;
        RECT 311.700 136.400 312.300 143.600 ;
        RECT 311.600 135.600 312.400 136.400 ;
        RECT 308.400 129.600 309.200 130.400 ;
        RECT 295.600 119.600 296.400 120.400 ;
        RECT 297.200 119.600 298.000 120.400 ;
        RECT 306.800 119.600 307.600 120.400 ;
        RECT 278.000 104.200 278.800 117.800 ;
        RECT 279.600 104.200 280.400 117.800 ;
        RECT 281.200 104.200 282.000 117.800 ;
        RECT 282.800 104.200 283.600 115.800 ;
        RECT 284.400 105.600 285.200 106.400 ;
        RECT 286.000 104.200 286.800 115.800 ;
        RECT 287.600 107.600 288.400 108.400 ;
        RECT 289.200 104.200 290.000 115.800 ;
        RECT 290.800 104.200 291.600 117.800 ;
        RECT 292.400 104.200 293.200 117.800 ;
        RECT 295.600 109.600 296.400 110.400 ;
        RECT 295.700 102.400 296.300 109.600 ;
        RECT 292.400 101.600 293.200 102.400 ;
        RECT 295.600 101.600 296.400 102.400 ;
        RECT 292.500 98.400 293.100 101.600 ;
        RECT 271.600 95.600 272.400 96.400 ;
        RECT 271.700 80.400 272.300 95.600 ;
        RECT 273.200 86.200 274.000 97.800 ;
        RECT 274.800 93.600 275.600 94.400 ;
        RECT 276.400 86.200 277.200 97.800 ;
        RECT 278.000 84.200 278.800 97.800 ;
        RECT 279.600 84.200 280.400 97.800 ;
        RECT 292.400 97.600 293.200 98.400 ;
        RECT 295.600 95.600 296.400 96.400 ;
        RECT 295.700 94.400 296.300 95.600 ;
        RECT 295.600 93.600 296.400 94.400 ;
        RECT 297.300 92.400 297.900 119.600 ;
        RECT 313.300 118.400 313.900 167.700 ;
        RECT 319.700 152.400 320.300 171.600 ;
        RECT 322.800 169.600 323.600 170.400 ;
        RECT 329.300 164.400 329.900 171.600 ;
        RECT 329.200 163.600 330.000 164.400 ;
        RECT 332.400 164.200 333.200 177.800 ;
        RECT 334.000 164.200 334.800 177.800 ;
        RECT 335.600 166.200 336.400 177.800 ;
        RECT 337.200 175.600 338.000 176.400 ;
        RECT 337.300 174.400 337.900 175.600 ;
        RECT 337.200 173.600 338.000 174.400 ;
        RECT 338.800 166.200 339.600 177.800 ;
        RECT 340.500 176.400 341.100 179.600 ;
        RECT 340.400 175.600 341.200 176.400 ;
        RECT 319.600 151.600 320.400 152.400 ;
        RECT 321.200 144.200 322.000 157.800 ;
        RECT 322.800 144.200 323.600 157.800 ;
        RECT 324.400 144.200 325.200 155.800 ;
        RECT 326.000 147.600 326.800 148.400 ;
        RECT 326.100 146.400 326.700 147.600 ;
        RECT 326.000 145.600 326.800 146.400 ;
        RECT 327.600 144.200 328.400 155.800 ;
        RECT 329.200 145.600 330.000 146.400 ;
        RECT 330.800 144.200 331.600 155.800 ;
        RECT 332.400 144.200 333.200 157.800 ;
        RECT 334.000 144.200 334.800 157.800 ;
        RECT 335.600 144.200 336.400 157.800 ;
        RECT 337.200 149.600 338.000 150.400 ;
        RECT 318.000 124.200 318.800 137.800 ;
        RECT 319.600 124.200 320.400 137.800 ;
        RECT 321.200 124.200 322.000 137.800 ;
        RECT 322.800 126.200 323.600 137.800 ;
        RECT 324.400 135.600 325.200 136.400 ;
        RECT 318.000 119.600 318.800 120.400 ;
        RECT 313.200 117.600 314.000 118.400 ;
        RECT 318.100 110.400 318.700 119.600 ;
        RECT 322.800 113.600 323.600 114.400 ;
        RECT 302.000 109.600 302.800 110.400 ;
        RECT 308.400 109.600 309.200 110.400 ;
        RECT 318.000 109.600 318.800 110.400 ;
        RECT 306.800 107.600 307.600 108.400 ;
        RECT 311.600 107.600 312.400 108.400 ;
        RECT 316.400 107.600 317.200 108.400 ;
        RECT 305.200 93.600 306.000 94.400 ;
        RECT 289.200 91.600 290.000 92.400 ;
        RECT 297.200 91.600 298.000 92.400 ;
        RECT 271.600 79.600 272.400 80.400 ;
        RECT 278.000 79.600 278.800 80.400 ;
        RECT 278.100 78.400 278.700 79.600 ;
        RECT 268.400 77.600 269.200 78.400 ;
        RECT 278.000 77.600 278.800 78.400 ;
        RECT 260.400 75.600 261.200 76.400 ;
        RECT 263.600 75.600 264.400 76.400 ;
        RECT 260.500 70.400 261.100 75.600 ;
        RECT 289.300 70.400 289.900 91.600 ;
        RECT 290.800 73.600 291.600 74.400 ;
        RECT 290.900 72.400 291.500 73.600 ;
        RECT 290.800 71.600 291.600 72.400 ;
        RECT 297.300 70.400 297.900 91.600 ;
        RECT 302.000 89.600 302.800 90.400 ;
        RECT 305.200 89.600 306.000 90.400 ;
        RECT 300.400 73.600 301.200 74.400 ;
        RECT 260.400 69.600 261.200 70.400 ;
        RECT 289.200 69.600 290.000 70.400 ;
        RECT 294.000 69.600 294.800 70.400 ;
        RECT 297.200 69.600 298.000 70.400 ;
        RECT 298.800 69.600 299.600 70.400 ;
        RECT 252.400 61.600 253.200 62.400 ;
        RECT 252.500 58.400 253.100 61.600 ;
        RECT 252.400 57.600 253.200 58.400 ;
        RECT 255.600 57.600 256.400 58.400 ;
        RECT 255.700 52.400 256.300 57.600 ;
        RECT 257.200 55.600 258.000 56.400 ;
        RECT 257.300 54.400 257.900 55.600 ;
        RECT 257.200 53.600 258.000 54.400 ;
        RECT 260.500 52.400 261.100 69.600 ;
        RECT 294.100 68.400 294.700 69.600 ;
        RECT 289.200 67.600 290.000 68.400 ;
        RECT 294.000 67.600 294.800 68.400 ;
        RECT 295.600 67.600 296.400 68.400 ;
        RECT 287.600 63.600 288.400 64.400 ;
        RECT 255.600 51.600 256.400 52.400 ;
        RECT 260.400 51.600 261.200 52.400 ;
        RECT 266.800 51.600 267.600 52.400 ;
        RECT 252.400 47.600 253.200 48.400 ;
        RECT 252.500 40.400 253.100 47.600 ;
        RECT 271.600 44.200 272.400 57.800 ;
        RECT 273.200 44.200 274.000 57.800 ;
        RECT 274.800 46.200 275.600 57.800 ;
        RECT 276.400 53.600 277.200 54.400 ;
        RECT 278.000 46.200 278.800 57.800 ;
        RECT 279.600 55.600 280.400 56.400 ;
        RECT 252.400 39.600 253.200 40.400 ;
        RECT 278.000 39.600 278.800 40.400 ;
        RECT 218.800 29.600 219.600 30.400 ;
        RECT 218.800 27.600 219.600 28.400 ;
        RECT 220.400 24.200 221.200 35.800 ;
        RECT 222.000 24.200 222.800 37.800 ;
        RECT 223.600 24.200 224.400 37.800 ;
        RECT 233.200 37.600 234.000 38.400 ;
        RECT 234.800 29.600 235.600 30.400 ;
        RECT 215.700 19.700 217.900 20.300 ;
        RECT 217.300 18.400 217.900 19.700 ;
        RECT 196.400 15.600 197.200 16.400 ;
        RECT 207.600 15.600 208.400 16.400 ;
        RECT 196.500 12.400 197.100 15.600 ;
        RECT 196.400 11.600 197.200 12.400 ;
        RECT 202.800 11.600 203.600 12.400 ;
        RECT 202.900 10.400 203.500 11.600 ;
        RECT 202.800 9.600 203.600 10.400 ;
        RECT 209.200 4.200 210.000 17.800 ;
        RECT 210.800 4.200 211.600 17.800 ;
        RECT 212.400 6.200 213.200 17.800 ;
        RECT 214.000 15.600 214.800 16.400 ;
        RECT 214.100 14.400 214.700 15.600 ;
        RECT 214.000 13.600 214.800 14.400 ;
        RECT 215.600 6.200 216.400 17.800 ;
        RECT 217.200 17.600 218.000 18.400 ;
        RECT 217.300 16.400 217.900 17.600 ;
        RECT 217.200 15.600 218.000 16.400 ;
        RECT 218.800 6.200 219.600 17.800 ;
        RECT 220.400 4.200 221.200 17.800 ;
        RECT 222.000 4.200 222.800 17.800 ;
        RECT 223.600 4.200 224.400 17.800 ;
        RECT 234.900 12.400 235.500 29.600 ;
        RECT 241.200 24.200 242.000 37.800 ;
        RECT 242.800 24.200 243.600 37.800 ;
        RECT 249.200 37.600 250.000 38.400 ;
        RECT 244.400 24.200 245.200 35.800 ;
        RECT 246.000 29.600 246.800 30.400 ;
        RECT 246.100 28.400 246.700 29.600 ;
        RECT 246.000 27.600 246.800 28.400 ;
        RECT 247.600 24.200 248.400 35.800 ;
        RECT 249.300 26.400 249.900 37.600 ;
        RECT 249.200 25.600 250.000 26.400 ;
        RECT 250.800 24.200 251.600 35.800 ;
        RECT 252.400 24.200 253.200 37.800 ;
        RECT 254.000 24.200 254.800 37.800 ;
        RECT 255.600 24.200 256.400 37.800 ;
        RECT 278.100 34.300 278.700 39.600 ;
        RECT 279.700 38.400 280.300 55.600 ;
        RECT 281.200 46.200 282.000 57.800 ;
        RECT 282.800 44.200 283.600 57.800 ;
        RECT 284.400 44.200 285.200 57.800 ;
        RECT 286.000 44.200 286.800 57.800 ;
        RECT 287.700 52.400 288.300 63.600 ;
        RECT 287.600 51.600 288.400 52.400 ;
        RECT 287.600 49.600 288.400 50.400 ;
        RECT 279.600 37.600 280.400 38.400 ;
        RECT 278.100 33.700 280.300 34.300 ;
        RECT 279.700 32.400 280.300 33.700 ;
        RECT 287.700 32.400 288.300 49.600 ;
        RECT 279.600 31.600 280.400 32.400 ;
        RECT 287.600 31.600 288.400 32.400 ;
        RECT 289.300 30.400 289.900 67.600 ;
        RECT 292.400 65.600 293.200 66.400 ;
        RECT 295.700 56.400 296.300 67.600 ;
        RECT 297.300 58.400 297.900 69.600 ;
        RECT 298.800 61.600 299.600 62.400 ;
        RECT 297.200 57.600 298.000 58.400 ;
        RECT 295.600 55.600 296.400 56.400 ;
        RECT 297.200 53.600 298.000 54.400 ;
        RECT 298.900 50.400 299.500 61.600 ;
        RECT 302.100 56.400 302.700 89.600 ;
        RECT 305.300 82.400 305.900 89.600 ;
        RECT 305.200 81.600 306.000 82.400 ;
        RECT 305.200 69.600 306.000 70.400 ;
        RECT 305.300 64.400 305.900 69.600 ;
        RECT 306.900 68.400 307.500 107.600 ;
        RECT 311.700 96.400 312.300 107.600 ;
        RECT 324.500 106.400 325.100 135.600 ;
        RECT 326.000 126.200 326.800 137.800 ;
        RECT 327.600 133.600 328.400 134.400 ;
        RECT 327.700 128.400 328.300 133.600 ;
        RECT 327.600 127.600 328.400 128.400 ;
        RECT 329.200 126.200 330.000 137.800 ;
        RECT 330.800 124.200 331.600 137.800 ;
        RECT 332.400 124.200 333.200 137.800 ;
        RECT 337.300 132.400 337.900 149.600 ;
        RECT 340.500 146.400 341.100 175.600 ;
        RECT 342.000 166.200 342.800 177.800 ;
        RECT 343.600 164.200 344.400 177.800 ;
        RECT 345.200 164.200 346.000 177.800 ;
        RECT 346.800 164.200 347.600 177.800 ;
        RECT 348.500 154.400 349.100 209.600 ;
        RECT 350.000 187.600 350.800 188.400 ;
        RECT 345.200 153.600 346.000 154.400 ;
        RECT 348.400 153.600 349.200 154.400 ;
        RECT 351.700 152.400 352.300 225.600 ;
        RECT 353.300 214.400 353.900 227.600 ;
        RECT 353.200 213.600 354.000 214.400 ;
        RECT 353.200 183.600 354.000 184.400 ;
        RECT 353.300 178.400 353.900 183.600 ;
        RECT 354.900 182.400 355.500 235.700 ;
        RECT 361.200 233.600 362.000 234.400 ;
        RECT 361.300 232.400 361.900 233.600 ;
        RECT 362.900 232.400 363.500 243.600 ;
        RECT 361.200 231.600 362.000 232.400 ;
        RECT 362.800 231.600 363.600 232.400 ;
        RECT 367.700 230.400 368.300 251.600 ;
        RECT 372.400 250.300 373.200 250.400 ;
        RECT 372.400 249.700 374.700 250.300 ;
        RECT 372.400 249.600 373.200 249.700 ;
        RECT 370.800 243.600 371.600 244.400 ;
        RECT 364.400 229.600 365.200 230.400 ;
        RECT 367.600 229.600 368.400 230.400 ;
        RECT 356.400 227.600 357.200 228.400 ;
        RECT 366.000 227.600 366.800 228.400 ;
        RECT 359.600 223.600 360.400 224.400 ;
        RECT 359.700 214.400 360.300 223.600 ;
        RECT 367.700 222.400 368.300 229.600 ;
        RECT 370.900 228.400 371.500 243.600 ;
        RECT 374.100 238.400 374.700 249.700 ;
        RECT 377.300 246.400 377.900 271.600 ;
        RECT 398.100 270.400 398.700 281.600 ;
        RECT 402.900 278.400 403.500 291.600 ;
        RECT 406.100 288.400 406.700 329.600 ;
        RECT 415.700 324.400 416.300 329.600 ;
        RECT 415.600 323.600 416.400 324.400 ;
        RECT 446.000 324.200 446.800 337.800 ;
        RECT 447.600 324.200 448.400 337.800 ;
        RECT 449.200 324.200 450.000 337.800 ;
        RECT 450.800 326.200 451.600 337.800 ;
        RECT 452.500 336.400 453.100 339.700 ;
        RECT 452.400 335.600 453.200 336.400 ;
        RECT 454.000 326.200 454.800 337.800 ;
        RECT 455.600 337.600 456.400 338.400 ;
        RECT 455.700 334.400 456.300 337.600 ;
        RECT 455.600 333.600 456.400 334.400 ;
        RECT 457.200 326.200 458.000 337.800 ;
        RECT 458.800 324.200 459.600 337.800 ;
        RECT 460.400 324.200 461.200 337.800 ;
        RECT 463.700 332.400 464.300 349.600 ;
        RECT 463.600 331.600 464.400 332.400 ;
        RECT 466.900 318.400 467.500 349.600 ;
        RECT 471.600 347.600 472.400 348.400 ;
        RECT 476.400 347.600 477.200 348.400 ;
        RECT 486.100 346.400 486.700 373.600 ;
        RECT 487.700 358.400 488.300 383.600 ;
        RECT 489.300 382.400 489.900 411.600 ;
        RECT 490.800 409.600 491.600 410.400 ;
        RECT 492.400 409.600 493.200 410.400 ;
        RECT 490.900 398.400 491.500 409.600 ;
        RECT 490.800 397.600 491.600 398.400 ;
        RECT 492.500 392.400 493.100 409.600 ;
        RECT 494.100 404.400 494.700 447.700 ;
        RECT 495.600 447.600 496.400 447.700 ;
        RECT 495.600 437.600 496.400 438.400 ;
        RECT 495.700 412.400 496.300 437.600 ;
        RECT 497.300 414.400 497.900 455.600 ;
        RECT 503.700 452.400 504.300 481.600 ;
        RECT 508.500 466.400 509.100 495.600 ;
        RECT 510.000 486.200 510.800 497.800 ;
        RECT 511.600 495.600 512.400 496.400 ;
        RECT 511.700 494.400 512.300 495.600 ;
        RECT 511.600 493.600 512.400 494.400 ;
        RECT 511.600 485.600 512.400 486.400 ;
        RECT 513.200 486.200 514.000 497.800 ;
        RECT 511.700 478.400 512.300 485.600 ;
        RECT 514.800 484.200 515.600 497.800 ;
        RECT 516.400 484.200 517.200 497.800 ;
        RECT 526.000 495.600 526.800 496.400 ;
        RECT 532.400 495.600 533.200 496.400 ;
        RECT 526.100 492.400 526.700 495.600 ;
        RECT 532.500 494.400 533.100 495.600 ;
        RECT 529.200 494.300 530.000 494.400 ;
        RECT 527.700 493.700 530.000 494.300 ;
        RECT 522.800 491.600 523.600 492.400 ;
        RECT 526.000 491.600 526.800 492.400 ;
        RECT 522.900 488.400 523.500 491.600 ;
        RECT 522.800 487.600 523.600 488.400 ;
        RECT 527.700 478.400 528.300 493.700 ;
        RECT 529.200 493.600 530.000 493.700 ;
        RECT 532.400 493.600 533.200 494.400 ;
        RECT 538.800 493.600 539.600 494.400 ;
        RECT 545.200 493.600 546.000 494.400 ;
        RECT 542.000 491.600 542.800 492.400 ;
        RECT 559.600 491.600 560.400 492.400 ;
        RECT 529.200 489.600 530.000 490.400 ;
        RECT 535.600 489.600 536.400 490.400 ;
        RECT 538.800 489.600 539.600 490.400 ;
        RECT 529.300 478.400 529.900 489.600 ;
        RECT 535.700 486.400 536.300 489.600 ;
        RECT 559.700 488.400 560.300 491.600 ;
        RECT 559.600 487.600 560.400 488.400 ;
        RECT 535.600 485.600 536.400 486.400 ;
        RECT 551.600 483.600 552.400 484.400 ;
        RECT 561.200 484.200 562.000 497.800 ;
        RECT 562.800 484.200 563.600 497.800 ;
        RECT 564.400 484.200 565.200 497.800 ;
        RECT 566.000 486.200 566.800 497.800 ;
        RECT 567.600 495.600 568.400 496.400 ;
        RECT 569.200 486.200 570.000 497.800 ;
        RECT 570.800 493.600 571.600 494.400 ;
        RECT 570.900 492.400 571.500 493.600 ;
        RECT 570.800 491.600 571.600 492.400 ;
        RECT 572.400 486.200 573.200 497.800 ;
        RECT 574.000 484.200 574.800 497.800 ;
        RECT 575.600 484.200 576.400 497.800 ;
        RECT 578.800 495.600 579.600 496.400 ;
        RECT 511.600 477.600 512.400 478.400 ;
        RECT 527.600 477.600 528.400 478.400 ;
        RECT 529.200 477.600 530.000 478.400 ;
        RECT 526.000 471.600 526.800 472.400 ;
        RECT 518.000 469.600 518.800 470.400 ;
        RECT 518.100 466.400 518.700 469.600 ;
        RECT 527.700 468.400 528.300 477.600 ;
        RECT 530.800 471.600 531.600 472.400 ;
        RECT 521.200 467.600 522.000 468.400 ;
        RECT 527.600 467.600 528.400 468.400 ;
        RECT 542.000 467.600 542.800 468.400 ;
        RECT 508.400 465.600 509.200 466.400 ;
        RECT 513.200 465.600 514.000 466.400 ;
        RECT 518.000 465.600 518.800 466.400 ;
        RECT 502.000 451.600 502.800 452.400 ;
        RECT 503.600 451.600 504.400 452.400 ;
        RECT 498.800 443.600 499.600 444.400 ;
        RECT 498.900 430.400 499.500 443.600 ;
        RECT 502.100 430.400 502.700 451.600 ;
        RECT 505.200 444.200 506.000 457.800 ;
        RECT 506.800 444.200 507.600 457.800 ;
        RECT 508.400 446.200 509.200 457.800 ;
        RECT 510.000 455.600 510.800 456.400 ;
        RECT 510.100 454.400 510.700 455.600 ;
        RECT 510.000 453.600 510.800 454.400 ;
        RECT 511.600 446.200 512.400 457.800 ;
        RECT 513.300 456.400 513.900 465.600 ;
        RECT 518.100 464.400 518.700 465.600 ;
        RECT 514.800 463.600 515.600 464.400 ;
        RECT 518.000 463.600 518.800 464.400 ;
        RECT 514.900 460.400 515.500 463.600 ;
        RECT 514.800 459.600 515.600 460.400 ;
        RECT 513.200 455.600 514.000 456.400 ;
        RECT 513.300 438.400 513.900 455.600 ;
        RECT 514.800 446.200 515.600 457.800 ;
        RECT 514.800 443.600 515.600 444.400 ;
        RECT 516.400 444.200 517.200 457.800 ;
        RECT 518.000 444.200 518.800 457.800 ;
        RECT 519.600 444.200 520.400 457.800 ;
        RECT 513.200 437.600 514.000 438.400 ;
        RECT 506.800 433.600 507.600 434.400 ;
        RECT 498.800 429.600 499.600 430.400 ;
        RECT 502.000 429.600 502.800 430.400 ;
        RECT 503.600 429.600 504.400 430.400 ;
        RECT 498.800 425.600 499.600 426.400 ;
        RECT 497.200 413.600 498.000 414.400 ;
        RECT 495.600 411.600 496.400 412.400 ;
        RECT 498.900 408.300 499.500 425.600 ;
        RECT 502.100 424.400 502.700 429.600 ;
        RECT 506.900 428.400 507.500 433.600 ;
        RECT 508.400 429.600 509.200 430.400 ;
        RECT 505.200 427.600 506.000 428.400 ;
        RECT 506.800 427.600 507.600 428.400 ;
        RECT 502.000 423.600 502.800 424.400 ;
        RECT 505.300 422.400 505.900 427.600 ;
        RECT 505.200 421.600 506.000 422.400 ;
        RECT 500.400 415.600 501.200 416.400 ;
        RECT 500.500 410.400 501.100 415.600 ;
        RECT 502.000 413.600 502.800 414.400 ;
        RECT 503.600 411.600 504.400 412.400 ;
        RECT 500.400 409.600 501.200 410.400 ;
        RECT 503.600 409.600 504.400 410.400 ;
        RECT 498.900 407.700 501.100 408.300 ;
        RECT 494.000 403.600 494.800 404.400 ;
        RECT 494.100 398.400 494.700 403.600 ;
        RECT 494.000 397.600 494.800 398.400 ;
        RECT 500.500 394.400 501.100 407.700 ;
        RECT 503.700 396.400 504.300 409.600 ;
        RECT 505.300 400.400 505.900 421.600 ;
        RECT 506.800 413.600 507.600 414.400 ;
        RECT 506.800 409.600 507.600 410.400 ;
        RECT 506.900 402.400 507.500 409.600 ;
        RECT 506.800 401.600 507.600 402.400 ;
        RECT 505.200 399.600 506.000 400.400 ;
        RECT 503.600 395.600 504.400 396.400 ;
        RECT 498.800 393.600 499.600 394.400 ;
        RECT 500.400 393.600 501.200 394.400 ;
        RECT 492.400 391.600 493.200 392.400 ;
        RECT 490.800 387.600 491.600 388.400 ;
        RECT 489.200 381.600 490.000 382.400 ;
        RECT 489.200 375.600 490.000 376.400 ;
        RECT 487.600 357.600 488.400 358.400 ;
        RECT 476.400 345.600 477.200 346.400 ;
        RECT 486.000 345.600 486.800 346.400 ;
        RECT 473.200 343.600 474.000 344.400 ;
        RECT 471.600 337.600 472.400 338.400 ;
        RECT 470.000 335.600 470.800 336.400 ;
        RECT 470.100 334.400 470.700 335.600 ;
        RECT 470.000 333.600 470.800 334.400 ;
        RECT 410.800 309.600 411.600 310.400 ;
        RECT 407.600 307.600 408.400 308.400 ;
        RECT 407.700 298.400 408.300 307.600 ;
        RECT 414.000 303.600 414.800 304.400 ;
        RECT 415.600 304.200 416.400 317.800 ;
        RECT 417.200 304.200 418.000 317.800 ;
        RECT 418.800 304.200 419.600 315.800 ;
        RECT 420.400 307.600 421.200 308.400 ;
        RECT 422.000 304.200 422.800 315.800 ;
        RECT 423.600 305.600 424.400 306.400 ;
        RECT 407.600 297.600 408.400 298.400 ;
        RECT 414.100 296.400 414.700 303.600 ;
        RECT 423.700 296.400 424.300 305.600 ;
        RECT 425.200 304.200 426.000 315.800 ;
        RECT 426.800 304.200 427.600 317.800 ;
        RECT 428.400 304.200 429.200 317.800 ;
        RECT 430.000 304.200 430.800 317.800 ;
        RECT 439.600 317.600 440.400 318.400 ;
        RECT 466.800 317.600 467.600 318.400 ;
        RECT 431.600 309.600 432.400 310.400 ;
        RECT 431.700 300.400 432.300 309.600 ;
        RECT 444.400 307.600 445.200 308.400 ;
        RECT 441.200 305.600 442.000 306.400 ;
        RECT 446.000 306.200 446.800 311.800 ;
        RECT 447.600 307.600 448.400 308.400 ;
        RECT 439.600 303.600 440.400 304.400 ;
        RECT 441.300 302.400 441.900 305.600 ;
        RECT 441.200 301.600 442.000 302.400 ;
        RECT 426.800 299.600 427.600 300.400 ;
        RECT 431.600 299.600 432.400 300.400 ;
        RECT 414.000 295.600 414.800 296.400 ;
        RECT 423.600 295.600 424.400 296.400 ;
        RECT 426.900 292.400 427.500 299.600 ;
        RECT 426.800 291.600 427.600 292.400 ;
        RECT 406.000 287.600 406.800 288.400 ;
        RECT 428.400 284.200 429.200 297.800 ;
        RECT 430.000 284.200 430.800 297.800 ;
        RECT 431.600 286.200 432.400 297.800 ;
        RECT 433.200 293.600 434.000 294.400 ;
        RECT 433.200 291.600 434.000 292.400 ;
        RECT 402.800 277.600 403.600 278.400 ;
        RECT 409.200 277.600 410.000 278.400 ;
        RECT 406.000 273.600 406.800 274.400 ;
        RECT 409.300 270.400 409.900 277.600 ;
        RECT 433.300 270.400 433.900 291.600 ;
        RECT 434.800 286.200 435.600 297.800 ;
        RECT 436.400 295.600 437.200 296.400 ;
        RECT 438.000 286.200 438.800 297.800 ;
        RECT 439.600 284.200 440.400 297.800 ;
        RECT 441.200 284.200 442.000 297.800 ;
        RECT 442.800 284.200 443.600 297.800 ;
        RECT 447.700 296.400 448.300 307.600 ;
        RECT 449.200 304.200 450.000 315.800 ;
        RECT 452.400 315.600 453.200 316.400 ;
        RECT 452.500 310.400 453.100 315.600 ;
        RECT 452.400 309.600 453.200 310.400 ;
        RECT 458.800 304.200 459.600 315.800 ;
        RECT 465.200 313.600 466.000 314.400 ;
        RECT 465.300 312.400 465.900 313.600 ;
        RECT 473.300 312.400 473.900 343.600 ;
        RECT 476.500 338.400 477.100 345.600 ;
        RECT 481.200 343.600 482.000 344.400 ;
        RECT 482.800 343.600 483.600 344.400 ;
        RECT 487.600 344.200 488.400 355.800 ;
        RECT 476.400 337.600 477.200 338.400 ;
        RECT 478.000 337.600 478.800 338.400 ;
        RECT 476.400 335.600 477.200 336.400 ;
        RECT 474.800 333.600 475.600 334.400 ;
        RECT 474.800 330.300 475.600 330.400 ;
        RECT 476.500 330.300 477.100 335.600 ;
        RECT 478.100 330.400 478.700 337.600 ;
        RECT 479.600 335.600 480.400 336.400 ;
        RECT 474.800 329.700 477.100 330.300 ;
        RECT 474.800 329.600 475.600 329.700 ;
        RECT 478.000 329.600 478.800 330.400 ;
        RECT 478.000 327.600 478.800 328.400 ;
        RECT 465.200 311.600 466.000 312.400 ;
        RECT 473.200 311.600 474.000 312.400 ;
        RECT 474.800 311.600 475.600 312.400 ;
        RECT 474.900 310.400 475.500 311.600 ;
        RECT 478.100 310.400 478.700 327.600 ;
        RECT 479.700 318.400 480.300 335.600 ;
        RECT 481.300 332.400 481.900 343.600 ;
        RECT 489.300 336.300 489.900 375.600 ;
        RECT 490.900 372.400 491.500 387.600 ;
        RECT 494.000 385.600 494.800 386.400 ;
        RECT 494.100 378.400 494.700 385.600 ;
        RECT 494.000 377.600 494.800 378.400 ;
        RECT 490.800 371.600 491.600 372.400 ;
        RECT 490.900 348.400 491.500 371.600 ;
        RECT 497.200 363.600 498.000 364.400 ;
        RECT 497.300 358.300 497.900 363.600 ;
        RECT 495.700 357.700 497.900 358.300 ;
        RECT 494.000 349.600 494.800 350.400 ;
        RECT 490.800 347.600 491.600 348.400 ;
        RECT 494.100 346.400 494.700 349.600 ;
        RECT 495.700 348.400 496.300 357.700 ;
        RECT 495.600 347.600 496.400 348.400 ;
        RECT 490.800 345.600 491.600 346.400 ;
        RECT 494.000 345.600 494.800 346.400 ;
        RECT 490.900 338.400 491.500 345.600 ;
        RECT 497.200 344.200 498.000 355.800 ;
        RECT 497.200 341.600 498.000 342.400 ;
        RECT 490.800 337.600 491.600 338.400 ;
        RECT 487.700 335.700 489.900 336.300 ;
        RECT 482.800 333.600 483.600 334.400 ;
        RECT 481.200 331.600 482.000 332.400 ;
        RECT 482.900 328.400 483.500 333.600 ;
        RECT 487.700 330.400 488.300 335.700 ;
        RECT 489.200 333.600 490.000 334.400 ;
        RECT 487.600 329.600 488.400 330.400 ;
        RECT 482.800 327.600 483.600 328.400 ;
        RECT 484.400 323.600 485.200 324.400 ;
        RECT 479.600 317.600 480.400 318.400 ;
        RECT 482.800 315.600 483.600 316.400 ;
        RECT 479.600 311.600 480.400 312.400 ;
        RECT 468.400 309.600 469.200 310.400 ;
        RECT 470.000 309.600 470.800 310.400 ;
        RECT 474.800 309.600 475.600 310.400 ;
        RECT 478.000 309.600 478.800 310.400 ;
        RECT 468.500 308.400 469.100 309.600 ;
        RECT 470.100 308.400 470.700 309.600 ;
        RECT 468.400 307.600 469.200 308.400 ;
        RECT 470.000 307.600 470.800 308.400 ;
        RECT 471.600 307.600 472.400 308.400 ;
        RECT 474.800 307.600 475.600 308.400 ;
        RECT 479.700 308.300 480.300 311.600 ;
        RECT 482.900 310.400 483.500 315.600 ;
        RECT 484.500 312.400 485.100 323.600 ;
        RECT 486.000 317.600 486.800 318.400 ;
        RECT 484.400 311.600 485.200 312.400 ;
        RECT 481.200 309.600 482.000 310.400 ;
        RECT 482.800 309.600 483.600 310.400 ;
        RECT 486.000 309.600 486.800 310.400 ;
        RECT 481.300 308.400 481.900 309.600 ;
        RECT 478.100 307.700 480.300 308.300 ;
        RECT 465.200 305.600 466.000 306.400 ;
        RECT 452.400 297.600 453.200 298.400 ;
        RECT 463.600 297.600 464.400 298.400 ;
        RECT 463.700 296.400 464.300 297.600 ;
        RECT 465.300 296.400 465.900 305.600 ;
        RECT 447.600 295.600 448.400 296.400 ;
        RECT 463.600 295.600 464.400 296.400 ;
        RECT 465.200 295.600 466.000 296.400 ;
        RECT 468.500 294.400 469.100 307.600 ;
        RECT 471.700 294.400 472.300 307.600 ;
        RECT 473.200 295.600 474.000 296.400 ;
        RECT 454.000 293.600 454.800 294.400 ;
        RECT 465.200 293.600 466.000 294.400 ;
        RECT 468.400 293.600 469.200 294.400 ;
        RECT 471.600 293.600 472.400 294.400 ;
        RECT 458.800 291.600 459.600 292.400 ;
        RECT 463.600 291.600 464.400 292.400 ;
        RECT 455.600 289.600 456.400 290.400 ;
        RECT 455.700 278.400 456.300 289.600 ;
        RECT 455.600 278.300 456.400 278.400 ;
        RECT 378.800 269.600 379.600 270.400 ;
        RECT 386.800 269.600 387.600 270.400 ;
        RECT 388.400 270.300 389.200 270.400 ;
        RECT 390.000 270.300 390.800 270.400 ;
        RECT 388.400 269.700 390.800 270.300 ;
        RECT 388.400 269.600 389.200 269.700 ;
        RECT 390.000 269.600 390.800 269.700 ;
        RECT 398.000 269.600 398.800 270.400 ;
        RECT 409.200 269.600 410.000 270.400 ;
        RECT 410.800 269.600 411.600 270.400 ;
        RECT 433.200 269.600 434.000 270.400 ;
        RECT 385.200 263.600 386.000 264.400 ;
        RECT 380.400 255.600 381.200 256.400 ;
        RECT 380.400 253.600 381.200 254.400 ;
        RECT 385.300 252.400 385.900 263.600 ;
        RECT 386.900 256.400 387.500 269.600 ;
        RECT 394.800 263.600 395.600 264.400 ;
        RECT 394.900 258.400 395.500 263.600 ;
        RECT 394.800 257.600 395.600 258.400 ;
        RECT 386.800 255.600 387.600 256.400 ;
        RECT 398.100 256.300 398.700 269.600 ;
        RECT 410.900 266.400 411.500 269.600 ;
        RECT 410.800 265.600 411.600 266.400 ;
        RECT 425.200 265.600 426.000 266.400 ;
        RECT 401.200 263.600 402.000 264.400 ;
        RECT 404.400 263.600 405.200 264.400 ;
        RECT 401.300 256.400 401.900 263.600 ;
        RECT 402.800 259.600 403.600 260.400 ;
        RECT 402.900 258.400 403.500 259.600 ;
        RECT 402.800 257.600 403.600 258.400 ;
        RECT 398.100 255.700 400.300 256.300 ;
        RECT 386.900 252.400 387.500 255.600 ;
        RECT 398.000 253.600 398.800 254.400 ;
        RECT 399.700 252.400 400.300 255.700 ;
        RECT 401.200 255.600 402.000 256.400 ;
        RECT 383.600 251.600 384.400 252.400 ;
        RECT 385.200 251.600 386.000 252.400 ;
        RECT 386.800 251.600 387.600 252.400 ;
        RECT 399.600 251.600 400.400 252.400 ;
        RECT 383.700 250.400 384.300 251.600 ;
        RECT 378.800 249.600 379.600 250.400 ;
        RECT 383.600 249.600 384.400 250.400 ;
        RECT 385.200 249.600 386.000 250.400 ;
        RECT 388.400 249.600 389.200 250.400 ;
        RECT 391.600 249.600 392.400 250.400 ;
        RECT 393.200 249.600 394.000 250.400 ;
        RECT 378.900 246.400 379.500 249.600 ;
        RECT 385.300 246.400 385.900 249.600 ;
        RECT 388.500 248.400 389.100 249.600 ;
        RECT 388.400 247.600 389.200 248.400 ;
        RECT 377.200 245.600 378.000 246.400 ;
        RECT 378.800 245.600 379.600 246.400 ;
        RECT 385.200 245.600 386.000 246.400 ;
        RECT 390.000 245.600 390.800 246.400 ;
        RECT 375.600 243.600 376.400 244.400 ;
        RECT 386.800 243.600 387.600 244.400 ;
        RECT 388.400 243.600 389.200 244.400 ;
        RECT 374.000 237.600 374.800 238.400 ;
        RECT 375.700 236.400 376.300 243.600 ;
        RECT 383.600 241.600 384.400 242.400 ;
        RECT 383.700 238.400 384.300 241.600 ;
        RECT 378.800 237.600 379.600 238.400 ;
        RECT 383.600 237.600 384.400 238.400 ;
        RECT 385.200 237.600 386.000 238.400 ;
        RECT 375.600 235.600 376.400 236.400 ;
        RECT 375.600 233.600 376.400 234.400 ;
        RECT 372.400 229.600 373.200 230.400 ;
        RECT 372.500 228.400 373.100 229.600 ;
        RECT 370.800 227.600 371.600 228.400 ;
        RECT 372.400 227.600 373.200 228.400 ;
        RECT 367.600 221.600 368.400 222.400 ;
        RECT 375.700 220.400 376.300 233.600 ;
        RECT 378.900 232.400 379.500 237.600 ;
        RECT 380.400 235.600 381.200 236.400 ;
        RECT 378.800 231.600 379.600 232.400 ;
        RECT 377.200 229.600 378.000 230.400 ;
        RECT 377.300 220.400 377.900 229.600 ;
        RECT 380.500 224.400 381.100 235.600 ;
        RECT 382.000 233.600 382.800 234.400 ;
        RECT 385.300 232.400 385.900 237.600 ;
        RECT 385.200 231.600 386.000 232.400 ;
        RECT 383.600 229.600 384.400 230.400 ;
        RECT 385.200 229.600 386.000 230.400 ;
        RECT 383.700 228.400 384.300 229.600 ;
        RECT 383.600 227.600 384.400 228.400 ;
        RECT 380.400 223.600 381.200 224.400 ;
        RECT 375.600 219.600 376.400 220.400 ;
        RECT 377.200 219.600 378.000 220.400 ;
        RECT 359.600 213.600 360.400 214.400 ;
        RECT 366.000 204.200 366.800 217.800 ;
        RECT 367.600 204.200 368.400 217.800 ;
        RECT 369.200 204.200 370.000 217.800 ;
        RECT 370.800 206.200 371.600 217.800 ;
        RECT 372.400 215.600 373.200 216.400 ;
        RECT 358.000 197.600 358.800 198.400 ;
        RECT 356.400 185.600 357.200 186.400 ;
        RECT 354.800 181.600 355.600 182.400 ;
        RECT 353.200 177.600 354.000 178.400 ;
        RECT 356.400 169.600 357.200 170.400 ;
        RECT 345.200 151.600 346.000 152.400 ;
        RECT 351.600 151.600 352.400 152.400 ;
        RECT 340.400 145.600 341.200 146.400 ;
        RECT 345.300 136.400 345.900 151.600 ;
        RECT 358.100 150.400 358.700 197.600 ;
        RECT 370.800 195.600 371.600 196.400 ;
        RECT 372.500 194.400 373.100 215.600 ;
        RECT 374.000 206.200 374.800 217.800 ;
        RECT 375.600 213.600 376.400 214.400 ;
        RECT 377.200 206.200 378.000 217.800 ;
        RECT 378.800 204.200 379.600 217.800 ;
        RECT 380.400 204.200 381.200 217.800 ;
        RECT 385.300 212.400 385.900 229.600 ;
        RECT 385.200 211.600 386.000 212.400 ;
        RECT 380.400 197.600 381.200 198.400 ;
        RECT 372.400 193.600 373.200 194.400 ;
        RECT 380.500 192.400 381.100 197.600 ;
        RECT 375.600 191.600 376.400 192.400 ;
        RECT 380.400 191.600 381.200 192.400 ;
        RECT 382.000 191.600 382.800 192.400 ;
        RECT 382.100 188.400 382.700 191.600 ;
        RECT 383.600 189.600 384.400 190.400 ;
        RECT 361.200 187.600 362.000 188.400 ;
        RECT 367.600 187.600 368.400 188.400 ;
        RECT 369.200 187.600 370.000 188.400 ;
        RECT 372.400 187.600 373.200 188.400 ;
        RECT 382.000 187.600 382.800 188.400 ;
        RECT 361.300 178.400 361.900 187.600 ;
        RECT 367.700 182.400 368.300 187.600 ;
        RECT 369.200 183.600 370.000 184.400 ;
        RECT 380.400 183.600 381.200 184.400 ;
        RECT 383.600 183.600 384.400 184.400 ;
        RECT 367.600 181.600 368.400 182.400 ;
        RECT 366.000 179.600 366.800 180.400 ;
        RECT 361.200 177.600 362.000 178.400 ;
        RECT 358.000 149.600 358.800 150.400 ;
        RECT 346.800 145.600 347.600 146.400 ;
        RECT 346.900 136.400 347.500 145.600 ;
        RECT 359.600 144.200 360.400 157.800 ;
        RECT 361.200 144.200 362.000 157.800 ;
        RECT 362.800 144.200 363.600 157.800 ;
        RECT 364.400 144.200 365.200 155.800 ;
        RECT 366.100 146.400 366.700 179.600 ;
        RECT 366.000 145.600 366.800 146.400 ;
        RECT 367.600 144.200 368.400 155.800 ;
        RECT 369.300 148.400 369.900 183.600 ;
        RECT 377.200 179.600 378.000 180.400 ;
        RECT 370.800 164.200 371.600 177.800 ;
        RECT 372.400 164.200 373.200 177.800 ;
        RECT 374.000 164.200 374.800 177.800 ;
        RECT 375.600 166.200 376.400 177.800 ;
        RECT 377.300 176.400 377.900 179.600 ;
        RECT 377.200 175.600 378.000 176.400 ;
        RECT 378.800 166.200 379.600 177.800 ;
        RECT 380.500 174.400 381.100 183.600 ;
        RECT 380.400 173.600 381.200 174.400 ;
        RECT 380.400 171.600 381.200 172.400 ;
        RECT 369.200 147.600 370.000 148.400 ;
        RECT 370.800 144.200 371.600 155.800 ;
        RECT 372.400 144.200 373.200 157.800 ;
        RECT 374.000 144.200 374.800 157.800 ;
        RECT 380.500 150.400 381.100 171.600 ;
        RECT 382.000 166.200 382.800 177.800 ;
        RECT 383.600 164.200 384.400 177.800 ;
        RECT 385.200 164.200 386.000 177.800 ;
        RECT 386.900 174.400 387.500 243.600 ;
        RECT 388.500 188.400 389.100 243.600 ;
        RECT 393.300 242.400 393.900 249.600 ;
        RECT 393.200 241.600 394.000 242.400 ;
        RECT 401.300 238.400 401.900 255.600 ;
        RECT 404.500 254.400 405.100 263.600 ;
        RECT 406.000 261.600 406.800 262.400 ;
        RECT 406.100 258.400 406.700 261.600 ;
        RECT 410.900 258.400 411.500 265.600 ;
        RECT 414.000 263.600 414.800 264.400 ;
        RECT 434.800 264.200 435.600 277.800 ;
        RECT 436.400 264.200 437.200 277.800 ;
        RECT 438.000 264.200 438.800 275.800 ;
        RECT 439.600 267.600 440.400 268.400 ;
        RECT 441.200 264.200 442.000 275.800 ;
        RECT 442.800 265.600 443.600 266.400 ;
        RECT 406.000 257.600 406.800 258.400 ;
        RECT 410.800 257.600 411.600 258.400 ;
        RECT 410.800 256.300 411.600 256.400 ;
        RECT 410.800 255.700 413.100 256.300 ;
        RECT 410.800 255.600 411.600 255.700 ;
        RECT 404.400 253.600 405.200 254.400 ;
        RECT 412.500 250.400 413.100 255.700 ;
        RECT 414.100 254.400 414.700 263.600 ;
        RECT 442.900 260.400 443.500 265.600 ;
        RECT 444.400 264.200 445.200 275.800 ;
        RECT 446.000 264.200 446.800 277.800 ;
        RECT 447.600 264.200 448.400 277.800 ;
        RECT 449.200 264.200 450.000 277.800 ;
        RECT 455.600 277.700 457.900 278.300 ;
        RECT 455.600 277.600 456.400 277.700 ;
        RECT 450.800 269.600 451.600 270.400 ;
        RECT 442.800 259.600 443.600 260.400 ;
        RECT 450.800 259.600 451.600 260.400 ;
        RECT 414.000 253.600 414.800 254.400 ;
        RECT 414.000 251.600 414.800 252.400 ;
        RECT 426.800 251.600 427.600 252.400 ;
        RECT 412.400 249.600 413.200 250.400 ;
        RECT 414.100 246.400 414.700 251.600 ;
        RECT 415.600 249.600 416.400 250.400 ;
        RECT 415.700 248.400 416.300 249.600 ;
        RECT 415.600 247.600 416.400 248.400 ;
        RECT 414.000 245.600 414.800 246.400 ;
        RECT 423.600 245.600 424.400 246.400 ;
        RECT 402.800 243.600 403.600 244.400 ;
        RECT 393.200 231.600 394.000 232.400 ;
        RECT 390.000 229.600 390.800 230.400 ;
        RECT 390.000 217.600 390.800 218.400 ;
        RECT 390.100 194.400 390.700 217.600 ;
        RECT 391.600 213.600 392.400 214.400 ;
        RECT 390.000 193.600 390.800 194.400 ;
        RECT 390.100 192.400 390.700 193.600 ;
        RECT 393.300 192.400 393.900 231.600 ;
        RECT 394.800 224.200 395.600 237.800 ;
        RECT 396.400 224.200 397.200 237.800 ;
        RECT 401.200 237.600 402.000 238.400 ;
        RECT 398.000 224.200 398.800 235.800 ;
        RECT 399.600 227.600 400.400 228.400 ;
        RECT 401.200 224.200 402.000 235.800 ;
        RECT 402.900 232.400 403.500 243.600 ;
        RECT 402.800 231.600 403.600 232.400 ;
        RECT 402.800 225.600 403.600 226.400 ;
        RECT 404.400 224.200 405.200 235.800 ;
        RECT 406.000 224.200 406.800 237.800 ;
        RECT 407.600 224.200 408.400 237.800 ;
        RECT 409.200 224.200 410.000 237.800 ;
        RECT 423.700 234.400 424.300 245.600 ;
        RECT 423.600 233.600 424.400 234.400 ;
        RECT 410.800 231.600 411.600 232.400 ;
        RECT 410.900 230.400 411.500 231.600 ;
        RECT 423.700 230.400 424.300 233.600 ;
        RECT 426.900 232.400 427.500 251.600 ;
        RECT 428.400 249.600 429.200 250.400 ;
        RECT 428.500 238.400 429.100 249.600 ;
        RECT 431.600 244.200 432.400 257.800 ;
        RECT 433.200 244.200 434.000 257.800 ;
        RECT 434.800 246.200 435.600 257.800 ;
        RECT 436.400 253.600 437.200 254.400 ;
        RECT 438.000 246.200 438.800 257.800 ;
        RECT 439.600 255.600 440.400 256.400 ;
        RECT 441.200 246.200 442.000 257.800 ;
        RECT 442.800 244.200 443.600 257.800 ;
        RECT 444.400 244.200 445.200 257.800 ;
        RECT 446.000 244.200 446.800 257.800 ;
        RECT 450.900 238.400 451.500 259.600 ;
        RECT 455.600 257.600 456.400 258.400 ;
        RECT 457.300 252.400 457.900 277.700 ;
        RECT 457.200 251.600 458.000 252.400 ;
        RECT 458.900 244.400 459.500 291.600 ;
        RECT 463.700 278.400 464.300 291.600 ;
        RECT 470.000 289.600 470.800 290.400 ;
        RECT 471.700 288.400 472.300 293.600 ;
        RECT 473.300 292.400 473.900 295.600 ;
        RECT 473.200 291.600 474.000 292.400 ;
        RECT 474.900 290.400 475.500 307.600 ;
        RECT 478.100 302.400 478.700 307.700 ;
        RECT 481.200 307.600 482.000 308.400 ;
        RECT 479.600 305.600 480.400 306.400 ;
        RECT 478.000 301.600 478.800 302.400 ;
        RECT 476.400 295.600 477.200 296.400 ;
        RECT 476.500 292.400 477.100 295.600 ;
        RECT 478.100 292.400 478.700 301.600 ;
        RECT 481.200 299.600 482.000 300.400 ;
        RECT 481.300 294.400 481.900 299.600 ;
        RECT 482.900 294.400 483.500 309.600 ;
        RECT 484.400 307.600 485.200 308.400 ;
        RECT 484.500 300.400 485.100 307.600 ;
        RECT 486.100 306.400 486.700 309.600 ;
        RECT 486.000 305.600 486.800 306.400 ;
        RECT 487.600 305.600 488.400 306.400 ;
        RECT 484.400 299.600 485.200 300.400 ;
        RECT 487.700 298.400 488.300 305.600 ;
        RECT 487.600 297.600 488.400 298.400 ;
        RECT 487.700 296.400 488.300 297.600 ;
        RECT 487.600 295.600 488.400 296.400 ;
        RECT 479.600 293.600 480.400 294.400 ;
        RECT 481.200 293.600 482.000 294.400 ;
        RECT 482.800 293.600 483.600 294.400 ;
        RECT 486.000 293.600 486.800 294.400 ;
        RECT 479.700 292.400 480.300 293.600 ;
        RECT 476.400 291.600 477.200 292.400 ;
        RECT 478.000 291.600 478.800 292.400 ;
        RECT 479.600 291.600 480.400 292.400 ;
        RECT 474.800 289.600 475.600 290.400 ;
        RECT 471.600 287.600 472.400 288.400 ;
        RECT 481.300 280.400 481.900 293.600 ;
        RECT 482.800 291.600 483.600 292.400 ;
        RECT 486.000 291.600 486.800 292.400 ;
        RECT 486.100 290.400 486.700 291.600 ;
        RECT 486.000 289.600 486.800 290.400 ;
        RECT 481.200 279.600 482.000 280.400 ;
        RECT 463.600 277.600 464.400 278.400 ;
        RECT 468.400 269.600 469.200 270.400 ;
        RECT 463.600 267.600 464.400 268.400 ;
        RECT 462.000 265.600 462.800 266.400 ;
        RECT 462.100 258.400 462.700 265.600 ;
        RECT 463.700 258.400 464.300 267.600 ;
        RECT 473.200 264.200 474.000 277.800 ;
        RECT 474.800 264.200 475.600 277.800 ;
        RECT 476.400 264.200 477.200 275.800 ;
        RECT 478.000 267.600 478.800 268.400 ;
        RECT 478.100 266.400 478.700 267.600 ;
        RECT 478.000 265.600 478.800 266.400 ;
        RECT 479.600 264.200 480.400 275.800 ;
        RECT 481.200 265.600 482.000 266.400 ;
        RECT 481.300 260.400 481.900 265.600 ;
        RECT 482.800 264.200 483.600 275.800 ;
        RECT 484.400 264.200 485.200 277.800 ;
        RECT 486.000 264.200 486.800 277.800 ;
        RECT 487.600 264.200 488.400 277.800 ;
        RECT 489.300 268.400 489.900 333.600 ;
        RECT 497.300 332.400 497.900 341.600 ;
        RECT 495.600 331.600 496.400 332.400 ;
        RECT 497.200 331.600 498.000 332.400 ;
        RECT 495.700 316.400 496.300 331.600 ;
        RECT 497.200 325.600 498.000 326.400 ;
        RECT 495.600 315.600 496.400 316.400 ;
        RECT 490.800 313.600 491.600 314.400 ;
        RECT 490.900 312.400 491.500 313.600 ;
        RECT 497.300 312.400 497.900 325.600 ;
        RECT 498.900 318.400 499.500 393.600 ;
        RECT 503.700 392.400 504.300 395.600 ;
        RECT 503.600 391.600 504.400 392.400 ;
        RECT 505.300 388.400 505.900 399.600 ;
        RECT 506.800 391.600 507.600 392.400 ;
        RECT 506.900 390.400 507.500 391.600 ;
        RECT 508.500 390.400 509.100 429.600 ;
        RECT 510.000 407.600 510.800 408.400 ;
        RECT 510.000 397.600 510.800 398.400 ;
        RECT 510.100 390.400 510.700 397.600 ;
        RECT 514.900 394.400 515.500 443.600 ;
        RECT 521.300 438.400 521.900 467.600 ;
        RECT 526.000 463.600 526.800 464.400 ;
        RECT 526.100 454.400 526.700 463.600 ;
        RECT 542.100 462.300 542.700 467.600 ;
        RECT 543.600 464.200 544.400 477.800 ;
        RECT 545.200 464.200 546.000 477.800 ;
        RECT 546.800 464.200 547.600 477.800 ;
        RECT 548.400 464.200 549.200 475.800 ;
        RECT 550.000 469.600 550.800 470.400 ;
        RECT 550.100 466.400 550.700 469.600 ;
        RECT 550.000 465.600 550.800 466.400 ;
        RECT 550.000 463.600 550.800 464.400 ;
        RECT 551.600 464.200 552.400 475.800 ;
        RECT 553.200 467.600 554.000 468.400 ;
        RECT 553.300 464.400 553.900 467.600 ;
        RECT 553.200 463.600 554.000 464.400 ;
        RECT 554.800 464.200 555.600 475.800 ;
        RECT 556.400 464.200 557.200 477.800 ;
        RECT 558.000 464.200 558.800 477.800 ;
        RECT 578.900 470.400 579.500 495.600 ;
        RECT 585.200 493.600 586.000 494.400 ;
        RECT 583.600 471.600 584.400 472.400 ;
        RECT 585.300 470.400 585.900 493.600 ;
        RECT 586.800 491.600 587.600 492.400 ;
        RECT 594.800 491.600 595.600 492.400 ;
        RECT 586.900 478.400 587.500 491.600 ;
        RECT 586.800 477.600 587.600 478.400 ;
        RECT 590.000 471.600 590.800 472.400 ;
        RECT 562.800 469.600 563.600 470.400 ;
        RECT 575.600 469.600 576.400 470.400 ;
        RECT 578.800 469.600 579.600 470.400 ;
        RECT 585.200 469.600 586.000 470.400 ;
        RECT 559.600 465.600 560.400 466.400 ;
        RECT 542.100 461.700 544.300 462.300 ;
        RECT 542.000 459.600 542.800 460.400 ;
        RECT 530.800 455.600 531.600 456.400 ;
        RECT 542.100 454.400 542.700 459.600 ;
        RECT 543.700 458.400 544.300 461.700 ;
        RECT 550.100 458.400 550.700 463.600 ;
        RECT 551.600 459.600 552.400 460.400 ;
        RECT 543.600 457.600 544.400 458.400 ;
        RECT 550.000 457.600 550.800 458.400 ;
        RECT 551.700 456.400 552.300 459.600 ;
        RECT 551.600 455.600 552.400 456.400 ;
        RECT 526.000 453.600 526.800 454.400 ;
        RECT 542.000 453.600 542.800 454.400 ;
        RECT 546.800 453.600 547.600 454.400 ;
        RECT 537.200 452.300 538.000 452.400 ;
        RECT 537.200 451.700 539.500 452.300 ;
        RECT 537.200 451.600 538.000 451.700 ;
        RECT 530.800 450.300 531.600 450.400 ;
        RECT 529.300 449.700 531.600 450.300 ;
        RECT 529.300 438.400 529.900 449.700 ;
        RECT 530.800 449.600 531.600 449.700 ;
        RECT 530.800 447.600 531.600 448.400 ;
        RECT 518.000 437.600 518.800 438.400 ;
        RECT 521.200 437.600 522.000 438.400 ;
        RECT 529.200 437.600 530.000 438.400 ;
        RECT 530.900 432.300 531.500 447.600 ;
        RECT 538.900 438.400 539.500 451.700 ;
        RECT 542.000 449.600 542.800 450.400 ;
        RECT 546.800 449.600 547.600 450.400 ;
        RECT 550.000 449.600 550.800 450.400 ;
        RECT 538.800 437.600 539.600 438.400 ;
        RECT 532.400 432.300 533.200 432.400 ;
        RECT 530.900 431.700 533.200 432.300 ;
        RECT 532.400 431.600 533.200 431.700 ;
        RECT 526.000 429.600 526.800 430.400 ;
        RECT 529.200 429.600 530.000 430.400 ;
        RECT 540.400 429.600 541.200 430.400 ;
        RECT 519.600 427.600 520.400 428.400 ;
        RECT 522.800 427.600 523.600 428.400 ;
        RECT 519.700 426.400 520.300 427.600 ;
        RECT 526.100 426.400 526.700 429.600 ;
        RECT 527.600 427.600 528.400 428.400 ;
        RECT 519.600 425.600 520.400 426.400 ;
        RECT 526.000 425.600 526.800 426.400 ;
        RECT 519.700 424.400 520.300 425.600 ;
        RECT 518.000 423.600 518.800 424.400 ;
        RECT 519.600 423.600 520.400 424.400 ;
        RECT 526.000 423.600 526.800 424.400 ;
        RECT 518.100 412.400 518.700 423.600 ;
        RECT 518.000 411.600 518.800 412.400 ;
        RECT 518.000 407.600 518.800 408.400 ;
        RECT 514.800 393.600 515.600 394.400 ;
        RECT 518.100 392.400 518.700 407.600 ;
        RECT 519.600 404.200 520.400 417.800 ;
        RECT 521.200 404.200 522.000 417.800 ;
        RECT 522.800 404.200 523.600 417.800 ;
        RECT 524.400 406.200 525.200 417.800 ;
        RECT 526.100 416.400 526.700 423.600 ;
        RECT 527.700 422.400 528.300 427.600 ;
        RECT 529.300 424.400 529.900 429.600 ;
        RECT 534.000 427.600 534.800 428.400 ;
        RECT 535.600 427.600 536.400 428.400 ;
        RECT 534.100 426.400 534.700 427.600 ;
        RECT 534.000 425.600 534.800 426.400 ;
        RECT 535.700 424.400 536.300 427.600 ;
        RECT 529.200 423.600 530.000 424.400 ;
        RECT 535.600 423.600 536.400 424.400 ;
        RECT 538.800 423.600 539.600 424.400 ;
        RECT 527.600 421.600 528.400 422.400 ;
        RECT 526.000 415.600 526.800 416.400 ;
        RECT 527.600 406.200 528.400 417.800 ;
        RECT 529.200 413.600 530.000 414.400 ;
        RECT 530.800 406.200 531.600 417.800 ;
        RECT 529.200 403.600 530.000 404.400 ;
        RECT 530.800 403.600 531.600 404.400 ;
        RECT 532.400 404.200 533.200 417.800 ;
        RECT 534.000 404.200 534.800 417.800 ;
        RECT 538.900 412.400 539.500 423.600 ;
        RECT 540.500 420.400 541.100 429.600 ;
        RECT 540.400 419.600 541.200 420.400 ;
        RECT 540.400 415.600 541.200 416.400 ;
        RECT 540.500 412.400 541.100 415.600 ;
        RECT 538.800 411.600 539.600 412.400 ;
        RECT 540.400 411.600 541.200 412.400 ;
        RECT 521.200 401.600 522.000 402.400 ;
        RECT 521.300 398.400 521.900 401.600 ;
        RECT 521.200 397.600 522.000 398.400 ;
        RECT 522.800 395.600 523.600 396.400 ;
        RECT 511.600 391.600 512.400 392.400 ;
        RECT 518.000 391.600 518.800 392.400 ;
        RECT 506.800 389.600 507.600 390.400 ;
        RECT 508.400 389.600 509.200 390.400 ;
        RECT 510.000 389.600 510.800 390.400 ;
        RECT 503.600 387.600 504.400 388.400 ;
        RECT 505.200 387.600 506.000 388.400 ;
        RECT 510.000 387.600 510.800 388.400 ;
        RECT 500.400 383.600 501.200 384.400 ;
        RECT 500.500 376.400 501.100 383.600 ;
        RECT 511.700 382.400 512.300 391.600 ;
        RECT 514.800 389.600 515.600 390.400 ;
        RECT 521.200 389.600 522.000 390.400 ;
        RECT 522.900 388.400 523.500 395.600 ;
        RECT 529.300 390.400 529.900 403.600 ;
        RECT 530.900 394.400 531.500 403.600 ;
        RECT 535.600 395.600 536.400 396.400 ;
        RECT 530.800 393.600 531.600 394.400 ;
        RECT 527.600 389.600 528.400 390.400 ;
        RECT 529.200 389.600 530.000 390.400 ;
        RECT 516.400 387.600 517.200 388.400 ;
        RECT 522.800 387.600 523.600 388.400 ;
        RECT 516.400 385.600 517.200 386.400 ;
        RECT 521.200 385.600 522.000 386.400 ;
        RECT 503.600 381.600 504.400 382.400 ;
        RECT 511.600 381.600 512.400 382.400 ;
        RECT 500.400 375.600 501.200 376.400 ;
        RECT 500.400 373.600 501.200 374.400 ;
        RECT 500.500 372.400 501.100 373.600 ;
        RECT 500.400 371.600 501.200 372.400 ;
        RECT 503.700 370.400 504.300 381.600 ;
        RECT 516.500 378.400 517.100 385.600 ;
        RECT 518.000 381.600 518.800 382.400 ;
        RECT 516.400 377.600 517.200 378.400 ;
        RECT 511.600 373.600 512.400 374.400 ;
        RECT 511.700 372.400 512.300 373.600 ;
        RECT 518.100 372.400 518.700 381.600 ;
        RECT 521.300 374.400 521.900 385.600 ;
        RECT 526.000 383.600 526.800 384.400 ;
        RECT 522.800 379.600 523.600 380.400 ;
        RECT 521.200 373.600 522.000 374.400 ;
        RECT 522.900 372.400 523.500 379.600 ;
        RECT 526.100 378.400 526.700 383.600 ;
        RECT 527.700 378.400 528.300 389.600 ;
        RECT 535.700 388.400 536.300 395.600 ;
        RECT 540.400 391.600 541.200 392.400 ;
        RECT 537.200 389.600 538.000 390.400 ;
        RECT 534.000 387.600 534.800 388.400 ;
        RECT 535.600 387.600 536.400 388.400 ;
        RECT 530.800 383.600 531.600 384.400 ;
        RECT 526.000 377.600 526.800 378.400 ;
        RECT 527.600 377.600 528.400 378.400 ;
        RECT 530.800 377.600 531.600 378.400 ;
        RECT 526.000 375.600 526.800 376.400 ;
        RECT 508.400 372.300 509.200 372.400 ;
        RECT 506.900 371.700 509.200 372.300 ;
        RECT 503.600 369.600 504.400 370.400 ;
        RECT 506.900 368.300 507.500 371.700 ;
        RECT 508.400 371.600 509.200 371.700 ;
        RECT 510.000 371.600 510.800 372.400 ;
        RECT 511.600 371.600 512.400 372.400 ;
        RECT 516.400 371.600 517.200 372.400 ;
        RECT 518.000 371.600 518.800 372.400 ;
        RECT 519.600 371.600 520.400 372.400 ;
        RECT 522.800 371.600 523.600 372.400 ;
        RECT 508.400 370.300 509.200 370.400 ;
        RECT 510.100 370.300 510.700 371.600 ;
        RECT 508.400 369.700 510.700 370.300 ;
        RECT 508.400 369.600 509.200 369.700 ;
        RECT 510.100 368.400 510.700 369.700 ;
        RECT 506.900 367.700 509.100 368.300 ;
        RECT 500.400 346.200 501.200 351.800 ;
        RECT 502.000 346.200 502.800 351.800 ;
        RECT 503.600 347.600 504.400 348.400 ;
        RECT 505.200 344.200 506.000 355.800 ;
        RECT 502.000 333.600 502.800 334.400 ;
        RECT 505.200 333.600 506.000 334.400 ;
        RECT 502.100 332.400 502.700 333.600 ;
        RECT 502.000 331.600 502.800 332.400 ;
        RECT 503.600 331.600 504.400 332.400 ;
        RECT 503.700 330.400 504.300 331.600 ;
        RECT 503.600 329.600 504.400 330.400 ;
        RECT 505.300 328.400 505.900 333.600 ;
        RECT 506.800 331.600 507.600 332.400 ;
        RECT 505.200 327.600 506.000 328.400 ;
        RECT 500.400 321.600 501.200 322.400 ;
        RECT 498.800 317.600 499.600 318.400 ;
        RECT 500.500 312.400 501.100 321.600 ;
        RECT 505.200 319.600 506.000 320.400 ;
        RECT 505.300 318.400 505.900 319.600 ;
        RECT 505.200 317.600 506.000 318.400 ;
        RECT 508.500 314.400 509.100 367.700 ;
        RECT 510.000 367.600 510.800 368.400 ;
        RECT 510.000 349.600 510.800 350.400 ;
        RECT 510.000 345.600 510.800 346.400 ;
        RECT 511.600 345.600 512.400 346.400 ;
        RECT 510.100 338.400 510.700 345.600 ;
        RECT 511.700 344.400 512.300 345.600 ;
        RECT 511.600 343.600 512.400 344.400 ;
        RECT 514.800 344.200 515.600 355.800 ;
        RECT 516.500 354.400 517.100 371.600 ;
        RECT 519.700 362.400 520.300 371.600 ;
        RECT 519.600 361.600 520.400 362.400 ;
        RECT 519.600 355.600 520.400 356.400 ;
        RECT 516.400 353.600 517.200 354.400 ;
        RECT 522.900 346.400 523.500 371.600 ;
        RECT 526.100 370.400 526.700 375.600 ;
        RECT 530.900 372.400 531.500 377.600 ;
        RECT 534.100 374.400 534.700 387.600 ;
        RECT 537.300 380.400 537.900 389.600 ;
        RECT 540.500 382.400 541.100 391.600 ;
        RECT 540.400 381.600 541.200 382.400 ;
        RECT 537.200 379.600 538.000 380.400 ;
        RECT 540.400 375.600 541.200 376.400 ;
        RECT 532.400 373.600 533.200 374.400 ;
        RECT 534.000 373.600 534.800 374.400 ;
        RECT 537.200 373.600 538.000 374.400 ;
        RECT 530.800 371.600 531.600 372.400 ;
        RECT 532.500 370.400 533.100 373.600 ;
        RECT 535.600 371.600 536.400 372.400 ;
        RECT 526.000 369.600 526.800 370.400 ;
        RECT 529.200 369.600 530.000 370.400 ;
        RECT 532.400 369.600 533.200 370.400 ;
        RECT 534.000 369.600 534.800 370.400 ;
        RECT 524.400 351.600 525.200 352.400 ;
        RECT 521.200 345.600 522.000 346.400 ;
        RECT 522.800 345.600 523.600 346.400 ;
        RECT 522.800 343.600 523.600 344.400 ;
        RECT 510.000 337.600 510.800 338.400 ;
        RECT 511.700 330.400 512.300 343.600 ;
        RECT 518.000 335.600 518.800 336.400 ;
        RECT 519.600 336.300 520.400 336.400 ;
        RECT 519.600 335.700 523.500 336.300 ;
        RECT 519.600 335.600 520.400 335.700 ;
        RECT 516.400 333.600 517.200 334.400 ;
        RECT 514.800 331.600 515.600 332.400 ;
        RECT 511.600 329.600 512.400 330.400 ;
        RECT 514.900 322.400 515.500 331.600 ;
        RECT 518.100 326.400 518.700 335.600 ;
        RECT 522.900 334.400 523.500 335.700 ;
        RECT 524.500 334.400 525.100 351.600 ;
        RECT 526.000 349.600 526.800 350.400 ;
        RECT 527.600 349.600 528.400 350.400 ;
        RECT 527.700 348.400 528.300 349.600 ;
        RECT 529.300 348.400 529.900 369.600 ;
        RECT 534.100 368.300 534.700 369.600 ;
        RECT 532.500 367.700 534.700 368.300 ;
        RECT 530.800 363.600 531.600 364.400 ;
        RECT 530.900 354.400 531.500 363.600 ;
        RECT 532.500 356.400 533.100 367.700 ;
        RECT 535.700 366.400 536.300 371.600 ;
        RECT 537.300 368.400 537.900 373.600 ;
        RECT 540.500 372.400 541.100 375.600 ;
        RECT 540.400 371.600 541.200 372.400 ;
        RECT 537.200 367.600 538.000 368.400 ;
        RECT 535.600 365.600 536.400 366.400 ;
        RECT 532.400 355.600 533.200 356.400 ;
        RECT 530.800 353.600 531.600 354.400 ;
        RECT 530.900 350.400 531.500 353.600 ;
        RECT 532.500 350.400 533.100 355.600 ;
        RECT 530.800 349.600 531.600 350.400 ;
        RECT 532.400 349.600 533.200 350.400 ;
        RECT 527.600 347.600 528.400 348.400 ;
        RECT 529.200 347.600 530.000 348.400 ;
        RECT 530.800 345.600 531.600 346.400 ;
        RECT 530.900 334.400 531.500 345.600 ;
        RECT 521.200 333.600 522.000 334.400 ;
        RECT 522.800 333.600 523.600 334.400 ;
        RECT 524.400 333.600 525.200 334.400 ;
        RECT 530.800 333.600 531.600 334.400 ;
        RECT 518.000 325.600 518.800 326.400 ;
        RECT 514.800 321.600 515.600 322.400 ;
        RECT 503.600 313.600 504.400 314.400 ;
        RECT 505.200 313.600 506.000 314.400 ;
        RECT 508.400 313.600 509.200 314.400 ;
        RECT 516.400 314.300 517.200 314.400 ;
        RECT 518.000 314.300 518.800 314.400 ;
        RECT 516.400 313.700 518.800 314.300 ;
        RECT 516.400 313.600 517.200 313.700 ;
        RECT 518.000 313.600 518.800 313.700 ;
        RECT 490.800 311.600 491.600 312.400 ;
        RECT 494.000 311.600 494.800 312.400 ;
        RECT 497.200 311.600 498.000 312.400 ;
        RECT 500.400 311.600 501.200 312.400 ;
        RECT 494.100 310.400 494.700 311.600 ;
        RECT 494.000 309.600 494.800 310.400 ;
        RECT 495.600 307.600 496.400 308.400 ;
        RECT 492.400 286.200 493.200 297.800 ;
        RECT 495.700 296.400 496.300 307.600 ;
        RECT 497.300 306.400 497.900 311.600 ;
        RECT 500.500 310.400 501.100 311.600 ;
        RECT 500.400 309.600 501.200 310.400 ;
        RECT 498.800 307.600 499.600 308.400 ;
        RECT 502.000 307.600 502.800 308.400 ;
        RECT 497.200 305.600 498.000 306.400 ;
        RECT 495.600 295.600 496.400 296.400 ;
        RECT 497.200 293.600 498.000 294.400 ;
        RECT 497.300 292.400 497.900 293.600 ;
        RECT 498.900 292.400 499.500 307.600 ;
        RECT 503.700 306.400 504.300 313.600 ;
        RECT 503.600 305.600 504.400 306.400 ;
        RECT 505.300 304.300 505.900 313.600 ;
        RECT 506.800 311.600 507.600 312.400 ;
        RECT 506.900 308.300 507.500 311.600 ;
        RECT 518.100 310.400 518.700 313.600 ;
        RECT 519.600 311.600 520.400 312.400 ;
        RECT 508.400 310.300 509.200 310.400 ;
        RECT 508.400 309.700 510.700 310.300 ;
        RECT 508.400 309.600 509.200 309.700 ;
        RECT 506.900 307.700 509.100 308.300 ;
        RECT 503.700 303.700 505.900 304.300 ;
        RECT 500.400 293.600 501.200 294.400 ;
        RECT 497.200 291.600 498.000 292.400 ;
        RECT 498.800 291.600 499.600 292.400 ;
        RECT 489.200 267.600 490.000 268.400 ;
        RECT 500.500 266.400 501.100 293.600 ;
        RECT 502.000 286.200 502.800 297.800 ;
        RECT 502.000 283.600 502.800 284.400 ;
        RECT 502.100 278.400 502.700 283.600 ;
        RECT 503.700 278.400 504.300 303.700 ;
        RECT 508.500 298.400 509.100 307.700 ;
        RECT 508.400 297.600 509.200 298.400 ;
        RECT 505.200 290.200 506.000 295.800 ;
        RECT 506.800 295.600 507.600 296.400 ;
        RECT 510.100 282.400 510.700 309.700 ;
        RECT 513.200 309.600 514.000 310.400 ;
        RECT 516.400 309.600 517.200 310.400 ;
        RECT 518.000 309.600 518.800 310.400 ;
        RECT 511.600 307.600 512.400 308.400 ;
        RECT 511.700 298.400 512.300 307.600 ;
        RECT 511.600 297.600 512.400 298.400 ;
        RECT 519.700 294.400 520.300 311.600 ;
        RECT 521.300 296.400 521.900 333.600 ;
        RECT 530.900 332.400 531.500 333.600 ;
        RECT 522.800 331.600 523.600 332.400 ;
        RECT 527.600 331.600 528.400 332.400 ;
        RECT 530.800 331.600 531.600 332.400 ;
        RECT 526.000 329.600 526.800 330.400 ;
        RECT 527.700 322.400 528.300 331.600 ;
        RECT 532.500 330.400 533.100 349.600 ;
        RECT 534.000 347.600 534.800 348.400 ;
        RECT 534.100 346.400 534.700 347.600 ;
        RECT 534.000 345.600 534.800 346.400 ;
        RECT 535.700 332.400 536.300 365.600 ;
        RECT 535.600 331.600 536.400 332.400 ;
        RECT 532.400 329.600 533.200 330.400 ;
        RECT 534.000 329.600 534.800 330.400 ;
        RECT 527.600 321.600 528.400 322.400 ;
        RECT 527.700 314.400 528.300 321.600 ;
        RECT 530.800 319.600 531.600 320.400 ;
        RECT 527.600 313.600 528.400 314.400 ;
        RECT 529.200 309.600 530.000 310.400 ;
        RECT 522.800 307.600 523.600 308.400 ;
        RECT 522.900 298.400 523.500 307.600 ;
        RECT 529.300 306.400 529.900 309.600 ;
        RECT 530.900 308.400 531.500 319.600 ;
        RECT 532.400 313.600 533.200 314.400 ;
        RECT 532.500 310.400 533.100 313.600 ;
        RECT 534.100 312.400 534.700 329.600 ;
        RECT 537.300 328.400 537.900 367.600 ;
        RECT 538.800 363.600 539.600 364.400 ;
        RECT 538.900 352.400 539.500 363.600 ;
        RECT 542.100 360.400 542.700 449.600 ;
        RECT 546.900 444.400 547.500 449.600 ;
        RECT 550.000 445.600 550.800 446.400 ;
        RECT 546.800 443.600 547.600 444.400 ;
        RECT 550.100 438.400 550.700 445.600 ;
        RECT 551.700 438.400 552.300 455.600 ;
        RECT 559.700 452.400 560.300 465.600 ;
        RECT 562.900 452.400 563.500 469.600 ;
        RECT 569.200 467.600 570.000 468.400 ;
        RECT 567.600 465.600 568.400 466.400 ;
        RECT 569.300 460.400 569.900 467.600 ;
        RECT 575.700 466.400 576.300 469.600 ;
        RECT 577.200 467.600 578.000 468.400 ;
        RECT 575.600 465.600 576.400 466.400 ;
        RECT 577.200 465.600 578.000 466.400 ;
        RECT 569.200 459.600 570.000 460.400 ;
        RECT 559.600 451.600 560.400 452.400 ;
        RECT 562.800 451.600 563.600 452.400 ;
        RECT 570.800 451.600 571.600 452.400 ;
        RECT 554.800 449.600 555.600 450.400 ;
        RECT 554.900 444.400 555.500 449.600 ;
        RECT 561.200 447.600 562.000 448.400 ;
        RECT 554.800 443.600 555.600 444.400 ;
        RECT 543.600 437.600 544.400 438.400 ;
        RECT 550.000 437.600 550.800 438.400 ;
        RECT 551.600 437.600 552.400 438.400 ;
        RECT 554.900 432.400 555.500 443.600 ;
        RECT 546.800 431.600 547.600 432.400 ;
        RECT 554.800 431.600 555.600 432.400 ;
        RECT 550.000 429.600 550.800 430.400 ;
        RECT 551.600 427.600 552.400 428.400 ;
        RECT 551.700 422.400 552.300 427.600 ;
        RECT 561.300 426.400 561.900 447.600 ;
        RECT 572.400 444.200 573.200 457.800 ;
        RECT 574.000 444.200 574.800 457.800 ;
        RECT 575.600 444.200 576.400 457.800 ;
        RECT 577.200 446.200 578.000 457.800 ;
        RECT 578.900 456.400 579.500 469.600 ;
        RECT 585.200 467.600 586.000 468.400 ;
        RECT 590.100 466.400 590.700 471.600 ;
        RECT 593.200 469.600 594.000 470.400 ;
        RECT 590.000 465.600 590.800 466.400 ;
        RECT 593.300 462.400 593.900 469.600 ;
        RECT 593.200 461.600 594.000 462.400 ;
        RECT 578.800 455.600 579.600 456.400 ;
        RECT 580.400 446.200 581.200 457.800 ;
        RECT 582.000 453.600 582.800 454.400 ;
        RECT 582.100 452.400 582.700 453.600 ;
        RECT 582.000 451.600 582.800 452.400 ;
        RECT 583.600 446.200 584.400 457.800 ;
        RECT 585.200 444.200 586.000 457.800 ;
        RECT 586.800 444.200 587.600 457.800 ;
        RECT 594.900 454.400 595.500 491.600 ;
        RECT 598.000 484.200 598.800 497.800 ;
        RECT 599.600 484.200 600.400 497.800 ;
        RECT 601.200 486.200 602.000 497.800 ;
        RECT 602.800 493.600 603.600 494.400 ;
        RECT 602.900 492.400 603.500 493.600 ;
        RECT 602.800 491.600 603.600 492.400 ;
        RECT 604.400 486.200 605.200 497.800 ;
        RECT 606.000 495.600 606.800 496.400 ;
        RECT 607.600 486.200 608.400 497.800 ;
        RECT 609.200 484.200 610.000 497.800 ;
        RECT 610.800 484.200 611.600 497.800 ;
        RECT 612.400 484.200 613.200 497.800 ;
        RECT 631.600 497.600 632.400 498.400 ;
        RECT 627.000 495.600 627.800 495.800 ;
        RECT 627.000 495.000 632.600 495.600 ;
        RECT 633.200 495.000 634.000 495.800 ;
        RECT 625.200 493.600 626.000 494.400 ;
        RECT 627.000 490.200 627.600 495.000 ;
        RECT 628.400 494.800 629.200 495.000 ;
        RECT 631.800 494.800 632.600 495.000 ;
        RECT 633.400 494.200 634.000 495.000 ;
        RECT 628.400 493.600 634.000 494.200 ;
        RECT 634.800 493.600 635.600 494.400 ;
        RECT 636.400 494.300 637.200 494.400 ;
        RECT 636.400 493.700 638.700 494.300 ;
        RECT 636.400 493.600 637.200 493.700 ;
        RECT 628.400 492.200 629.000 493.600 ;
        RECT 628.200 491.400 629.000 492.200 ;
        RECT 633.400 490.200 634.000 493.600 ;
        RECT 627.000 489.400 627.800 490.200 ;
        RECT 633.200 489.400 634.000 490.200 ;
        RECT 634.900 484.400 635.500 493.600 ;
        RECT 622.000 483.600 622.800 484.400 ;
        RECT 634.800 483.600 635.600 484.400 ;
        RECT 601.200 471.600 602.000 472.400 ;
        RECT 606.000 471.600 606.800 472.400 ;
        RECT 609.200 471.600 610.000 472.400 ;
        RECT 617.200 471.600 618.000 472.400 ;
        RECT 599.600 469.600 600.400 470.400 ;
        RECT 601.300 468.400 601.900 471.600 ;
        RECT 606.100 470.400 606.700 471.600 ;
        RECT 609.300 470.400 609.900 471.600 ;
        RECT 606.000 469.600 606.800 470.400 ;
        RECT 609.200 469.600 610.000 470.400 ;
        RECT 612.400 469.600 613.200 470.400 ;
        RECT 612.500 468.400 613.100 469.600 ;
        RECT 596.400 467.600 597.200 468.400 ;
        RECT 601.200 467.600 602.000 468.400 ;
        RECT 609.200 467.600 610.000 468.400 ;
        RECT 610.800 467.600 611.600 468.400 ;
        RECT 612.400 467.600 613.200 468.400 ;
        RECT 596.500 458.400 597.100 467.600 ;
        RECT 602.800 463.600 603.600 464.400 ;
        RECT 596.400 457.600 597.200 458.400 ;
        RECT 591.600 453.600 592.400 454.400 ;
        RECT 594.800 453.600 595.600 454.400 ;
        RECT 601.200 454.300 602.000 454.400 ;
        RECT 602.900 454.300 603.500 463.600 ;
        RECT 606.000 457.600 606.800 458.400 ;
        RECT 606.100 454.400 606.700 457.600 ;
        RECT 609.300 456.400 609.900 467.600 ;
        RECT 610.900 466.400 611.500 467.600 ;
        RECT 610.800 465.600 611.600 466.400 ;
        RECT 610.800 461.600 611.600 462.400 ;
        RECT 610.900 458.400 611.500 461.600 ;
        RECT 610.800 457.600 611.600 458.400 ;
        RECT 612.500 456.400 613.100 467.600 ;
        RECT 614.000 463.600 614.800 464.400 ;
        RECT 609.200 455.600 610.000 456.400 ;
        RECT 612.400 455.600 613.200 456.400 ;
        RECT 609.300 454.400 609.900 455.600 ;
        RECT 601.200 453.700 603.500 454.300 ;
        RECT 601.200 453.600 602.000 453.700 ;
        RECT 606.000 453.600 606.800 454.400 ;
        RECT 609.200 453.600 610.000 454.400 ;
        RECT 612.400 453.600 613.200 454.400 ;
        RECT 591.700 452.400 592.300 453.600 ;
        RECT 591.600 451.600 592.400 452.400 ;
        RECT 599.600 451.600 600.400 452.400 ;
        RECT 602.800 451.600 603.600 452.400 ;
        RECT 599.700 450.400 600.300 451.600 ;
        RECT 596.400 449.600 597.200 450.400 ;
        RECT 599.600 449.600 600.400 450.400 ;
        RECT 593.200 447.600 594.000 448.400 ;
        RECT 561.200 425.600 562.000 426.400 ;
        RECT 554.800 423.600 555.600 424.400 ;
        RECT 562.800 423.600 563.600 424.400 ;
        RECT 564.400 424.200 565.200 437.800 ;
        RECT 566.000 424.200 566.800 437.800 ;
        RECT 567.600 424.200 568.400 437.800 ;
        RECT 569.200 424.200 570.000 435.800 ;
        RECT 570.800 425.600 571.600 426.400 ;
        RECT 572.400 424.200 573.200 435.800 ;
        RECT 574.000 427.600 574.800 428.400 ;
        RECT 575.600 424.200 576.400 435.800 ;
        RECT 577.200 424.200 578.000 437.800 ;
        RECT 578.800 424.200 579.600 437.800 ;
        RECT 583.600 431.600 584.400 432.400 ;
        RECT 593.300 430.400 593.900 447.600 ;
        RECT 596.400 431.600 597.200 432.400 ;
        RECT 583.600 429.600 584.400 430.400 ;
        RECT 593.200 429.600 594.000 430.400 ;
        RECT 551.600 421.600 552.400 422.400 ;
        RECT 554.900 420.400 555.500 423.600 ;
        RECT 554.800 419.600 555.600 420.400 ;
        RECT 554.800 417.600 555.600 418.400 ;
        RECT 558.000 415.600 558.800 416.400 ;
        RECT 550.000 413.600 550.800 414.400 ;
        RECT 548.400 411.600 549.200 412.400 ;
        RECT 548.500 410.400 549.100 411.600 ;
        RECT 550.100 410.400 550.700 413.600 ;
        RECT 551.600 411.600 552.400 412.400 ;
        RECT 554.800 411.600 555.600 412.400 ;
        RECT 554.900 410.400 555.500 411.600 ;
        RECT 548.400 409.600 549.200 410.400 ;
        RECT 550.000 409.600 550.800 410.400 ;
        RECT 554.800 409.600 555.600 410.400 ;
        RECT 556.400 409.600 557.200 410.400 ;
        RECT 558.100 410.300 558.700 415.600 ;
        RECT 559.600 413.600 560.400 414.400 ;
        RECT 559.700 412.400 560.300 413.600 ;
        RECT 562.900 412.400 563.500 423.600 ;
        RECT 569.200 421.600 570.000 422.400 ;
        RECT 569.300 414.400 569.900 421.600 ;
        RECT 564.400 413.600 565.200 414.400 ;
        RECT 566.000 413.600 566.800 414.400 ;
        RECT 569.200 413.600 570.000 414.400 ;
        RECT 559.600 411.600 560.400 412.400 ;
        RECT 562.800 411.600 563.600 412.400 ;
        RECT 559.600 410.300 560.400 410.400 ;
        RECT 558.100 409.700 560.400 410.300 ;
        RECT 559.600 409.600 560.400 409.700 ;
        RECT 545.200 403.600 546.000 404.400 ;
        RECT 545.300 396.400 545.900 403.600 ;
        RECT 545.200 395.600 546.000 396.400 ;
        RECT 546.800 393.600 547.600 394.400 ;
        RECT 545.200 391.600 546.000 392.400 ;
        RECT 546.900 390.400 547.500 393.600 ;
        RECT 546.800 389.600 547.600 390.400 ;
        RECT 546.800 388.300 547.600 388.400 ;
        RECT 545.300 387.700 547.600 388.300 ;
        RECT 543.600 377.600 544.400 378.400 ;
        RECT 545.300 370.400 545.900 387.700 ;
        RECT 546.800 387.600 547.600 387.700 ;
        RECT 548.400 386.200 549.200 391.800 ;
        RECT 551.600 384.200 552.400 395.800 ;
        RECT 554.800 391.600 555.600 392.400 ;
        RECT 554.900 390.400 555.500 391.600 ;
        RECT 554.800 389.600 555.600 390.400 ;
        RECT 556.400 387.600 557.200 388.400 ;
        RECT 556.500 386.400 557.100 387.600 ;
        RECT 556.400 385.600 557.200 386.400 ;
        RECT 546.800 371.600 547.600 372.400 ;
        RECT 548.400 371.600 549.200 372.400 ;
        RECT 545.200 369.600 546.000 370.400 ;
        RECT 546.900 368.400 547.500 371.600 ;
        RECT 546.800 367.600 547.600 368.400 ;
        RECT 543.600 361.600 544.400 362.400 ;
        RECT 542.000 359.600 542.800 360.400 ;
        RECT 542.000 353.600 542.800 354.400 ;
        RECT 538.800 351.600 539.600 352.400 ;
        RECT 542.100 350.400 542.700 353.600 ;
        RECT 538.800 349.600 539.600 350.400 ;
        RECT 542.000 349.600 542.800 350.400 ;
        RECT 538.900 346.400 539.500 349.600 ;
        RECT 540.400 347.600 541.200 348.400 ;
        RECT 538.800 345.600 539.600 346.400 ;
        RECT 538.900 342.400 539.500 345.600 ;
        RECT 540.500 344.400 541.100 347.600 ;
        RECT 540.400 343.600 541.200 344.400 ;
        RECT 538.800 341.600 539.600 342.400 ;
        RECT 538.800 339.600 539.600 340.400 ;
        RECT 537.200 327.600 538.000 328.400 ;
        RECT 538.900 324.400 539.500 339.600 ;
        RECT 540.400 333.600 541.200 334.400 ;
        RECT 542.100 332.400 542.700 349.600 ;
        RECT 543.700 344.400 544.300 361.600 ;
        RECT 546.900 358.400 547.500 367.600 ;
        RECT 548.500 360.400 549.100 371.600 ;
        RECT 554.800 366.200 555.600 377.800 ;
        RECT 556.500 372.400 557.100 385.600 ;
        RECT 561.200 384.200 562.000 395.800 ;
        RECT 562.900 392.400 563.500 411.600 ;
        RECT 564.500 396.400 565.100 413.600 ;
        RECT 567.600 412.300 568.400 412.400 ;
        RECT 566.100 411.700 568.400 412.300 ;
        RECT 564.400 395.600 565.200 396.400 ;
        RECT 562.800 391.600 563.600 392.400 ;
        RECT 564.400 387.600 565.200 388.400 ;
        RECT 564.500 382.400 565.100 387.600 ;
        RECT 564.400 381.600 565.200 382.400 ;
        RECT 556.400 371.600 557.200 372.400 ;
        RECT 562.800 371.800 563.600 372.600 ;
        RECT 562.900 368.400 563.500 371.800 ;
        RECT 562.800 367.600 563.600 368.400 ;
        RECT 564.400 366.200 565.200 377.800 ;
        RECT 550.000 363.600 550.800 364.400 ;
        RECT 548.400 359.600 549.200 360.400 ;
        RECT 546.800 357.600 547.600 358.400 ;
        RECT 550.100 356.400 550.700 363.600 ;
        RECT 550.000 355.600 550.800 356.400 ;
        RECT 561.200 355.600 562.000 356.400 ;
        RECT 545.200 351.600 546.000 352.400 ;
        RECT 548.400 351.600 549.200 352.400 ;
        RECT 551.600 351.600 552.400 352.400 ;
        RECT 553.200 351.600 554.000 352.400 ;
        RECT 558.000 351.600 558.800 352.400 ;
        RECT 548.400 349.600 549.200 350.400 ;
        RECT 551.600 349.600 552.400 350.400 ;
        RECT 553.300 348.400 553.900 351.600 ;
        RECT 556.400 349.600 557.200 350.400 ;
        RECT 553.200 347.600 554.000 348.400 ;
        RECT 543.600 343.600 544.400 344.400 ;
        RECT 556.500 342.400 557.100 349.600 ;
        RECT 556.400 341.600 557.200 342.400 ;
        RECT 556.400 335.600 557.200 336.400 ;
        RECT 556.500 334.400 557.100 335.600 ;
        RECT 545.200 333.600 546.000 334.400 ;
        RECT 553.200 333.600 554.000 334.400 ;
        RECT 556.400 333.600 557.200 334.400 ;
        RECT 542.000 331.600 542.800 332.400 ;
        RECT 548.400 331.600 549.200 332.400 ;
        RECT 554.800 331.600 555.600 332.400 ;
        RECT 535.600 323.600 536.400 324.400 ;
        RECT 538.800 323.600 539.600 324.400 ;
        RECT 535.700 312.400 536.300 323.600 ;
        RECT 538.900 318.400 539.500 323.600 ;
        RECT 538.800 317.600 539.600 318.400 ;
        RECT 542.100 314.400 542.700 331.600 ;
        RECT 543.600 329.600 544.400 330.400 ;
        RECT 545.200 329.600 546.000 330.400 ;
        RECT 548.400 329.600 549.200 330.400 ;
        RECT 551.600 329.600 552.400 330.400 ;
        RECT 542.000 313.600 542.800 314.400 ;
        RECT 534.000 311.600 534.800 312.400 ;
        RECT 535.600 311.600 536.400 312.400 ;
        RECT 542.000 311.600 542.800 312.400 ;
        RECT 543.700 310.400 544.300 329.600 ;
        RECT 546.800 325.600 547.600 326.400 ;
        RECT 546.900 318.400 547.500 325.600 ;
        RECT 546.800 317.600 547.600 318.400 ;
        RECT 532.400 309.600 533.200 310.400 ;
        RECT 538.800 309.600 539.600 310.400 ;
        RECT 543.600 309.600 544.400 310.400 ;
        RECT 538.900 308.400 539.500 309.600 ;
        RECT 530.800 307.600 531.600 308.400 ;
        RECT 538.800 307.600 539.600 308.400 ;
        RECT 542.000 307.600 542.800 308.400 ;
        RECT 529.200 305.600 530.000 306.400 ;
        RECT 526.000 303.600 526.800 304.400 ;
        RECT 522.800 297.600 523.600 298.400 ;
        RECT 521.200 295.600 522.000 296.400 ;
        RECT 516.400 293.600 517.200 294.400 ;
        RECT 519.600 293.600 520.400 294.400 ;
        RECT 516.500 292.400 517.100 293.600 ;
        RECT 511.600 291.600 512.400 292.400 ;
        RECT 516.400 291.600 517.200 292.400 ;
        RECT 518.000 291.600 518.800 292.400 ;
        RECT 511.700 288.400 512.300 291.600 ;
        RECT 519.700 290.400 520.300 293.600 ;
        RECT 522.900 292.400 523.500 297.600 ;
        RECT 526.100 296.400 526.700 303.600 ;
        RECT 538.800 301.600 539.600 302.400 ;
        RECT 526.000 295.600 526.800 296.400 ;
        RECT 526.100 294.400 526.700 295.600 ;
        RECT 526.000 293.600 526.800 294.400 ;
        RECT 530.800 293.600 531.600 294.400 ;
        RECT 534.000 293.600 534.800 294.400 ;
        RECT 521.200 291.600 522.000 292.400 ;
        RECT 522.800 291.600 523.600 292.400 ;
        RECT 519.600 289.600 520.400 290.400 ;
        RECT 511.600 287.600 512.400 288.400 ;
        RECT 514.800 283.600 515.600 284.400 ;
        RECT 510.000 281.600 510.800 282.400 ;
        RECT 502.000 277.600 502.800 278.400 ;
        RECT 503.600 277.600 504.400 278.400 ;
        RECT 514.900 270.400 515.500 283.600 ;
        RECT 519.700 274.400 520.300 289.600 ;
        RECT 519.600 273.600 520.400 274.400 ;
        RECT 521.300 272.400 521.900 291.600 ;
        RECT 530.900 290.400 531.500 293.600 ;
        RECT 534.100 292.400 534.700 293.600 ;
        RECT 538.900 292.400 539.500 301.600 ;
        RECT 542.100 298.400 542.700 307.600 ;
        RECT 543.700 306.400 544.300 309.600 ;
        RECT 543.600 305.600 544.400 306.400 ;
        RECT 542.000 297.600 542.800 298.400 ;
        RECT 532.400 291.600 533.200 292.400 ;
        RECT 534.000 291.600 534.800 292.400 ;
        RECT 538.800 291.600 539.600 292.400 ;
        RECT 545.200 291.600 546.000 292.400 ;
        RECT 530.800 289.600 531.600 290.400 ;
        RECT 527.600 283.600 528.400 284.400 ;
        RECT 527.700 272.400 528.300 283.600 ;
        RECT 532.400 281.600 533.200 282.400 ;
        RECT 529.200 279.600 530.000 280.400 ;
        RECT 529.300 278.400 529.900 279.600 ;
        RECT 529.200 277.600 530.000 278.400 ;
        RECT 521.200 271.600 522.000 272.400 ;
        RECT 527.600 271.600 528.400 272.400 ;
        RECT 532.500 270.400 533.100 281.600 ;
        RECT 534.100 278.400 534.700 291.600 ;
        RECT 542.000 289.600 542.800 290.400 ;
        RECT 535.600 283.600 536.400 284.400 ;
        RECT 534.000 277.600 534.800 278.400 ;
        RECT 535.700 270.400 536.300 283.600 ;
        RECT 542.100 280.400 542.700 289.600 ;
        RECT 542.000 279.600 542.800 280.400 ;
        RECT 548.500 278.400 549.100 329.600 ;
        RECT 550.000 327.600 550.800 328.400 ;
        RECT 554.900 318.400 555.500 331.600 ;
        RECT 558.100 330.400 558.700 351.600 ;
        RECT 561.300 346.400 561.900 355.600 ;
        RECT 566.100 354.400 566.700 411.700 ;
        RECT 567.600 411.600 568.400 411.700 ;
        RECT 570.800 409.600 571.600 410.400 ;
        RECT 575.600 409.600 576.400 410.400 ;
        RECT 570.900 408.400 571.500 409.600 ;
        RECT 575.700 408.400 576.300 409.600 ;
        RECT 567.600 407.600 568.400 408.400 ;
        RECT 570.800 407.600 571.600 408.400 ;
        RECT 575.600 407.600 576.400 408.400 ;
        RECT 567.700 398.400 568.300 407.600 ;
        RECT 567.600 397.600 568.400 398.400 ;
        RECT 575.700 394.400 576.300 407.600 ;
        RECT 583.700 398.400 584.300 429.600 ;
        RECT 599.700 428.400 600.300 449.600 ;
        RECT 602.900 448.400 603.500 451.600 ;
        RECT 602.800 447.600 603.600 448.400 ;
        RECT 612.500 446.400 613.100 453.600 ;
        RECT 614.100 452.400 614.700 463.600 ;
        RECT 617.300 462.400 617.900 471.600 ;
        RECT 622.100 470.400 622.700 483.600 ;
        RECT 623.600 471.800 624.400 472.600 ;
        RECT 629.800 471.800 630.600 472.600 ;
        RECT 634.900 472.400 635.500 483.600 ;
        RECT 622.000 469.600 622.800 470.400 ;
        RECT 623.600 468.400 624.200 471.800 ;
        RECT 626.800 469.600 627.600 470.400 ;
        RECT 628.600 469.800 629.400 470.600 ;
        RECT 628.600 468.400 629.200 469.800 ;
        RECT 620.400 467.600 621.200 468.400 ;
        RECT 622.000 467.600 622.800 468.400 ;
        RECT 623.600 467.800 629.200 468.400 ;
        RECT 620.500 466.400 621.100 467.600 ;
        RECT 620.400 465.600 621.200 466.400 ;
        RECT 622.100 462.400 622.700 467.600 ;
        RECT 623.600 467.000 624.200 467.800 ;
        RECT 625.000 467.000 625.800 467.200 ;
        RECT 628.400 467.000 629.200 467.200 ;
        RECT 630.000 467.000 630.600 471.800 ;
        RECT 634.800 471.600 635.600 472.400 ;
        RECT 633.200 469.600 634.000 470.400 ;
        RECT 634.800 469.600 635.600 470.400 ;
        RECT 631.600 467.600 632.400 468.400 ;
        RECT 623.600 466.200 624.400 467.000 ;
        RECT 625.000 466.400 630.600 467.000 ;
        RECT 631.700 466.400 632.300 467.600 ;
        RECT 629.800 466.200 630.600 466.400 ;
        RECT 631.600 465.600 632.400 466.400 ;
        RECT 617.200 461.600 618.000 462.400 ;
        RECT 622.000 461.600 622.800 462.400 ;
        RECT 631.600 461.600 632.400 462.400 ;
        RECT 615.600 455.600 616.400 456.400 ;
        RECT 625.200 455.600 626.000 456.400 ;
        RECT 631.700 452.400 632.300 461.600 ;
        RECT 633.300 454.400 633.900 469.600 ;
        RECT 636.400 465.600 637.200 466.400 ;
        RECT 634.800 463.600 635.600 464.400 ;
        RECT 633.200 453.600 634.000 454.400 ;
        RECT 614.000 451.600 614.800 452.400 ;
        RECT 620.400 451.600 621.200 452.400 ;
        RECT 622.000 451.600 622.800 452.400 ;
        RECT 631.600 451.600 632.400 452.400 ;
        RECT 620.500 450.400 621.100 451.600 ;
        RECT 617.200 449.600 618.000 450.400 ;
        RECT 620.400 449.600 621.200 450.400 ;
        RECT 631.700 448.400 632.300 451.600 ;
        RECT 633.200 449.600 634.000 450.400 ;
        RECT 626.800 447.600 627.600 448.400 ;
        RECT 630.000 447.600 630.800 448.400 ;
        RECT 631.600 447.600 632.400 448.400 ;
        RECT 612.400 445.600 613.200 446.400 ;
        RECT 628.400 445.600 629.200 446.400 ;
        RECT 609.200 431.600 610.000 432.400 ;
        RECT 609.300 430.400 609.900 431.600 ;
        RECT 609.200 429.600 610.000 430.400 ;
        RECT 599.600 427.600 600.400 428.400 ;
        RECT 594.800 425.600 595.600 426.400 ;
        RECT 586.800 415.600 587.600 416.400 ;
        RECT 586.900 412.400 587.500 415.600 ;
        RECT 586.800 411.600 587.600 412.400 ;
        RECT 588.400 404.200 589.200 417.800 ;
        RECT 590.000 404.200 590.800 417.800 ;
        RECT 591.600 404.200 592.400 417.800 ;
        RECT 593.200 406.200 594.000 417.800 ;
        RECT 594.900 416.400 595.500 425.600 ;
        RECT 601.200 423.600 602.000 424.400 ;
        RECT 607.600 423.600 608.400 424.400 ;
        RECT 610.800 424.200 611.600 437.800 ;
        RECT 612.400 424.200 613.200 437.800 ;
        RECT 614.000 424.200 614.800 437.800 ;
        RECT 615.600 424.200 616.400 435.800 ;
        RECT 617.200 425.600 618.000 426.400 ;
        RECT 618.800 424.200 619.600 435.800 ;
        RECT 620.400 427.600 621.200 428.400 ;
        RECT 594.800 415.600 595.600 416.400 ;
        RECT 596.400 406.200 597.200 417.800 ;
        RECT 598.000 417.600 598.800 418.400 ;
        RECT 598.100 414.400 598.700 417.600 ;
        RECT 598.000 413.600 598.800 414.400 ;
        RECT 599.600 406.200 600.400 417.800 ;
        RECT 601.200 404.200 602.000 417.800 ;
        RECT 602.800 404.200 603.600 417.800 ;
        RECT 606.000 407.600 606.800 408.400 ;
        RECT 606.100 398.400 606.700 407.600 ;
        RECT 607.700 400.400 608.300 423.600 ;
        RECT 620.500 422.300 621.100 427.600 ;
        RECT 622.000 424.200 622.800 435.800 ;
        RECT 623.600 424.200 624.400 437.800 ;
        RECT 625.200 424.200 626.000 437.800 ;
        RECT 630.000 429.600 630.800 430.400 ;
        RECT 631.600 429.600 632.400 430.400 ;
        RECT 618.900 421.700 621.100 422.300 ;
        RECT 618.900 418.400 619.500 421.700 ;
        RECT 618.800 417.600 619.600 418.400 ;
        RECT 612.400 415.600 613.200 416.400 ;
        RECT 612.500 414.400 613.100 415.600 ;
        RECT 613.800 415.000 614.600 415.800 ;
        RECT 615.600 415.000 619.800 415.600 ;
        RECT 620.400 415.000 621.200 415.800 ;
        RECT 612.400 413.600 613.200 414.400 ;
        RECT 609.200 411.600 610.000 412.400 ;
        RECT 607.600 399.600 608.400 400.400 ;
        RECT 583.600 397.600 584.400 398.400 ;
        RECT 606.000 397.600 606.800 398.400 ;
        RECT 569.200 393.600 570.000 394.400 ;
        RECT 575.600 393.600 576.400 394.400 ;
        RECT 569.300 386.400 569.900 393.600 ;
        RECT 580.400 391.600 581.200 392.400 ;
        RECT 578.800 387.600 579.600 388.400 ;
        RECT 569.200 385.600 570.000 386.400 ;
        RECT 569.300 376.400 569.900 385.600 ;
        RECT 570.800 383.600 571.600 384.400 ;
        RECT 580.500 378.400 581.100 391.600 ;
        RECT 583.600 389.600 584.400 390.400 ;
        RECT 583.700 384.400 584.300 389.600 ;
        RECT 585.200 387.600 586.000 388.400 ;
        RECT 583.600 383.600 584.400 384.400 ;
        RECT 585.300 382.400 585.900 387.600 ;
        RECT 586.800 386.200 587.600 391.800 ;
        RECT 588.400 387.600 589.200 388.400 ;
        RECT 588.500 386.400 589.100 387.600 ;
        RECT 588.400 385.600 589.200 386.400 ;
        RECT 590.000 384.200 590.800 395.800 ;
        RECT 591.600 389.400 592.400 390.400 ;
        RECT 596.400 387.600 597.200 388.400 ;
        RECT 585.200 381.600 586.000 382.400 ;
        RECT 570.800 377.600 571.600 378.400 ;
        RECT 577.200 377.600 578.000 378.400 ;
        RECT 580.400 377.600 581.200 378.400 ;
        RECT 567.600 370.200 568.400 375.800 ;
        RECT 569.200 375.600 570.000 376.400 ;
        RECT 569.200 374.300 570.000 374.400 ;
        RECT 570.900 374.300 571.500 377.600 ;
        RECT 572.400 375.600 573.200 376.400 ;
        RECT 582.000 375.600 582.800 376.400 ;
        RECT 590.000 375.600 590.800 376.400 ;
        RECT 569.200 373.700 571.500 374.300 ;
        RECT 569.200 373.600 570.000 373.700 ;
        RECT 569.200 371.600 570.000 372.400 ;
        RECT 572.500 372.300 573.100 375.600 ;
        RECT 582.100 374.400 582.700 375.600 ;
        RECT 590.100 374.400 590.700 375.600 ;
        RECT 578.800 373.600 579.600 374.400 ;
        RECT 582.000 373.600 582.800 374.400 ;
        RECT 590.000 373.600 590.800 374.400 ;
        RECT 591.600 373.600 592.400 374.400 ;
        RECT 578.900 372.400 579.500 373.600 ;
        RECT 591.700 372.400 592.300 373.600 ;
        RECT 570.900 371.700 573.100 372.300 ;
        RECT 566.000 354.300 566.800 354.400 ;
        RECT 566.000 353.700 568.300 354.300 ;
        RECT 566.000 353.600 566.800 353.700 ;
        RECT 562.800 351.600 563.600 352.400 ;
        RECT 562.800 347.600 563.600 348.400 ;
        RECT 566.000 347.600 566.800 348.400 ;
        RECT 561.200 345.600 562.000 346.400 ;
        RECT 566.100 344.400 566.700 347.600 ;
        RECT 559.600 343.600 560.400 344.400 ;
        RECT 566.000 343.600 566.800 344.400 ;
        RECT 559.700 338.400 560.300 343.600 ;
        RECT 559.600 337.600 560.400 338.400 ;
        RECT 558.000 329.600 558.800 330.400 ;
        RECT 556.400 323.600 557.200 324.400 ;
        RECT 553.200 317.600 554.000 318.400 ;
        RECT 554.800 317.600 555.600 318.400 ;
        RECT 556.500 316.400 557.100 323.600 ;
        RECT 556.400 315.600 557.200 316.400 ;
        RECT 558.100 312.400 558.700 329.600 ;
        RECT 562.800 327.600 563.600 328.400 ;
        RECT 561.200 313.600 562.000 314.400 ;
        RECT 561.300 312.400 561.900 313.600 ;
        RECT 562.900 312.400 563.500 327.600 ;
        RECT 564.400 326.200 565.200 337.800 ;
        RECT 567.700 316.400 568.300 353.700 ;
        RECT 569.300 334.400 569.900 371.600 ;
        RECT 570.900 368.400 571.500 371.700 ;
        RECT 577.200 371.600 578.000 372.400 ;
        RECT 578.800 371.600 579.600 372.400 ;
        RECT 582.000 371.600 582.800 372.400 ;
        RECT 588.400 371.600 589.200 372.400 ;
        RECT 591.600 371.600 592.400 372.400 ;
        RECT 572.400 369.600 573.200 370.400 ;
        RECT 572.500 368.400 573.100 369.600 ;
        RECT 570.800 367.600 571.600 368.400 ;
        RECT 572.400 367.600 573.200 368.400 ;
        RECT 572.500 352.400 573.100 367.600 ;
        RECT 577.300 358.400 577.900 371.600 ;
        RECT 577.200 357.600 578.000 358.400 ;
        RECT 578.800 355.600 579.600 356.400 ;
        RECT 578.900 352.400 579.500 355.600 ;
        RECT 580.400 353.600 581.200 354.400 ;
        RECT 572.400 351.600 573.200 352.400 ;
        RECT 578.800 351.600 579.600 352.400 ;
        RECT 578.900 350.400 579.500 351.600 ;
        RECT 580.500 350.400 581.100 353.600 ;
        RECT 574.000 349.600 574.800 350.400 ;
        RECT 578.800 349.600 579.600 350.400 ;
        RECT 580.400 349.600 581.200 350.400 ;
        RECT 574.100 346.400 574.700 349.600 ;
        RECT 582.100 348.400 582.700 371.600 ;
        RECT 585.200 369.600 586.000 370.400 ;
        RECT 585.300 352.400 585.900 369.600 ;
        RECT 588.500 368.400 589.100 371.600 ;
        RECT 588.400 367.600 589.200 368.400 ;
        RECT 593.200 367.600 594.000 368.400 ;
        RECT 590.000 359.600 590.800 360.400 ;
        RECT 585.200 351.600 586.000 352.400 ;
        RECT 590.100 350.400 590.700 359.600 ;
        RECT 583.600 349.600 584.400 350.400 ;
        RECT 588.400 349.600 589.200 350.400 ;
        RECT 590.000 349.600 590.800 350.400 ;
        RECT 582.000 347.600 582.800 348.400 ;
        RECT 574.000 345.600 574.800 346.400 ;
        RECT 569.200 333.600 570.000 334.400 ;
        RECT 572.400 331.600 573.200 332.600 ;
        RECT 574.000 326.200 574.800 337.800 ;
        RECT 577.200 330.200 578.000 335.800 ;
        RECT 582.100 334.400 582.700 347.600 ;
        RECT 583.700 346.400 584.300 349.600 ;
        RECT 583.600 345.600 584.400 346.400 ;
        RECT 588.500 344.400 589.100 349.600 ;
        RECT 585.200 343.600 586.000 344.400 ;
        RECT 588.400 343.600 589.200 344.400 ;
        RECT 582.000 333.600 582.800 334.400 ;
        RECT 585.300 332.400 585.900 343.600 ;
        RECT 588.500 332.400 589.100 343.600 ;
        RECT 590.100 336.400 590.700 349.600 ;
        RECT 591.600 346.200 592.400 351.800 ;
        RECT 593.300 336.400 593.900 367.600 ;
        RECT 594.800 344.200 595.600 355.800 ;
        RECT 596.500 348.400 597.100 387.600 ;
        RECT 599.600 384.200 600.400 395.800 ;
        RECT 607.700 394.400 608.300 399.600 ;
        RECT 609.300 394.400 609.900 411.600 ;
        RECT 613.800 410.200 614.400 415.000 ;
        RECT 615.600 414.800 616.400 415.000 ;
        RECT 619.000 414.800 619.800 415.000 ;
        RECT 620.600 414.200 621.200 415.000 ;
        RECT 616.400 413.600 621.200 414.200 ;
        RECT 622.000 413.600 622.800 414.400 ;
        RECT 623.600 413.600 624.400 414.400 ;
        RECT 626.800 413.600 627.600 414.400 ;
        RECT 628.400 413.600 629.200 414.400 ;
        RECT 616.400 413.400 617.200 413.600 ;
        RECT 620.600 410.200 621.200 413.600 ;
        RECT 622.000 411.600 622.800 412.400 ;
        RECT 623.700 410.400 624.300 413.600 ;
        RECT 626.900 410.400 627.500 413.600 ;
        RECT 613.800 409.400 614.600 410.200 ;
        RECT 620.400 409.400 621.200 410.200 ;
        RECT 623.600 409.600 624.400 410.400 ;
        RECT 626.800 409.600 627.600 410.400 ;
        RECT 612.400 395.600 613.200 396.400 ;
        RECT 620.400 395.600 621.200 396.400 ;
        RECT 622.000 395.600 622.800 396.400 ;
        RECT 604.400 393.600 605.200 394.400 ;
        RECT 607.600 393.600 608.400 394.400 ;
        RECT 609.200 393.600 610.000 394.400 ;
        RECT 604.400 381.600 605.200 382.400 ;
        RECT 604.500 378.400 605.100 381.600 ;
        RECT 604.400 377.600 605.200 378.400 ;
        RECT 599.600 375.600 600.400 376.400 ;
        RECT 606.000 375.600 606.800 376.400 ;
        RECT 598.000 371.600 598.800 372.400 ;
        RECT 602.800 371.600 603.600 372.400 ;
        RECT 598.000 365.600 598.800 366.400 ;
        RECT 596.400 347.600 597.200 348.400 ;
        RECT 598.100 342.400 598.700 365.600 ;
        RECT 599.600 349.600 600.400 350.400 ;
        RECT 598.000 341.600 598.800 342.400 ;
        RECT 590.000 336.300 590.800 336.400 ;
        RECT 590.000 335.700 592.300 336.300 ;
        RECT 590.000 335.600 590.800 335.700 ;
        RECT 590.000 333.600 590.800 334.400 ;
        RECT 585.200 331.600 586.000 332.400 ;
        RECT 586.800 331.600 587.600 332.400 ;
        RECT 588.400 331.600 589.200 332.400 ;
        RECT 588.400 330.300 589.200 330.400 ;
        RECT 590.100 330.300 590.700 333.600 ;
        RECT 588.400 329.700 590.700 330.300 ;
        RECT 588.400 329.600 589.200 329.700 ;
        RECT 582.000 323.600 582.800 324.400 ;
        RECT 567.600 315.600 568.400 316.400 ;
        RECT 550.000 311.600 550.800 312.400 ;
        RECT 558.000 311.600 558.800 312.400 ;
        RECT 561.200 311.600 562.000 312.400 ;
        RECT 562.800 311.600 563.600 312.400 ;
        RECT 567.700 310.400 568.300 315.600 ;
        RECT 553.200 309.600 554.000 310.400 ;
        RECT 556.400 309.600 557.200 310.400 ;
        RECT 558.000 309.600 558.800 310.400 ;
        RECT 567.600 309.600 568.400 310.400 ;
        RECT 551.600 305.600 552.400 306.400 ;
        RECT 550.000 295.600 550.800 296.400 ;
        RECT 548.400 277.600 549.200 278.400 ;
        RECT 538.800 271.600 539.600 272.400 ;
        RECT 514.800 269.600 515.600 270.400 ;
        RECT 524.400 269.600 525.200 270.400 ;
        RECT 532.400 269.600 533.200 270.400 ;
        RECT 535.600 269.600 536.400 270.400 ;
        RECT 538.800 269.600 539.600 270.400 ;
        RECT 506.800 267.600 507.600 268.400 ;
        RECT 519.600 267.600 520.400 268.400 ;
        RECT 529.200 267.600 530.000 268.400 ;
        RECT 534.000 267.600 534.800 268.400 ;
        RECT 519.700 266.400 520.300 267.600 ;
        RECT 489.200 265.600 490.000 266.400 ;
        RECT 500.400 265.600 501.200 266.400 ;
        RECT 505.200 265.600 506.000 266.400 ;
        RECT 519.600 265.600 520.400 266.400 ;
        RECT 481.200 259.600 482.000 260.400 ;
        RECT 489.300 258.400 489.900 265.600 ;
        RECT 497.200 263.600 498.000 264.400 ;
        RECT 462.000 257.600 462.800 258.400 ;
        RECT 463.600 257.600 464.400 258.400 ;
        RECT 470.000 257.600 470.800 258.400 ;
        RECT 489.200 257.600 490.000 258.400 ;
        RECT 470.100 256.400 470.700 257.600 ;
        RECT 497.300 256.400 497.900 263.600 ;
        RECT 505.300 256.400 505.900 265.600 ;
        RECT 521.200 263.600 522.000 264.400 ;
        RECT 521.300 262.400 521.900 263.600 ;
        RECT 521.200 261.600 522.000 262.400 ;
        RECT 534.100 260.400 534.700 267.600 ;
        RECT 540.400 266.200 541.200 271.800 ;
        RECT 542.000 267.600 542.800 268.400 ;
        RECT 542.100 266.400 542.700 267.600 ;
        RECT 542.000 265.600 542.800 266.400 ;
        RECT 543.600 264.200 544.400 275.800 ;
        RECT 546.800 273.600 547.600 274.400 ;
        RECT 545.200 269.400 546.000 270.400 ;
        RECT 527.600 259.600 528.400 260.400 ;
        RECT 534.000 259.600 534.800 260.400 ;
        RECT 470.000 255.600 470.800 256.400 ;
        RECT 471.600 255.600 472.400 256.400 ;
        RECT 497.200 255.600 498.000 256.400 ;
        RECT 505.200 255.600 506.000 256.400 ;
        RECT 510.000 255.600 510.800 256.400 ;
        RECT 471.700 254.400 472.300 255.600 ;
        RECT 471.600 253.600 472.400 254.400 ;
        RECT 481.200 253.600 482.000 254.400 ;
        RECT 484.400 253.600 485.200 254.400 ;
        RECT 506.800 253.600 507.600 254.400 ;
        RECT 460.400 251.600 461.200 252.400 ;
        RECT 460.500 250.400 461.100 251.600 ;
        RECT 460.400 249.600 461.200 250.400 ;
        RECT 478.000 249.600 478.800 250.400 ;
        RECT 458.800 243.600 459.600 244.400 ;
        RECT 428.400 237.600 429.200 238.400 ;
        RECT 450.800 237.600 451.600 238.400 ;
        RECT 426.800 231.600 427.600 232.400 ;
        RECT 428.500 230.400 429.100 237.600 ;
        RECT 457.200 231.600 458.000 232.400 ;
        RECT 457.300 230.400 457.900 231.600 ;
        RECT 410.800 229.600 411.600 230.400 ;
        RECT 423.600 229.600 424.400 230.400 ;
        RECT 428.400 229.600 429.200 230.400 ;
        RECT 431.600 229.600 432.400 230.400 ;
        RECT 457.200 229.600 458.000 230.400 ;
        RECT 394.800 221.600 395.600 222.400 ;
        RECT 390.000 191.600 390.800 192.400 ;
        RECT 393.200 191.600 394.000 192.400 ;
        RECT 393.300 188.400 393.900 191.600 ;
        RECT 388.400 187.600 389.200 188.400 ;
        RECT 393.200 187.600 394.000 188.400 ;
        RECT 394.900 184.300 395.500 221.600 ;
        RECT 401.200 219.600 402.000 220.400 ;
        RECT 396.400 213.600 397.200 214.400 ;
        RECT 396.400 211.600 397.200 212.400 ;
        RECT 398.000 212.300 398.800 212.400 ;
        RECT 398.000 211.700 400.300 212.300 ;
        RECT 398.000 211.600 398.800 211.700 ;
        RECT 396.400 205.600 397.200 206.400 ;
        RECT 396.500 198.400 397.100 205.600 ;
        RECT 396.400 197.600 397.200 198.400 ;
        RECT 398.000 193.600 398.800 194.400 ;
        RECT 396.400 189.600 397.200 190.400 ;
        RECT 396.500 186.400 397.100 189.600 ;
        RECT 396.400 185.600 397.200 186.400 ;
        RECT 394.900 183.700 397.100 184.300 ;
        RECT 386.800 173.600 387.600 174.400 ;
        RECT 394.800 173.600 395.600 174.400 ;
        RECT 394.900 172.400 395.500 173.600 ;
        RECT 396.500 172.400 397.100 183.700 ;
        RECT 394.800 171.600 395.600 172.400 ;
        RECT 396.400 171.600 397.200 172.400 ;
        RECT 398.000 163.600 398.800 164.400 ;
        RECT 398.100 158.300 398.700 163.600 ;
        RECT 399.700 158.400 400.300 211.700 ;
        RECT 401.300 210.400 401.900 219.600 ;
        RECT 410.900 212.400 411.500 229.600 ;
        RECT 431.700 228.400 432.300 229.600 ;
        RECT 431.600 227.600 432.400 228.400 ;
        RECT 439.600 227.600 440.400 228.400 ;
        RECT 423.600 225.600 424.400 226.400 ;
        RECT 425.200 225.600 426.000 226.400 ;
        RECT 436.400 225.600 437.200 226.400 ;
        RECT 406.000 211.600 406.800 212.400 ;
        RECT 410.800 211.600 411.600 212.400 ;
        RECT 401.200 209.600 402.000 210.400 ;
        RECT 401.300 208.400 401.900 209.600 ;
        RECT 401.200 207.600 402.000 208.400 ;
        RECT 402.800 203.600 403.600 204.400 ;
        RECT 402.900 198.400 403.500 203.600 ;
        RECT 402.800 197.600 403.600 198.400 ;
        RECT 404.400 193.600 405.200 194.400 ;
        RECT 401.200 191.600 402.000 192.400 ;
        RECT 402.800 189.600 403.600 190.400 ;
        RECT 406.100 176.400 406.700 211.600 ;
        RECT 415.600 204.200 416.400 217.800 ;
        RECT 417.200 204.200 418.000 217.800 ;
        RECT 418.800 206.200 419.600 217.800 ;
        RECT 420.400 213.600 421.200 214.400 ;
        RECT 422.000 206.200 422.800 217.800 ;
        RECT 423.700 216.400 424.300 225.600 ;
        RECT 423.600 215.600 424.400 216.400 ;
        RECT 425.200 206.200 426.000 217.800 ;
        RECT 426.800 204.200 427.600 217.800 ;
        RECT 428.400 204.200 429.200 217.800 ;
        RECT 430.000 204.200 430.800 217.800 ;
        RECT 417.200 197.600 418.000 198.400 ;
        RECT 428.400 197.600 429.200 198.400 ;
        RECT 417.300 190.400 417.900 197.600 ;
        RECT 436.500 192.400 437.100 225.600 ;
        RECT 439.700 208.400 440.300 227.600 ;
        RECT 450.800 223.600 451.600 224.400 ;
        RECT 450.900 216.400 451.500 223.600 ;
        RECT 450.800 215.600 451.600 216.400 ;
        RECT 442.800 211.600 443.600 212.400 ;
        RECT 450.600 211.600 451.600 212.400 ;
        RECT 439.600 207.600 440.400 208.400 ;
        RECT 439.600 203.600 440.400 204.400 ;
        RECT 446.000 203.600 446.800 204.400 ;
        RECT 439.700 202.400 440.300 203.600 ;
        RECT 439.600 201.600 440.400 202.400 ;
        RECT 446.100 198.400 446.700 203.600 ;
        RECT 436.400 191.600 437.200 192.400 ;
        RECT 417.200 189.600 418.000 190.400 ;
        RECT 407.600 187.600 408.400 188.400 ;
        RECT 407.700 182.400 408.300 187.600 ;
        RECT 409.200 183.600 410.000 184.400 ;
        RECT 412.400 183.600 413.200 184.400 ;
        RECT 407.600 181.600 408.400 182.400 ;
        RECT 407.700 178.400 408.300 181.600 ;
        RECT 409.300 180.400 409.900 183.600 ;
        RECT 409.200 179.600 410.000 180.400 ;
        RECT 412.500 178.400 413.100 183.600 ;
        RECT 417.300 178.400 417.900 189.600 ;
        RECT 420.400 187.600 421.200 188.400 ;
        RECT 433.200 185.600 434.000 186.400 ;
        RECT 407.600 177.600 408.400 178.400 ;
        RECT 412.400 177.600 413.200 178.400 ;
        RECT 417.200 177.600 418.000 178.400 ;
        RECT 406.000 175.600 406.800 176.400 ;
        RECT 401.200 171.600 402.000 172.400 ;
        RECT 425.200 171.600 426.000 172.400 ;
        RECT 401.300 168.400 401.900 171.600 ;
        RECT 401.200 167.600 402.000 168.400 ;
        RECT 422.000 167.600 422.800 168.400 ;
        RECT 425.300 168.300 425.900 171.600 ;
        RECT 423.700 167.700 425.900 168.300 ;
        RECT 422.100 158.400 422.700 167.600 ;
        RECT 380.400 149.600 381.200 150.400 ;
        RECT 386.800 149.600 387.600 150.400 ;
        RECT 391.600 144.200 392.400 157.800 ;
        RECT 393.200 144.200 394.000 157.800 ;
        RECT 396.500 157.700 398.700 158.300 ;
        RECT 394.800 144.200 395.600 155.800 ;
        RECT 396.500 148.400 397.100 157.700 ;
        RECT 399.600 157.600 400.400 158.400 ;
        RECT 396.400 147.600 397.200 148.400 ;
        RECT 398.000 144.200 398.800 155.800 ;
        RECT 399.600 145.600 400.400 146.400 ;
        RECT 399.700 142.400 400.300 145.600 ;
        RECT 401.200 144.200 402.000 155.800 ;
        RECT 402.800 144.200 403.600 157.800 ;
        RECT 404.400 144.200 405.200 157.800 ;
        RECT 406.000 144.200 406.800 157.800 ;
        RECT 422.000 157.600 422.800 158.400 ;
        RECT 407.600 149.600 408.400 150.400 ;
        RECT 415.600 145.600 416.400 146.400 ;
        RECT 367.600 141.600 368.400 142.400 ;
        RECT 399.600 141.600 400.400 142.400 ;
        RECT 410.800 141.600 411.600 142.400 ;
        RECT 345.200 135.600 346.000 136.400 ;
        RECT 346.800 135.600 347.600 136.400 ;
        RECT 337.200 131.600 338.000 132.400 ;
        RECT 342.000 131.600 342.800 132.400 ;
        RECT 350.000 131.600 350.800 132.400 ;
        RECT 335.600 125.600 336.400 126.400 ;
        RECT 329.200 113.600 330.000 114.400 ;
        RECT 326.000 111.600 326.800 112.400 ;
        RECT 327.600 107.600 328.400 108.400 ;
        RECT 314.800 105.600 315.600 106.400 ;
        RECT 324.400 105.600 325.200 106.400 ;
        RECT 311.600 95.600 312.400 96.400 ;
        RECT 308.400 89.600 309.200 90.400 ;
        RECT 306.800 67.600 307.600 68.400 ;
        RECT 305.200 63.600 306.000 64.400 ;
        RECT 306.900 60.300 307.500 67.600 ;
        RECT 310.000 64.200 310.800 77.800 ;
        RECT 311.600 64.200 312.400 77.800 ;
        RECT 313.200 64.200 314.000 75.800 ;
        RECT 314.900 74.400 315.500 105.600 ;
        RECT 316.400 101.600 317.200 102.400 ;
        RECT 316.500 92.400 317.100 101.600 ;
        RECT 316.400 91.600 317.200 92.400 ;
        RECT 318.000 84.200 318.800 97.800 ;
        RECT 319.600 84.200 320.400 97.800 ;
        RECT 321.200 84.200 322.000 97.800 ;
        RECT 322.800 86.200 323.600 97.800 ;
        RECT 324.500 96.400 325.100 105.600 ;
        RECT 324.400 95.600 325.200 96.400 ;
        RECT 326.000 86.200 326.800 97.800 ;
        RECT 327.600 93.600 328.400 94.400 ;
        RECT 329.200 86.200 330.000 97.800 ;
        RECT 330.800 84.200 331.600 97.800 ;
        RECT 332.400 84.200 333.200 97.800 ;
        RECT 314.800 73.600 315.600 74.400 ;
        RECT 314.800 67.600 315.600 68.400 ;
        RECT 314.900 66.400 315.500 67.600 ;
        RECT 314.800 65.600 315.600 66.400 ;
        RECT 316.400 64.200 317.200 75.800 ;
        RECT 318.000 65.600 318.800 66.400 ;
        RECT 306.900 59.700 309.100 60.300 ;
        RECT 306.800 57.600 307.600 58.400 ;
        RECT 302.000 55.600 302.800 56.400 ;
        RECT 306.900 52.400 307.500 57.600 ;
        RECT 308.500 54.400 309.100 59.700 ;
        RECT 310.000 55.600 310.800 56.400 ;
        RECT 310.100 54.400 310.700 55.600 ;
        RECT 308.400 53.600 309.200 54.400 ;
        RECT 310.000 53.600 310.800 54.400 ;
        RECT 306.800 51.600 307.600 52.400 ;
        RECT 295.600 49.600 296.400 50.400 ;
        RECT 298.800 49.600 299.600 50.400 ;
        RECT 302.000 49.600 302.800 50.400 ;
        RECT 313.200 47.600 314.000 48.400 ;
        RECT 311.600 43.600 312.400 44.400 ;
        RECT 290.800 37.600 291.600 38.400 ;
        RECT 302.000 33.600 302.800 34.400 ;
        RECT 302.100 30.400 302.700 33.600 ;
        RECT 311.700 32.400 312.300 43.600 ;
        RECT 308.400 31.600 309.200 32.400 ;
        RECT 311.600 31.600 312.400 32.400 ;
        RECT 257.200 29.600 258.000 30.400 ;
        RECT 271.600 29.600 272.400 30.400 ;
        RECT 276.400 29.600 277.200 30.400 ;
        RECT 289.200 29.600 290.000 30.400 ;
        RECT 302.000 29.600 302.800 30.400 ;
        RECT 305.200 29.600 306.000 30.400 ;
        RECT 308.400 29.600 309.200 30.400 ;
        RECT 257.300 26.400 257.900 29.600 ;
        RECT 257.200 25.600 258.000 26.400 ;
        RECT 260.400 23.600 261.200 24.400 ;
        RECT 265.200 23.600 266.000 24.400 ;
        RECT 260.500 16.400 261.100 23.600 ;
        RECT 271.700 18.400 272.300 29.600 ;
        RECT 302.100 28.400 302.700 29.600 ;
        RECT 313.300 28.400 313.900 47.600 ;
        RECT 273.200 27.600 274.000 28.400 ;
        RECT 276.400 27.600 277.200 28.400 ;
        RECT 284.400 27.600 285.200 28.400 ;
        RECT 302.000 27.600 302.800 28.400 ;
        RECT 303.600 27.600 304.400 28.400 ;
        RECT 313.200 27.600 314.000 28.400 ;
        RECT 266.800 17.600 267.600 18.400 ;
        RECT 271.600 17.600 272.400 18.400 ;
        RECT 276.500 16.400 277.100 27.600 ;
        RECT 292.400 25.600 293.200 26.400 ;
        RECT 308.400 25.600 309.200 26.400 ;
        RECT 286.000 23.600 286.800 24.400 ;
        RECT 290.800 23.600 291.600 24.400 ;
        RECT 236.400 15.600 237.200 16.400 ;
        RECT 244.400 15.600 245.200 16.400 ;
        RECT 250.800 15.600 251.600 16.400 ;
        RECT 260.400 15.600 261.200 16.400 ;
        RECT 273.200 15.600 274.000 16.400 ;
        RECT 276.400 15.600 277.200 16.400 ;
        RECT 282.800 15.600 283.600 16.400 ;
        RECT 236.500 14.400 237.100 15.600 ;
        RECT 250.900 14.400 251.500 15.600 ;
        RECT 236.400 13.600 237.200 14.400 ;
        RECT 239.600 13.600 240.400 14.400 ;
        RECT 250.800 13.600 251.600 14.400 ;
        RECT 239.700 12.400 240.300 13.600 ;
        RECT 260.500 12.400 261.100 15.600 ;
        RECT 273.300 14.400 273.900 15.600 ;
        RECT 276.500 14.400 277.100 15.600 ;
        RECT 273.200 13.600 274.000 14.400 ;
        RECT 276.400 13.600 277.200 14.400 ;
        RECT 282.800 13.600 283.600 14.400 ;
        RECT 273.300 12.400 273.900 13.600 ;
        RECT 225.200 11.600 226.000 12.400 ;
        RECT 234.800 11.600 235.600 12.400 ;
        RECT 238.000 11.600 238.800 12.400 ;
        RECT 239.600 11.600 240.400 12.400 ;
        RECT 247.600 11.600 248.400 12.400 ;
        RECT 260.400 11.600 261.200 12.400 ;
        RECT 273.200 11.600 274.000 12.400 ;
        RECT 286.100 10.400 286.700 23.600 ;
        RECT 290.900 18.400 291.500 23.600 ;
        RECT 290.800 17.600 291.600 18.400 ;
        RECT 292.500 12.400 293.100 25.600 ;
        RECT 314.800 23.600 315.600 24.400 ;
        RECT 318.100 18.400 318.700 65.600 ;
        RECT 319.600 64.200 320.400 75.800 ;
        RECT 321.200 64.200 322.000 77.800 ;
        RECT 322.800 64.200 323.600 77.800 ;
        RECT 324.400 64.200 325.200 77.800 ;
        RECT 334.000 73.600 334.800 74.400 ;
        RECT 335.700 64.400 336.300 125.600 ;
        RECT 337.300 110.400 337.900 131.600 ;
        RECT 342.100 126.400 342.700 131.600 ;
        RECT 342.000 125.600 342.800 126.400 ;
        RECT 350.100 126.300 350.700 131.600 ;
        RECT 350.100 125.700 352.300 126.300 ;
        RECT 342.000 123.600 342.800 124.400 ;
        RECT 350.000 123.600 350.800 124.400 ;
        RECT 342.100 120.400 342.700 123.600 ;
        RECT 342.000 119.600 342.800 120.400 ;
        RECT 350.100 118.400 350.700 123.600 ;
        RECT 351.700 120.400 352.300 125.700 ;
        RECT 359.600 124.200 360.400 137.800 ;
        RECT 361.200 124.200 362.000 137.800 ;
        RECT 362.800 126.200 363.600 137.800 ;
        RECT 364.400 133.600 365.200 134.400 ;
        RECT 364.500 122.400 365.100 133.600 ;
        RECT 366.000 126.200 366.800 137.800 ;
        RECT 367.700 136.400 368.300 141.600 ;
        RECT 367.600 135.600 368.400 136.400 ;
        RECT 369.200 126.200 370.000 137.800 ;
        RECT 370.800 124.200 371.600 137.800 ;
        RECT 372.400 124.200 373.200 137.800 ;
        RECT 374.000 124.200 374.800 137.800 ;
        RECT 394.800 137.600 395.600 138.400 ;
        RECT 391.600 133.600 392.400 134.400 ;
        RECT 391.700 132.400 392.300 133.600 ;
        RECT 375.600 131.600 376.400 132.400 ;
        RECT 391.600 131.600 392.400 132.400 ;
        RECT 402.800 131.600 403.600 132.400 ;
        RECT 383.600 123.600 384.400 124.400 ;
        RECT 388.400 123.600 389.200 124.400 ;
        RECT 401.200 123.600 402.000 124.400 ;
        RECT 404.400 124.200 405.200 137.800 ;
        RECT 406.000 124.200 406.800 137.800 ;
        RECT 407.600 124.200 408.400 137.800 ;
        RECT 409.200 126.200 410.000 137.800 ;
        RECT 410.900 136.400 411.500 141.600 ;
        RECT 414.000 139.600 414.800 140.400 ;
        RECT 410.800 135.600 411.600 136.400 ;
        RECT 412.400 126.200 413.200 137.800 ;
        RECT 414.100 134.400 414.700 139.600 ;
        RECT 414.000 133.600 414.800 134.400 ;
        RECT 415.600 126.200 416.400 137.800 ;
        RECT 417.200 124.200 418.000 137.800 ;
        RECT 418.800 124.200 419.600 137.800 ;
        RECT 423.700 132.400 424.300 167.700 ;
        RECT 426.800 164.200 427.600 177.800 ;
        RECT 428.400 164.200 429.200 177.800 ;
        RECT 430.000 164.200 430.800 177.800 ;
        RECT 431.600 166.200 432.400 177.800 ;
        RECT 433.300 176.400 433.900 185.600 ;
        RECT 438.000 184.200 438.800 197.800 ;
        RECT 439.600 184.200 440.400 197.800 ;
        RECT 441.200 184.200 442.000 197.800 ;
        RECT 446.000 197.600 446.800 198.400 ;
        RECT 442.800 184.200 443.600 195.800 ;
        RECT 444.400 185.600 445.200 186.400 ;
        RECT 446.000 184.200 446.800 195.800 ;
        RECT 447.600 187.600 448.400 188.400 ;
        RECT 447.700 182.400 448.300 187.600 ;
        RECT 449.200 184.200 450.000 195.800 ;
        RECT 450.800 184.200 451.600 197.800 ;
        RECT 452.400 184.200 453.200 197.800 ;
        RECT 455.600 191.600 456.400 192.400 ;
        RECT 447.600 181.600 448.400 182.400 ;
        RECT 452.400 181.600 453.200 182.400 ;
        RECT 452.500 178.400 453.100 181.600 ;
        RECT 433.200 175.600 434.000 176.400 ;
        RECT 428.400 157.600 429.200 158.400 ;
        RECT 428.500 150.400 429.100 157.600 ;
        RECT 431.600 151.600 432.400 152.400 ;
        RECT 428.400 149.600 429.200 150.400 ;
        RECT 426.800 147.600 427.600 148.400 ;
        RECT 425.200 145.600 426.000 146.400 ;
        RECT 425.300 136.400 425.900 145.600 ;
        RECT 425.200 135.600 426.000 136.400 ;
        RECT 423.600 131.600 424.400 132.400 ;
        RECT 423.700 126.400 424.300 131.600 ;
        RECT 423.600 125.600 424.400 126.400 ;
        RECT 364.400 121.600 365.200 122.400 ;
        RECT 388.500 120.400 389.100 123.600 ;
        RECT 351.600 119.600 352.400 120.400 ;
        RECT 364.400 119.600 365.200 120.400 ;
        RECT 388.400 119.600 389.200 120.400 ;
        RECT 391.600 119.600 392.400 120.400 ;
        RECT 399.600 119.600 400.400 120.400 ;
        RECT 364.500 118.400 365.100 119.600 ;
        RECT 337.200 109.600 338.000 110.400 ;
        RECT 337.300 92.400 337.900 109.600 ;
        RECT 338.800 104.200 339.600 117.800 ;
        RECT 340.400 104.200 341.200 117.800 ;
        RECT 342.000 104.200 342.800 117.800 ;
        RECT 350.000 117.600 350.800 118.400 ;
        RECT 343.600 104.200 344.400 115.800 ;
        RECT 345.200 105.600 346.000 106.400 ;
        RECT 346.800 104.200 347.600 115.800 ;
        RECT 348.400 107.600 349.200 108.400 ;
        RECT 350.000 104.200 350.800 115.800 ;
        RECT 351.600 104.200 352.400 117.800 ;
        RECT 353.200 104.200 354.000 117.800 ;
        RECT 364.400 117.600 365.200 118.400 ;
        RECT 369.200 109.600 370.000 110.400 ;
        RECT 372.400 109.600 373.200 110.400 ;
        RECT 361.200 105.600 362.000 106.400 ;
        RECT 358.000 99.600 358.800 100.400 ;
        RECT 342.000 95.600 342.800 96.400 ;
        RECT 337.200 91.600 338.000 92.400 ;
        RECT 343.600 83.600 344.400 84.400 ;
        RECT 353.200 84.200 354.000 97.800 ;
        RECT 354.800 84.200 355.600 97.800 ;
        RECT 356.400 86.200 357.200 97.800 ;
        RECT 358.100 94.400 358.700 99.600 ;
        RECT 358.000 93.600 358.800 94.400 ;
        RECT 359.600 86.200 360.400 97.800 ;
        RECT 361.300 96.400 361.900 105.600 ;
        RECT 364.400 103.600 365.200 104.400 ;
        RECT 364.500 100.400 365.100 103.600 ;
        RECT 364.400 99.600 365.200 100.400 ;
        RECT 361.200 95.600 362.000 96.400 ;
        RECT 343.700 72.400 344.300 83.600 ;
        RECT 343.600 71.600 344.400 72.400 ;
        RECT 343.600 69.600 344.400 70.400 ;
        RECT 335.600 63.600 336.400 64.400 ;
        RECT 326.000 44.200 326.800 57.800 ;
        RECT 327.600 44.200 328.400 57.800 ;
        RECT 329.200 44.200 330.000 57.800 ;
        RECT 330.800 46.200 331.600 57.800 ;
        RECT 332.400 55.600 333.200 56.400 ;
        RECT 334.000 46.200 334.800 57.800 ;
        RECT 335.700 54.400 336.300 63.600 ;
        RECT 335.600 53.600 336.400 54.400 ;
        RECT 337.200 46.200 338.000 57.800 ;
        RECT 338.800 44.200 339.600 57.800 ;
        RECT 340.400 44.200 341.200 57.800 ;
        RECT 343.700 52.400 344.300 69.600 ;
        RECT 345.200 64.200 346.000 77.800 ;
        RECT 346.800 64.200 347.600 77.800 ;
        RECT 348.400 64.200 349.200 75.800 ;
        RECT 350.000 71.600 350.800 72.400 ;
        RECT 350.100 68.400 350.700 71.600 ;
        RECT 350.000 67.600 350.800 68.400 ;
        RECT 351.600 64.200 352.400 75.800 ;
        RECT 353.200 73.600 354.000 74.400 ;
        RECT 353.300 66.400 353.900 73.600 ;
        RECT 353.200 65.600 354.000 66.400 ;
        RECT 354.800 64.200 355.600 75.800 ;
        RECT 356.400 64.200 357.200 77.800 ;
        RECT 358.000 64.200 358.800 77.800 ;
        RECT 359.600 64.200 360.400 77.800 ;
        RECT 361.300 74.400 361.900 95.600 ;
        RECT 362.800 86.200 363.600 97.800 ;
        RECT 364.400 84.200 365.200 97.800 ;
        RECT 366.000 84.200 366.800 97.800 ;
        RECT 367.600 84.200 368.400 97.800 ;
        RECT 369.300 92.400 369.900 109.600 ;
        RECT 374.000 104.200 374.800 117.800 ;
        RECT 375.600 104.200 376.400 117.800 ;
        RECT 377.200 104.200 378.000 117.800 ;
        RECT 378.800 104.200 379.600 115.800 ;
        RECT 380.400 105.600 381.200 106.400 ;
        RECT 382.000 104.200 382.800 115.800 ;
        RECT 383.600 107.600 384.400 108.400 ;
        RECT 383.600 105.600 384.400 106.400 ;
        RECT 380.400 93.600 381.200 94.400 ;
        RECT 369.200 91.600 370.000 92.400 ;
        RECT 382.000 91.600 382.800 92.400 ;
        RECT 369.300 80.300 369.900 91.600 ;
        RECT 377.200 83.600 378.000 84.400 ;
        RECT 367.700 79.700 369.900 80.300 ;
        RECT 361.200 73.600 362.000 74.400 ;
        RECT 348.400 61.600 349.200 62.400 ;
        RECT 343.600 51.600 344.400 52.400 ;
        RECT 322.800 29.600 323.600 30.400 ;
        RECT 321.200 23.600 322.000 24.400 ;
        RECT 292.400 11.600 293.200 12.400 ;
        RECT 244.400 9.600 245.200 10.400 ;
        RECT 250.800 9.600 251.600 10.400 ;
        RECT 254.000 9.600 254.800 10.400 ;
        RECT 281.200 9.600 282.000 10.400 ;
        RECT 286.000 9.600 286.800 10.400 ;
        RECT 294.000 4.200 294.800 17.800 ;
        RECT 295.600 4.200 296.400 17.800 ;
        RECT 297.200 4.200 298.000 17.800 ;
        RECT 298.800 6.200 299.600 17.800 ;
        RECT 300.400 17.600 301.200 18.400 ;
        RECT 300.500 16.400 301.100 17.600 ;
        RECT 300.400 15.600 301.200 16.400 ;
        RECT 302.000 6.200 302.800 17.800 ;
        RECT 303.600 15.600 304.400 16.400 ;
        RECT 303.700 14.400 304.300 15.600 ;
        RECT 303.600 13.600 304.400 14.400 ;
        RECT 305.200 6.200 306.000 17.800 ;
        RECT 306.800 4.200 307.600 17.800 ;
        RECT 308.400 4.200 309.200 17.800 ;
        RECT 318.000 17.600 318.800 18.400 ;
        RECT 321.300 12.400 321.900 23.600 ;
        RECT 322.900 22.300 323.500 29.600 ;
        RECT 324.400 24.200 325.200 37.800 ;
        RECT 326.000 24.200 326.800 37.800 ;
        RECT 327.600 24.200 328.400 37.800 ;
        RECT 329.200 24.200 330.000 35.800 ;
        RECT 330.800 25.600 331.600 26.400 ;
        RECT 322.900 21.700 325.100 22.300 ;
        RECT 324.500 18.400 325.100 21.700 ;
        RECT 330.900 18.400 331.500 25.600 ;
        RECT 332.400 24.200 333.200 35.800 ;
        RECT 334.000 27.600 334.800 28.400 ;
        RECT 334.100 26.400 334.700 27.600 ;
        RECT 334.000 25.600 334.800 26.400 ;
        RECT 335.600 24.200 336.400 35.800 ;
        RECT 337.200 24.200 338.000 37.800 ;
        RECT 338.800 24.200 339.600 37.800 ;
        RECT 343.700 30.400 344.300 51.600 ;
        RECT 348.500 34.400 349.100 61.600 ;
        RECT 359.600 57.600 360.400 58.400 ;
        RECT 367.700 52.400 368.300 79.700 ;
        RECT 377.300 74.400 377.900 83.600 ;
        RECT 383.700 78.400 384.300 105.600 ;
        RECT 385.200 104.200 386.000 115.800 ;
        RECT 386.800 104.200 387.600 117.800 ;
        RECT 388.400 104.200 389.200 117.800 ;
        RECT 390.000 95.600 390.800 96.400 ;
        RECT 391.700 94.400 392.300 119.600 ;
        RECT 393.200 117.600 394.000 118.400 ;
        RECT 391.600 93.600 392.400 94.400 ;
        RECT 393.300 92.400 393.900 117.600 ;
        RECT 399.700 110.400 400.300 119.600 ;
        RECT 401.300 114.400 401.900 123.600 ;
        RECT 409.200 121.600 410.000 122.400 ;
        RECT 409.300 118.400 409.900 121.600 ;
        RECT 404.400 117.600 405.200 118.400 ;
        RECT 409.200 117.600 410.000 118.400 ;
        RECT 415.600 117.600 416.400 118.400 ;
        RECT 401.200 113.600 402.000 114.400 ;
        RECT 404.500 110.400 405.100 117.600 ;
        RECT 412.400 115.600 413.200 116.400 ;
        RECT 412.500 114.400 413.100 115.600 ;
        RECT 410.800 113.600 411.600 114.400 ;
        RECT 412.400 113.600 413.200 114.400 ;
        RECT 410.900 112.400 411.500 113.600 ;
        RECT 410.800 111.600 411.600 112.400 ;
        RECT 415.700 110.400 416.300 117.600 ;
        RECT 425.200 115.600 426.000 116.400 ;
        RECT 426.900 110.400 427.500 147.600 ;
        RECT 428.500 118.400 429.100 149.600 ;
        RECT 431.700 138.400 432.300 151.600 ;
        RECT 433.300 142.400 433.900 175.600 ;
        RECT 434.800 166.200 435.600 177.800 ;
        RECT 436.400 177.600 437.200 178.400 ;
        RECT 436.500 174.400 437.100 177.600 ;
        RECT 436.400 173.600 437.200 174.400 ;
        RECT 438.000 166.200 438.800 177.800 ;
        RECT 439.600 164.200 440.400 177.800 ;
        RECT 441.200 164.200 442.000 177.800 ;
        RECT 452.400 177.600 453.200 178.400 ;
        RECT 455.700 176.400 456.300 191.600 ;
        RECT 457.200 189.600 458.000 190.400 ;
        RECT 450.800 175.600 451.600 176.400 ;
        RECT 455.600 175.600 456.400 176.400 ;
        RECT 450.900 174.400 451.500 175.600 ;
        RECT 450.800 173.600 451.600 174.400 ;
        RECT 457.300 172.400 457.900 189.600 ;
        RECT 458.900 182.400 459.500 243.600 ;
        RECT 462.000 224.200 462.800 237.800 ;
        RECT 463.600 224.200 464.400 237.800 ;
        RECT 465.200 224.200 466.000 235.800 ;
        RECT 466.800 227.600 467.600 228.400 ;
        RECT 468.400 224.200 469.200 235.800 ;
        RECT 470.000 225.600 470.800 226.400 ;
        RECT 470.100 218.400 470.700 225.600 ;
        RECT 471.600 224.200 472.400 235.800 ;
        RECT 473.200 224.200 474.000 237.800 ;
        RECT 474.800 224.200 475.600 237.800 ;
        RECT 476.400 224.200 477.200 237.800 ;
        RECT 478.100 230.400 478.700 249.600 ;
        RECT 478.000 229.600 478.800 230.400 ;
        RECT 460.400 204.200 461.200 217.800 ;
        RECT 462.000 204.200 462.800 217.800 ;
        RECT 463.600 204.200 464.400 217.800 ;
        RECT 465.200 206.200 466.000 217.800 ;
        RECT 466.800 215.600 467.600 216.400 ;
        RECT 468.400 206.200 469.200 217.800 ;
        RECT 470.000 217.600 470.800 218.400 ;
        RECT 470.000 215.600 470.800 216.400 ;
        RECT 470.100 214.400 470.700 215.600 ;
        RECT 470.000 213.600 470.800 214.400 ;
        RECT 471.600 206.200 472.400 217.800 ;
        RECT 473.200 204.200 474.000 217.800 ;
        RECT 474.800 204.200 475.600 217.800 ;
        RECT 476.400 213.600 477.200 214.400 ;
        RECT 466.800 197.600 467.600 198.400 ;
        RECT 466.900 196.400 467.500 197.600 ;
        RECT 465.200 195.600 466.000 196.400 ;
        RECT 466.800 195.600 467.600 196.400 ;
        RECT 465.300 192.400 465.900 195.600 ;
        RECT 462.000 191.600 462.800 192.400 ;
        RECT 465.200 191.600 466.000 192.400 ;
        RECT 462.100 190.400 462.700 191.600 ;
        RECT 462.000 189.600 462.800 190.400 ;
        RECT 465.200 189.600 466.000 190.400 ;
        RECT 466.900 188.400 467.500 195.600 ;
        RECT 476.500 190.400 477.100 213.600 ;
        RECT 479.600 209.600 480.400 210.400 ;
        RECT 481.300 194.400 481.900 253.600 ;
        RECT 486.000 251.600 486.800 252.400 ;
        RECT 487.600 251.600 488.400 252.400 ;
        RECT 498.800 251.600 499.600 252.400 ;
        RECT 500.400 251.600 501.200 252.400 ;
        RECT 514.800 251.600 515.600 252.400 ;
        RECT 482.800 233.600 483.600 234.400 ;
        RECT 481.200 193.600 482.000 194.400 ;
        RECT 468.400 189.600 469.200 190.400 ;
        RECT 476.400 189.600 477.200 190.400 ;
        RECT 468.500 188.400 469.100 189.600 ;
        RECT 481.300 188.400 481.900 193.600 ;
        RECT 482.900 190.400 483.500 233.600 ;
        RECT 486.000 225.600 486.800 226.400 ;
        RECT 486.100 224.400 486.700 225.600 ;
        RECT 486.000 224.300 486.800 224.400 ;
        RECT 484.500 223.700 486.800 224.300 ;
        RECT 484.500 216.400 485.100 223.700 ;
        RECT 486.000 223.600 486.800 223.700 ;
        RECT 484.400 215.600 485.200 216.400 ;
        RECT 486.000 203.600 486.800 204.400 ;
        RECT 484.400 191.600 485.200 192.400 ;
        RECT 484.500 190.400 485.100 191.600 ;
        RECT 482.800 189.600 483.600 190.400 ;
        RECT 484.400 189.600 485.200 190.400 ;
        RECT 465.200 187.600 466.000 188.400 ;
        RECT 466.800 187.600 467.600 188.400 ;
        RECT 468.400 187.600 469.200 188.400 ;
        RECT 481.200 187.600 482.000 188.400 ;
        RECT 462.000 183.600 462.800 184.400 ;
        RECT 458.800 181.600 459.600 182.400 ;
        RECT 458.800 177.600 459.600 178.400 ;
        RECT 462.100 174.400 462.700 183.600 ;
        RECT 458.800 173.600 459.600 174.400 ;
        RECT 462.000 173.600 462.800 174.400 ;
        RECT 447.600 171.600 448.400 172.400 ;
        RECT 457.200 171.600 458.000 172.400 ;
        RECT 458.900 170.400 459.500 173.600 ;
        RECT 465.300 172.400 465.900 187.600 ;
        RECT 463.600 171.600 464.400 172.400 ;
        RECT 465.200 171.600 466.000 172.400 ;
        RECT 454.000 169.600 454.800 170.400 ;
        RECT 458.800 169.600 459.600 170.400 ;
        RECT 454.100 164.400 454.700 169.600 ;
        RECT 454.000 163.600 454.800 164.400 ;
        RECT 457.200 163.600 458.000 164.400 ;
        RECT 465.200 163.600 466.000 164.400 ;
        RECT 466.800 163.600 467.600 164.400 ;
        RECT 457.300 160.400 457.900 163.600 ;
        RECT 457.200 159.600 458.000 160.400 ;
        RECT 436.400 153.600 437.200 154.400 ;
        RECT 436.500 152.400 437.100 153.600 ;
        RECT 436.400 151.600 437.200 152.400 ;
        RECT 441.200 149.600 442.000 150.400 ;
        RECT 434.800 143.600 435.600 144.400 ;
        RECT 433.200 141.600 434.000 142.400 ;
        RECT 434.900 140.400 435.500 143.600 ;
        RECT 434.800 139.600 435.600 140.400 ;
        RECT 431.600 137.600 432.400 138.400 ;
        RECT 438.000 135.600 438.800 136.400 ;
        RECT 441.300 132.400 441.900 149.600 ;
        RECT 446.000 144.200 446.800 157.800 ;
        RECT 447.600 144.200 448.400 157.800 ;
        RECT 449.200 144.200 450.000 155.800 ;
        RECT 450.800 147.600 451.600 148.400 ;
        RECT 452.400 144.200 453.200 155.800 ;
        RECT 454.000 145.600 454.800 146.400 ;
        RECT 454.100 142.400 454.700 145.600 ;
        RECT 455.600 144.200 456.400 155.800 ;
        RECT 457.200 144.200 458.000 157.800 ;
        RECT 458.800 144.200 459.600 157.800 ;
        RECT 460.400 144.200 461.200 157.800 ;
        RECT 462.000 149.600 462.800 150.400 ;
        RECT 454.000 141.600 454.800 142.400 ;
        RECT 457.200 141.600 458.000 142.400 ;
        RECT 436.400 131.600 437.200 132.400 ;
        RECT 441.200 131.600 442.000 132.400 ;
        RECT 444.400 131.600 445.200 132.400 ;
        RECT 433.200 125.600 434.000 126.400 ;
        RECT 430.000 123.600 430.800 124.400 ;
        RECT 428.400 117.600 429.200 118.400 ;
        RECT 399.600 109.600 400.400 110.400 ;
        RECT 404.400 109.600 405.200 110.400 ;
        RECT 406.000 109.600 406.800 110.400 ;
        RECT 415.600 109.600 416.400 110.400 ;
        RECT 426.800 109.600 427.600 110.400 ;
        RECT 398.000 107.600 398.800 108.400 ;
        RECT 399.700 106.400 400.300 109.600 ;
        RECT 406.100 108.400 406.700 109.600 ;
        RECT 402.800 107.600 403.600 108.400 ;
        RECT 406.000 107.600 406.800 108.400 ;
        RECT 407.600 107.600 408.400 108.400 ;
        RECT 417.200 107.600 418.000 108.400 ;
        RECT 399.600 105.600 400.400 106.400 ;
        RECT 425.200 105.600 426.000 106.400 ;
        RECT 412.400 103.600 413.200 104.400 ;
        RECT 412.500 94.400 413.100 103.600 ;
        RECT 412.400 93.600 413.200 94.400 ;
        RECT 393.200 91.600 394.000 92.400 ;
        RECT 394.800 91.600 395.600 92.400 ;
        RECT 401.200 91.600 402.000 92.400 ;
        RECT 386.800 89.600 387.600 90.400 ;
        RECT 390.000 90.300 390.800 90.400 ;
        RECT 394.900 90.300 395.500 91.600 ;
        RECT 401.300 90.400 401.900 91.600 ;
        RECT 390.000 89.700 395.500 90.300 ;
        RECT 390.000 89.600 390.800 89.700 ;
        RECT 401.200 89.600 402.000 90.400 ;
        RECT 409.200 89.600 410.000 90.400 ;
        RECT 398.000 87.600 398.800 88.400 ;
        RECT 383.600 77.600 384.400 78.400 ;
        RECT 377.200 73.600 378.000 74.400 ;
        RECT 390.000 73.600 390.800 74.400 ;
        RECT 396.400 73.600 397.200 74.400 ;
        RECT 390.100 68.400 390.700 73.600 ;
        RECT 396.500 72.400 397.100 73.600 ;
        RECT 398.100 72.400 398.700 87.600 ;
        RECT 399.600 83.600 400.400 84.400 ;
        RECT 418.800 84.200 419.600 97.800 ;
        RECT 420.400 84.200 421.200 97.800 ;
        RECT 422.000 84.200 422.800 97.800 ;
        RECT 423.600 86.200 424.400 97.800 ;
        RECT 425.300 96.400 425.900 105.600 ;
        RECT 428.500 98.400 429.100 117.600 ;
        RECT 430.100 108.400 430.700 123.600 ;
        RECT 433.300 110.400 433.900 125.600 ;
        RECT 439.600 123.600 440.400 124.400 ;
        RECT 449.200 124.200 450.000 137.800 ;
        RECT 450.800 124.200 451.600 137.800 ;
        RECT 452.400 126.200 453.200 137.800 ;
        RECT 454.000 133.600 454.800 134.400 ;
        RECT 455.600 126.200 456.400 137.800 ;
        RECT 457.300 136.400 457.900 141.600 ;
        RECT 457.200 135.600 458.000 136.400 ;
        RECT 439.700 118.400 440.300 123.600 ;
        RECT 433.200 109.600 434.000 110.400 ;
        RECT 430.000 107.600 430.800 108.400 ;
        RECT 430.100 100.400 430.700 107.600 ;
        RECT 434.800 104.200 435.600 117.800 ;
        RECT 436.400 104.200 437.200 117.800 ;
        RECT 438.000 104.200 438.800 117.800 ;
        RECT 439.600 117.600 440.400 118.400 ;
        RECT 439.600 104.200 440.400 115.800 ;
        RECT 441.200 105.600 442.000 106.400 ;
        RECT 442.800 104.200 443.600 115.800 ;
        RECT 444.400 107.600 445.200 108.400 ;
        RECT 430.000 99.600 430.800 100.400 ;
        RECT 444.500 98.400 445.100 107.600 ;
        RECT 446.000 104.200 446.800 115.800 ;
        RECT 447.600 104.200 448.400 117.800 ;
        RECT 449.200 104.200 450.000 117.800 ;
        RECT 454.000 109.600 454.800 110.400 ;
        RECT 450.800 107.600 451.600 108.400 ;
        RECT 450.900 98.400 451.500 107.600 ;
        RECT 457.300 106.400 457.900 135.600 ;
        RECT 458.800 126.200 459.600 137.800 ;
        RECT 460.400 124.200 461.200 137.800 ;
        RECT 462.000 124.200 462.800 137.800 ;
        RECT 463.600 124.200 464.400 137.800 ;
        RECT 465.300 118.400 465.900 163.600 ;
        RECT 466.900 148.400 467.500 163.600 ;
        RECT 466.800 147.600 467.600 148.400 ;
        RECT 465.200 117.600 466.000 118.400 ;
        RECT 463.600 112.300 464.400 112.400 ;
        RECT 462.100 111.700 464.400 112.300 ;
        RECT 458.800 109.600 459.600 110.400 ;
        RECT 458.900 108.400 459.500 109.600 ;
        RECT 458.800 107.600 459.600 108.400 ;
        RECT 457.200 105.600 458.000 106.400 ;
        RECT 452.400 99.600 453.200 100.400 ;
        RECT 460.400 99.600 461.200 100.400 ;
        RECT 425.200 95.600 426.000 96.400 ;
        RECT 426.800 86.200 427.600 97.800 ;
        RECT 428.400 97.600 429.200 98.400 ;
        RECT 428.400 95.600 429.200 96.400 ;
        RECT 428.500 94.400 429.100 95.600 ;
        RECT 428.400 93.600 429.200 94.400 ;
        RECT 430.000 86.200 430.800 97.800 ;
        RECT 431.600 84.200 432.400 97.800 ;
        RECT 433.200 84.200 434.000 97.800 ;
        RECT 444.400 97.600 445.200 98.400 ;
        RECT 450.800 97.600 451.600 98.400 ;
        RECT 442.800 93.600 443.600 94.400 ;
        RECT 450.900 92.400 451.500 97.600 ;
        RECT 452.500 94.400 453.100 99.600 ;
        RECT 457.200 95.600 458.000 96.400 ;
        RECT 452.400 93.600 453.200 94.400 ;
        RECT 457.300 92.400 457.900 95.600 ;
        RECT 460.500 94.400 461.100 99.600 ;
        RECT 458.800 93.600 459.600 94.400 ;
        RECT 460.400 93.600 461.200 94.400 ;
        RECT 438.000 91.600 438.800 92.400 ;
        RECT 449.200 91.600 450.000 92.400 ;
        RECT 450.800 91.600 451.600 92.400 ;
        RECT 457.200 91.600 458.000 92.400 ;
        RECT 438.100 88.400 438.700 91.600 ;
        RECT 446.000 89.600 446.800 90.400 ;
        RECT 438.000 87.600 438.800 88.400 ;
        RECT 439.600 87.600 440.400 88.400 ;
        RECT 396.400 71.600 397.200 72.400 ;
        RECT 398.000 71.600 398.800 72.400 ;
        RECT 399.700 70.400 400.300 83.600 ;
        RECT 404.400 71.600 405.200 72.400 ;
        RECT 399.600 69.600 400.400 70.400 ;
        RECT 372.400 67.600 373.200 68.400 ;
        RECT 390.000 67.600 390.800 68.400 ;
        RECT 401.200 67.600 402.000 68.400 ;
        RECT 369.200 63.600 370.000 64.400 ;
        RECT 372.500 62.400 373.100 67.600 ;
        RECT 386.800 65.600 387.600 66.400 ;
        RECT 372.400 61.600 373.200 62.400 ;
        RECT 378.800 59.600 379.600 60.400 ;
        RECT 358.000 51.600 358.800 52.400 ;
        RECT 367.600 51.600 368.400 52.400 ;
        RECT 359.600 43.600 360.400 44.400 ;
        RECT 369.200 44.200 370.000 57.800 ;
        RECT 370.800 44.200 371.600 57.800 ;
        RECT 372.400 44.200 373.200 57.800 ;
        RECT 374.000 46.200 374.800 57.800 ;
        RECT 375.600 55.600 376.400 56.400 ;
        RECT 375.700 44.300 376.300 55.600 ;
        RECT 377.200 46.200 378.000 57.800 ;
        RECT 378.900 54.400 379.500 59.600 ;
        RECT 386.900 58.400 387.500 65.600 ;
        RECT 378.800 53.600 379.600 54.400 ;
        RECT 378.800 51.600 379.600 52.400 ;
        RECT 375.700 43.700 377.900 44.300 ;
        RECT 348.400 33.600 349.200 34.400 ;
        RECT 343.600 29.600 344.400 30.400 ;
        RECT 348.500 28.400 349.100 33.600 ;
        RECT 359.700 30.400 360.300 43.600 ;
        RECT 370.800 39.600 371.600 40.400 ;
        RECT 370.900 32.400 371.500 39.600 ;
        RECT 370.800 31.600 371.600 32.400 ;
        RECT 359.600 29.600 360.400 30.400 ;
        RECT 370.800 29.600 371.600 30.400 ;
        RECT 348.400 27.600 349.200 28.400 ;
        RECT 366.000 27.600 366.800 28.400 ;
        RECT 369.200 27.600 370.000 28.400 ;
        RECT 362.800 25.600 363.600 26.400 ;
        RECT 359.600 23.600 360.400 24.400 ;
        RECT 337.200 21.600 338.000 22.400 ;
        RECT 337.300 18.400 337.900 21.600 ;
        RECT 359.700 20.400 360.300 23.600 ;
        RECT 362.900 22.400 363.500 25.600 ;
        RECT 362.800 21.600 363.600 22.400 ;
        RECT 353.200 19.600 354.000 20.400 ;
        RECT 359.600 19.600 360.400 20.400 ;
        RECT 324.400 17.600 325.200 18.400 ;
        RECT 330.800 17.600 331.600 18.400 ;
        RECT 337.200 17.600 338.000 18.400 ;
        RECT 324.500 12.400 325.100 17.600 ;
        RECT 313.200 11.600 314.000 12.400 ;
        RECT 321.200 11.600 322.000 12.400 ;
        RECT 324.400 11.600 325.200 12.400 ;
        RECT 346.800 4.200 347.600 17.800 ;
        RECT 348.400 4.200 349.200 17.800 ;
        RECT 350.000 4.200 350.800 17.800 ;
        RECT 351.600 6.200 352.400 17.800 ;
        RECT 353.300 16.400 353.900 19.600 ;
        RECT 353.200 15.600 354.000 16.400 ;
        RECT 354.800 6.200 355.600 17.800 ;
        RECT 356.400 13.600 357.200 14.400 ;
        RECT 358.000 6.200 358.800 17.800 ;
        RECT 359.600 4.200 360.400 17.800 ;
        RECT 361.200 4.200 362.000 17.800 ;
        RECT 369.300 14.400 369.900 27.600 ;
        RECT 369.200 13.600 370.000 14.400 ;
        RECT 370.900 12.400 371.500 29.600 ;
        RECT 375.600 23.600 376.400 24.400 ;
        RECT 375.700 12.400 376.300 23.600 ;
        RECT 377.300 20.400 377.900 43.700 ;
        RECT 378.900 30.400 379.500 51.600 ;
        RECT 380.400 46.200 381.200 57.800 ;
        RECT 382.000 44.200 382.800 57.800 ;
        RECT 383.600 44.200 384.400 57.800 ;
        RECT 386.800 57.600 387.600 58.400 ;
        RECT 390.100 54.400 390.700 67.600 ;
        RECT 394.800 63.600 395.600 64.400 ;
        RECT 394.900 60.400 395.500 63.600 ;
        RECT 394.800 59.600 395.600 60.400 ;
        RECT 399.600 57.600 400.400 58.400 ;
        RECT 401.300 54.400 401.900 67.600 ;
        RECT 407.600 63.600 408.400 64.400 ;
        RECT 422.000 64.200 422.800 77.800 ;
        RECT 423.600 64.200 424.400 77.800 ;
        RECT 425.200 64.200 426.000 77.800 ;
        RECT 426.800 64.200 427.600 75.800 ;
        RECT 428.400 65.600 429.200 66.400 ;
        RECT 390.000 53.600 390.800 54.400 ;
        RECT 393.200 53.600 394.000 54.400 ;
        RECT 401.200 53.600 402.000 54.400 ;
        RECT 394.800 43.600 395.600 44.400 ;
        RECT 394.900 40.400 395.500 43.600 ;
        RECT 394.800 39.600 395.600 40.400 ;
        RECT 378.800 29.600 379.600 30.400 ;
        RECT 377.200 19.600 378.000 20.400 ;
        RECT 378.900 12.400 379.500 29.600 ;
        RECT 380.400 24.200 381.200 37.800 ;
        RECT 382.000 24.200 382.800 37.800 ;
        RECT 383.600 24.200 384.400 35.800 ;
        RECT 385.200 33.600 386.000 34.400 ;
        RECT 385.300 28.400 385.900 33.600 ;
        RECT 385.200 27.600 386.000 28.400 ;
        RECT 386.800 24.200 387.600 35.800 ;
        RECT 388.400 25.600 389.200 26.400 ;
        RECT 388.500 20.400 389.100 25.600 ;
        RECT 390.000 24.200 390.800 35.800 ;
        RECT 391.600 24.200 392.400 37.800 ;
        RECT 393.200 24.200 394.000 37.800 ;
        RECT 394.800 24.200 395.600 37.800 ;
        RECT 401.300 28.400 401.900 53.600 ;
        RECT 407.700 36.400 408.300 63.600 ;
        RECT 418.800 59.600 419.600 60.400 ;
        RECT 409.200 44.200 410.000 57.800 ;
        RECT 410.800 44.200 411.600 57.800 ;
        RECT 412.400 44.200 413.200 57.800 ;
        RECT 414.000 46.200 414.800 57.800 ;
        RECT 415.600 55.600 416.400 56.400 ;
        RECT 417.200 46.200 418.000 57.800 ;
        RECT 418.900 54.400 419.500 59.600 ;
        RECT 418.800 53.600 419.600 54.400 ;
        RECT 420.400 46.200 421.200 57.800 ;
        RECT 422.000 44.200 422.800 57.800 ;
        RECT 423.600 44.200 424.400 57.800 ;
        RECT 428.500 56.400 429.100 65.600 ;
        RECT 430.000 64.200 430.800 75.800 ;
        RECT 431.600 69.600 432.400 70.400 ;
        RECT 431.700 68.400 432.300 69.600 ;
        RECT 431.600 67.600 432.400 68.400 ;
        RECT 433.200 64.200 434.000 75.800 ;
        RECT 434.800 64.200 435.600 77.800 ;
        RECT 436.400 64.200 437.200 77.800 ;
        RECT 439.700 70.400 440.300 87.600 ;
        RECT 446.100 82.400 446.700 89.600 ;
        RECT 447.600 87.600 448.400 88.400 ;
        RECT 446.000 81.600 446.800 82.400 ;
        RECT 446.100 72.400 446.700 81.600 ;
        RECT 446.000 71.600 446.800 72.400 ;
        RECT 439.600 69.600 440.400 70.400 ;
        RECT 428.400 55.600 429.200 56.400 ;
        RECT 439.700 52.400 440.300 69.600 ;
        RECT 446.000 63.600 446.800 64.400 ;
        RECT 446.100 60.400 446.700 63.600 ;
        RECT 446.000 59.600 446.800 60.400 ;
        RECT 447.700 58.400 448.300 87.600 ;
        RECT 449.300 68.400 449.900 91.600 ;
        RECT 454.000 90.300 454.800 90.400 ;
        RECT 454.000 89.700 456.300 90.300 ;
        RECT 454.000 89.600 454.800 89.700 ;
        RECT 450.800 72.300 451.600 72.400 ;
        RECT 450.800 71.700 453.100 72.300 ;
        RECT 450.800 71.600 451.600 71.700 ;
        RECT 449.200 67.600 450.000 68.400 ;
        RECT 450.800 63.600 451.600 64.400 ;
        RECT 450.900 62.400 451.500 63.600 ;
        RECT 450.800 61.600 451.600 62.400 ;
        RECT 452.500 58.400 453.100 71.700 ;
        RECT 454.000 69.600 454.800 70.400 ;
        RECT 455.700 58.400 456.300 89.700 ;
        RECT 457.200 83.600 458.000 84.400 ;
        RECT 457.200 68.300 458.000 68.400 ;
        RECT 458.900 68.300 459.500 93.600 ;
        RECT 460.400 91.600 461.200 92.400 ;
        RECT 462.100 78.400 462.700 111.700 ;
        RECT 463.600 111.600 464.400 111.700 ;
        RECT 463.700 110.400 464.300 111.600 ;
        RECT 463.600 109.600 464.400 110.400 ;
        RECT 466.800 109.600 467.600 110.400 ;
        RECT 466.900 108.400 467.500 109.600 ;
        RECT 465.200 107.600 466.000 108.400 ;
        RECT 466.800 108.300 467.600 108.400 ;
        RECT 468.500 108.300 469.100 187.600 ;
        RECT 470.000 185.600 470.800 186.400 ;
        RECT 474.800 183.600 475.600 184.400 ;
        RECT 474.900 172.400 475.500 183.600 ;
        RECT 482.900 172.400 483.500 189.600 ;
        RECT 484.400 175.600 485.200 176.400 ;
        RECT 471.600 171.600 472.400 172.400 ;
        RECT 473.200 171.600 474.000 172.400 ;
        RECT 474.800 171.600 475.600 172.400 ;
        RECT 482.800 171.600 483.600 172.400 ;
        RECT 471.700 170.300 472.300 171.600 ;
        RECT 482.900 170.300 483.500 171.600 ;
        RECT 484.400 170.300 485.200 170.400 ;
        RECT 471.700 169.700 473.900 170.300 ;
        RECT 482.900 169.700 485.200 170.300 ;
        RECT 473.300 158.400 473.900 169.700 ;
        RECT 484.400 169.600 485.200 169.700 ;
        RECT 486.100 164.400 486.700 203.600 ;
        RECT 487.700 192.400 488.300 251.600 ;
        RECT 500.500 248.400 501.100 251.600 ;
        RECT 514.900 250.400 515.500 251.600 ;
        RECT 514.800 249.600 515.600 250.400 ;
        RECT 490.800 247.600 491.600 248.400 ;
        RECT 500.400 247.600 501.200 248.400 ;
        RECT 489.200 233.600 490.000 234.400 ;
        RECT 489.300 230.400 489.900 233.600 ;
        RECT 490.900 230.400 491.500 247.600 ;
        RECT 519.600 244.200 520.400 257.800 ;
        RECT 521.200 244.200 522.000 257.800 ;
        RECT 522.800 246.200 523.600 257.800 ;
        RECT 524.400 253.600 525.200 254.400 ;
        RECT 526.000 246.200 526.800 257.800 ;
        RECT 527.700 256.400 528.300 259.600 ;
        RECT 546.900 258.400 547.500 273.600 ;
        RECT 550.100 264.400 550.700 295.600 ;
        RECT 551.700 292.400 552.300 305.600 ;
        RECT 553.300 296.400 553.900 309.600 ;
        RECT 556.500 308.400 557.100 309.600 ;
        RECT 554.800 307.600 555.600 308.400 ;
        RECT 556.400 307.600 557.200 308.400 ;
        RECT 558.100 306.300 558.700 309.600 ;
        RECT 559.600 307.600 560.400 308.400 ;
        RECT 562.800 307.600 563.600 308.400 ;
        RECT 569.200 307.600 570.000 308.400 ;
        RECT 556.500 305.700 558.700 306.300 ;
        RECT 553.200 295.600 554.000 296.400 ;
        RECT 551.600 291.600 552.400 292.400 ;
        RECT 556.500 284.400 557.100 305.700 ;
        RECT 559.700 298.400 560.300 307.600 ;
        RECT 569.300 302.400 569.900 307.600 ;
        RECT 570.800 305.600 571.600 306.400 ;
        RECT 577.200 306.200 578.000 311.800 ;
        RECT 578.800 307.600 579.600 308.400 ;
        RECT 570.900 304.400 571.500 305.600 ;
        RECT 570.800 303.600 571.600 304.400 ;
        RECT 569.200 301.600 570.000 302.400 ;
        RECT 559.600 297.600 560.400 298.400 ;
        RECT 558.000 290.200 558.800 295.800 ;
        RECT 561.200 286.200 562.000 297.800 ;
        RECT 569.200 293.600 570.000 294.400 ;
        RECT 569.300 292.400 569.900 293.600 ;
        RECT 564.400 291.600 565.200 292.400 ;
        RECT 569.200 291.600 570.000 292.400 ;
        RECT 562.800 287.600 563.600 288.400 ;
        RECT 554.800 283.600 555.600 284.400 ;
        RECT 556.400 283.600 557.200 284.400 ;
        RECT 550.000 263.600 550.800 264.400 ;
        RECT 553.200 264.200 554.000 275.800 ;
        RECT 527.600 255.600 528.400 256.400 ;
        RECT 529.200 246.200 530.000 257.800 ;
        RECT 530.800 244.200 531.600 257.800 ;
        RECT 532.400 244.200 533.200 257.800 ;
        RECT 534.000 244.200 534.800 257.800 ;
        RECT 546.800 257.600 547.600 258.400 ;
        RECT 543.600 255.600 544.400 256.400 ;
        RECT 551.600 246.200 552.400 257.800 ;
        RECT 553.200 257.600 554.000 258.400 ;
        RECT 489.200 229.600 490.000 230.400 ;
        RECT 490.800 229.600 491.600 230.400 ;
        RECT 506.800 229.600 507.600 230.400 ;
        RECT 492.400 227.600 493.200 228.400 ;
        RECT 492.500 226.400 493.100 227.600 ;
        RECT 492.400 225.600 493.200 226.400 ;
        RECT 500.400 225.600 501.200 226.400 ;
        RECT 506.900 222.400 507.500 229.600 ;
        RECT 510.000 224.200 510.800 237.800 ;
        RECT 511.600 224.200 512.400 237.800 ;
        RECT 513.200 224.200 514.000 235.800 ;
        RECT 514.800 227.600 515.600 228.400 ;
        RECT 516.400 224.200 517.200 235.800 ;
        RECT 518.000 225.600 518.800 226.400 ;
        RECT 506.800 221.600 507.600 222.400 ;
        RECT 511.600 221.600 512.400 222.400 ;
        RECT 489.200 211.600 490.000 212.400 ;
        RECT 489.300 210.400 489.900 211.600 ;
        RECT 489.200 209.600 490.000 210.400 ;
        RECT 495.600 204.200 496.400 217.800 ;
        RECT 497.200 204.200 498.000 217.800 ;
        RECT 498.800 206.200 499.600 217.800 ;
        RECT 500.400 213.600 501.200 214.400 ;
        RECT 500.400 211.600 501.200 212.400 ;
        RECT 494.000 201.600 494.800 202.400 ;
        RECT 487.600 191.600 488.400 192.400 ;
        RECT 487.600 189.600 488.400 190.400 ;
        RECT 494.100 186.400 494.700 201.600 ;
        RECT 495.600 193.600 496.400 194.400 ;
        RECT 495.700 188.400 496.300 193.600 ;
        RECT 495.600 187.600 496.400 188.400 ;
        RECT 494.000 186.300 494.800 186.400 ;
        RECT 494.000 185.700 496.300 186.300 ;
        RECT 494.000 185.600 494.800 185.700 ;
        RECT 489.200 181.600 490.000 182.400 ;
        RECT 489.300 172.400 489.900 181.600 ;
        RECT 495.700 176.400 496.300 185.700 ;
        RECT 494.000 175.600 494.800 176.400 ;
        RECT 495.600 175.600 496.400 176.400 ;
        RECT 489.200 171.600 490.000 172.400 ;
        RECT 476.400 163.600 477.200 164.400 ;
        RECT 486.000 163.600 486.800 164.400 ;
        RECT 489.200 163.600 490.000 164.400 ;
        RECT 473.200 157.600 474.000 158.400 ;
        RECT 473.200 155.600 474.000 156.400 ;
        RECT 470.000 145.600 470.800 146.400 ;
        RECT 473.300 138.400 473.900 155.600 ;
        RECT 474.800 145.600 475.600 146.400 ;
        RECT 473.200 137.600 474.000 138.400 ;
        RECT 476.500 134.400 477.100 163.600 ;
        RECT 479.600 149.600 480.400 150.400 ;
        RECT 484.400 144.200 485.200 157.800 ;
        RECT 486.000 144.200 486.800 157.800 ;
        RECT 487.600 144.200 488.400 155.800 ;
        RECT 489.300 148.400 489.900 163.600 ;
        RECT 494.100 160.400 494.700 175.600 ;
        RECT 500.500 174.400 501.100 211.600 ;
        RECT 502.000 206.200 502.800 217.800 ;
        RECT 503.600 217.600 504.400 218.400 ;
        RECT 503.700 216.400 504.300 217.600 ;
        RECT 503.600 215.600 504.400 216.400 ;
        RECT 503.700 202.400 504.300 215.600 ;
        RECT 505.200 206.200 506.000 217.800 ;
        RECT 506.800 204.200 507.600 217.800 ;
        RECT 508.400 204.200 509.200 217.800 ;
        RECT 510.000 204.200 510.800 217.800 ;
        RECT 511.700 212.400 512.300 221.600 ;
        RECT 518.100 218.400 518.700 225.600 ;
        RECT 519.600 224.200 520.400 235.800 ;
        RECT 521.200 224.200 522.000 237.800 ;
        RECT 522.800 224.200 523.600 237.800 ;
        RECT 524.400 224.200 525.200 237.800 ;
        RECT 538.800 231.600 539.600 232.400 ;
        RECT 529.200 227.600 530.000 228.400 ;
        RECT 529.300 218.400 529.900 227.600 ;
        RECT 538.900 226.400 539.500 231.600 ;
        RECT 553.300 230.400 553.900 257.600 ;
        RECT 554.900 254.400 555.500 283.600 ;
        RECT 561.200 279.600 562.000 280.400 ;
        RECT 561.300 278.400 561.900 279.600 ;
        RECT 558.000 277.600 558.800 278.400 ;
        RECT 561.200 277.600 562.000 278.400 ;
        RECT 559.600 271.600 560.400 272.400 ;
        RECT 562.900 270.400 563.500 287.600 ;
        RECT 564.500 286.400 565.100 291.600 ;
        RECT 564.400 285.600 565.200 286.400 ;
        RECT 562.800 269.600 563.600 270.400 ;
        RECT 562.800 267.600 563.600 268.400 ;
        RECT 569.300 266.400 569.900 291.600 ;
        RECT 570.800 286.200 571.600 297.800 ;
        RECT 578.900 294.400 579.500 307.600 ;
        RECT 580.400 304.200 581.200 315.800 ;
        RECT 582.100 312.400 582.700 323.600 ;
        RECT 582.000 311.600 582.800 312.400 ;
        RECT 580.400 297.600 581.200 298.400 ;
        RECT 580.500 294.400 581.100 297.600 ;
        RECT 578.800 293.600 579.600 294.400 ;
        RECT 580.400 293.600 581.200 294.400 ;
        RECT 582.100 292.400 582.700 311.600 ;
        RECT 583.600 309.600 584.400 310.400 ;
        RECT 583.700 300.400 584.300 309.600 ;
        RECT 588.400 303.600 589.200 304.400 ;
        RECT 590.000 304.200 590.800 315.800 ;
        RECT 583.600 299.600 584.400 300.400 ;
        RECT 588.500 292.400 589.100 303.600 ;
        RECT 591.700 292.400 592.300 335.700 ;
        RECT 593.200 335.600 594.000 336.400 ;
        RECT 593.300 332.400 593.900 335.600 ;
        RECT 594.800 333.600 595.600 334.400 ;
        RECT 593.200 331.600 594.000 332.400 ;
        RECT 594.900 326.400 595.500 333.600 ;
        RECT 598.100 332.400 598.700 341.600 ;
        RECT 599.600 339.600 600.400 340.400 ;
        RECT 598.000 331.600 598.800 332.400 ;
        RECT 598.000 329.600 598.800 330.400 ;
        RECT 596.400 327.600 597.200 328.400 ;
        RECT 594.800 326.300 595.600 326.400 ;
        RECT 594.800 325.700 597.100 326.300 ;
        RECT 594.800 325.600 595.600 325.700 ;
        RECT 594.800 313.600 595.600 314.400 ;
        RECT 596.500 308.400 597.100 325.700 ;
        RECT 598.100 314.400 598.700 329.600 ;
        RECT 599.700 328.400 600.300 339.600 ;
        RECT 602.900 332.400 603.500 371.600 ;
        RECT 604.400 344.200 605.200 355.800 ;
        RECT 606.100 352.400 606.700 375.600 ;
        RECT 607.700 374.400 608.300 393.600 ;
        RECT 610.800 391.600 611.600 392.400 ;
        RECT 610.900 390.400 611.500 391.600 ;
        RECT 609.200 389.600 610.000 390.400 ;
        RECT 610.800 389.600 611.600 390.400 ;
        RECT 609.300 386.400 609.900 389.600 ;
        RECT 612.500 388.400 613.100 395.600 ;
        RECT 618.800 391.600 619.600 392.400 ;
        RECT 614.000 389.600 614.800 390.400 ;
        RECT 614.100 388.400 614.700 389.600 ;
        RECT 612.400 387.600 613.200 388.400 ;
        RECT 614.000 387.600 614.800 388.400 ;
        RECT 618.800 387.600 619.600 388.400 ;
        RECT 609.200 385.600 610.000 386.400 ;
        RECT 610.800 385.600 611.600 386.400 ;
        RECT 610.900 376.400 611.500 385.600 ;
        RECT 615.600 383.600 616.400 384.400 ;
        RECT 615.700 378.400 616.300 383.600 ;
        RECT 615.600 377.600 616.400 378.400 ;
        RECT 610.800 375.600 611.600 376.400 ;
        RECT 612.400 375.600 613.200 376.400 ;
        RECT 607.600 373.600 608.400 374.400 ;
        RECT 607.700 372.400 608.300 373.600 ;
        RECT 607.600 371.600 608.400 372.400 ;
        RECT 606.000 351.600 606.800 352.400 ;
        RECT 607.700 340.400 608.300 371.600 ;
        RECT 609.200 369.600 610.000 370.400 ;
        RECT 612.500 366.400 613.100 375.600 ;
        RECT 620.500 374.400 621.100 395.600 ;
        RECT 622.100 388.400 622.700 395.600 ;
        RECT 623.600 389.600 624.400 390.400 ;
        RECT 622.000 387.600 622.800 388.400 ;
        RECT 623.700 384.400 624.300 389.600 ;
        RECT 626.900 386.400 627.500 409.600 ;
        RECT 628.500 400.400 629.100 413.600 ;
        RECT 628.400 399.600 629.200 400.400 ;
        RECT 626.800 385.600 627.600 386.400 ;
        RECT 623.600 383.600 624.400 384.400 ;
        RECT 628.400 384.200 629.200 395.800 ;
        RECT 618.800 373.600 619.600 374.400 ;
        RECT 620.400 373.600 621.200 374.400 ;
        RECT 620.400 371.600 621.200 372.400 ;
        RECT 618.800 369.600 619.600 370.400 ;
        RECT 612.400 365.600 613.200 366.400 ;
        RECT 617.200 351.600 618.000 352.400 ;
        RECT 612.400 349.600 613.200 350.400 ;
        RECT 614.000 349.600 614.800 350.400 ;
        RECT 610.800 347.600 611.600 348.400 ;
        RECT 609.200 345.600 610.000 346.400 ;
        RECT 609.300 344.400 609.900 345.600 ;
        RECT 612.500 344.400 613.100 349.600 ;
        RECT 617.300 346.400 617.900 351.600 ;
        RECT 617.200 345.600 618.000 346.400 ;
        RECT 609.200 343.600 610.000 344.400 ;
        RECT 612.400 343.600 613.200 344.400 ;
        RECT 607.600 339.600 608.400 340.400 ;
        RECT 609.200 337.600 610.000 338.400 ;
        RECT 607.600 333.600 608.400 334.400 ;
        RECT 614.000 333.600 614.800 334.400 ;
        RECT 602.800 331.600 603.600 332.400 ;
        RECT 599.600 327.600 600.400 328.400 ;
        RECT 598.000 313.600 598.800 314.400 ;
        RECT 601.200 313.600 602.000 314.400 ;
        RECT 601.300 312.400 601.900 313.600 ;
        RECT 601.200 311.600 602.000 312.400 ;
        RECT 601.300 310.400 601.900 311.600 ;
        RECT 598.000 309.600 598.800 310.400 ;
        RECT 601.200 309.600 602.000 310.400 ;
        RECT 602.900 308.400 603.500 331.600 ;
        RECT 607.700 326.400 608.300 333.600 ;
        RECT 614.000 331.600 614.800 332.400 ;
        RECT 615.600 331.600 616.400 332.400 ;
        RECT 609.200 329.600 610.000 330.400 ;
        RECT 607.600 325.600 608.400 326.400 ;
        RECT 606.000 309.600 606.800 310.400 ;
        RECT 606.100 308.400 606.700 309.600 ;
        RECT 607.700 308.400 608.300 325.600 ;
        RECT 609.200 319.600 610.000 320.400 ;
        RECT 609.300 310.400 609.900 319.600 ;
        RECT 609.200 309.600 610.000 310.400 ;
        RECT 610.800 309.600 611.600 310.400 ;
        RECT 596.400 307.600 597.200 308.400 ;
        RECT 598.000 307.600 598.800 308.400 ;
        RECT 599.600 307.600 600.400 308.400 ;
        RECT 602.800 307.600 603.600 308.400 ;
        RECT 606.000 307.600 606.800 308.400 ;
        RECT 607.600 307.600 608.400 308.400 ;
        RECT 612.400 307.600 613.200 308.400 ;
        RECT 596.500 302.400 597.100 307.600 ;
        RECT 598.100 304.400 598.700 307.600 ;
        RECT 598.000 303.600 598.800 304.400 ;
        RECT 596.400 301.600 597.200 302.400 ;
        RECT 593.200 293.600 594.000 294.400 ;
        RECT 593.300 292.400 593.900 293.600 ;
        RECT 598.100 292.400 598.700 303.600 ;
        RECT 582.000 291.600 582.800 292.400 ;
        RECT 583.600 291.600 584.400 292.400 ;
        RECT 588.400 291.600 589.200 292.400 ;
        RECT 591.600 291.600 592.400 292.400 ;
        RECT 593.200 291.600 594.000 292.400 ;
        RECT 598.000 291.600 598.800 292.400 ;
        RECT 583.700 290.400 584.300 291.600 ;
        RECT 583.600 289.600 584.400 290.400 ;
        RECT 586.800 287.600 587.600 288.400 ;
        RECT 586.800 279.600 587.600 280.400 ;
        RECT 572.400 277.600 573.200 278.400 ;
        RECT 572.500 270.400 573.100 277.600 ;
        RECT 583.600 275.600 584.400 276.400 ;
        RECT 586.900 270.400 587.500 279.600 ;
        RECT 588.500 272.400 589.100 291.600 ;
        RECT 591.700 280.400 592.300 291.600 ;
        RECT 598.000 287.600 598.800 288.400 ;
        RECT 596.400 283.600 597.200 284.400 ;
        RECT 591.600 279.600 592.400 280.400 ;
        RECT 588.400 271.600 589.200 272.400 ;
        RECT 591.600 272.300 592.400 272.400 ;
        RECT 594.800 272.300 595.600 272.400 ;
        RECT 591.600 271.700 595.600 272.300 ;
        RECT 591.600 271.600 592.400 271.700 ;
        RECT 594.800 271.600 595.600 271.700 ;
        RECT 570.800 269.600 571.600 270.400 ;
        RECT 572.400 269.600 573.200 270.400 ;
        RECT 580.400 269.600 581.200 270.400 ;
        RECT 585.200 269.600 586.000 270.400 ;
        RECT 586.800 269.600 587.600 270.400 ;
        RECT 559.600 265.600 560.400 266.400 ;
        RECT 569.200 265.600 570.000 266.400 ;
        RECT 559.700 256.400 560.300 265.600 ;
        RECT 567.600 263.600 568.400 264.400 ;
        RECT 566.000 259.600 566.800 260.400 ;
        RECT 559.600 255.600 560.400 256.400 ;
        RECT 554.800 253.600 555.600 254.400 ;
        RECT 558.000 251.600 558.800 252.400 ;
        RECT 561.200 246.200 562.000 257.800 ;
        RECT 564.400 250.200 565.200 255.800 ;
        RECT 566.100 254.400 566.700 259.600 ;
        RECT 566.000 253.600 566.800 254.400 ;
        RECT 567.700 252.400 568.300 263.600 ;
        RECT 569.300 256.400 569.900 265.600 ;
        RECT 570.900 264.400 571.500 269.600 ;
        RECT 585.300 268.400 585.900 269.600 ;
        RECT 585.200 267.600 586.000 268.400 ;
        RECT 570.800 263.600 571.600 264.400 ;
        RECT 578.800 263.600 579.600 264.400 ;
        RECT 569.200 255.600 570.000 256.400 ;
        RECT 575.600 253.600 576.400 254.400 ;
        RECT 575.700 252.400 576.300 253.600 ;
        RECT 567.600 251.600 568.400 252.400 ;
        RECT 575.600 251.600 576.400 252.400 ;
        RECT 577.200 250.300 578.000 250.400 ;
        RECT 578.900 250.300 579.500 263.600 ;
        RECT 580.400 259.600 581.200 260.400 ;
        RECT 580.500 252.400 581.100 259.600 ;
        RECT 588.500 258.400 589.100 271.600 ;
        RECT 593.200 269.600 594.000 270.400 ;
        RECT 594.800 270.300 595.600 270.400 ;
        RECT 596.500 270.300 597.100 283.600 ;
        RECT 598.100 270.400 598.700 287.600 ;
        RECT 599.700 282.400 600.300 307.600 ;
        RECT 607.700 306.400 608.300 307.600 ;
        RECT 612.500 306.400 613.100 307.600 ;
        RECT 601.200 305.600 602.000 306.400 ;
        RECT 607.600 305.600 608.400 306.400 ;
        RECT 612.400 305.600 613.200 306.400 ;
        RECT 601.300 294.400 601.900 305.600 ;
        RECT 602.800 303.600 603.600 304.400 ;
        RECT 602.900 300.400 603.500 303.600 ;
        RECT 607.600 301.600 608.400 302.400 ;
        RECT 602.800 299.600 603.600 300.400 ;
        RECT 604.400 297.600 605.200 298.400 ;
        RECT 601.200 293.600 602.000 294.400 ;
        RECT 602.800 285.600 603.600 286.400 ;
        RECT 599.600 281.600 600.400 282.400 ;
        RECT 599.700 270.400 600.300 281.600 ;
        RECT 604.500 274.400 605.100 297.600 ;
        RECT 607.700 294.400 608.300 301.600 ;
        RECT 612.400 299.600 613.200 300.400 ;
        RECT 612.500 294.400 613.100 299.600 ;
        RECT 614.100 298.400 614.700 331.600 ;
        RECT 615.700 322.400 616.300 331.600 ;
        RECT 618.900 324.400 619.500 369.600 ;
        RECT 620.500 352.400 621.100 371.600 ;
        RECT 623.700 370.300 624.300 383.600 ;
        RECT 626.800 371.600 627.600 372.400 ;
        RECT 628.400 371.600 629.200 372.400 ;
        RECT 625.200 370.300 626.000 370.400 ;
        RECT 623.700 369.700 626.000 370.300 ;
        RECT 625.200 369.600 626.000 369.700 ;
        RECT 622.000 367.600 622.800 368.400 ;
        RECT 626.900 364.400 627.500 371.600 ;
        RECT 628.500 370.400 629.100 371.600 ;
        RECT 628.400 369.600 629.200 370.400 ;
        RECT 626.800 363.600 627.600 364.400 ;
        RECT 626.900 354.400 627.500 363.600 ;
        RECT 623.600 353.600 624.400 354.400 ;
        RECT 626.800 353.600 627.600 354.400 ;
        RECT 620.400 351.600 621.200 352.400 ;
        RECT 620.500 350.400 621.100 351.600 ;
        RECT 623.700 350.400 624.300 353.600 ;
        RECT 620.400 349.600 621.200 350.400 ;
        RECT 623.600 349.600 624.400 350.400 ;
        RECT 625.200 349.600 626.000 350.400 ;
        RECT 620.500 336.400 621.100 349.600 ;
        RECT 622.000 347.600 622.800 348.400 ;
        RECT 625.300 346.400 625.900 349.600 ;
        RECT 625.200 345.600 626.000 346.400 ;
        RECT 626.800 343.600 627.600 344.400 ;
        RECT 620.400 335.600 621.200 336.400 ;
        RECT 622.000 335.600 622.800 336.400 ;
        RECT 620.500 334.400 621.100 335.600 ;
        RECT 622.100 334.400 622.700 335.600 ;
        RECT 620.400 333.600 621.200 334.400 ;
        RECT 622.000 333.600 622.800 334.400 ;
        RECT 625.200 333.600 626.000 334.400 ;
        RECT 626.800 333.600 627.600 334.400 ;
        RECT 623.600 331.600 624.400 332.400 ;
        RECT 618.800 323.600 619.600 324.400 ;
        RECT 615.600 321.600 616.400 322.400 ;
        RECT 618.800 321.600 619.600 322.400 ;
        RECT 618.900 310.400 619.500 321.600 ;
        RECT 623.700 316.400 624.300 331.600 ;
        RECT 623.600 315.600 624.400 316.400 ;
        RECT 626.900 312.400 627.500 333.600 ;
        RECT 630.100 330.300 630.700 429.600 ;
        RECT 631.700 428.400 632.300 429.600 ;
        RECT 631.600 427.600 632.400 428.400 ;
        RECT 633.300 424.400 633.900 449.600 ;
        RECT 633.200 423.600 634.000 424.400 ;
        RECT 631.600 413.600 632.400 414.400 ;
        RECT 633.200 412.300 634.000 412.400 ;
        RECT 634.900 412.300 635.500 463.600 ;
        RECT 636.500 458.400 637.100 465.600 ;
        RECT 636.400 457.600 637.200 458.400 ;
        RECT 636.400 447.600 637.200 448.400 ;
        RECT 636.500 438.400 637.100 447.600 ;
        RECT 636.400 437.600 637.200 438.400 ;
        RECT 638.100 434.400 638.700 493.700 ;
        RECT 660.400 491.600 661.200 492.400 ;
        RECT 647.600 483.600 648.400 484.400 ;
        RECT 652.400 483.600 653.200 484.400 ;
        RECT 647.700 474.400 648.300 483.600 ;
        RECT 660.500 482.300 661.100 491.600 ;
        RECT 662.000 484.200 662.800 497.800 ;
        RECT 663.600 484.200 664.400 497.800 ;
        RECT 665.200 484.200 666.000 497.800 ;
        RECT 666.800 486.200 667.600 497.800 ;
        RECT 668.400 495.600 669.200 496.400 ;
        RECT 660.500 481.700 662.700 482.300 ;
        RECT 647.600 473.600 648.400 474.400 ;
        RECT 652.400 471.600 653.200 472.400 ;
        RECT 639.600 469.600 640.400 470.400 ;
        RECT 642.800 469.600 643.600 470.400 ;
        RECT 644.400 469.600 645.200 470.400 ;
        RECT 649.200 469.600 650.000 470.400 ;
        RECT 655.600 469.600 656.400 470.400 ;
        RECT 639.700 466.400 640.300 469.600 ;
        RECT 641.200 467.600 642.000 468.400 ;
        RECT 641.300 466.400 641.900 467.600 ;
        RECT 639.600 465.600 640.400 466.400 ;
        RECT 641.200 465.600 642.000 466.400 ;
        RECT 642.900 464.400 643.500 469.600 ;
        RECT 644.500 468.400 645.100 469.600 ;
        RECT 644.400 467.600 645.200 468.400 ;
        RECT 649.300 466.400 649.900 469.600 ;
        RECT 657.200 467.600 658.000 468.400 ;
        RECT 649.200 465.600 650.000 466.400 ;
        RECT 642.800 463.600 643.600 464.400 ;
        RECT 647.600 463.600 648.400 464.400 ;
        RECT 652.400 463.600 653.200 464.400 ;
        RECT 658.800 463.600 659.600 464.400 ;
        RECT 647.700 460.400 648.300 463.600 ;
        RECT 647.600 459.600 648.400 460.400 ;
        RECT 652.500 458.400 653.100 463.600 ;
        RECT 655.600 459.600 656.400 460.400 ;
        RECT 644.400 457.600 645.200 458.400 ;
        RECT 641.200 453.600 642.000 454.400 ;
        RECT 638.000 433.600 638.800 434.400 ;
        RECT 639.400 415.000 640.200 415.800 ;
        RECT 641.300 415.600 641.900 453.600 ;
        RECT 644.500 452.400 645.100 457.600 ;
        RECT 644.400 451.600 645.200 452.400 ;
        RECT 646.000 444.200 646.800 457.800 ;
        RECT 647.600 444.200 648.400 457.800 ;
        RECT 649.200 444.200 650.000 457.800 ;
        RECT 650.800 446.200 651.600 457.800 ;
        RECT 652.400 457.600 653.200 458.400 ;
        RECT 652.400 455.600 653.200 456.400 ;
        RECT 652.500 448.400 653.100 455.600 ;
        RECT 652.400 447.600 653.200 448.400 ;
        RECT 654.000 446.200 654.800 457.800 ;
        RECT 655.700 454.400 656.300 459.600 ;
        RECT 655.600 453.600 656.400 454.400 ;
        RECT 657.200 446.200 658.000 457.800 ;
        RECT 658.800 444.200 659.600 457.800 ;
        RECT 660.400 444.200 661.200 457.800 ;
        RECT 662.100 452.400 662.700 481.700 ;
        RECT 663.600 464.200 664.400 475.800 ;
        RECT 666.800 473.600 667.600 474.400 ;
        RECT 662.000 451.600 662.800 452.400 ;
        RECT 649.200 441.600 650.000 442.400 ;
        RECT 647.600 433.600 648.400 434.400 ;
        RECT 647.700 428.400 648.300 433.600 ;
        RECT 647.600 427.600 648.400 428.400 ;
        RECT 647.600 423.600 648.400 424.400 ;
        RECT 644.400 421.600 645.200 422.400 ;
        RECT 644.500 418.400 645.100 421.600 ;
        RECT 644.400 417.600 645.200 418.400 ;
        RECT 641.200 415.000 645.400 415.600 ;
        RECT 646.000 415.000 646.800 415.800 ;
        RECT 638.000 413.600 638.800 414.400 ;
        RECT 633.200 411.700 635.500 412.300 ;
        RECT 633.200 411.600 634.000 411.700 ;
        RECT 633.200 403.600 634.000 404.400 ;
        RECT 633.300 374.300 633.900 403.600 ;
        RECT 634.900 378.400 635.500 411.700 ;
        RECT 636.400 409.600 637.200 410.400 ;
        RECT 638.100 402.400 638.700 413.600 ;
        RECT 639.400 410.200 640.000 415.000 ;
        RECT 641.200 414.800 642.000 415.000 ;
        RECT 644.600 414.800 645.400 415.000 ;
        RECT 646.200 414.200 646.800 415.000 ;
        RECT 647.700 414.400 648.300 423.600 ;
        RECT 642.000 413.600 646.800 414.200 ;
        RECT 647.600 413.600 648.400 414.400 ;
        RECT 642.000 413.400 642.800 413.600 ;
        RECT 646.200 410.200 646.800 413.600 ;
        RECT 639.400 409.400 640.200 410.200 ;
        RECT 646.000 409.400 646.800 410.200 ;
        RECT 647.700 408.400 648.300 413.600 ;
        RECT 647.600 407.600 648.400 408.400 ;
        RECT 638.000 401.600 638.800 402.400 ;
        RECT 636.400 389.400 637.200 390.200 ;
        RECT 636.500 378.400 637.100 389.400 ;
        RECT 638.000 384.200 638.800 395.800 ;
        RECT 642.800 392.300 643.600 392.400 ;
        RECT 639.600 387.600 640.400 388.400 ;
        RECT 639.700 380.400 640.300 387.600 ;
        RECT 641.200 386.200 642.000 391.800 ;
        RECT 642.800 391.700 645.100 392.300 ;
        RECT 642.800 391.600 643.600 391.700 ;
        RECT 642.800 383.600 643.600 384.400 ;
        RECT 639.600 379.600 640.400 380.400 ;
        RECT 642.900 378.400 643.500 383.600 ;
        RECT 634.800 377.600 635.600 378.400 ;
        RECT 636.400 377.600 637.200 378.400 ;
        RECT 638.000 377.600 638.800 378.400 ;
        RECT 642.800 377.600 643.600 378.400 ;
        RECT 631.700 373.700 633.900 374.300 ;
        RECT 631.700 356.400 632.300 373.700 ;
        RECT 634.800 373.600 635.600 374.400 ;
        RECT 634.900 372.400 635.500 373.600 ;
        RECT 633.200 371.600 634.000 372.400 ;
        RECT 634.800 371.600 635.600 372.400 ;
        RECT 633.300 358.400 633.900 371.600 ;
        RECT 636.400 369.600 637.200 370.400 ;
        RECT 636.500 368.400 637.100 369.600 ;
        RECT 636.400 367.600 637.200 368.400 ;
        RECT 633.200 357.600 634.000 358.400 ;
        RECT 631.600 355.600 632.400 356.400 ;
        RECT 633.300 350.400 633.900 357.600 ;
        RECT 638.100 354.400 638.700 377.600 ;
        RECT 641.200 375.600 642.000 376.400 ;
        RECT 641.300 374.400 641.900 375.600 ;
        RECT 641.200 373.600 642.000 374.400 ;
        RECT 642.800 373.600 643.600 374.400 ;
        RECT 639.600 371.600 640.400 372.400 ;
        RECT 644.500 370.400 645.100 391.700 ;
        RECT 646.000 389.600 646.800 390.400 ;
        RECT 647.600 387.600 648.400 388.400 ;
        RECT 647.700 386.400 648.300 387.600 ;
        RECT 647.600 385.600 648.400 386.400 ;
        RECT 647.600 375.600 648.400 376.400 ;
        RECT 647.700 374.400 648.300 375.600 ;
        RECT 647.600 373.600 648.400 374.400 ;
        RECT 639.600 369.600 640.400 370.400 ;
        RECT 644.400 369.600 645.200 370.400 ;
        RECT 646.000 369.600 646.800 370.400 ;
        RECT 636.400 353.600 637.200 354.400 ;
        RECT 638.000 353.600 638.800 354.400 ;
        RECT 634.800 351.600 635.600 352.400 ;
        RECT 634.900 350.400 635.500 351.600 ;
        RECT 633.200 349.600 634.000 350.400 ;
        RECT 634.800 349.600 635.600 350.400 ;
        RECT 633.200 347.600 634.000 348.400 ;
        RECT 633.200 345.600 634.000 346.400 ;
        RECT 631.600 341.600 632.400 342.400 ;
        RECT 631.700 332.400 632.300 341.600 ;
        RECT 633.300 332.400 633.900 345.600 ;
        RECT 634.900 340.400 635.500 349.600 ;
        RECT 636.500 342.300 637.100 353.600 ;
        RECT 638.000 351.600 638.800 352.400 ;
        RECT 638.100 344.300 638.700 351.600 ;
        RECT 639.700 346.300 640.300 369.600 ;
        RECT 644.400 363.600 645.200 364.400 ;
        RECT 642.800 349.600 643.600 350.400 ;
        RECT 641.200 347.600 642.000 348.400 ;
        RECT 639.700 345.700 641.900 346.300 ;
        RECT 638.100 343.700 640.300 344.300 ;
        RECT 638.000 342.300 638.800 342.400 ;
        RECT 636.500 341.700 638.800 342.300 ;
        RECT 638.000 341.600 638.800 341.700 ;
        RECT 634.800 339.600 635.600 340.400 ;
        RECT 636.400 337.600 637.200 338.400 ;
        RECT 636.500 336.400 637.100 337.600 ;
        RECT 634.800 335.600 635.600 336.400 ;
        RECT 636.400 335.600 637.200 336.400 ;
        RECT 638.100 332.400 638.700 341.600 ;
        RECT 639.700 332.400 640.300 343.700 ;
        RECT 631.600 331.600 632.400 332.400 ;
        RECT 633.200 331.600 634.000 332.400 ;
        RECT 636.400 331.600 637.200 332.400 ;
        RECT 638.000 331.600 638.800 332.400 ;
        RECT 639.600 331.600 640.400 332.400 ;
        RECT 630.100 329.700 632.300 330.300 ;
        RECT 631.700 328.400 632.300 329.700 ;
        RECT 633.200 329.600 634.000 330.400 ;
        RECT 630.000 327.600 630.800 328.400 ;
        RECT 631.600 327.600 632.400 328.400 ;
        RECT 628.400 323.600 629.200 324.400 ;
        RECT 628.500 312.400 629.100 323.600 ;
        RECT 636.500 318.400 637.100 331.600 ;
        RECT 638.100 320.400 638.700 331.600 ;
        RECT 639.700 330.400 640.300 331.600 ;
        RECT 639.600 329.600 640.400 330.400 ;
        RECT 639.600 327.600 640.400 328.400 ;
        RECT 638.000 319.600 638.800 320.400 ;
        RECT 633.200 317.600 634.000 318.400 ;
        RECT 636.400 317.600 637.200 318.400 ;
        RECT 638.000 315.600 638.800 316.400 ;
        RECT 626.800 311.600 627.600 312.400 ;
        RECT 628.400 311.600 629.200 312.400 ;
        RECT 615.600 309.600 616.400 310.400 ;
        RECT 618.800 309.600 619.600 310.400 ;
        RECT 623.600 309.600 624.400 310.400 ;
        RECT 614.000 297.600 614.800 298.400 ;
        RECT 607.600 293.600 608.400 294.400 ;
        RECT 610.800 293.600 611.600 294.400 ;
        RECT 612.400 293.600 613.200 294.400 ;
        RECT 607.700 290.400 608.300 293.600 ;
        RECT 610.900 292.400 611.500 293.600 ;
        RECT 610.800 291.600 611.600 292.400 ;
        RECT 615.700 290.400 616.300 309.600 ;
        RECT 622.000 303.600 622.800 304.400 ;
        RECT 620.400 295.600 621.200 296.400 ;
        RECT 622.100 294.400 622.700 303.600 ;
        RECT 618.800 293.600 619.600 294.400 ;
        RECT 622.000 293.600 622.800 294.400 ;
        RECT 617.200 291.600 618.000 292.400 ;
        RECT 607.600 289.600 608.400 290.400 ;
        RECT 614.000 289.600 614.800 290.400 ;
        RECT 615.600 289.600 616.400 290.400 ;
        RECT 614.100 286.400 614.700 289.600 ;
        RECT 618.900 288.300 619.500 293.600 ;
        RECT 623.700 292.400 624.300 309.600 ;
        RECT 625.200 307.600 626.000 308.400 ;
        RECT 625.300 302.400 625.900 307.600 ;
        RECT 625.200 301.600 626.000 302.400 ;
        RECT 625.200 295.600 626.000 296.400 ;
        RECT 625.300 294.400 625.900 295.600 ;
        RECT 625.200 293.600 626.000 294.400 ;
        RECT 623.600 291.600 624.400 292.400 ;
        RECT 625.200 291.600 626.000 292.400 ;
        RECT 625.300 290.400 625.900 291.600 ;
        RECT 620.400 289.600 621.200 290.400 ;
        RECT 625.200 289.600 626.000 290.400 ;
        RECT 626.800 290.300 627.600 290.400 ;
        RECT 628.500 290.300 629.100 311.600 ;
        RECT 633.200 309.600 634.000 310.400 ;
        RECT 634.800 309.600 635.600 310.400 ;
        RECT 634.900 308.400 635.500 309.600 ;
        RECT 634.800 307.600 635.600 308.400 ;
        RECT 634.800 297.600 635.600 298.400 ;
        RECT 631.600 295.600 632.400 296.400 ;
        RECT 633.200 295.600 634.000 296.400 ;
        RECT 630.000 293.600 630.800 294.400 ;
        RECT 626.800 289.700 629.100 290.300 ;
        RECT 626.800 289.600 627.600 289.700 ;
        RECT 618.900 287.700 621.100 288.300 ;
        RECT 614.000 285.600 614.800 286.400 ;
        RECT 609.200 283.600 610.000 284.400 ;
        RECT 604.400 273.600 605.200 274.400 ;
        RECT 609.300 270.400 609.900 283.600 ;
        RECT 620.500 278.400 621.100 287.700 ;
        RECT 625.200 285.600 626.000 286.400 ;
        RECT 625.300 278.400 625.900 285.600 ;
        RECT 620.400 277.600 621.200 278.400 ;
        RECT 625.200 277.600 626.000 278.400 ;
        RECT 617.200 275.600 618.000 276.400 ;
        RECT 612.400 271.600 613.200 272.400 ;
        RECT 594.800 269.700 597.100 270.300 ;
        RECT 594.800 269.600 595.600 269.700 ;
        RECT 593.300 268.400 593.900 269.600 ;
        RECT 593.200 267.600 594.000 268.400 ;
        RECT 582.000 253.600 582.800 254.400 ;
        RECT 580.400 251.600 581.200 252.400 ;
        RECT 577.200 249.700 579.500 250.300 ;
        RECT 583.600 250.200 584.400 255.800 ;
        RECT 577.200 249.600 578.000 249.700 ;
        RECT 586.800 246.200 587.600 257.800 ;
        RECT 588.400 257.600 589.200 258.400 ;
        RECT 588.400 255.600 589.200 256.400 ;
        RECT 593.300 254.400 593.900 267.600 ;
        RECT 594.800 263.600 595.600 264.400 ;
        RECT 593.200 253.600 594.000 254.400 ;
        RECT 588.400 251.600 589.200 252.600 ;
        RECT 594.900 252.400 595.500 263.600 ;
        RECT 596.500 260.400 597.100 269.700 ;
        RECT 598.000 269.600 598.800 270.400 ;
        RECT 599.600 269.600 600.400 270.400 ;
        RECT 607.600 269.600 608.400 270.400 ;
        RECT 609.200 269.600 610.000 270.400 ;
        RECT 607.700 268.400 608.300 269.600 ;
        RECT 599.600 267.600 600.400 268.400 ;
        RECT 604.400 267.600 605.200 268.400 ;
        RECT 607.600 267.600 608.400 268.400 ;
        RECT 612.500 266.400 613.100 271.600 ;
        RECT 617.300 270.400 617.900 275.600 ;
        RECT 626.900 272.400 627.500 289.600 ;
        RECT 628.400 283.600 629.200 284.400 ;
        RECT 628.500 278.400 629.100 283.600 ;
        RECT 628.400 277.600 629.200 278.400 ;
        RECT 623.600 271.600 624.400 272.400 ;
        RECT 626.800 271.600 627.600 272.400 ;
        RECT 628.500 270.400 629.100 277.600 ;
        RECT 630.100 276.400 630.700 293.600 ;
        RECT 634.900 292.400 635.500 297.600 ;
        RECT 636.400 295.600 637.200 296.400 ;
        RECT 636.500 292.400 637.100 295.600 ;
        RECT 634.800 291.600 635.600 292.400 ;
        RECT 636.400 291.600 637.200 292.400 ;
        RECT 634.900 284.400 635.500 291.600 ;
        RECT 634.800 283.600 635.600 284.400 ;
        RECT 630.000 275.600 630.800 276.400 ;
        RECT 638.100 274.400 638.700 315.600 ;
        RECT 639.700 308.400 640.300 327.600 ;
        RECT 641.300 324.400 641.900 345.700 ;
        RECT 642.900 338.400 643.500 349.600 ;
        RECT 642.800 337.600 643.600 338.400 ;
        RECT 642.800 335.600 643.600 336.400 ;
        RECT 641.200 323.600 642.000 324.400 ;
        RECT 642.900 318.400 643.500 335.600 ;
        RECT 644.500 334.400 645.100 363.600 ;
        RECT 646.100 352.400 646.700 369.600 ;
        RECT 647.700 362.400 648.300 373.600 ;
        RECT 649.300 368.400 649.900 441.600 ;
        RECT 655.600 433.600 656.400 434.400 ;
        RECT 650.800 423.600 651.600 424.400 ;
        RECT 650.800 409.600 651.600 410.400 ;
        RECT 650.800 407.600 651.600 408.400 ;
        RECT 650.900 372.400 651.500 407.600 ;
        RECT 654.000 393.600 654.800 394.400 ;
        RECT 654.100 390.400 654.700 393.600 ;
        RECT 654.000 389.600 654.800 390.400 ;
        RECT 650.800 371.600 651.600 372.400 ;
        RECT 650.900 368.400 651.500 371.600 ;
        RECT 649.200 367.600 650.000 368.400 ;
        RECT 650.800 367.600 651.600 368.400 ;
        RECT 650.800 363.600 651.600 364.400 ;
        RECT 654.000 363.600 654.800 364.400 ;
        RECT 647.600 361.600 648.400 362.400 ;
        RECT 649.200 361.600 650.000 362.400 ;
        RECT 646.000 351.600 646.800 352.400 ;
        RECT 646.100 350.400 646.700 351.600 ;
        RECT 646.000 349.600 646.800 350.400 ;
        RECT 647.600 349.600 648.400 350.400 ;
        RECT 646.000 347.600 646.800 348.400 ;
        RECT 644.400 333.600 645.200 334.400 ;
        RECT 644.400 331.600 645.200 332.400 ;
        RECT 642.800 317.600 643.600 318.400 ;
        RECT 644.500 316.400 645.100 331.600 ;
        RECT 646.100 326.400 646.700 347.600 ;
        RECT 649.300 346.400 649.900 361.600 ;
        RECT 650.900 360.400 651.500 363.600 ;
        RECT 654.100 362.400 654.700 363.600 ;
        RECT 654.000 361.600 654.800 362.400 ;
        RECT 650.800 359.600 651.600 360.400 ;
        RECT 655.700 358.400 656.300 433.600 ;
        RECT 658.800 429.600 659.600 430.400 ;
        RECT 658.900 428.400 659.500 429.600 ;
        RECT 658.800 427.600 659.600 428.400 ;
        RECT 658.900 412.400 659.500 427.600 ;
        RECT 660.400 424.200 661.200 437.800 ;
        RECT 662.000 424.200 662.800 437.800 ;
        RECT 663.600 424.200 664.400 437.800 ;
        RECT 665.200 424.200 666.000 435.800 ;
        RECT 666.900 426.400 667.500 473.600 ;
        RECT 668.500 448.400 669.100 495.600 ;
        RECT 670.000 486.200 670.800 497.800 ;
        RECT 671.600 497.600 672.400 498.400 ;
        RECT 671.700 494.400 672.300 497.600 ;
        RECT 671.600 493.600 672.400 494.400 ;
        RECT 673.200 486.200 674.000 497.800 ;
        RECT 674.800 484.200 675.600 497.800 ;
        RECT 676.400 484.200 677.200 497.800 ;
        RECT 670.000 469.600 670.800 470.400 ;
        RECT 673.200 464.200 674.000 475.800 ;
        RECT 674.800 467.600 675.600 468.400 ;
        RECT 676.400 466.200 677.200 471.800 ;
        RECT 678.000 469.600 678.800 470.400 ;
        RECT 670.000 453.600 670.800 454.400 ;
        RECT 670.100 450.400 670.700 453.600 ;
        RECT 670.000 449.600 670.800 450.400 ;
        RECT 668.400 447.600 669.200 448.400 ;
        RECT 666.800 425.600 667.600 426.400 ;
        RECT 658.800 411.600 659.600 412.400 ;
        RECT 660.400 404.200 661.200 417.800 ;
        RECT 662.000 404.200 662.800 417.800 ;
        RECT 663.600 404.200 664.400 417.800 ;
        RECT 665.200 406.200 666.000 417.800 ;
        RECT 666.900 416.400 667.500 425.600 ;
        RECT 668.400 424.200 669.200 435.800 ;
        RECT 670.000 427.600 670.800 428.400 ;
        RECT 670.100 422.400 670.700 427.600 ;
        RECT 671.600 424.200 672.400 435.800 ;
        RECT 673.200 424.200 674.000 437.800 ;
        RECT 674.800 424.200 675.600 437.800 ;
        RECT 670.000 421.600 670.800 422.400 ;
        RECT 666.800 415.600 667.600 416.400 ;
        RECT 666.900 398.300 667.500 415.600 ;
        RECT 668.400 406.200 669.200 417.800 ;
        RECT 670.000 413.600 670.800 414.400 ;
        RECT 671.600 406.200 672.400 417.800 ;
        RECT 673.200 404.200 674.000 417.800 ;
        RECT 674.800 404.200 675.600 417.800 ;
        RECT 678.100 398.400 678.700 469.600 ;
        RECT 681.200 467.600 682.000 468.400 ;
        RECT 681.300 458.400 681.900 467.600 ;
        RECT 681.200 457.600 682.000 458.400 ;
        RECT 681.200 443.600 682.000 444.400 ;
        RECT 679.600 411.600 680.400 412.400 ;
        RECT 657.200 384.200 658.000 397.800 ;
        RECT 658.800 384.200 659.600 397.800 ;
        RECT 665.300 397.700 667.500 398.300 ;
        RECT 660.400 384.200 661.200 395.800 ;
        RECT 662.000 387.600 662.800 388.400 ;
        RECT 663.600 384.200 664.400 395.800 ;
        RECT 665.300 386.400 665.900 397.700 ;
        RECT 665.200 385.600 666.000 386.400 ;
        RECT 666.800 384.200 667.600 395.800 ;
        RECT 668.400 384.200 669.200 397.800 ;
        RECT 670.000 384.200 670.800 397.800 ;
        RECT 671.600 384.200 672.400 397.800 ;
        RECT 678.000 397.600 678.800 398.400 ;
        RECT 678.100 392.400 678.700 397.600 ;
        RECT 678.000 391.600 678.800 392.400 ;
        RECT 670.000 379.600 670.800 380.400 ;
        RECT 658.800 373.600 659.600 374.400 ;
        RECT 655.600 357.600 656.400 358.400 ;
        RECT 647.600 345.600 648.400 346.400 ;
        RECT 649.200 345.600 650.000 346.400 ;
        RECT 647.700 334.400 648.300 345.600 ;
        RECT 650.800 343.600 651.600 344.400 ;
        RECT 655.600 344.200 656.400 355.800 ;
        RECT 649.200 339.600 650.000 340.400 ;
        RECT 647.600 333.600 648.400 334.400 ;
        RECT 646.000 325.600 646.800 326.400 ;
        RECT 644.400 315.600 645.200 316.400 ;
        RECT 644.400 311.600 645.200 312.400 ;
        RECT 642.800 309.600 643.600 310.400 ;
        RECT 639.600 307.600 640.400 308.400 ;
        RECT 641.200 307.600 642.000 308.400 ;
        RECT 641.300 306.400 641.900 307.600 ;
        RECT 644.500 306.400 645.100 311.600 ;
        RECT 646.000 309.600 646.800 310.400 ;
        RECT 639.600 305.600 640.400 306.400 ;
        RECT 641.200 305.600 642.000 306.400 ;
        RECT 644.400 305.600 645.200 306.400 ;
        RECT 639.700 298.400 640.300 305.600 ;
        RECT 646.100 304.400 646.700 309.600 ;
        RECT 646.000 303.600 646.800 304.400 ;
        RECT 647.700 300.400 648.300 333.600 ;
        RECT 649.300 332.400 649.900 339.600 ;
        RECT 649.200 331.600 650.000 332.400 ;
        RECT 650.900 330.400 651.500 343.600 ;
        RECT 652.400 337.600 653.200 338.400 ;
        RECT 652.500 330.400 653.100 337.600 ;
        RECT 654.000 333.600 654.800 334.400 ;
        RECT 654.100 332.400 654.700 333.600 ;
        RECT 654.000 331.600 654.800 332.400 ;
        RECT 655.600 331.600 656.400 332.400 ;
        RECT 657.200 331.600 658.000 332.400 ;
        RECT 650.800 329.600 651.600 330.400 ;
        RECT 652.400 329.600 653.200 330.400 ;
        RECT 657.300 328.400 657.900 331.600 ;
        RECT 649.200 327.600 650.000 328.400 ;
        RECT 657.200 327.600 658.000 328.400 ;
        RECT 649.200 323.600 650.000 324.400 ;
        RECT 647.600 299.600 648.400 300.400 ;
        RECT 649.300 298.400 649.900 323.600 ;
        RECT 655.600 313.600 656.400 314.400 ;
        RECT 652.400 311.600 653.200 312.400 ;
        RECT 652.500 310.400 653.100 311.600 ;
        RECT 652.400 309.600 653.200 310.400 ;
        RECT 654.000 310.300 654.800 310.400 ;
        RECT 655.700 310.300 656.300 313.600 ;
        RECT 654.000 309.700 656.300 310.300 ;
        RECT 654.000 309.600 654.800 309.700 ;
        RECT 657.200 309.600 658.000 310.400 ;
        RECT 650.800 307.600 651.600 308.400 ;
        RECT 650.900 306.400 651.500 307.600 ;
        RECT 650.800 305.600 651.600 306.400 ;
        RECT 654.100 298.400 654.700 309.600 ;
        RECT 655.600 307.600 656.400 308.400 ;
        RECT 655.700 300.400 656.300 307.600 ;
        RECT 655.600 299.600 656.400 300.400 ;
        RECT 639.600 297.600 640.400 298.400 ;
        RECT 649.200 297.600 650.000 298.400 ;
        RECT 650.800 297.600 651.600 298.400 ;
        RECT 654.000 297.600 654.800 298.400 ;
        RECT 650.900 296.400 651.500 297.600 ;
        RECT 650.800 295.600 651.600 296.400 ;
        RECT 639.600 293.600 640.400 294.400 ;
        RECT 644.400 293.600 645.200 294.400 ;
        RECT 646.000 293.600 646.800 294.400 ;
        RECT 634.800 273.600 635.600 274.400 ;
        RECT 638.000 273.600 638.800 274.400 ;
        RECT 634.900 270.400 635.500 273.600 ;
        RECT 639.700 272.400 640.300 293.600 ;
        RECT 641.200 291.600 642.000 292.400 ;
        RECT 641.300 288.400 641.900 291.600 ;
        RECT 641.200 287.600 642.000 288.400 ;
        RECT 639.600 271.600 640.400 272.400 ;
        RECT 642.800 271.600 643.600 272.400 ;
        RECT 639.700 270.400 640.300 271.600 ;
        RECT 617.200 269.600 618.000 270.400 ;
        RECT 628.400 269.600 629.200 270.400 ;
        RECT 630.000 269.600 630.800 270.400 ;
        RECT 634.800 269.600 635.600 270.400 ;
        RECT 636.400 269.600 637.200 270.400 ;
        RECT 639.600 269.600 640.400 270.400 ;
        RECT 618.800 267.600 619.600 268.400 ;
        RECT 626.800 267.600 627.600 268.400 ;
        RECT 612.400 265.600 613.200 266.400 ;
        RECT 622.000 265.600 622.800 266.400 ;
        RECT 601.200 263.600 602.000 264.400 ;
        RECT 596.400 259.600 597.200 260.400 ;
        RECT 601.300 258.400 601.900 263.600 ;
        RECT 612.500 258.400 613.100 265.600 ;
        RECT 626.900 264.400 627.500 267.600 ;
        RECT 630.100 266.400 630.700 269.600 ;
        RECT 630.000 265.600 630.800 266.400 ;
        RECT 614.000 263.600 614.800 264.400 ;
        RECT 626.800 263.600 627.600 264.400 ;
        RECT 594.800 251.600 595.600 252.400 ;
        RECT 596.400 246.200 597.200 257.800 ;
        RECT 601.200 257.600 602.000 258.400 ;
        RECT 602.800 257.600 603.600 258.400 ;
        RECT 607.600 246.200 608.400 257.800 ;
        RECT 612.400 257.600 613.200 258.400 ;
        RECT 614.100 252.400 614.700 263.600 ;
        RECT 612.400 251.600 613.200 252.400 ;
        RECT 614.000 251.600 614.800 252.400 ;
        RECT 617.200 246.200 618.000 257.800 ;
        RECT 622.000 257.600 622.800 258.400 ;
        RECT 618.800 253.600 619.600 254.400 ;
        RECT 554.800 231.600 555.600 232.400 ;
        RECT 556.400 231.600 557.200 232.400 ;
        RECT 558.000 231.600 558.800 232.400 ;
        RECT 566.000 231.600 566.800 232.400 ;
        RECT 572.400 231.600 573.200 232.400 ;
        RECT 542.000 229.600 542.800 230.400 ;
        RECT 550.000 229.600 550.800 230.400 ;
        RECT 553.200 229.600 554.000 230.400 ;
        RECT 540.400 227.600 541.200 228.400 ;
        RECT 542.100 226.400 542.700 229.600 ;
        RECT 534.000 225.600 534.800 226.400 ;
        RECT 538.800 225.600 539.600 226.400 ;
        RECT 542.000 226.300 542.800 226.400 ;
        RECT 540.500 225.700 542.800 226.300 ;
        RECT 537.200 223.600 538.000 224.400 ;
        RECT 518.000 217.600 518.800 218.400 ;
        RECT 527.600 217.600 528.400 218.400 ;
        RECT 529.200 217.600 530.000 218.400 ;
        RECT 537.300 218.300 537.900 223.600 ;
        RECT 537.300 217.700 539.500 218.300 ;
        RECT 537.200 215.600 538.000 216.400 ;
        RECT 522.800 213.600 523.600 214.400 ;
        RECT 511.600 211.600 512.400 212.400 ;
        RECT 519.600 203.600 520.400 204.400 ;
        RECT 503.600 201.600 504.400 202.400 ;
        RECT 506.800 201.600 507.600 202.400 ;
        RECT 506.900 198.400 507.500 201.600 ;
        RECT 506.800 197.600 507.600 198.400 ;
        RECT 518.000 195.600 518.800 196.400 ;
        RECT 518.100 188.400 518.700 195.600 ;
        RECT 519.700 188.400 520.300 203.600 ;
        RECT 522.900 196.400 523.500 213.600 ;
        RECT 537.300 212.400 537.900 215.600 ;
        RECT 538.900 214.400 539.500 217.700 ;
        RECT 540.500 216.400 541.100 225.700 ;
        RECT 542.000 225.600 542.800 225.700 ;
        RECT 546.800 225.600 547.600 226.400 ;
        RECT 545.200 223.600 546.000 224.400 ;
        RECT 548.400 223.600 549.200 224.400 ;
        RECT 540.400 215.600 541.200 216.400 ;
        RECT 545.300 214.400 545.900 223.600 ;
        RECT 548.500 216.400 549.100 223.600 ;
        RECT 548.400 215.600 549.200 216.400 ;
        RECT 538.800 213.600 539.600 214.400 ;
        RECT 543.600 213.600 544.400 214.400 ;
        RECT 545.200 213.600 546.000 214.400 ;
        RECT 548.400 213.600 549.200 214.400 ;
        RECT 524.400 211.600 525.200 212.400 ;
        RECT 537.200 211.600 538.000 212.400 ;
        RECT 545.200 211.600 546.000 212.400 ;
        RECT 522.800 195.600 523.600 196.400 ;
        RECT 516.400 187.600 517.200 188.400 ;
        RECT 518.000 187.600 518.800 188.400 ;
        RECT 519.600 187.600 520.400 188.400 ;
        RECT 516.500 186.400 517.100 187.600 ;
        RECT 522.900 186.400 523.500 195.600 ;
        RECT 524.500 186.400 525.100 211.600 ;
        RECT 527.600 209.600 528.400 210.400 ;
        RECT 529.200 209.600 530.000 210.400 ;
        RECT 534.000 209.600 534.800 210.400 ;
        RECT 529.300 208.400 529.900 209.600 ;
        RECT 529.200 207.600 530.000 208.400 ;
        RECT 534.100 206.400 534.700 209.600 ;
        RECT 526.000 205.600 526.800 206.400 ;
        RECT 534.000 205.600 534.800 206.400 ;
        RECT 526.100 198.400 526.700 205.600 ;
        RECT 526.000 197.600 526.800 198.400 ;
        RECT 529.000 191.800 529.800 192.600 ;
        RECT 535.600 191.800 536.400 192.600 ;
        RECT 526.000 189.600 526.800 190.400 ;
        RECT 526.100 186.400 526.700 189.600 ;
        RECT 529.000 187.000 529.600 191.800 ;
        RECT 531.600 188.400 532.400 188.600 ;
        RECT 535.800 188.400 536.400 191.800 ;
        RECT 531.600 187.800 536.400 188.400 ;
        RECT 530.800 187.000 531.600 187.200 ;
        RECT 534.200 187.000 535.000 187.200 ;
        RECT 535.800 187.000 536.400 187.800 ;
        RECT 537.200 187.600 538.000 188.400 ;
        RECT 516.400 185.600 517.200 186.400 ;
        RECT 522.800 185.600 523.600 186.400 ;
        RECT 524.400 185.600 525.200 186.400 ;
        RECT 526.000 185.600 526.800 186.400 ;
        RECT 529.000 186.200 529.800 187.000 ;
        RECT 530.800 186.400 535.000 187.000 ;
        RECT 506.800 183.600 507.600 184.400 ;
        RECT 513.200 183.600 514.000 184.400 ;
        RECT 518.000 183.600 518.800 184.400 ;
        RECT 521.200 183.600 522.000 184.400 ;
        RECT 530.800 183.600 531.600 184.400 ;
        RECT 532.400 183.600 533.200 184.400 ;
        RECT 506.900 178.400 507.500 183.600 ;
        RECT 513.300 180.400 513.900 183.600 ;
        RECT 513.200 179.600 514.000 180.400 ;
        RECT 506.800 177.600 507.600 178.400 ;
        RECT 500.400 173.600 501.200 174.400 ;
        RECT 500.500 172.400 501.100 173.600 ;
        RECT 500.400 171.600 501.200 172.400 ;
        RECT 503.600 171.600 504.400 172.400 ;
        RECT 497.200 163.600 498.000 164.400 ;
        RECT 497.300 162.400 497.900 163.600 ;
        RECT 497.200 161.600 498.000 162.400 ;
        RECT 494.000 159.600 494.800 160.400 ;
        RECT 489.200 147.600 490.000 148.400 ;
        RECT 490.800 144.200 491.600 155.800 ;
        RECT 492.400 145.600 493.200 146.400 ;
        RECT 492.500 142.400 493.100 145.600 ;
        RECT 494.000 144.200 494.800 155.800 ;
        RECT 495.600 144.200 496.400 157.800 ;
        RECT 497.200 144.200 498.000 157.800 ;
        RECT 498.800 144.200 499.600 157.800 ;
        RECT 492.400 141.600 493.200 142.400 ;
        RECT 476.400 133.600 477.200 134.400 ;
        RECT 473.200 123.600 474.000 124.400 ;
        RECT 484.400 124.200 485.200 137.800 ;
        RECT 486.000 124.200 486.800 137.800 ;
        RECT 487.600 126.200 488.400 137.800 ;
        RECT 489.200 133.600 490.000 134.400 ;
        RECT 490.800 126.200 491.600 137.800 ;
        RECT 492.400 135.600 493.200 136.400 ;
        RECT 494.000 126.200 494.800 137.800 ;
        RECT 495.600 124.200 496.400 137.800 ;
        RECT 497.200 124.200 498.000 137.800 ;
        RECT 498.800 124.200 499.600 137.800 ;
        RECT 500.500 132.400 501.100 171.600 ;
        RECT 503.700 168.400 504.300 171.600 ;
        RECT 503.600 167.600 504.400 168.400 ;
        RECT 506.900 136.400 507.500 177.600 ;
        RECT 508.400 171.600 509.200 172.400 ;
        RECT 513.200 164.200 514.000 177.800 ;
        RECT 514.800 164.200 515.600 177.800 ;
        RECT 516.400 166.200 517.200 177.800 ;
        RECT 518.100 174.400 518.700 183.600 ;
        RECT 521.300 182.400 521.900 183.600 ;
        RECT 521.200 181.600 522.000 182.400 ;
        RECT 530.800 181.600 531.600 182.400 ;
        RECT 518.000 173.600 518.800 174.400 ;
        RECT 518.000 165.600 518.800 166.400 ;
        RECT 519.600 166.200 520.400 177.800 ;
        RECT 521.200 177.600 522.000 178.400 ;
        RECT 521.300 176.400 521.900 177.600 ;
        RECT 521.200 175.600 522.000 176.400 ;
        RECT 522.800 166.200 523.600 177.800 ;
        RECT 508.400 159.600 509.200 160.400 ;
        RECT 508.500 158.400 509.100 159.600 ;
        RECT 518.100 158.400 518.700 165.600 ;
        RECT 524.400 164.200 525.200 177.800 ;
        RECT 526.000 164.200 526.800 177.800 ;
        RECT 527.600 164.200 528.400 177.800 ;
        RECT 508.400 157.600 509.200 158.400 ;
        RECT 511.600 157.600 512.400 158.400 ;
        RECT 518.000 157.600 518.800 158.400 ;
        RECT 508.400 147.600 509.200 148.400 ;
        RECT 508.500 138.400 509.100 147.600 ;
        RECT 510.000 145.600 510.800 146.400 ;
        RECT 511.700 138.400 512.300 157.600 ;
        RECT 530.900 152.400 531.500 181.600 ;
        RECT 514.800 152.300 515.600 152.400 ;
        RECT 513.300 151.700 515.600 152.300 ;
        RECT 508.400 137.600 509.200 138.400 ;
        RECT 511.600 137.600 512.400 138.400 ;
        RECT 506.800 135.600 507.600 136.400 ;
        RECT 500.400 131.600 501.200 132.400 ;
        RECT 510.000 129.600 510.800 130.400 ;
        RECT 471.600 115.600 472.400 116.400 ;
        RECT 471.700 114.400 472.300 115.600 ;
        RECT 471.600 113.600 472.400 114.400 ;
        RECT 466.800 107.700 469.100 108.300 ;
        RECT 466.800 107.600 467.600 107.700 ;
        RECT 470.000 107.600 470.800 108.400 ;
        RECT 471.600 107.600 472.400 108.400 ;
        RECT 465.300 100.400 465.900 107.600 ;
        RECT 465.200 99.600 466.000 100.400 ;
        RECT 471.700 98.400 472.300 107.600 ;
        RECT 473.300 98.400 473.900 123.600 ;
        RECT 474.800 117.600 475.600 118.400 ;
        RECT 474.900 112.400 475.500 117.600 ;
        RECT 482.800 115.600 483.600 116.400 ;
        RECT 479.600 113.600 480.400 114.400 ;
        RECT 479.700 112.400 480.300 113.600 ;
        RECT 474.800 111.600 475.600 112.400 ;
        RECT 479.600 111.600 480.400 112.400 ;
        RECT 490.800 109.600 491.600 110.400 ;
        RECT 476.400 107.600 477.200 108.400 ;
        RECT 481.200 107.600 482.000 108.400 ;
        RECT 484.400 105.600 485.200 106.400 ;
        RECT 474.800 103.600 475.600 104.400 ;
        RECT 465.200 97.600 466.000 98.400 ;
        RECT 471.600 97.600 472.400 98.400 ;
        RECT 473.200 97.600 474.000 98.400 ;
        RECT 474.900 96.400 475.500 103.600 ;
        RECT 474.800 95.600 475.600 96.400 ;
        RECT 476.400 91.600 477.200 92.400 ;
        RECT 476.500 88.400 477.100 91.600 ;
        RECT 465.200 87.600 466.000 88.400 ;
        RECT 476.400 87.600 477.200 88.400 ;
        RECT 462.000 77.600 462.800 78.400 ;
        RECT 465.300 74.400 465.900 87.600 ;
        RECT 478.000 84.200 478.800 97.800 ;
        RECT 479.600 84.200 480.400 97.800 ;
        RECT 481.200 84.200 482.000 97.800 ;
        RECT 482.800 86.200 483.600 97.800 ;
        RECT 484.500 96.400 485.100 105.600 ;
        RECT 490.900 100.400 491.500 109.600 ;
        RECT 492.400 104.200 493.200 117.800 ;
        RECT 494.000 104.200 494.800 117.800 ;
        RECT 495.600 104.200 496.400 117.800 ;
        RECT 497.200 104.200 498.000 115.800 ;
        RECT 498.800 105.600 499.600 106.400 ;
        RECT 500.400 104.200 501.200 115.800 ;
        RECT 502.000 107.600 502.800 108.400 ;
        RECT 503.600 104.200 504.400 115.800 ;
        RECT 505.200 104.200 506.000 117.800 ;
        RECT 506.800 104.200 507.600 117.800 ;
        RECT 506.800 101.600 507.600 102.400 ;
        RECT 490.800 99.600 491.600 100.400 ;
        RECT 495.600 99.600 496.400 100.400 ;
        RECT 484.400 95.600 485.200 96.400 ;
        RECT 486.000 86.200 486.800 97.800 ;
        RECT 487.600 95.600 488.400 96.400 ;
        RECT 487.700 94.400 488.300 95.600 ;
        RECT 487.600 93.600 488.400 94.400 ;
        RECT 489.200 86.200 490.000 97.800 ;
        RECT 490.800 84.200 491.600 97.800 ;
        RECT 492.400 84.200 493.200 97.800 ;
        RECT 495.700 92.400 496.300 99.600 ;
        RECT 506.900 98.400 507.500 101.600 ;
        RECT 510.100 98.400 510.700 129.600 ;
        RECT 511.600 109.600 512.400 110.400 ;
        RECT 513.300 98.400 513.900 151.700 ;
        RECT 514.800 151.600 515.600 151.700 ;
        RECT 521.200 151.600 522.000 152.400 ;
        RECT 527.600 151.600 528.400 152.400 ;
        RECT 530.800 151.600 531.600 152.400 ;
        RECT 514.800 149.600 515.600 150.400 ;
        RECT 518.000 149.600 518.800 150.400 ;
        RECT 519.600 149.600 520.400 150.400 ;
        RECT 519.700 148.400 520.300 149.600 ;
        RECT 521.300 148.400 521.900 151.600 ;
        RECT 522.800 149.600 523.600 150.400 ;
        RECT 519.600 147.600 520.400 148.400 ;
        RECT 521.200 147.600 522.000 148.400 ;
        RECT 519.700 136.400 520.300 147.600 ;
        RECT 522.900 146.300 523.500 149.600 ;
        RECT 527.700 148.400 528.300 151.600 ;
        RECT 530.900 150.400 531.500 151.600 ;
        RECT 530.800 149.600 531.600 150.400 ;
        RECT 532.500 148.400 533.100 183.600 ;
        RECT 534.100 170.400 534.700 186.400 ;
        RECT 535.600 186.200 536.400 187.000 ;
        RECT 537.300 184.400 537.900 187.600 ;
        RECT 538.800 186.200 539.600 191.800 ;
        RECT 540.400 187.600 541.200 188.400 ;
        RECT 537.200 183.600 538.000 184.400 ;
        RECT 540.500 178.400 541.100 187.600 ;
        RECT 542.000 184.200 542.800 195.800 ;
        RECT 545.200 189.600 546.000 190.400 ;
        RECT 545.200 187.600 546.000 188.400 ;
        RECT 540.400 177.600 541.200 178.400 ;
        RECT 542.000 175.600 542.800 176.400 ;
        RECT 545.300 172.400 545.900 187.600 ;
        RECT 550.100 178.400 550.700 229.600 ;
        RECT 554.900 226.400 555.500 231.600 ;
        RECT 556.500 230.400 557.100 231.600 ;
        RECT 558.100 230.400 558.700 231.600 ;
        RECT 556.400 229.600 557.200 230.400 ;
        RECT 558.000 229.600 558.800 230.400 ;
        RECT 556.400 227.600 557.200 228.400 ;
        RECT 559.600 227.600 560.400 228.400 ;
        RECT 561.200 227.600 562.000 228.400 ;
        RECT 554.800 225.600 555.600 226.400 ;
        RECT 556.500 216.400 557.100 227.600 ;
        RECT 561.300 226.400 561.900 227.600 ;
        RECT 561.200 225.600 562.000 226.400 ;
        RECT 562.800 223.600 563.600 224.400 ;
        RECT 556.400 215.600 557.200 216.400 ;
        RECT 551.600 213.600 552.400 214.400 ;
        RECT 554.800 213.600 555.600 214.400 ;
        RECT 551.700 212.400 552.300 213.600 ;
        RECT 554.900 212.400 555.500 213.600 ;
        RECT 551.600 211.600 552.400 212.400 ;
        RECT 554.800 211.600 555.600 212.400 ;
        RECT 556.500 210.400 557.100 215.600 ;
        RECT 561.200 212.300 562.000 212.400 ;
        RECT 562.900 212.300 563.500 223.600 ;
        RECT 564.400 215.600 565.200 216.400 ;
        RECT 561.200 211.700 563.500 212.300 ;
        RECT 561.200 211.600 562.000 211.700 ;
        RECT 554.800 209.600 555.600 210.400 ;
        RECT 556.400 209.600 557.200 210.400 ;
        RECT 554.900 208.400 555.500 209.600 ;
        RECT 551.600 207.600 552.400 208.400 ;
        RECT 554.800 207.600 555.600 208.400 ;
        RECT 551.600 184.200 552.400 195.800 ;
        RECT 554.900 182.400 555.500 207.600 ;
        RECT 556.500 188.300 557.100 209.600 ;
        RECT 564.500 208.400 565.100 215.600 ;
        RECT 566.100 214.400 566.700 231.600 ;
        RECT 572.500 230.400 573.100 231.600 ;
        RECT 572.400 229.600 573.200 230.400 ;
        RECT 585.200 229.600 586.000 230.400 ;
        RECT 567.600 228.300 568.400 228.400 ;
        RECT 569.200 228.300 570.000 228.400 ;
        RECT 567.600 227.700 570.000 228.300 ;
        RECT 567.600 227.600 568.400 227.700 ;
        RECT 569.200 227.600 570.000 227.700 ;
        RECT 566.000 213.600 566.800 214.400 ;
        RECT 566.100 212.400 566.700 213.600 ;
        RECT 566.000 211.600 566.800 212.400 ;
        RECT 564.400 207.600 565.200 208.400 ;
        RECT 559.600 193.600 560.400 194.400 ;
        RECT 559.700 190.400 560.300 193.600 ;
        RECT 564.400 191.600 565.200 192.400 ;
        RECT 564.500 190.400 565.100 191.600 ;
        RECT 559.600 189.600 560.400 190.400 ;
        RECT 561.200 189.600 562.000 190.400 ;
        RECT 564.400 190.300 565.200 190.400 ;
        RECT 562.900 189.700 565.200 190.300 ;
        RECT 558.000 188.300 558.800 188.400 ;
        RECT 556.500 187.700 558.800 188.300 ;
        RECT 558.000 187.600 558.800 187.700 ;
        RECT 558.100 186.400 558.700 187.600 ;
        RECT 558.000 185.600 558.800 186.400 ;
        RECT 556.400 183.600 557.200 184.400 ;
        RECT 554.800 181.600 555.600 182.400 ;
        RECT 550.000 177.600 550.800 178.400 ;
        RECT 554.800 175.600 555.600 176.400 ;
        RECT 554.800 173.600 555.600 174.400 ;
        RECT 545.200 171.600 546.000 172.400 ;
        RECT 546.800 171.600 547.600 172.400 ;
        RECT 534.000 169.600 534.800 170.400 ;
        RECT 545.300 164.400 545.900 171.600 ;
        RECT 546.900 168.400 547.500 171.600 ;
        RECT 556.400 169.600 557.200 170.400 ;
        RECT 546.800 167.600 547.600 168.400 ;
        RECT 537.200 163.600 538.000 164.400 ;
        RECT 542.000 163.600 542.800 164.400 ;
        RECT 545.200 163.600 546.000 164.400 ;
        RECT 553.200 163.600 554.000 164.400 ;
        RECT 534.000 159.600 534.800 160.400 ;
        RECT 527.600 147.600 528.400 148.400 ;
        RECT 532.400 147.600 533.200 148.400 ;
        RECT 532.500 146.400 533.100 147.600 ;
        RECT 534.100 146.400 534.700 159.600 ;
        RECT 537.300 156.400 537.900 163.600 ;
        RECT 540.400 161.600 541.200 162.400 ;
        RECT 540.500 158.400 541.100 161.600 ;
        RECT 540.400 157.600 541.200 158.400 ;
        RECT 537.200 155.600 538.000 156.400 ;
        RECT 542.100 152.400 542.700 163.600 ;
        RECT 546.800 161.600 547.600 162.400 ;
        RECT 543.600 159.600 544.400 160.400 ;
        RECT 537.200 151.600 538.000 152.400 ;
        RECT 542.000 151.600 542.800 152.400 ;
        RECT 522.900 145.700 525.100 146.300 ;
        RECT 516.400 135.600 517.200 136.400 ;
        RECT 519.600 135.600 520.400 136.400 ;
        RECT 516.500 134.400 517.100 135.600 ;
        RECT 516.400 133.600 517.200 134.400 ;
        RECT 514.800 131.600 515.600 132.400 ;
        RECT 518.000 127.600 518.800 128.400 ;
        RECT 516.400 109.600 517.200 110.400 ;
        RECT 516.500 108.400 517.100 109.600 ;
        RECT 516.400 107.600 517.200 108.400 ;
        RECT 506.800 97.600 507.600 98.400 ;
        RECT 510.000 97.600 510.800 98.400 ;
        RECT 513.200 97.600 514.000 98.400 ;
        RECT 518.000 97.600 518.800 98.400 ;
        RECT 518.100 96.400 518.700 97.600 ;
        RECT 503.600 95.600 504.400 96.400 ;
        RECT 518.000 95.600 518.800 96.400 ;
        RECT 502.000 93.600 502.800 94.400 ;
        RECT 503.700 92.400 504.300 95.600 ;
        RECT 508.400 93.600 509.200 94.400 ;
        RECT 510.000 93.600 510.800 94.400 ;
        RECT 518.000 94.300 518.800 94.400 ;
        RECT 519.700 94.300 520.300 135.600 ;
        RECT 522.800 126.200 523.600 137.800 ;
        RECT 522.800 115.600 523.600 116.400 ;
        RECT 522.900 112.400 523.500 115.600 ;
        RECT 521.200 111.600 522.000 112.400 ;
        RECT 522.800 111.600 523.600 112.400 ;
        RECT 521.300 110.400 521.900 111.600 ;
        RECT 521.200 109.600 522.000 110.400 ;
        RECT 524.500 104.400 525.100 145.700 ;
        RECT 532.400 145.600 533.200 146.400 ;
        RECT 534.000 145.600 534.800 146.400 ;
        RECT 537.300 146.300 537.900 151.600 ;
        RECT 538.800 149.600 539.600 150.400 ;
        RECT 542.000 149.600 542.800 150.400 ;
        RECT 542.000 148.300 542.800 148.400 ;
        RECT 543.700 148.300 544.300 159.600 ;
        RECT 546.900 152.400 547.500 161.600 ;
        RECT 550.000 155.600 550.800 156.400 ;
        RECT 546.800 151.600 547.600 152.400 ;
        RECT 550.100 148.400 550.700 155.600 ;
        RECT 542.000 147.700 544.300 148.300 ;
        RECT 542.000 147.600 542.800 147.700 ;
        RECT 550.000 147.600 550.800 148.400 ;
        RECT 538.800 146.300 539.600 146.400 ;
        RECT 537.300 145.700 539.600 146.300 ;
        RECT 538.800 145.600 539.600 145.700 ;
        RECT 548.400 145.600 549.200 146.400 ;
        RECT 526.000 143.600 526.800 144.400 ;
        RECT 535.600 144.300 536.400 144.400 ;
        RECT 535.600 143.700 537.900 144.300 ;
        RECT 535.600 143.600 536.400 143.700 ;
        RECT 526.100 134.400 526.700 143.600 ;
        RECT 526.000 133.600 526.800 134.400 ;
        RECT 530.800 131.600 531.600 132.600 ;
        RECT 532.400 126.200 533.200 137.800 ;
        RECT 534.000 133.600 534.800 134.400 ;
        RECT 534.100 130.400 534.700 133.600 ;
        RECT 534.000 129.600 534.800 130.400 ;
        RECT 535.600 130.200 536.400 135.800 ;
        RECT 537.300 132.400 537.900 143.700 ;
        RECT 537.200 131.600 538.000 132.400 ;
        RECT 537.300 124.400 537.900 131.600 ;
        RECT 537.200 123.600 538.000 124.400 ;
        RECT 530.800 119.600 531.600 120.400 ;
        RECT 526.000 113.600 526.800 114.400 ;
        RECT 526.000 111.600 526.800 112.400 ;
        RECT 526.100 110.400 526.700 111.600 ;
        RECT 526.000 109.600 526.800 110.400 ;
        RECT 527.600 107.600 528.400 108.400 ;
        RECT 529.200 107.600 530.000 108.400 ;
        RECT 524.400 103.600 525.200 104.400 ;
        RECT 527.700 98.400 528.300 107.600 ;
        RECT 529.300 106.400 529.900 107.600 ;
        RECT 529.200 105.600 530.000 106.400 ;
        RECT 527.600 97.600 528.400 98.400 ;
        RECT 521.200 94.300 522.000 94.400 ;
        RECT 518.000 93.700 522.000 94.300 ;
        RECT 518.000 93.600 518.800 93.700 ;
        RECT 521.200 93.600 522.000 93.700 ;
        RECT 495.600 91.600 496.400 92.400 ;
        RECT 503.600 91.600 504.400 92.400 ;
        RECT 506.800 89.600 507.600 90.400 ;
        RECT 465.200 73.600 466.000 74.400 ;
        RECT 468.400 69.600 469.200 70.400 ;
        RECT 457.200 67.700 459.500 68.300 ;
        RECT 457.200 67.600 458.000 67.700 ;
        RECT 447.600 57.600 448.400 58.400 ;
        RECT 452.400 57.600 453.200 58.400 ;
        RECT 455.600 57.600 456.400 58.400 ;
        RECT 442.800 55.600 443.600 56.400 ;
        RECT 441.200 53.600 442.000 54.400 ;
        RECT 428.400 51.600 429.200 52.400 ;
        RECT 434.800 51.600 435.600 52.400 ;
        RECT 439.600 51.600 440.400 52.400 ;
        RECT 433.200 47.600 434.000 48.400 ;
        RECT 433.300 38.400 433.900 47.600 ;
        RECT 426.800 37.600 427.600 38.400 ;
        RECT 433.200 37.600 434.000 38.400 ;
        RECT 407.600 35.600 408.400 36.400 ;
        RECT 422.000 35.600 422.800 36.400 ;
        RECT 414.000 33.600 414.800 34.400 ;
        RECT 422.100 32.400 422.700 35.600 ;
        RECT 410.800 31.600 411.600 32.400 ;
        RECT 422.000 31.600 422.800 32.400 ;
        RECT 410.800 29.600 411.600 30.400 ;
        RECT 414.000 29.600 414.800 30.400 ;
        RECT 426.900 28.400 427.500 37.600 ;
        RECT 434.900 32.400 435.500 51.600 ;
        RECT 442.900 40.400 443.500 55.600 ;
        RECT 457.300 54.400 457.900 67.600 ;
        RECT 468.500 66.400 469.100 69.600 ;
        RECT 462.000 65.600 462.800 66.400 ;
        RECT 468.400 65.600 469.200 66.400 ;
        RECT 444.400 53.600 445.200 54.400 ;
        RECT 449.200 53.600 450.000 54.400 ;
        RECT 454.000 53.600 454.800 54.400 ;
        RECT 457.200 54.300 458.000 54.400 ;
        RECT 457.200 53.700 459.500 54.300 ;
        RECT 457.200 53.600 458.000 53.700 ;
        RECT 442.800 39.600 443.600 40.400 ;
        RECT 434.800 31.600 435.600 32.400 ;
        RECT 428.400 29.600 429.200 30.400 ;
        RECT 434.800 29.600 435.600 30.400 ;
        RECT 401.200 27.600 402.000 28.400 ;
        RECT 415.600 27.600 416.400 28.400 ;
        RECT 426.800 27.600 427.600 28.400 ;
        RECT 404.400 23.600 405.200 24.400 ;
        RECT 417.200 23.600 418.000 24.400 ;
        RECT 388.400 19.600 389.200 20.400 ;
        RECT 396.400 19.600 397.200 20.400 ;
        RECT 366.000 11.600 366.800 12.400 ;
        RECT 370.800 11.600 371.600 12.400 ;
        RECT 375.600 11.600 376.400 12.400 ;
        RECT 378.800 11.600 379.600 12.400 ;
        RECT 383.600 11.600 384.400 12.400 ;
        RECT 388.400 4.200 389.200 17.800 ;
        RECT 390.000 4.200 390.800 17.800 ;
        RECT 391.600 6.200 392.400 17.800 ;
        RECT 393.200 15.600 394.000 16.400 ;
        RECT 393.300 14.400 393.900 15.600 ;
        RECT 393.200 13.600 394.000 14.400 ;
        RECT 394.800 6.200 395.600 17.800 ;
        RECT 396.500 16.400 397.100 19.600 ;
        RECT 396.400 15.600 397.200 16.400 ;
        RECT 398.000 6.200 398.800 17.800 ;
        RECT 399.600 4.200 400.400 17.800 ;
        RECT 401.200 4.200 402.000 17.800 ;
        RECT 402.800 4.200 403.600 17.800 ;
        RECT 417.300 16.400 417.900 23.600 ;
        RECT 417.200 15.600 418.000 16.400 ;
        RECT 412.400 13.600 413.400 14.400 ;
        RECT 418.800 13.600 419.600 14.400 ;
        RECT 418.900 12.400 419.500 13.600 ;
        RECT 428.500 12.400 429.100 29.600 ;
        RECT 430.000 25.600 430.800 26.400 ;
        RECT 430.100 14.400 430.700 25.600 ;
        RECT 439.600 24.200 440.400 37.800 ;
        RECT 441.200 24.200 442.000 37.800 ;
        RECT 442.800 24.200 443.600 35.800 ;
        RECT 444.500 30.400 445.100 53.600 ;
        RECT 455.600 51.600 456.400 52.400 ;
        RECT 454.000 47.600 454.800 48.400 ;
        RECT 447.600 43.600 448.400 44.400 ;
        RECT 444.400 29.600 445.200 30.400 ;
        RECT 444.400 27.600 445.200 28.400 ;
        RECT 446.000 24.200 446.800 35.800 ;
        RECT 447.700 32.400 448.300 43.600 ;
        RECT 454.100 42.400 454.700 47.600 ;
        RECT 454.000 41.600 454.800 42.400 ;
        RECT 447.600 31.600 448.400 32.400 ;
        RECT 447.600 25.600 448.400 26.400 ;
        RECT 447.700 20.400 448.300 25.600 ;
        RECT 449.200 24.200 450.000 35.800 ;
        RECT 450.800 24.200 451.600 37.800 ;
        RECT 452.400 24.200 453.200 37.800 ;
        RECT 454.000 24.200 454.800 37.800 ;
        RECT 455.700 30.400 456.300 51.600 ;
        RECT 457.200 47.600 458.000 48.400 ;
        RECT 457.300 38.400 457.900 47.600 ;
        RECT 457.200 37.600 458.000 38.400 ;
        RECT 455.600 29.600 456.400 30.400 ;
        RECT 441.200 19.600 442.000 20.400 ;
        RECT 447.600 19.600 448.400 20.400 ;
        RECT 430.000 13.600 430.800 14.400 ;
        RECT 404.400 11.600 405.200 12.400 ;
        RECT 418.800 11.600 419.600 12.400 ;
        RECT 428.400 11.600 429.200 12.400 ;
        RECT 433.200 4.200 434.000 17.800 ;
        RECT 434.800 4.200 435.600 17.800 ;
        RECT 436.400 6.200 437.200 17.800 ;
        RECT 438.000 13.600 438.800 14.400 ;
        RECT 439.600 6.200 440.400 17.800 ;
        RECT 441.300 16.400 441.900 19.600 ;
        RECT 441.200 15.600 442.000 16.400 ;
        RECT 442.800 6.200 443.600 17.800 ;
        RECT 444.400 4.200 445.200 17.800 ;
        RECT 446.000 4.200 446.800 17.800 ;
        RECT 447.600 4.200 448.400 17.800 ;
        RECT 458.900 16.400 459.500 53.700 ;
        RECT 462.100 52.400 462.700 65.600 ;
        RECT 473.200 64.200 474.000 77.800 ;
        RECT 474.800 64.200 475.600 77.800 ;
        RECT 476.400 64.200 477.200 75.800 ;
        RECT 478.000 71.600 478.800 72.400 ;
        RECT 478.100 68.400 478.700 71.600 ;
        RECT 478.000 67.600 478.800 68.400 ;
        RECT 479.600 64.200 480.400 75.800 ;
        RECT 481.200 65.600 482.000 66.400 ;
        RECT 481.300 60.400 481.900 65.600 ;
        RECT 482.800 64.200 483.600 75.800 ;
        RECT 484.400 64.200 485.200 77.800 ;
        RECT 486.000 64.200 486.800 77.800 ;
        RECT 487.600 64.200 488.400 77.800 ;
        RECT 502.000 73.600 502.800 74.400 ;
        RECT 502.100 66.400 502.700 73.600 ;
        RECT 497.200 65.600 498.000 66.400 ;
        RECT 498.800 65.600 499.600 66.400 ;
        RECT 502.000 65.600 502.800 66.400 ;
        RECT 503.600 65.600 504.400 66.400 ;
        RECT 474.800 59.600 475.600 60.400 ;
        RECT 481.200 59.600 482.000 60.400 ;
        RECT 462.000 51.600 462.800 52.400 ;
        RECT 466.800 44.200 467.600 57.800 ;
        RECT 468.400 44.200 469.200 57.800 ;
        RECT 470.000 46.200 470.800 57.800 ;
        RECT 471.600 53.600 472.400 54.400 ;
        RECT 473.200 46.200 474.000 57.800 ;
        RECT 474.900 56.400 475.500 59.600 ;
        RECT 474.800 55.600 475.600 56.400 ;
        RECT 468.400 41.600 469.200 42.400 ;
        RECT 463.600 37.600 464.400 38.400 ;
        RECT 462.000 31.600 462.800 32.400 ;
        RECT 466.800 31.600 467.600 32.400 ;
        RECT 462.100 16.400 462.700 31.600 ;
        RECT 466.900 30.400 467.500 31.600 ;
        RECT 466.800 29.600 467.600 30.400 ;
        RECT 465.200 27.600 466.000 28.400 ;
        RECT 465.300 18.400 465.900 27.600 ;
        RECT 466.900 26.400 467.500 29.600 ;
        RECT 466.800 25.600 467.600 26.400 ;
        RECT 468.500 18.400 469.100 41.600 ;
        RECT 473.200 37.600 474.000 38.400 ;
        RECT 473.300 32.400 473.900 37.600 ;
        RECT 473.200 31.600 474.000 32.400 ;
        RECT 470.000 27.600 470.800 28.400 ;
        RECT 474.900 20.400 475.500 55.600 ;
        RECT 476.400 46.200 477.200 57.800 ;
        RECT 478.000 44.200 478.800 57.800 ;
        RECT 479.600 44.200 480.400 57.800 ;
        RECT 481.200 44.200 482.000 57.800 ;
        RECT 490.800 57.600 491.600 58.400 ;
        RECT 498.900 54.400 499.500 65.600 ;
        RECT 502.100 58.400 502.700 65.600 ;
        RECT 506.900 58.400 507.500 89.600 ;
        RECT 508.400 71.600 509.200 72.400 ;
        RECT 508.400 69.600 509.200 70.400 ;
        RECT 502.000 57.600 502.800 58.400 ;
        RECT 506.800 57.600 507.600 58.400 ;
        RECT 492.400 53.600 493.200 54.400 ;
        RECT 498.800 53.600 499.600 54.400 ;
        RECT 500.400 53.600 501.200 54.400 ;
        RECT 500.500 52.400 501.100 53.600 ;
        RECT 494.000 51.600 494.800 52.400 ;
        RECT 498.800 51.600 499.600 52.400 ;
        RECT 500.400 51.600 501.200 52.400 ;
        RECT 494.100 50.400 494.700 51.600 ;
        RECT 498.900 50.400 499.500 51.600 ;
        RECT 494.000 49.600 494.800 50.400 ;
        RECT 498.800 49.600 499.600 50.400 ;
        RECT 500.400 50.300 501.200 50.400 ;
        RECT 502.100 50.300 502.700 57.600 ;
        RECT 505.200 55.600 506.000 56.400 ;
        RECT 505.300 54.400 505.900 55.600 ;
        RECT 505.200 53.600 506.000 54.400 ;
        RECT 503.600 51.600 504.400 52.400 ;
        RECT 500.400 49.700 502.700 50.300 ;
        RECT 500.400 49.600 501.200 49.700 ;
        RECT 497.200 47.600 498.000 48.400 ;
        RECT 479.600 41.600 480.400 42.400 ;
        RECT 478.000 39.600 478.800 40.400 ;
        RECT 478.100 34.400 478.700 39.600 ;
        RECT 478.000 33.600 478.800 34.400 ;
        RECT 476.400 29.600 477.200 30.400 ;
        RECT 478.100 28.400 478.700 33.600 ;
        RECT 479.700 32.400 480.300 41.600 ;
        RECT 497.300 38.400 497.900 47.600 ;
        RECT 497.200 37.600 498.000 38.400 ;
        RECT 484.400 33.600 485.200 34.400 ;
        RECT 479.600 31.600 480.400 32.400 ;
        RECT 482.800 31.600 483.600 32.400 ;
        RECT 482.800 29.600 483.600 30.400 ;
        RECT 484.500 28.400 485.100 33.600 ;
        RECT 486.000 31.600 486.800 32.400 ;
        RECT 489.200 29.600 490.000 30.400 ;
        RECT 478.000 27.600 478.800 28.400 ;
        RECT 484.400 27.600 485.200 28.400 ;
        RECT 487.600 27.600 488.400 28.400 ;
        RECT 474.800 19.600 475.600 20.400 ;
        RECT 484.400 19.600 485.200 20.400 ;
        RECT 465.200 17.600 466.000 18.400 ;
        RECT 468.400 17.600 469.200 18.400 ;
        RECT 458.800 15.600 459.600 16.400 ;
        RECT 462.000 15.600 462.800 16.400 ;
        RECT 458.800 13.600 459.600 14.400 ;
        RECT 449.200 11.600 450.000 12.400 ;
        RECT 476.400 11.600 477.200 12.400 ;
        RECT 478.000 4.200 478.800 17.800 ;
        RECT 479.600 4.200 480.400 17.800 ;
        RECT 481.200 4.200 482.000 17.800 ;
        RECT 482.800 6.200 483.600 17.800 ;
        RECT 484.500 16.400 485.100 19.600 ;
        RECT 484.400 15.600 485.200 16.400 ;
        RECT 486.000 6.200 486.800 17.800 ;
        RECT 487.700 14.400 488.300 27.600 ;
        RECT 489.300 26.400 489.900 29.600 ;
        RECT 498.900 26.400 499.500 49.600 ;
        RECT 503.700 30.400 504.300 51.600 ;
        RECT 505.300 34.400 505.900 53.600 ;
        RECT 508.500 50.400 509.100 69.600 ;
        RECT 510.100 54.400 510.700 93.600 ;
        RECT 530.900 92.400 531.500 119.600 ;
        RECT 537.200 115.600 538.000 116.400 ;
        RECT 537.300 110.400 537.900 115.600 ;
        RECT 537.200 109.600 538.000 110.400 ;
        RECT 532.400 107.600 533.200 108.400 ;
        RECT 530.800 91.600 531.600 92.400 ;
        RECT 526.000 89.600 526.800 90.400 ;
        RECT 527.600 89.600 528.400 90.400 ;
        RECT 511.600 87.600 512.400 88.400 ;
        RECT 513.200 87.600 514.000 88.400 ;
        RECT 511.700 72.300 512.300 87.600 ;
        RECT 513.300 74.400 513.900 87.600 ;
        RECT 522.800 85.600 523.600 86.400 ;
        RECT 513.200 73.600 514.000 74.400 ;
        RECT 513.200 72.300 514.000 72.400 ;
        RECT 511.700 71.700 514.000 72.300 ;
        RECT 511.700 66.400 512.300 71.700 ;
        RECT 513.200 71.600 514.000 71.700 ;
        RECT 518.000 71.600 518.800 72.400 ;
        RECT 516.400 69.600 517.200 70.400 ;
        RECT 511.600 65.600 512.400 66.400 ;
        RECT 510.000 53.600 510.800 54.400 ;
        RECT 514.800 52.300 515.600 52.400 ;
        RECT 516.500 52.300 517.100 69.600 ;
        RECT 518.100 68.400 518.700 71.600 ;
        RECT 518.000 67.600 518.800 68.400 ;
        RECT 518.100 56.400 518.700 67.600 ;
        RECT 521.200 63.600 522.000 64.400 ;
        RECT 518.000 55.600 518.800 56.400 ;
        RECT 519.600 55.600 520.400 56.400 ;
        RECT 514.800 51.700 517.100 52.300 ;
        RECT 514.800 51.600 515.600 51.700 ;
        RECT 508.400 49.600 509.200 50.400 ;
        RECT 511.600 49.600 512.400 50.400 ;
        RECT 511.700 48.400 512.300 49.600 ;
        RECT 506.800 47.600 507.600 48.400 ;
        RECT 511.600 47.600 512.400 48.400 ;
        RECT 514.900 46.400 515.500 51.600 ;
        RECT 514.800 45.600 515.600 46.400 ;
        RECT 514.800 43.600 515.600 44.400 ;
        RECT 513.200 39.600 514.000 40.400 ;
        RECT 505.200 33.600 506.000 34.400 ;
        RECT 503.600 29.600 504.400 30.400 ;
        RECT 505.200 29.600 506.000 30.400 ;
        RECT 503.600 27.600 504.400 28.400 ;
        RECT 489.200 25.600 490.000 26.400 ;
        RECT 498.800 25.600 499.600 26.400 ;
        RECT 503.700 18.400 504.300 27.600 ;
        RECT 487.600 13.600 488.400 14.400 ;
        RECT 489.200 6.200 490.000 17.800 ;
        RECT 490.800 4.200 491.600 17.800 ;
        RECT 492.400 4.200 493.200 17.800 ;
        RECT 503.600 17.600 504.400 18.400 ;
        RECT 505.300 12.400 505.900 29.600 ;
        RECT 506.800 24.200 507.600 37.800 ;
        RECT 508.400 24.200 509.200 37.800 ;
        RECT 510.000 24.200 510.800 37.800 ;
        RECT 511.600 24.200 512.400 35.800 ;
        RECT 513.300 26.400 513.900 39.600 ;
        RECT 514.900 38.400 515.500 43.600 ;
        RECT 521.300 40.400 521.900 63.600 ;
        RECT 526.100 58.400 526.700 89.600 ;
        RECT 527.700 88.400 528.300 89.600 ;
        RECT 527.600 87.600 528.400 88.400 ;
        RECT 532.500 68.400 533.100 107.600 ;
        RECT 535.600 95.600 536.400 96.400 ;
        RECT 535.600 91.600 536.400 92.400 ;
        RECT 535.700 90.400 536.300 91.600 ;
        RECT 537.300 90.400 537.900 109.600 ;
        RECT 535.600 89.600 536.400 90.400 ;
        RECT 537.200 89.600 538.000 90.400 ;
        RECT 532.400 67.600 533.200 68.400 ;
        RECT 534.000 66.200 534.800 71.800 ;
        RECT 535.600 69.600 536.400 70.400 ;
        RECT 535.700 58.400 536.300 69.600 ;
        RECT 537.200 64.200 538.000 75.800 ;
        RECT 538.900 72.400 539.500 145.600 ;
        RECT 546.800 143.600 547.600 144.400 ;
        RECT 546.900 138.400 547.500 143.600 ;
        RECT 548.400 139.600 549.200 140.400 ;
        RECT 546.800 137.600 547.600 138.400 ;
        RECT 540.400 135.600 541.200 136.400 ;
        RECT 543.600 133.600 544.400 134.400 ;
        RECT 545.200 131.600 546.000 132.400 ;
        RECT 546.800 131.600 547.600 132.400 ;
        RECT 540.400 129.600 541.200 130.400 ;
        RECT 538.800 71.600 539.600 72.400 ;
        RECT 540.500 72.300 541.100 129.600 ;
        RECT 542.000 111.600 542.800 112.400 ;
        RECT 543.600 111.600 544.400 112.400 ;
        RECT 542.100 110.400 542.700 111.600 ;
        RECT 542.000 109.600 542.800 110.400 ;
        RECT 545.300 108.400 545.900 131.600 ;
        RECT 546.800 109.600 547.600 110.400 ;
        RECT 542.000 107.600 542.800 108.400 ;
        RECT 545.200 107.600 546.000 108.400 ;
        RECT 546.900 104.400 547.500 109.600 ;
        RECT 548.500 108.400 549.100 139.600 ;
        RECT 550.100 132.400 550.700 147.600 ;
        RECT 551.600 143.600 552.400 144.400 ;
        RECT 550.000 131.600 550.800 132.400 ;
        RECT 550.000 129.600 550.800 130.400 ;
        RECT 550.100 128.400 550.700 129.600 ;
        RECT 550.000 127.600 550.800 128.400 ;
        RECT 550.100 114.400 550.700 127.600 ;
        RECT 551.700 120.400 552.300 143.600 ;
        RECT 553.300 140.400 553.900 163.600 ;
        RECT 558.100 158.400 558.700 185.600 ;
        RECT 562.900 184.400 563.500 189.700 ;
        RECT 564.400 189.600 565.200 189.700 ;
        RECT 562.800 183.600 563.600 184.400 ;
        RECT 562.900 174.400 563.500 183.600 ;
        RECT 561.200 173.600 562.000 174.400 ;
        RECT 562.800 173.600 563.600 174.400 ;
        RECT 559.600 171.600 560.400 172.400 ;
        RECT 561.300 160.400 561.900 173.600 ;
        RECT 566.100 172.400 566.700 211.600 ;
        RECT 567.700 210.400 568.300 227.600 ;
        RECT 586.800 224.200 587.600 237.800 ;
        RECT 588.400 224.200 589.200 237.800 ;
        RECT 590.000 224.200 590.800 237.800 ;
        RECT 591.600 224.200 592.400 235.800 ;
        RECT 593.200 225.600 594.000 226.400 ;
        RECT 593.300 224.400 593.900 225.600 ;
        RECT 593.200 223.600 594.000 224.400 ;
        RECT 594.800 224.200 595.600 235.800 ;
        RECT 596.400 227.600 597.200 228.400 ;
        RECT 596.500 222.400 597.100 227.600 ;
        RECT 598.000 224.200 598.800 235.800 ;
        RECT 599.600 224.200 600.400 237.800 ;
        RECT 601.200 224.200 602.000 237.800 ;
        RECT 610.800 237.600 611.600 238.400 ;
        RECT 607.600 229.600 608.400 230.400 ;
        RECT 615.600 224.200 616.400 235.800 ;
        RECT 618.900 230.400 619.500 253.600 ;
        RECT 620.400 250.200 621.200 255.800 ;
        RECT 626.800 246.200 627.600 257.800 ;
        RECT 630.100 254.400 630.700 265.600 ;
        RECT 631.600 263.600 632.400 264.400 ;
        RECT 628.400 253.600 629.200 254.400 ;
        RECT 630.000 253.600 630.800 254.400 ;
        RECT 628.500 252.400 629.100 253.600 ;
        RECT 628.400 251.600 629.200 252.400 ;
        RECT 630.100 238.400 630.700 253.600 ;
        RECT 631.700 250.400 632.300 263.600 ;
        RECT 634.900 256.400 635.500 269.600 ;
        RECT 636.500 268.400 637.100 269.600 ;
        RECT 636.400 267.600 637.200 268.400 ;
        RECT 641.200 267.600 642.000 268.400 ;
        RECT 641.300 260.400 641.900 267.600 ;
        RECT 642.900 264.400 643.500 271.600 ;
        RECT 644.500 270.400 645.100 293.600 ;
        RECT 646.100 292.400 646.700 293.600 ;
        RECT 646.000 291.600 646.800 292.400 ;
        RECT 652.400 287.600 653.200 288.400 ;
        RECT 650.800 281.600 651.600 282.400 ;
        RECT 646.000 273.600 646.800 274.400 ;
        RECT 646.000 271.600 646.800 272.400 ;
        RECT 649.200 271.600 650.000 272.400 ;
        RECT 646.100 270.400 646.700 271.600 ;
        RECT 649.300 270.400 649.900 271.600 ;
        RECT 644.400 269.600 645.200 270.400 ;
        RECT 646.000 269.600 646.800 270.400 ;
        RECT 649.200 269.600 650.000 270.400 ;
        RECT 644.500 268.400 645.100 269.600 ;
        RECT 644.400 267.600 645.200 268.400 ;
        RECT 642.800 263.600 643.600 264.400 ;
        RECT 641.200 259.600 642.000 260.400 ;
        RECT 642.900 258.400 643.500 263.600 ;
        RECT 634.800 255.600 635.600 256.400 ;
        RECT 633.200 251.600 634.000 252.400 ;
        RECT 631.600 249.600 632.400 250.400 ;
        RECT 636.400 246.200 637.200 257.800 ;
        RECT 642.800 257.600 643.600 258.400 ;
        RECT 639.600 250.200 640.400 255.800 ;
        RECT 641.200 253.600 642.000 254.400 ;
        RECT 644.500 254.300 645.100 267.600 ;
        RECT 646.000 254.300 646.800 254.400 ;
        RECT 644.500 253.700 646.800 254.300 ;
        RECT 646.000 253.600 646.800 253.700 ;
        RECT 641.300 250.400 641.900 253.600 ;
        RECT 644.400 251.600 645.200 252.400 ;
        RECT 646.000 251.600 646.800 252.400 ;
        RECT 641.200 249.600 642.000 250.400 ;
        RECT 644.400 247.600 645.200 248.400 ;
        RECT 630.000 237.600 630.800 238.400 ;
        RECT 623.600 231.600 624.400 232.400 ;
        RECT 618.800 229.600 619.600 230.400 ;
        RECT 620.400 229.600 621.200 230.400 ;
        RECT 623.700 230.200 624.300 231.600 ;
        RECT 586.800 221.600 587.600 222.400 ;
        RECT 596.400 221.600 597.200 222.400 ;
        RECT 586.900 218.400 587.500 221.600 ;
        RECT 580.400 217.600 581.200 218.400 ;
        RECT 586.800 217.600 587.600 218.400 ;
        RECT 578.800 215.600 579.600 216.400 ;
        RECT 577.200 213.600 578.000 214.400 ;
        RECT 578.900 212.400 579.500 215.600 ;
        RECT 580.500 214.400 581.100 217.600 ;
        RECT 582.200 215.600 583.000 215.800 ;
        RECT 582.200 215.000 587.800 215.600 ;
        RECT 588.400 215.000 589.200 215.800 ;
        RECT 580.400 213.600 581.200 214.400 ;
        RECT 569.200 211.600 570.000 212.400 ;
        RECT 578.800 211.600 579.600 212.400 ;
        RECT 578.900 210.400 579.500 211.600 ;
        RECT 567.600 209.600 568.400 210.400 ;
        RECT 578.800 209.600 579.600 210.400 ;
        RECT 582.200 210.200 582.800 215.000 ;
        RECT 583.600 214.800 584.400 215.000 ;
        RECT 587.000 214.800 587.800 215.000 ;
        RECT 588.600 214.200 589.200 215.000 ;
        RECT 583.600 213.600 589.200 214.200 ;
        RECT 590.000 213.600 590.800 214.400 ;
        RECT 599.600 213.600 600.400 214.400 ;
        RECT 607.600 213.600 608.400 214.400 ;
        RECT 610.800 213.600 611.600 214.400 ;
        RECT 583.600 212.200 584.200 213.600 ;
        RECT 583.400 211.400 584.200 212.200 ;
        RECT 588.600 210.200 589.200 213.600 ;
        RECT 607.700 212.400 608.300 213.600 ;
        RECT 620.500 212.400 621.100 229.600 ;
        RECT 623.600 229.400 624.400 230.200 ;
        RECT 625.200 224.200 626.000 235.800 ;
        RECT 626.800 227.600 627.600 228.400 ;
        RECT 626.900 224.400 627.500 227.600 ;
        RECT 628.400 226.200 629.200 231.800 ;
        RECT 633.200 229.600 634.000 230.400 ;
        RECT 626.800 223.600 627.600 224.400 ;
        RECT 628.400 223.600 629.200 224.400 ;
        RECT 638.000 224.200 638.800 237.800 ;
        RECT 639.600 224.200 640.400 237.800 ;
        RECT 641.200 224.200 642.000 235.800 ;
        RECT 642.800 227.600 643.600 228.400 ;
        RECT 590.000 211.600 590.800 212.400 ;
        RECT 593.200 211.600 594.000 212.400 ;
        RECT 598.000 211.600 598.800 212.400 ;
        RECT 601.200 211.600 602.000 212.400 ;
        RECT 602.800 211.600 603.600 212.400 ;
        RECT 607.600 211.600 608.400 212.400 ;
        RECT 612.200 211.600 613.200 212.400 ;
        RECT 620.400 211.600 621.200 212.400 ;
        RECT 582.200 209.400 583.000 210.200 ;
        RECT 588.400 209.400 589.200 210.200 ;
        RECT 582.000 195.600 582.800 196.400 ;
        RECT 578.800 193.600 579.600 194.400 ;
        RECT 575.600 191.600 576.400 192.400 ;
        RECT 575.700 190.400 576.300 191.600 ;
        RECT 582.100 190.400 582.700 195.600 ;
        RECT 567.600 189.600 568.400 190.400 ;
        RECT 575.600 189.600 576.400 190.400 ;
        RECT 577.200 189.600 578.000 190.400 ;
        RECT 582.000 189.600 582.800 190.400 ;
        RECT 586.800 189.600 587.600 190.400 ;
        RECT 588.400 189.600 589.200 190.400 ;
        RECT 566.000 171.600 566.800 172.400 ;
        RECT 562.800 169.600 563.600 170.400 ;
        RECT 566.000 169.600 566.800 170.400 ;
        RECT 561.200 159.600 562.000 160.400 ;
        RECT 558.000 157.600 558.800 158.400 ;
        RECT 558.000 155.600 558.800 156.400 ;
        RECT 556.400 147.600 557.200 148.400 ;
        RECT 554.800 145.600 555.600 146.400 ;
        RECT 553.200 139.600 554.000 140.400 ;
        RECT 553.200 135.600 554.000 136.400 ;
        RECT 553.300 132.400 553.900 135.600 ;
        RECT 554.900 134.400 555.500 145.600 ;
        RECT 556.500 136.400 557.100 147.600 ;
        RECT 556.400 135.600 557.200 136.400 ;
        RECT 554.800 133.600 555.600 134.400 ;
        RECT 553.200 131.600 554.000 132.400 ;
        RECT 556.500 128.400 557.100 135.600 ;
        RECT 556.400 127.600 557.200 128.400 ;
        RECT 558.100 126.300 558.700 155.600 ;
        RECT 562.900 152.400 563.500 169.600 ;
        RECT 564.400 163.600 565.200 164.400 ;
        RECT 564.500 152.400 565.100 163.600 ;
        RECT 562.800 151.600 563.600 152.400 ;
        RECT 564.400 151.600 565.200 152.400 ;
        RECT 561.200 149.600 562.000 150.400 ;
        RECT 562.800 149.600 563.600 150.400 ;
        RECT 561.300 138.400 561.900 149.600 ;
        RECT 561.200 137.600 562.000 138.400 ;
        RECT 559.600 131.600 560.400 132.400 ;
        RECT 556.500 125.700 558.700 126.300 ;
        RECT 551.600 119.600 552.400 120.400 ;
        RECT 550.000 113.600 550.800 114.400 ;
        RECT 550.100 108.400 550.700 113.600 ;
        RECT 551.600 111.600 552.400 112.400 ;
        RECT 553.200 111.600 554.000 112.400 ;
        RECT 556.500 110.400 557.100 125.700 ;
        RECT 558.000 123.600 558.800 124.400 ;
        RECT 558.100 116.400 558.700 123.600 ;
        RECT 558.000 115.600 558.800 116.400 ;
        RECT 558.100 112.400 558.700 115.600 ;
        RECT 558.000 111.600 558.800 112.400 ;
        RECT 556.400 109.600 557.200 110.400 ;
        RECT 548.400 107.600 549.200 108.400 ;
        RECT 550.000 107.600 550.800 108.400 ;
        RECT 553.200 107.600 554.000 108.400 ;
        RECT 554.800 107.600 555.600 108.400 ;
        RECT 546.800 103.600 547.600 104.400 ;
        RECT 542.000 93.600 542.800 94.400 ;
        RECT 542.100 76.400 542.700 93.600 ;
        RECT 546.900 92.400 547.500 103.600 ;
        RECT 548.400 101.600 549.200 102.400 ;
        RECT 546.800 91.600 547.600 92.400 ;
        RECT 543.600 89.600 544.400 90.400 ;
        RECT 542.000 75.600 542.800 76.400 ;
        RECT 543.700 72.400 544.300 89.600 ;
        RECT 540.500 71.700 542.700 72.300 ;
        RECT 538.800 69.400 539.600 70.400 ;
        RECT 540.400 69.600 541.200 70.400 ;
        RECT 526.000 57.600 526.800 58.400 ;
        RECT 535.600 57.600 536.400 58.400 ;
        RECT 540.500 56.400 541.100 69.600 ;
        RECT 542.100 68.400 542.700 71.700 ;
        RECT 543.600 71.600 544.400 72.400 ;
        RECT 542.000 67.600 542.800 68.400 ;
        RECT 542.000 63.600 542.800 64.400 ;
        RECT 546.800 64.200 547.600 75.800 ;
        RECT 529.200 55.600 530.000 56.400 ;
        RECT 540.400 55.600 541.200 56.400 ;
        RECT 529.300 54.400 529.900 55.600 ;
        RECT 540.500 54.400 541.100 55.600 ;
        RECT 524.400 53.600 525.200 54.400 ;
        RECT 529.200 53.600 530.000 54.400 ;
        RECT 538.800 53.600 539.600 54.400 ;
        RECT 540.400 53.600 541.200 54.400 ;
        RECT 522.800 51.600 523.600 52.400 ;
        RECT 521.200 39.600 522.000 40.400 ;
        RECT 514.800 37.600 515.600 38.400 ;
        RECT 513.200 25.600 514.000 26.400 ;
        RECT 513.300 20.400 513.900 25.600 ;
        RECT 514.800 24.200 515.600 35.800 ;
        RECT 516.400 29.600 517.200 30.400 ;
        RECT 516.500 28.400 517.100 29.600 ;
        RECT 516.400 27.600 517.200 28.400 ;
        RECT 518.000 24.200 518.800 35.800 ;
        RECT 519.600 24.200 520.400 37.800 ;
        RECT 521.200 24.200 522.000 37.800 ;
        RECT 524.500 32.400 525.100 53.600 ;
        RECT 538.900 52.400 539.500 53.600 ;
        RECT 542.100 52.400 542.700 63.600 ;
        RECT 543.600 53.600 544.400 54.400 ;
        RECT 548.500 52.400 549.100 101.600 ;
        RECT 551.600 95.600 552.400 96.400 ;
        RECT 551.700 92.400 552.300 95.600 ;
        RECT 551.600 91.600 552.400 92.400 ;
        RECT 553.200 89.600 554.000 90.400 ;
        RECT 553.200 87.600 554.000 88.400 ;
        RECT 553.300 78.400 553.900 87.600 ;
        RECT 553.200 77.600 554.000 78.400 ;
        RECT 554.900 74.400 555.500 107.600 ;
        RECT 556.500 102.400 557.100 109.600 ;
        RECT 559.700 108.400 560.300 131.600 ;
        RECT 561.200 130.200 562.000 135.800 ;
        RECT 564.400 126.200 565.200 137.800 ;
        RECT 564.400 123.600 565.200 124.400 ;
        RECT 561.200 113.600 562.000 114.400 ;
        RECT 561.300 110.400 561.900 113.600 ;
        RECT 562.800 111.600 563.600 112.400 ;
        RECT 562.900 110.400 563.500 111.600 ;
        RECT 564.500 110.400 565.100 123.600 ;
        RECT 566.100 116.400 566.700 169.600 ;
        RECT 567.700 150.400 568.300 189.600 ;
        RECT 569.200 187.600 570.000 188.400 ;
        RECT 567.600 149.600 568.400 150.400 ;
        RECT 569.300 148.400 569.900 187.600 ;
        RECT 582.100 184.400 582.700 189.600 ;
        RECT 585.200 187.600 586.000 188.400 ;
        RECT 585.300 186.400 585.900 187.600 ;
        RECT 585.200 185.600 586.000 186.400 ;
        RECT 582.000 183.600 582.800 184.400 ;
        RECT 586.900 178.400 587.500 189.600 ;
        RECT 590.100 186.400 590.700 211.600 ;
        RECT 593.300 210.400 593.900 211.600 ;
        RECT 593.200 209.600 594.000 210.400 ;
        RECT 591.600 191.600 592.400 192.400 ;
        RECT 590.000 185.600 590.800 186.400 ;
        RECT 591.700 184.400 592.300 191.600 ;
        RECT 591.600 183.600 592.400 184.400 ;
        RECT 577.200 177.600 578.000 178.400 ;
        RECT 586.800 177.600 587.600 178.400 ;
        RECT 591.600 177.600 592.400 178.400 ;
        RECT 578.800 175.600 579.600 176.400 ;
        RECT 578.900 172.400 579.500 175.600 ;
        RECT 570.800 171.600 571.600 172.400 ;
        RECT 574.000 171.600 574.800 172.400 ;
        RECT 578.800 171.600 579.600 172.400 ;
        RECT 580.400 171.600 581.200 172.400 ;
        RECT 582.000 171.600 582.800 172.400 ;
        RECT 585.200 171.600 586.000 172.400 ;
        RECT 567.600 147.600 568.400 148.400 ;
        RECT 569.200 147.600 570.000 148.400 ;
        RECT 567.700 144.400 568.300 147.600 ;
        RECT 567.600 143.600 568.400 144.400 ;
        RECT 570.900 144.300 571.500 171.600 ;
        RECT 574.100 156.400 574.700 171.600 ;
        RECT 580.500 166.400 581.100 171.600 ;
        RECT 582.000 169.600 582.800 170.400 ;
        RECT 580.400 165.600 581.200 166.400 ;
        RECT 582.000 163.600 582.800 164.400 ;
        RECT 577.200 161.600 578.000 162.400 ;
        RECT 574.000 155.600 574.800 156.400 ;
        RECT 574.000 151.600 574.800 152.400 ;
        RECT 577.300 150.400 577.900 161.600 ;
        RECT 578.800 155.600 579.600 156.400 ;
        RECT 577.200 149.600 578.000 150.400 ;
        RECT 577.300 146.300 577.900 149.600 ;
        RECT 578.900 148.400 579.500 155.600 ;
        RECT 582.100 150.400 582.700 163.600 ;
        RECT 585.300 162.400 585.900 171.600 ;
        RECT 591.700 170.400 592.300 177.600 ;
        RECT 591.600 169.600 592.400 170.400 ;
        RECT 585.200 161.600 586.000 162.400 ;
        RECT 593.300 160.400 593.900 209.600 ;
        RECT 601.300 208.400 601.900 211.600 ;
        RECT 602.900 210.400 603.500 211.600 ;
        RECT 602.800 209.600 603.600 210.400 ;
        RECT 601.200 207.600 602.000 208.400 ;
        RECT 622.000 204.200 622.800 217.800 ;
        RECT 623.600 204.200 624.400 217.800 ;
        RECT 625.200 204.200 626.000 217.800 ;
        RECT 626.800 206.200 627.600 217.800 ;
        RECT 628.500 216.400 629.100 223.600 ;
        RECT 642.900 222.400 643.500 227.600 ;
        RECT 644.400 224.200 645.200 235.800 ;
        RECT 646.100 232.400 646.700 251.600 ;
        RECT 647.600 249.600 648.400 250.400 ;
        RECT 647.700 248.400 648.300 249.600 ;
        RECT 647.600 247.600 648.400 248.400 ;
        RECT 650.900 240.400 651.500 281.600 ;
        RECT 652.500 270.400 653.100 287.600 ;
        RECT 655.600 286.200 656.400 297.800 ;
        RECT 657.300 294.400 657.900 309.600 ;
        RECT 657.200 293.600 658.000 294.400 ;
        RECT 658.900 282.400 659.500 373.600 ;
        RECT 663.600 364.200 664.400 377.800 ;
        RECT 665.200 364.200 666.000 377.800 ;
        RECT 666.800 364.200 667.600 377.800 ;
        RECT 668.400 366.200 669.200 377.800 ;
        RECT 670.100 376.400 670.700 379.600 ;
        RECT 670.000 375.600 670.800 376.400 ;
        RECT 670.100 360.400 670.700 375.600 ;
        RECT 671.600 366.200 672.400 377.800 ;
        RECT 673.200 373.600 674.000 374.400 ;
        RECT 674.800 366.200 675.600 377.800 ;
        RECT 676.400 364.200 677.200 377.800 ;
        RECT 678.000 364.200 678.800 377.800 ;
        RECT 679.700 374.300 680.300 411.600 ;
        RECT 681.300 400.400 681.900 443.600 ;
        RECT 681.200 399.600 682.000 400.400 ;
        RECT 681.200 397.600 682.000 398.400 ;
        RECT 679.700 373.700 681.900 374.300 ;
        RECT 681.300 372.400 681.900 373.700 ;
        RECT 681.200 371.600 682.000 372.400 ;
        RECT 679.600 361.600 680.400 362.400 ;
        RECT 666.800 359.600 667.600 360.400 ;
        RECT 670.000 359.600 670.800 360.400 ;
        RECT 660.400 349.600 661.200 350.400 ;
        RECT 662.000 349.600 662.800 350.400 ;
        RECT 660.500 314.400 661.100 349.600 ;
        RECT 662.100 348.400 662.700 349.600 ;
        RECT 662.000 347.600 662.800 348.400 ;
        RECT 665.200 344.200 666.000 355.800 ;
        RECT 666.900 348.400 667.500 359.600 ;
        RECT 666.800 347.600 667.600 348.400 ;
        RECT 666.900 334.400 667.500 347.600 ;
        RECT 668.400 346.200 669.200 351.800 ;
        RECT 670.000 349.600 670.800 350.400 ;
        RECT 673.200 349.600 674.000 350.400 ;
        RECT 670.100 344.300 670.700 349.600 ;
        RECT 673.300 346.400 673.900 349.600 ;
        RECT 679.700 346.400 680.300 361.600 ;
        RECT 673.200 345.600 674.000 346.400 ;
        RECT 678.000 345.600 678.800 346.400 ;
        RECT 679.600 345.600 680.400 346.400 ;
        RECT 668.500 343.700 670.700 344.300 ;
        RECT 668.500 334.400 669.100 343.700 ;
        RECT 671.600 343.600 672.400 344.400 ;
        RECT 676.400 343.600 677.200 344.400 ;
        RECT 671.700 336.400 672.300 343.600 ;
        RECT 676.500 342.400 677.100 343.600 ;
        RECT 676.400 341.600 677.200 342.400 ;
        RECT 666.800 333.600 667.600 334.400 ;
        RECT 668.400 333.600 669.200 334.400 ;
        RECT 662.000 331.600 662.800 332.400 ;
        RECT 666.800 331.600 667.600 332.400 ;
        RECT 662.100 330.400 662.700 331.600 ;
        RECT 662.000 329.600 662.800 330.400 ;
        RECT 663.600 329.600 664.400 330.400 ;
        RECT 663.700 328.400 664.300 329.600 ;
        RECT 663.600 327.600 664.400 328.400 ;
        RECT 666.800 327.600 667.600 328.400 ;
        RECT 668.500 326.400 669.100 333.600 ;
        RECT 670.000 330.200 670.800 335.800 ;
        RECT 671.600 335.600 672.400 336.400 ;
        RECT 671.600 333.600 672.400 334.400 ;
        RECT 666.800 325.600 667.600 326.400 ;
        RECT 668.400 325.600 669.200 326.400 ;
        RECT 673.200 326.200 674.000 337.800 ;
        RECT 674.800 331.800 675.600 332.600 ;
        RECT 674.900 328.400 675.500 331.800 ;
        RECT 674.800 327.600 675.600 328.400 ;
        RECT 662.000 317.600 662.800 318.400 ;
        RECT 660.400 313.600 661.200 314.400 ;
        RECT 660.400 311.600 661.200 312.400 ;
        RECT 662.100 292.400 662.700 317.600 ;
        RECT 663.600 309.600 664.400 310.400 ;
        RECT 665.200 309.600 666.000 310.400 ;
        RECT 665.300 308.400 665.900 309.600 ;
        RECT 666.900 308.400 667.500 325.600 ;
        RECT 676.400 319.600 677.200 320.400 ;
        RECT 665.200 307.600 666.000 308.400 ;
        RECT 666.800 307.600 667.600 308.400 ;
        RECT 668.400 306.200 669.200 311.800 ;
        RECT 671.600 304.200 672.400 315.800 ;
        RECT 673.200 309.400 674.000 310.400 ;
        RECT 676.500 308.400 677.100 319.600 ;
        RECT 676.400 307.600 677.200 308.400 ;
        RECT 676.500 302.400 677.100 307.600 ;
        RECT 666.800 301.600 667.600 302.400 ;
        RECT 673.200 301.600 674.000 302.400 ;
        RECT 676.400 301.600 677.200 302.400 ;
        RECT 662.000 291.600 662.800 292.400 ;
        RECT 665.200 286.200 666.000 297.800 ;
        RECT 666.900 294.400 667.500 301.600 ;
        RECT 666.800 293.600 667.600 294.400 ;
        RECT 668.400 290.200 669.200 295.800 ;
        RECT 670.000 293.600 670.800 294.400 ;
        RECT 658.800 281.600 659.600 282.400 ;
        RECT 658.800 279.600 659.600 280.400 ;
        RECT 657.200 275.600 658.000 276.400 ;
        RECT 654.000 271.600 654.800 272.400 ;
        RECT 657.300 270.400 657.900 275.600 ;
        RECT 658.900 270.400 659.500 279.600 ;
        RECT 666.800 275.600 667.600 276.400 ;
        RECT 660.400 273.600 661.200 274.400 ;
        RECT 663.600 273.600 664.400 274.400 ;
        RECT 660.500 272.400 661.100 273.600 ;
        RECT 660.400 271.600 661.200 272.400 ;
        RECT 663.600 271.600 664.400 272.400 ;
        RECT 663.700 270.400 664.300 271.600 ;
        RECT 652.400 269.600 653.200 270.400 ;
        RECT 657.200 269.600 658.000 270.400 ;
        RECT 658.800 269.600 659.600 270.400 ;
        RECT 663.600 269.600 664.400 270.400 ;
        RECT 666.800 269.600 667.600 270.400 ;
        RECT 652.400 267.600 653.200 268.400 ;
        RECT 652.500 254.400 653.100 267.600 ;
        RECT 658.900 256.400 659.500 269.600 ;
        RECT 663.600 267.600 664.400 268.400 ;
        RECT 665.200 267.600 666.000 268.400 ;
        RECT 660.400 257.600 661.200 258.400 ;
        RECT 655.600 255.600 656.400 256.400 ;
        RECT 658.800 255.600 659.600 256.400 ;
        RECT 652.400 253.600 653.200 254.400 ;
        RECT 655.700 252.400 656.300 255.600 ;
        RECT 658.800 253.600 659.600 254.400 ;
        RECT 652.400 251.600 653.200 252.400 ;
        RECT 655.600 251.600 656.400 252.400 ;
        RECT 657.200 251.600 658.000 252.400 ;
        RECT 652.500 250.400 653.100 251.600 ;
        RECT 652.400 249.600 653.200 250.400 ;
        RECT 650.800 239.600 651.600 240.400 ;
        RECT 646.000 231.600 646.800 232.400 ;
        RECT 646.000 225.600 646.800 226.400 ;
        RECT 646.100 224.400 646.700 225.600 ;
        RECT 646.000 223.600 646.800 224.400 ;
        RECT 647.600 224.200 648.400 235.800 ;
        RECT 649.200 224.200 650.000 237.800 ;
        RECT 650.800 224.200 651.600 237.800 ;
        RECT 652.400 224.200 653.200 237.800 ;
        RECT 642.800 221.600 643.600 222.400 ;
        RECT 649.200 221.600 650.000 222.400 ;
        RECT 649.300 218.400 649.900 221.600 ;
        RECT 628.400 215.600 629.200 216.400 ;
        RECT 630.000 206.200 630.800 217.800 ;
        RECT 631.600 213.600 632.400 214.400 ;
        RECT 633.200 206.200 634.000 217.800 ;
        RECT 634.800 204.200 635.600 217.800 ;
        RECT 636.400 204.200 637.200 217.800 ;
        RECT 649.200 217.600 650.000 218.400 ;
        RECT 647.400 215.000 648.200 215.800 ;
        RECT 649.200 215.000 653.400 215.600 ;
        RECT 654.000 215.000 654.800 215.800 ;
        RECT 655.600 215.600 656.400 216.400 ;
        RECT 646.000 213.600 646.800 214.400 ;
        RECT 642.800 211.600 643.600 212.400 ;
        RECT 598.000 191.600 598.800 192.400 ;
        RECT 594.800 189.600 595.600 190.400 ;
        RECT 594.900 172.400 595.500 189.600 ;
        RECT 596.400 187.600 597.200 188.400 ;
        RECT 598.100 186.400 598.700 191.600 ;
        RECT 598.000 185.600 598.800 186.400 ;
        RECT 598.000 183.600 598.800 184.400 ;
        RECT 602.800 184.200 603.600 195.800 ;
        RECT 609.200 189.600 610.000 190.400 ;
        RECT 607.600 187.600 608.400 188.400 ;
        RECT 594.800 171.600 595.600 172.400 ;
        RECT 594.900 164.400 595.500 171.600 ;
        RECT 596.400 166.200 597.200 177.800 ;
        RECT 598.100 176.400 598.700 183.600 ;
        RECT 598.000 175.600 598.800 176.400 ;
        RECT 604.400 171.800 605.200 172.600 ;
        RECT 604.500 168.400 605.100 171.800 ;
        RECT 604.400 167.600 605.200 168.400 ;
        RECT 602.800 165.600 603.600 166.400 ;
        RECT 606.000 166.200 606.800 177.800 ;
        RECT 607.700 174.400 608.300 187.600 ;
        RECT 612.400 184.200 613.200 195.800 ;
        RECT 636.400 195.600 637.200 196.400 ;
        RECT 622.000 193.600 622.800 194.400 ;
        RECT 631.600 193.600 632.400 194.400 ;
        RECT 622.100 192.400 622.700 193.600 ;
        RECT 615.600 186.200 616.400 191.800 ;
        RECT 620.400 191.600 621.200 192.400 ;
        RECT 622.000 191.600 622.800 192.400 ;
        RECT 628.400 191.600 629.200 192.400 ;
        RECT 630.000 191.600 630.800 192.400 ;
        RECT 620.500 190.400 621.100 191.600 ;
        RECT 618.800 189.600 619.600 190.400 ;
        RECT 620.400 189.600 621.200 190.400 ;
        RECT 617.200 187.600 618.000 188.400 ;
        RECT 615.600 183.600 616.400 184.400 ;
        RECT 612.400 181.600 613.200 182.400 ;
        RECT 612.500 176.400 613.100 181.600 ;
        RECT 607.600 173.600 608.400 174.400 ;
        RECT 609.200 170.200 610.000 175.800 ;
        RECT 612.400 175.600 613.200 176.400 ;
        RECT 614.000 175.600 614.800 176.400 ;
        RECT 614.100 174.400 614.700 175.600 ;
        RECT 614.000 173.600 614.800 174.400 ;
        RECT 615.700 172.400 616.300 183.600 ;
        RECT 617.300 176.400 617.900 187.600 ;
        RECT 618.900 184.400 619.500 189.600 ;
        RECT 618.800 183.600 619.600 184.400 ;
        RECT 622.100 182.400 622.700 191.600 ;
        RECT 630.100 190.400 630.700 191.600 ;
        RECT 631.700 190.400 632.300 193.600 ;
        RECT 636.500 190.400 637.100 195.600 ;
        RECT 639.600 193.600 640.400 194.400 ;
        RECT 623.600 189.600 624.400 190.400 ;
        RECT 625.200 189.600 626.000 190.400 ;
        RECT 630.000 189.600 630.800 190.400 ;
        RECT 631.600 189.600 632.400 190.400 ;
        RECT 636.400 189.600 637.200 190.400 ;
        RECT 638.000 189.600 638.800 190.400 ;
        RECT 623.700 188.400 624.300 189.600 ;
        RECT 625.300 188.400 625.900 189.600 ;
        RECT 623.600 187.600 624.400 188.400 ;
        RECT 625.200 187.600 626.000 188.400 ;
        RECT 630.000 187.600 630.800 188.400 ;
        RECT 631.600 187.600 632.400 188.400 ;
        RECT 622.000 181.600 622.800 182.400 ;
        RECT 623.700 180.300 624.300 187.600 ;
        RECT 623.700 179.700 625.900 180.300 ;
        RECT 617.200 175.600 618.000 176.400 ;
        RECT 623.600 175.600 624.400 176.400 ;
        RECT 615.600 171.600 616.400 172.400 ;
        RECT 594.800 163.600 595.600 164.400 ;
        RECT 588.400 159.600 589.200 160.400 ;
        RECT 593.200 159.600 594.000 160.400 ;
        RECT 585.200 154.300 586.000 154.400 ;
        RECT 583.700 153.700 586.000 154.300 ;
        RECT 582.000 149.600 582.800 150.400 ;
        RECT 578.800 147.600 579.600 148.400 ;
        RECT 580.400 147.600 581.200 148.400 ;
        RECT 577.300 145.700 579.500 146.300 ;
        RECT 569.300 143.700 571.500 144.300 ;
        RECT 567.600 131.600 568.400 132.400 ;
        RECT 566.000 115.600 566.800 116.400 ;
        RECT 561.200 109.600 562.000 110.400 ;
        RECT 562.800 109.600 563.600 110.400 ;
        RECT 564.400 109.600 565.200 110.400 ;
        RECT 559.600 107.600 560.400 108.400 ;
        RECT 562.800 103.600 563.600 104.400 ;
        RECT 567.600 103.600 568.400 104.400 ;
        RECT 556.400 101.600 557.200 102.400 ;
        RECT 558.000 93.600 558.800 94.400 ;
        RECT 561.200 93.600 562.000 94.400 ;
        RECT 556.400 83.600 557.200 84.400 ;
        RECT 556.500 82.400 557.100 83.600 ;
        RECT 556.400 81.600 557.200 82.400 ;
        RECT 558.100 80.400 558.700 93.600 ;
        RECT 559.600 89.600 560.400 90.400 ;
        RECT 558.000 79.600 558.800 80.400 ;
        RECT 556.400 77.600 557.200 78.400 ;
        RECT 554.800 73.600 555.600 74.400 ;
        RECT 556.500 70.400 557.100 77.600 ;
        RECT 558.000 71.600 558.800 72.400 ;
        RECT 553.200 69.600 554.000 70.400 ;
        RECT 556.400 69.600 557.200 70.400 ;
        RECT 551.600 63.600 552.400 64.400 ;
        RECT 551.600 57.600 552.400 58.400 ;
        RECT 551.700 54.400 552.300 57.600 ;
        RECT 551.600 53.600 552.400 54.400 ;
        RECT 530.800 51.600 531.600 52.400 ;
        RECT 538.800 51.600 539.600 52.400 ;
        RECT 540.400 51.600 541.200 52.400 ;
        RECT 542.000 51.600 542.800 52.400 ;
        RECT 548.400 51.600 549.200 52.400 ;
        RECT 550.000 51.600 550.800 52.400 ;
        RECT 540.500 50.400 541.100 51.600 ;
        RECT 534.000 49.600 534.800 50.400 ;
        RECT 540.400 49.600 541.200 50.400 ;
        RECT 527.600 47.600 528.400 48.400 ;
        RECT 527.700 34.400 528.300 47.600 ;
        RECT 548.500 46.400 549.100 51.600 ;
        RECT 546.800 45.600 547.600 46.400 ;
        RECT 548.400 45.600 549.200 46.400 ;
        RECT 530.800 37.600 531.600 38.400 ;
        RECT 527.600 33.600 528.400 34.400 ;
        RECT 530.900 32.400 531.500 37.600 ;
        RECT 538.800 33.600 539.600 34.400 ;
        RECT 543.600 33.600 544.400 34.400 ;
        RECT 524.400 31.600 525.200 32.400 ;
        RECT 530.800 31.600 531.600 32.400 ;
        RECT 530.800 29.600 531.600 30.400 ;
        RECT 534.000 29.600 534.800 30.400 ;
        RECT 534.100 26.400 534.700 29.600 ;
        RECT 535.600 27.600 536.400 28.400 ;
        RECT 537.200 27.600 538.000 28.400 ;
        RECT 535.700 26.400 536.300 27.600 ;
        RECT 534.000 25.600 534.800 26.400 ;
        RECT 535.600 25.600 536.400 26.400 ;
        RECT 513.200 19.600 514.000 20.400 ;
        RECT 521.200 19.600 522.000 20.400 ;
        RECT 498.800 11.600 499.600 12.400 ;
        RECT 505.200 11.600 506.000 12.400 ;
        RECT 508.400 11.600 509.200 12.400 ;
        RECT 513.200 4.200 514.000 17.800 ;
        RECT 514.800 4.200 515.600 17.800 ;
        RECT 516.400 6.200 517.200 17.800 ;
        RECT 518.000 13.600 518.800 14.400 ;
        RECT 519.600 6.200 520.400 17.800 ;
        RECT 521.300 16.400 521.900 19.600 ;
        RECT 521.200 15.600 522.000 16.400 ;
        RECT 522.800 6.200 523.600 17.800 ;
        RECT 524.400 4.200 525.200 17.800 ;
        RECT 526.000 4.200 526.800 17.800 ;
        RECT 527.600 4.200 528.400 17.800 ;
        RECT 538.900 16.400 539.500 33.600 ;
        RECT 543.700 32.400 544.300 33.600 ;
        RECT 543.600 31.600 544.400 32.400 ;
        RECT 546.900 30.400 547.500 45.600 ;
        RECT 550.100 36.400 550.700 51.600 ;
        RECT 550.000 35.600 550.800 36.400 ;
        RECT 551.700 34.300 552.300 53.600 ;
        RECT 553.300 52.400 553.900 69.600 ;
        RECT 558.100 66.400 558.700 71.600 ;
        RECT 561.300 70.400 561.900 93.600 ;
        RECT 562.900 92.400 563.500 103.600 ;
        RECT 564.400 95.600 565.200 96.400 ;
        RECT 564.500 94.400 565.100 95.600 ;
        RECT 567.700 94.400 568.300 103.600 ;
        RECT 564.400 93.600 565.200 94.400 ;
        RECT 567.600 93.600 568.400 94.400 ;
        RECT 562.800 91.600 563.600 92.400 ;
        RECT 564.400 91.600 565.200 92.400 ;
        RECT 567.600 91.600 568.400 92.400 ;
        RECT 562.800 89.600 563.600 90.400 ;
        RECT 561.200 69.600 562.000 70.400 ;
        RECT 559.600 67.600 560.400 68.400 ;
        RECT 562.900 68.300 563.500 89.600 ;
        RECT 564.500 72.400 565.100 91.600 ;
        RECT 567.700 86.400 568.300 91.600 ;
        RECT 567.600 85.600 568.400 86.400 ;
        RECT 564.400 71.600 565.200 72.400 ;
        RECT 561.300 67.700 563.500 68.300 ;
        RECT 558.000 65.600 558.800 66.400 ;
        RECT 559.700 64.300 560.300 67.600 ;
        RECT 558.100 63.700 560.300 64.300 ;
        RECT 558.100 58.400 558.700 63.700 ;
        RECT 559.600 61.600 560.400 62.400 ;
        RECT 558.000 57.600 558.800 58.400 ;
        RECT 558.000 53.600 558.800 54.400 ;
        RECT 553.200 51.600 554.000 52.400 ;
        RECT 554.800 51.600 555.600 52.400 ;
        RECT 550.100 33.700 552.300 34.300 ;
        RECT 546.800 29.600 547.600 30.400 ;
        RECT 540.400 27.600 541.200 28.400 ;
        RECT 540.400 25.600 541.200 26.400 ;
        RECT 540.500 18.400 541.100 25.600 ;
        RECT 546.900 18.400 547.500 29.600 ;
        RECT 550.100 28.400 550.700 33.700 ;
        RECT 553.300 32.400 553.900 51.600 ;
        RECT 554.900 50.400 555.500 51.600 ;
        RECT 554.800 49.600 555.600 50.400 ;
        RECT 556.400 50.300 557.200 50.400 ;
        RECT 558.100 50.300 558.700 53.600 ;
        RECT 556.400 49.700 558.700 50.300 ;
        RECT 556.400 49.600 557.200 49.700 ;
        RECT 556.500 34.400 557.100 49.600 ;
        RECT 559.700 38.400 560.300 61.600 ;
        RECT 561.300 58.400 561.900 67.700 ;
        RECT 567.700 66.400 568.300 85.600 ;
        RECT 569.300 82.400 569.900 143.700 ;
        RECT 572.400 131.600 573.200 132.400 ;
        RECT 572.500 130.400 573.100 131.600 ;
        RECT 572.400 129.600 573.200 130.400 ;
        RECT 572.500 122.400 573.100 129.600 ;
        RECT 574.000 126.200 574.800 137.800 ;
        RECT 578.900 132.300 579.500 145.700 ;
        RECT 583.700 138.400 584.300 153.700 ;
        RECT 585.200 153.600 586.000 153.700 ;
        RECT 585.300 152.400 585.900 153.600 ;
        RECT 585.200 151.600 586.000 152.400 ;
        RECT 585.200 149.600 586.000 150.400 ;
        RECT 585.300 138.400 585.900 149.600 ;
        RECT 586.800 143.600 587.600 144.400 ;
        RECT 583.600 137.600 584.400 138.400 ;
        RECT 585.200 137.600 586.000 138.400 ;
        RECT 586.900 132.400 587.500 143.600 ;
        RECT 588.500 140.400 589.100 159.600 ;
        RECT 599.600 157.600 600.400 158.400 ;
        RECT 594.800 153.600 595.600 154.400 ;
        RECT 593.200 151.600 594.000 152.400 ;
        RECT 593.300 150.400 593.900 151.600 ;
        RECT 594.900 150.400 595.500 153.600 ;
        RECT 599.700 150.400 600.300 157.600 ;
        RECT 590.000 149.600 590.800 150.400 ;
        RECT 593.200 149.600 594.000 150.400 ;
        RECT 594.800 149.600 595.600 150.400 ;
        RECT 599.600 149.600 600.400 150.400 ;
        RECT 601.200 149.600 602.000 150.400 ;
        RECT 590.100 144.400 590.700 149.600 ;
        RECT 591.600 147.600 592.400 148.400 ;
        RECT 591.600 145.600 592.400 146.400 ;
        RECT 590.000 143.600 590.800 144.400 ;
        RECT 588.400 139.600 589.200 140.400 ;
        RECT 588.400 137.600 589.200 138.400 ;
        RECT 588.500 134.400 589.100 137.600 ;
        RECT 588.400 133.600 589.200 134.400 ;
        RECT 577.300 131.700 579.500 132.300 ;
        RECT 572.400 121.600 573.200 122.400 ;
        RECT 577.300 118.400 577.900 131.700 ;
        RECT 586.800 131.600 587.600 132.400 ;
        RECT 585.200 129.600 586.000 130.400 ;
        RECT 590.000 129.600 590.800 130.400 ;
        RECT 591.700 130.300 592.300 145.600 ;
        RECT 593.200 131.600 594.000 132.400 ;
        RECT 594.900 130.400 595.500 149.600 ;
        RECT 596.400 143.600 597.200 144.400 ;
        RECT 599.700 140.400 600.300 149.600 ;
        RECT 596.400 139.600 597.200 140.400 ;
        RECT 599.600 139.600 600.400 140.400 ;
        RECT 596.500 138.400 597.100 139.600 ;
        RECT 596.400 137.600 597.200 138.400 ;
        RECT 601.300 136.400 601.900 149.600 ;
        RECT 601.200 135.600 602.000 136.400 ;
        RECT 601.200 134.300 602.000 134.400 ;
        RECT 598.100 133.700 602.000 134.300 ;
        RECT 591.700 129.700 593.900 130.300 ;
        RECT 582.000 127.600 582.800 128.400 ;
        RECT 578.800 119.600 579.600 120.400 ;
        RECT 577.200 117.600 578.000 118.400 ;
        RECT 574.000 107.600 574.800 108.400 ;
        RECT 577.200 103.600 578.000 104.400 ;
        RECT 575.600 95.600 576.400 96.400 ;
        RECT 572.400 91.600 573.200 92.400 ;
        RECT 574.000 91.600 574.800 92.400 ;
        RECT 570.800 83.600 571.600 84.400 ;
        RECT 569.200 81.600 570.000 82.400 ;
        RECT 569.200 71.600 570.000 72.400 ;
        RECT 570.900 70.400 571.500 83.600 ;
        RECT 572.500 82.400 573.100 91.600 ;
        RECT 572.400 81.600 573.200 82.400 ;
        RECT 577.200 73.600 578.000 74.400 ;
        RECT 577.300 72.400 577.900 73.600 ;
        RECT 577.200 71.600 578.000 72.400 ;
        RECT 570.800 69.600 571.600 70.400 ;
        RECT 578.900 70.300 579.500 119.600 ;
        RECT 580.400 111.600 581.200 112.400 ;
        RECT 580.500 96.400 581.100 111.600 ;
        RECT 582.100 106.400 582.700 127.600 ;
        RECT 585.300 116.400 585.900 129.600 ;
        RECT 586.800 117.600 587.600 118.400 ;
        RECT 585.200 115.600 586.000 116.400 ;
        RECT 590.000 113.600 590.800 114.400 ;
        RECT 583.600 111.600 584.400 112.400 ;
        RECT 583.700 110.400 584.300 111.600 ;
        RECT 590.100 110.400 590.700 113.600 ;
        RECT 591.600 111.600 592.400 112.400 ;
        RECT 591.700 110.400 592.300 111.600 ;
        RECT 583.600 109.600 584.400 110.400 ;
        RECT 586.800 109.600 587.600 110.400 ;
        RECT 590.000 109.600 590.800 110.400 ;
        RECT 591.600 109.600 592.400 110.400 ;
        RECT 585.200 107.600 586.000 108.400 ;
        RECT 588.400 107.600 589.200 108.400 ;
        RECT 590.000 107.600 590.800 108.400 ;
        RECT 582.000 105.600 582.800 106.400 ;
        RECT 580.400 95.600 581.200 96.400 ;
        RECT 582.100 78.400 582.700 105.600 ;
        RECT 583.600 97.600 584.400 98.400 ;
        RECT 582.000 77.600 582.800 78.400 ;
        RECT 582.100 76.400 582.700 77.600 ;
        RECT 580.400 75.600 581.200 76.400 ;
        RECT 582.000 75.600 582.800 76.400 ;
        RECT 585.300 74.400 585.900 107.600 ;
        RECT 588.500 106.400 589.100 107.600 ;
        RECT 588.400 105.600 589.200 106.400 ;
        RECT 590.100 104.400 590.700 107.600 ;
        RECT 590.000 103.600 590.800 104.400 ;
        RECT 588.400 86.200 589.200 97.800 ;
        RECT 590.000 81.600 590.800 82.400 ;
        RECT 590.100 78.400 590.700 81.600 ;
        RECT 590.000 77.600 590.800 78.400 ;
        RECT 586.800 75.600 587.600 76.400 ;
        RECT 583.600 73.600 584.400 74.400 ;
        RECT 585.200 73.600 586.000 74.400 ;
        RECT 586.900 70.400 587.500 75.600 ;
        RECT 588.400 71.600 589.200 72.400 ;
        RECT 580.400 70.300 581.200 70.400 ;
        RECT 578.900 69.700 581.200 70.300 ;
        RECT 580.400 69.600 581.200 69.700 ;
        RECT 585.200 69.600 586.000 70.400 ;
        RECT 586.800 69.600 587.600 70.400 ;
        RECT 570.800 67.600 571.600 68.400 ;
        RECT 582.000 67.600 582.800 68.400 ;
        RECT 567.600 65.600 568.400 66.400 ;
        RECT 570.900 64.300 571.500 67.600 ;
        RECT 567.700 63.700 571.500 64.300 ;
        RECT 561.200 57.600 562.000 58.400 ;
        RECT 567.700 56.400 568.300 63.700 ;
        RECT 569.200 59.600 570.000 60.400 ;
        RECT 580.400 59.600 581.200 60.400 ;
        RECT 567.600 55.600 568.400 56.400 ;
        RECT 567.700 54.400 568.300 55.600 ;
        RECT 569.300 54.400 569.900 59.600 ;
        RECT 580.500 58.400 581.100 59.600 ;
        RECT 582.100 58.400 582.700 67.600 ;
        RECT 583.600 61.600 584.400 62.400 ;
        RECT 580.400 57.600 581.200 58.400 ;
        RECT 582.000 57.600 582.800 58.400 ;
        RECT 575.600 55.000 576.400 55.800 ;
        RECT 581.800 55.600 582.600 55.800 ;
        RECT 577.000 55.000 582.600 55.600 ;
        RECT 561.200 53.600 562.000 54.400 ;
        RECT 567.600 53.600 568.400 54.400 ;
        RECT 569.200 53.600 570.000 54.400 ;
        RECT 575.600 54.200 576.200 55.000 ;
        RECT 577.000 54.800 577.800 55.000 ;
        RECT 580.400 54.800 581.200 55.000 ;
        RECT 575.600 53.600 581.200 54.200 ;
        RECT 561.300 50.400 561.900 53.600 ;
        RECT 566.000 52.300 566.800 52.400 ;
        RECT 564.500 51.700 566.800 52.300 ;
        RECT 561.200 49.600 562.000 50.400 ;
        RECT 562.800 49.600 563.600 50.400 ;
        RECT 564.500 38.400 565.100 51.700 ;
        RECT 566.000 51.600 566.800 51.700 ;
        RECT 575.600 50.200 576.200 53.600 ;
        RECT 580.600 52.200 581.200 53.600 ;
        RECT 580.600 51.400 581.400 52.200 ;
        RECT 582.000 50.200 582.600 55.000 ;
        RECT 583.700 54.400 584.300 61.600 ;
        RECT 585.300 58.400 585.900 69.600 ;
        RECT 588.500 58.400 589.100 71.600 ;
        RECT 593.300 60.400 593.900 129.700 ;
        RECT 594.800 129.600 595.600 130.400 ;
        RECT 596.400 129.600 597.200 130.400 ;
        RECT 598.100 128.400 598.700 133.700 ;
        RECT 601.200 133.600 602.000 133.700 ;
        RECT 599.600 131.600 600.400 132.400 ;
        RECT 601.200 131.600 602.000 132.400 ;
        RECT 599.700 130.400 600.300 131.600 ;
        RECT 599.600 129.600 600.400 130.400 ;
        RECT 594.800 127.600 595.600 128.400 ;
        RECT 598.000 127.600 598.800 128.400 ;
        RECT 594.900 126.400 595.500 127.600 ;
        RECT 594.800 125.600 595.600 126.400 ;
        RECT 594.900 108.400 595.500 125.600 ;
        RECT 599.700 120.400 600.300 129.600 ;
        RECT 599.600 119.600 600.400 120.400 ;
        RECT 596.400 115.600 597.200 116.400 ;
        RECT 596.500 112.400 597.100 115.600 ;
        RECT 601.300 112.400 601.900 131.600 ;
        RECT 596.400 111.600 597.200 112.400 ;
        RECT 601.200 111.600 602.000 112.400 ;
        RECT 594.800 107.600 595.600 108.400 ;
        RECT 599.600 107.600 600.400 108.400 ;
        RECT 601.200 103.600 602.000 104.400 ;
        RECT 596.400 91.800 597.200 92.600 ;
        RECT 596.500 90.400 597.100 91.800 ;
        RECT 596.400 89.600 597.200 90.400 ;
        RECT 598.000 86.200 598.800 97.800 ;
        RECT 599.600 95.600 600.400 96.400 ;
        RECT 599.700 94.400 600.300 95.600 ;
        RECT 599.600 93.600 600.400 94.400 ;
        RECT 601.200 90.200 602.000 95.800 ;
        RECT 602.900 92.400 603.500 165.600 ;
        RECT 610.800 163.600 611.600 164.400 ;
        RECT 610.900 152.300 611.500 163.600 ;
        RECT 617.300 158.400 617.900 175.600 ;
        RECT 623.700 172.400 624.300 175.600 ;
        RECT 625.300 174.400 625.900 179.700 ;
        RECT 630.000 175.600 630.800 176.400 ;
        RECT 625.200 173.600 626.000 174.400 ;
        RECT 623.600 171.600 624.400 172.400 ;
        RECT 626.800 171.600 627.600 172.400 ;
        RECT 628.400 171.600 629.200 172.400 ;
        RECT 618.800 169.600 619.600 170.400 ;
        RECT 623.600 167.600 624.400 168.400 ;
        RECT 626.900 166.400 627.500 171.600 ;
        RECT 628.500 170.400 629.100 171.600 ;
        RECT 628.400 169.600 629.200 170.400 ;
        RECT 626.800 165.600 627.600 166.400 ;
        RECT 626.800 159.600 627.600 160.400 ;
        RECT 617.200 157.600 618.000 158.400 ;
        RECT 614.000 153.600 614.800 154.400 ;
        RECT 622.000 153.600 622.800 154.400 ;
        RECT 623.600 153.600 624.400 154.400 ;
        RECT 614.100 152.400 614.700 153.600 ;
        RECT 609.300 151.700 611.500 152.300 ;
        RECT 609.300 148.400 609.900 151.700 ;
        RECT 614.000 151.600 614.800 152.400 ;
        RECT 610.800 149.600 611.600 150.400 ;
        RECT 620.400 149.600 621.200 150.400 ;
        RECT 606.000 147.600 606.800 148.400 ;
        RECT 609.200 147.600 610.000 148.400 ;
        RECT 606.100 144.400 606.700 147.600 ;
        RECT 606.000 143.600 606.800 144.400 ;
        RECT 604.400 137.600 605.200 138.400 ;
        RECT 604.500 132.400 605.100 137.600 ;
        RECT 606.100 134.400 606.700 143.600 ;
        RECT 609.200 139.600 610.000 140.400 ;
        RECT 606.000 133.600 606.800 134.400 ;
        RECT 609.300 132.400 609.900 139.600 ;
        RECT 604.400 131.600 605.200 132.400 ;
        RECT 609.200 131.600 610.000 132.400 ;
        RECT 610.900 130.400 611.500 149.600 ;
        RECT 614.000 143.600 614.800 144.400 ;
        RECT 617.200 143.600 618.000 144.400 ;
        RECT 614.100 142.400 614.700 143.600 ;
        RECT 614.000 141.600 614.800 142.400 ;
        RECT 617.300 136.300 617.900 143.600 ;
        RECT 617.300 135.700 619.500 136.300 ;
        RECT 618.900 134.400 619.500 135.700 ;
        RECT 612.400 133.600 613.200 134.400 ;
        RECT 617.200 133.600 618.000 134.400 ;
        RECT 618.800 133.600 619.600 134.400 ;
        RECT 620.400 131.600 621.200 132.400 ;
        RECT 610.800 129.600 611.600 130.400 ;
        RECT 617.200 129.600 618.000 130.400 ;
        RECT 620.400 129.600 621.200 130.400 ;
        RECT 604.400 115.600 605.200 116.400 ;
        RECT 607.600 113.600 608.400 114.400 ;
        RECT 604.400 97.600 605.200 98.400 ;
        RECT 604.500 92.400 605.100 97.600 ;
        RECT 602.800 91.600 603.600 92.400 ;
        RECT 604.400 91.600 605.200 92.400 ;
        RECT 594.800 64.200 595.600 75.800 ;
        RECT 601.200 71.600 602.000 72.400 ;
        RECT 601.300 70.400 601.900 71.600 ;
        RECT 601.200 69.600 602.000 70.400 ;
        RECT 602.800 65.600 603.600 66.400 ;
        RECT 593.200 59.600 594.000 60.400 ;
        RECT 585.200 57.600 586.000 58.400 ;
        RECT 588.400 57.600 589.200 58.400 ;
        RECT 599.600 57.600 600.400 58.400 ;
        RECT 594.800 55.600 595.600 56.400 ;
        RECT 583.600 53.600 584.400 54.400 ;
        RECT 585.200 53.600 586.000 54.400 ;
        RECT 588.400 53.600 589.200 54.400 ;
        RECT 585.300 50.400 585.900 53.600 ;
        RECT 575.600 49.400 576.400 50.200 ;
        RECT 581.800 49.400 582.600 50.200 ;
        RECT 585.200 49.600 586.000 50.400 ;
        RECT 588.500 48.400 589.100 53.600 ;
        RECT 591.600 51.600 592.400 52.400 ;
        RECT 569.200 47.600 570.000 48.400 ;
        RECT 588.400 47.600 589.200 48.400 ;
        RECT 566.000 43.600 566.800 44.400 ;
        RECT 559.600 37.600 560.400 38.400 ;
        RECT 564.400 37.600 565.200 38.400 ;
        RECT 556.400 33.600 557.200 34.400 ;
        RECT 551.600 31.600 552.400 32.400 ;
        RECT 553.200 31.600 554.000 32.400 ;
        RECT 556.400 31.600 557.200 32.400 ;
        RECT 551.700 30.400 552.300 31.600 ;
        RECT 556.500 30.400 557.100 31.600 ;
        RECT 559.700 30.400 560.300 37.600 ;
        RECT 566.100 30.400 566.700 43.600 ;
        RECT 567.600 33.600 568.400 34.400 ;
        RECT 567.700 30.400 568.300 33.600 ;
        RECT 569.300 30.400 569.900 47.600 ;
        RECT 591.700 46.400 592.300 51.600 ;
        RECT 591.600 45.600 592.400 46.400 ;
        RECT 593.200 43.600 594.000 44.400 ;
        RECT 572.400 33.600 573.200 34.400 ;
        RECT 551.600 29.600 552.400 30.400 ;
        RECT 556.400 29.600 557.200 30.400 ;
        RECT 559.600 29.600 560.400 30.400 ;
        RECT 566.000 29.600 566.800 30.400 ;
        RECT 567.600 29.600 568.400 30.400 ;
        RECT 569.200 29.600 570.000 30.400 ;
        RECT 550.000 27.600 550.800 28.400 ;
        RECT 559.600 27.600 560.400 28.400 ;
        RECT 554.800 23.600 555.600 24.400 ;
        RECT 580.400 24.200 581.200 35.800 ;
        RECT 583.600 29.600 584.400 30.400 ;
        RECT 582.000 27.600 582.800 28.400 ;
        RECT 554.900 20.300 555.500 23.600 ;
        RECT 554.900 19.700 557.100 20.300 ;
        RECT 540.400 17.600 541.200 18.400 ;
        RECT 546.800 17.600 547.600 18.400 ;
        RECT 538.800 15.600 539.600 16.400 ;
        RECT 529.200 11.600 530.000 12.400 ;
        RECT 546.800 11.600 547.600 12.400 ;
        RECT 551.600 4.200 552.400 17.800 ;
        RECT 553.200 4.200 554.000 17.800 ;
        RECT 554.800 6.200 555.600 17.800 ;
        RECT 556.500 14.400 557.100 19.700 ;
        RECT 556.400 13.600 557.200 14.400 ;
        RECT 558.000 6.200 558.800 17.800 ;
        RECT 559.600 15.600 560.400 16.400 ;
        RECT 561.200 6.200 562.000 17.800 ;
        RECT 562.800 4.200 563.600 17.800 ;
        RECT 564.400 4.200 565.200 17.800 ;
        RECT 566.000 4.200 566.800 17.800 ;
        RECT 575.600 17.600 576.400 18.400 ;
        RECT 582.100 16.400 582.700 27.600 ;
        RECT 590.000 24.200 590.800 35.800 ;
        RECT 593.300 34.400 593.900 43.600 ;
        RECT 594.900 38.400 595.500 55.600 ;
        RECT 598.000 53.600 598.800 54.400 ;
        RECT 598.100 52.400 598.700 53.600 ;
        RECT 596.400 51.600 597.200 52.400 ;
        RECT 598.000 51.600 598.800 52.400 ;
        RECT 594.800 37.600 595.600 38.400 ;
        RECT 593.200 33.600 594.000 34.400 ;
        RECT 591.600 27.600 592.400 28.400 ;
        RECT 593.200 26.200 594.000 31.800 ;
        RECT 596.500 18.400 597.100 51.600 ;
        RECT 599.700 50.400 600.300 57.600 ;
        RECT 602.900 52.400 603.500 65.600 ;
        RECT 604.400 64.200 605.200 75.800 ;
        RECT 607.700 74.300 608.300 113.600 ;
        RECT 609.200 104.200 610.000 115.800 ;
        RECT 610.900 102.400 611.500 129.600 ;
        RECT 623.700 126.400 624.300 153.600 ;
        RECT 626.900 152.400 627.500 159.600 ;
        RECT 631.700 158.400 632.300 187.600 ;
        RECT 636.500 182.400 637.100 189.600 ;
        RECT 636.400 181.600 637.200 182.400 ;
        RECT 638.100 180.300 638.700 189.600 ;
        RECT 636.500 179.700 638.700 180.300 ;
        RECT 636.500 178.400 637.100 179.700 ;
        RECT 641.200 179.600 642.000 180.400 ;
        RECT 636.400 177.600 637.200 178.400 ;
        RECT 641.300 176.400 641.900 179.600 ;
        RECT 641.200 175.600 642.000 176.400 ;
        RECT 642.900 172.400 643.500 211.600 ;
        RECT 647.400 210.200 648.000 215.000 ;
        RECT 649.200 214.800 650.000 215.000 ;
        RECT 652.600 214.800 653.400 215.000 ;
        RECT 654.200 214.200 654.800 215.000 ;
        RECT 655.700 214.400 656.300 215.600 ;
        RECT 650.000 213.600 654.800 214.200 ;
        RECT 655.600 213.600 656.400 214.400 ;
        RECT 650.000 213.400 650.800 213.600 ;
        RECT 654.200 210.200 654.800 213.600 ;
        RECT 658.900 212.400 659.500 253.600 ;
        RECT 660.500 252.400 661.100 257.600 ;
        RECT 662.000 255.600 662.800 256.400 ;
        RECT 662.100 252.400 662.700 255.600 ;
        RECT 663.700 254.400 664.300 267.600 ;
        RECT 663.600 253.600 664.400 254.400 ;
        RECT 660.400 251.600 661.200 252.400 ;
        RECT 662.000 251.600 662.800 252.400 ;
        RECT 665.200 251.600 666.000 252.400 ;
        RECT 663.600 249.600 664.400 250.400 ;
        RECT 663.700 226.400 664.300 249.600 ;
        RECT 666.900 238.400 667.500 269.600 ;
        RECT 671.600 264.200 672.400 275.800 ;
        RECT 673.300 270.400 673.900 301.600 ;
        RECT 676.400 273.600 677.200 274.400 ;
        RECT 676.500 270.400 677.100 273.600 ;
        RECT 673.200 269.600 674.000 270.400 ;
        RECT 676.400 269.600 677.200 270.400 ;
        RECT 668.400 251.600 669.200 252.400 ;
        RECT 668.400 249.600 669.200 250.400 ;
        RECT 670.000 250.200 670.800 255.800 ;
        RECT 671.600 253.600 672.400 254.400 ;
        RECT 671.700 248.300 672.300 253.600 ;
        RECT 670.100 247.700 672.300 248.300 ;
        RECT 666.800 237.600 667.600 238.400 ;
        RECT 663.600 225.600 664.400 226.400 ;
        RECT 668.400 226.200 669.200 231.800 ;
        RECT 662.000 223.600 662.800 224.400 ;
        RECT 668.400 224.300 669.200 224.400 ;
        RECT 670.100 224.300 670.700 247.700 ;
        RECT 673.200 246.200 674.000 257.800 ;
        RECT 674.800 251.600 675.600 252.600 ;
        RECT 673.200 243.600 674.000 244.400 ;
        RECT 668.400 223.700 670.700 224.300 ;
        RECT 671.600 224.200 672.400 235.800 ;
        RECT 668.400 223.600 669.200 223.700 ;
        RECT 662.100 216.400 662.700 223.600 ;
        RECT 668.500 218.400 669.100 223.600 ;
        RECT 668.400 217.600 669.200 218.400 ;
        RECT 662.000 215.600 662.800 216.400 ;
        RECT 655.600 211.600 656.400 212.400 ;
        RECT 658.800 211.600 659.600 212.400 ;
        RECT 647.400 209.400 648.200 210.200 ;
        RECT 654.000 209.400 654.800 210.200 ;
        RECT 652.400 197.600 653.200 198.400 ;
        RECT 644.400 184.200 645.200 195.800 ;
        RECT 647.600 195.600 648.400 196.400 ;
        RECT 646.000 177.600 646.800 178.400 ;
        RECT 646.100 172.400 646.700 177.600 ;
        RECT 633.200 171.600 634.000 172.400 ;
        RECT 639.600 171.600 640.400 172.400 ;
        RECT 642.800 171.600 643.600 172.400 ;
        RECT 646.000 171.600 646.800 172.400 ;
        RECT 633.300 158.400 633.900 171.600 ;
        RECT 646.100 170.400 646.700 171.600 ;
        RECT 636.400 169.600 637.200 170.400 ;
        RECT 646.000 169.600 646.800 170.400 ;
        RECT 638.000 167.600 638.800 168.400 ;
        RECT 639.600 167.600 640.400 168.400 ;
        RECT 638.100 158.400 638.700 167.600 ;
        RECT 631.600 157.600 632.400 158.400 ;
        RECT 633.200 157.600 634.000 158.400 ;
        RECT 638.000 157.600 638.800 158.400 ;
        RECT 626.800 151.600 627.600 152.400 ;
        RECT 630.000 151.600 630.800 152.400 ;
        RECT 625.200 149.600 626.000 150.400 ;
        RECT 628.400 149.600 629.200 150.400 ;
        RECT 625.300 146.400 625.900 149.600 ;
        RECT 625.200 145.600 626.000 146.400 ;
        RECT 630.100 140.300 630.700 151.600 ;
        RECT 634.800 149.600 635.600 150.400 ;
        RECT 631.600 143.600 632.400 144.400 ;
        RECT 628.500 139.700 630.700 140.300 ;
        RECT 625.200 137.600 626.000 138.400 ;
        RECT 623.600 125.600 624.400 126.400 ;
        RECT 620.400 121.600 621.200 122.400 ;
        RECT 617.200 113.600 618.000 114.400 ;
        RECT 617.300 110.200 617.900 113.600 ;
        RECT 617.200 109.400 618.000 110.200 ;
        RECT 612.400 105.600 613.200 106.400 ;
        RECT 610.800 101.600 611.600 102.400 ;
        RECT 612.500 98.400 613.100 105.600 ;
        RECT 618.800 104.200 619.600 115.800 ;
        RECT 620.500 108.400 621.100 121.600 ;
        RECT 626.800 117.600 627.600 118.400 ;
        RECT 625.200 113.600 626.000 114.400 ;
        RECT 620.400 107.600 621.200 108.400 ;
        RECT 622.000 106.200 622.800 111.800 ;
        RECT 625.200 110.300 626.000 110.400 ;
        RECT 626.900 110.300 627.500 117.600 ;
        RECT 625.200 109.700 627.500 110.300 ;
        RECT 625.200 109.600 626.000 109.700 ;
        RECT 623.600 107.600 624.400 108.400 ;
        RECT 623.700 106.400 624.300 107.600 ;
        RECT 623.600 105.600 624.400 106.400 ;
        RECT 615.600 101.600 616.400 102.400 ;
        RECT 612.400 97.600 613.200 98.400 ;
        RECT 610.800 93.600 611.600 94.400 ;
        RECT 610.900 92.400 611.500 93.600 ;
        RECT 615.700 92.400 616.300 101.600 ;
        RECT 622.000 99.600 622.800 100.400 ;
        RECT 617.200 93.600 618.000 94.400 ;
        RECT 618.800 93.600 619.600 94.400 ;
        RECT 609.200 91.600 610.000 92.400 ;
        RECT 610.800 91.600 611.600 92.400 ;
        RECT 615.600 91.600 616.400 92.400 ;
        RECT 606.100 73.700 608.300 74.300 ;
        RECT 606.100 68.400 606.700 73.700 ;
        RECT 606.000 67.600 606.800 68.400 ;
        RECT 607.600 66.200 608.400 71.800 ;
        RECT 609.300 64.400 609.900 91.600 ;
        RECT 612.400 89.600 613.200 90.400 ;
        RECT 612.500 78.400 613.100 89.600 ;
        RECT 612.400 77.600 613.200 78.400 ;
        RECT 612.400 75.600 613.200 76.400 ;
        RECT 610.800 73.600 611.600 74.400 ;
        RECT 612.500 70.400 613.100 75.600 ;
        RECT 614.000 71.600 614.800 72.400 ;
        RECT 612.400 69.600 613.200 70.400 ;
        RECT 609.200 63.600 610.000 64.400 ;
        RECT 602.800 51.600 603.600 52.400 ;
        RECT 599.600 49.600 600.400 50.400 ;
        RECT 604.400 46.200 605.200 57.800 ;
        RECT 609.300 38.400 609.900 63.600 ;
        RECT 614.100 62.400 614.700 71.600 ;
        RECT 615.700 70.400 616.300 91.600 ;
        RECT 617.300 88.400 617.900 93.600 ;
        RECT 620.400 91.600 621.200 92.400 ;
        RECT 620.400 89.600 621.200 90.400 ;
        RECT 617.200 87.600 618.000 88.400 ;
        RECT 617.200 79.600 618.000 80.400 ;
        RECT 617.300 78.400 617.900 79.600 ;
        RECT 617.200 77.600 618.000 78.400 ;
        RECT 615.600 69.600 616.400 70.400 ;
        RECT 615.600 67.600 616.400 68.400 ;
        RECT 614.000 61.600 614.800 62.400 ;
        RECT 612.400 59.600 613.200 60.400 ;
        RECT 612.500 56.400 613.100 59.600 ;
        RECT 612.400 55.600 613.200 56.400 ;
        RECT 612.400 51.800 613.200 52.600 ;
        RECT 612.500 48.400 613.100 51.800 ;
        RECT 612.400 47.600 613.200 48.400 ;
        RECT 614.000 46.200 614.800 57.800 ;
        RECT 615.700 44.400 616.300 67.600 ;
        RECT 617.200 50.200 618.000 55.800 ;
        RECT 618.800 53.600 619.600 54.400 ;
        RECT 618.900 52.400 619.500 53.600 ;
        RECT 618.800 51.600 619.600 52.400 ;
        RECT 620.400 51.600 621.200 52.400 ;
        RECT 620.500 50.400 621.100 51.600 ;
        RECT 620.400 49.600 621.200 50.400 ;
        RECT 615.600 43.600 616.400 44.400 ;
        RECT 609.200 37.600 610.000 38.400 ;
        RECT 598.000 33.600 598.800 34.400 ;
        RECT 598.100 30.400 598.700 33.600 ;
        RECT 598.000 29.600 598.800 30.400 ;
        RECT 602.800 24.200 603.600 35.800 ;
        RECT 609.200 33.600 610.000 34.400 ;
        RECT 610.800 33.600 611.600 34.400 ;
        RECT 604.400 27.600 605.200 28.400 ;
        RECT 588.400 17.600 589.200 18.400 ;
        RECT 582.000 15.600 582.800 16.400 ;
        RECT 593.200 6.200 594.000 17.800 ;
        RECT 596.400 17.600 597.200 18.400 ;
        RECT 601.200 11.800 602.000 12.600 ;
        RECT 601.300 10.400 601.900 11.800 ;
        RECT 601.200 9.600 602.000 10.400 ;
        RECT 602.800 6.200 603.600 17.800 ;
        RECT 604.500 14.400 605.100 27.600 ;
        RECT 604.400 13.600 605.200 14.400 ;
        RECT 606.000 10.200 606.800 15.800 ;
        RECT 607.600 15.600 608.400 16.400 ;
        RECT 607.700 14.400 608.300 15.600 ;
        RECT 607.600 13.600 608.400 14.400 ;
        RECT 609.300 12.400 609.900 33.600 ;
        RECT 610.900 30.200 611.500 33.600 ;
        RECT 610.800 29.400 611.600 30.200 ;
        RECT 612.400 24.200 613.200 35.800 ;
        RECT 622.100 34.300 622.700 99.600 ;
        RECT 623.700 94.400 624.300 105.600 ;
        RECT 625.200 97.600 626.000 98.400 ;
        RECT 623.600 93.600 624.400 94.400 ;
        RECT 625.300 90.400 625.900 97.600 ;
        RECT 625.200 89.600 626.000 90.400 ;
        RECT 625.200 75.600 626.000 76.400 ;
        RECT 623.600 73.600 624.400 74.400 ;
        RECT 625.300 70.400 625.900 75.600 ;
        RECT 626.800 71.600 627.600 72.400 ;
        RECT 628.500 70.400 629.100 139.700 ;
        RECT 630.000 126.200 630.800 137.800 ;
        RECT 631.700 126.300 632.300 143.600 ;
        RECT 633.200 133.600 634.000 134.400 ;
        RECT 633.300 132.400 633.900 133.600 ;
        RECT 633.200 131.600 634.000 132.400 ;
        RECT 631.700 125.700 633.900 126.300 ;
        RECT 631.600 123.600 632.400 124.400 ;
        RECT 630.000 115.600 630.800 116.400 ;
        RECT 630.100 112.400 630.700 115.600 ;
        RECT 630.000 111.600 630.800 112.400 ;
        RECT 630.000 107.600 630.800 108.400 ;
        RECT 630.100 104.400 630.700 107.600 ;
        RECT 630.000 103.600 630.800 104.400 ;
        RECT 630.000 93.600 630.800 94.400 ;
        RECT 631.700 92.400 632.300 123.600 ;
        RECT 633.300 108.300 633.900 125.700 ;
        RECT 634.900 124.400 635.500 149.600 ;
        RECT 638.000 143.600 638.800 144.400 ;
        RECT 636.400 139.600 637.200 140.400 ;
        RECT 634.800 123.600 635.600 124.400 ;
        RECT 634.800 119.600 635.600 120.400 ;
        RECT 634.900 110.400 635.500 119.600 ;
        RECT 636.500 110.400 637.100 139.600 ;
        RECT 638.100 132.400 638.700 143.600 ;
        RECT 639.700 142.400 640.300 167.600 ;
        RECT 644.400 163.600 645.200 164.400 ;
        RECT 646.000 163.600 646.800 164.400 ;
        RECT 641.200 155.600 642.000 156.400 ;
        RECT 644.500 150.400 645.100 163.600 ;
        RECT 646.100 154.400 646.700 163.600 ;
        RECT 647.700 156.400 648.300 195.600 ;
        RECT 650.800 193.600 651.600 194.400 ;
        RECT 649.200 191.600 650.000 192.400 ;
        RECT 649.300 168.400 649.900 191.600 ;
        RECT 650.900 190.400 651.500 193.600 ;
        RECT 650.800 189.600 651.600 190.400 ;
        RECT 652.500 188.400 653.100 197.600 ;
        RECT 652.400 187.600 653.200 188.400 ;
        RECT 650.800 183.600 651.600 184.400 ;
        RECT 650.900 178.400 651.500 183.600 ;
        RECT 650.800 177.600 651.600 178.400 ;
        RECT 652.500 174.400 653.100 187.600 ;
        RECT 654.000 184.200 654.800 195.800 ;
        RECT 655.700 184.300 656.300 211.600 ;
        RECT 657.200 186.200 658.000 191.800 ;
        RECT 662.100 190.400 662.700 215.600 ;
        RECT 665.200 213.600 666.000 214.400 ;
        RECT 671.600 213.600 672.400 214.400 ;
        RECT 663.600 195.600 664.400 196.400 ;
        RECT 662.000 189.600 662.800 190.400 ;
        RECT 662.100 186.400 662.700 189.600 ;
        RECT 658.800 185.600 659.600 186.400 ;
        RECT 660.400 185.600 661.200 186.400 ;
        RECT 662.000 185.600 662.800 186.400 ;
        RECT 655.700 183.700 657.900 184.300 ;
        RECT 655.600 179.600 656.400 180.400 ;
        RECT 655.700 178.400 656.300 179.600 ;
        RECT 655.600 177.600 656.400 178.400 ;
        RECT 652.400 173.600 653.200 174.400 ;
        RECT 649.200 167.600 650.000 168.400 ;
        RECT 655.600 159.600 656.400 160.400 ;
        RECT 649.200 157.600 650.000 158.400 ;
        RECT 647.600 155.600 648.400 156.400 ;
        RECT 646.000 153.600 646.800 154.400 ;
        RECT 644.400 149.600 645.200 150.400 ;
        RECT 646.000 149.600 646.800 150.400 ;
        RECT 642.800 145.600 643.600 146.400 ;
        RECT 639.600 141.600 640.400 142.400 ;
        RECT 644.500 140.400 645.100 149.600 ;
        RECT 646.100 146.400 646.700 149.600 ;
        RECT 646.000 145.600 646.800 146.400 ;
        RECT 647.600 141.600 648.400 142.400 ;
        RECT 644.400 139.600 645.200 140.400 ;
        RECT 638.000 131.600 638.800 132.400 ;
        RECT 638.100 120.400 638.700 131.600 ;
        RECT 639.600 126.200 640.400 137.800 ;
        RECT 641.200 133.600 642.000 134.400 ;
        RECT 641.300 130.400 641.900 133.600 ;
        RECT 641.200 129.600 642.000 130.400 ;
        RECT 642.800 130.200 643.600 135.800 ;
        RECT 646.000 135.600 646.800 136.400 ;
        RECT 646.100 134.400 646.700 135.600 ;
        RECT 646.000 133.600 646.800 134.400 ;
        RECT 647.700 132.400 648.300 141.600 ;
        RECT 649.300 132.400 649.900 157.600 ;
        RECT 655.700 154.400 656.300 159.600 ;
        RECT 654.000 153.600 654.800 154.400 ;
        RECT 655.600 153.600 656.400 154.400 ;
        RECT 654.100 150.400 654.700 153.600 ;
        RECT 655.700 150.400 656.300 153.600 ;
        RECT 650.800 149.600 651.600 150.400 ;
        RECT 654.000 149.600 654.800 150.400 ;
        RECT 655.600 149.600 656.400 150.400 ;
        RECT 652.400 147.600 653.200 148.400 ;
        RECT 650.800 133.600 651.600 134.400 ;
        RECT 647.600 131.600 648.400 132.400 ;
        RECT 649.200 131.600 650.000 132.400 ;
        RECT 641.300 122.400 641.900 129.600 ;
        RECT 644.400 127.600 645.200 128.400 ;
        RECT 641.200 121.600 642.000 122.400 ;
        RECT 638.000 119.600 638.800 120.400 ;
        RECT 639.600 117.600 640.400 118.400 ;
        RECT 638.000 115.600 638.800 116.400 ;
        RECT 638.100 110.400 638.700 115.600 ;
        RECT 647.700 110.400 648.300 131.600 ;
        RECT 634.800 109.600 635.600 110.400 ;
        RECT 636.400 109.600 637.200 110.400 ;
        RECT 638.000 109.600 638.800 110.400 ;
        RECT 642.800 109.600 643.600 110.400 ;
        RECT 647.600 109.600 648.400 110.400 ;
        RECT 634.800 108.300 635.600 108.400 ;
        RECT 633.300 107.700 635.600 108.300 ;
        RECT 634.800 107.600 635.600 107.700 ;
        RECT 634.900 96.300 635.500 107.600 ;
        RECT 638.000 105.600 638.800 106.400 ;
        RECT 634.900 95.700 637.100 96.300 ;
        RECT 636.500 94.400 637.100 95.700 ;
        RECT 634.800 93.600 635.600 94.400 ;
        RECT 636.400 93.600 637.200 94.400 ;
        RECT 630.000 91.600 630.800 92.400 ;
        RECT 631.600 91.600 632.400 92.400 ;
        RECT 634.900 92.300 635.500 93.600 ;
        RECT 636.400 92.300 637.200 92.400 ;
        RECT 634.900 91.700 637.200 92.300 ;
        RECT 636.400 91.600 637.200 91.700 ;
        RECT 633.200 77.600 634.000 78.400 ;
        RECT 630.000 71.600 630.800 72.400 ;
        RECT 630.100 70.400 630.700 71.600 ;
        RECT 625.200 69.600 626.000 70.400 ;
        RECT 628.400 69.600 629.200 70.400 ;
        RECT 630.000 69.600 630.800 70.400 ;
        RECT 626.800 55.600 627.600 56.400 ;
        RECT 626.900 54.400 627.500 55.600 ;
        RECT 628.500 54.400 629.100 69.600 ;
        RECT 626.800 53.600 627.600 54.400 ;
        RECT 628.400 53.600 629.200 54.400 ;
        RECT 633.300 52.400 633.900 77.600 ;
        RECT 634.800 69.600 635.600 70.400 ;
        RECT 636.400 69.600 637.200 70.400 ;
        RECT 634.900 68.400 635.500 69.600 ;
        RECT 634.800 67.600 635.600 68.400 ;
        RECT 636.500 64.400 637.100 69.600 ;
        RECT 638.100 68.400 638.700 105.600 ;
        RECT 642.900 100.400 643.500 109.600 ;
        RECT 647.600 105.600 648.400 106.400 ;
        RECT 642.800 99.600 643.600 100.400 ;
        RECT 650.900 98.400 651.500 133.600 ;
        RECT 652.500 132.400 653.100 147.600 ;
        RECT 657.300 138.400 657.900 183.700 ;
        RECT 658.900 180.400 659.500 185.600 ;
        RECT 660.400 181.600 661.200 182.400 ;
        RECT 662.000 181.600 662.800 182.400 ;
        RECT 658.800 179.600 659.600 180.400 ;
        RECT 658.800 175.600 659.600 176.400 ;
        RECT 657.200 137.600 658.000 138.400 ;
        RECT 657.200 135.600 658.000 136.400 ;
        RECT 654.000 133.600 654.800 134.400 ;
        RECT 654.100 132.400 654.700 133.600 ;
        RECT 657.300 132.400 657.900 135.600 ;
        RECT 652.400 131.600 653.200 132.400 ;
        RECT 654.000 131.600 654.800 132.400 ;
        RECT 657.200 131.600 658.000 132.400 ;
        RECT 652.400 123.600 653.200 124.400 ;
        RECT 652.500 116.400 653.100 123.600 ;
        RECT 652.400 115.600 653.200 116.400 ;
        RECT 657.300 114.400 657.900 131.600 ;
        RECT 652.400 113.600 653.200 114.400 ;
        RECT 657.200 113.600 658.000 114.400 ;
        RECT 652.500 110.400 653.100 113.600 ;
        RECT 657.300 110.400 657.900 113.600 ;
        RECT 652.400 109.600 653.200 110.400 ;
        RECT 657.200 109.600 658.000 110.400 ;
        RECT 654.000 103.600 654.800 104.400 ;
        RECT 650.800 97.600 651.600 98.400 ;
        RECT 644.400 93.600 645.200 94.400 ;
        RECT 641.200 91.600 642.000 92.400 ;
        RECT 646.000 92.300 646.800 92.400 ;
        RECT 646.000 91.700 648.300 92.300 ;
        RECT 646.000 91.600 646.800 91.700 ;
        RECT 641.300 72.300 641.900 91.600 ;
        RECT 642.800 89.600 643.600 90.400 ;
        RECT 642.900 74.400 643.500 89.600 ;
        RECT 646.000 83.600 646.800 84.400 ;
        RECT 642.800 73.600 643.600 74.400 ;
        RECT 644.400 73.600 645.200 74.400 ;
        RECT 646.100 72.400 646.700 83.600 ;
        RECT 642.800 72.300 643.600 72.400 ;
        RECT 641.300 71.700 643.600 72.300 ;
        RECT 642.800 71.600 643.600 71.700 ;
        RECT 646.000 71.600 646.800 72.400 ;
        RECT 639.600 69.600 640.400 70.400 ;
        RECT 642.800 69.600 643.600 70.400 ;
        RECT 638.000 67.600 638.800 68.400 ;
        RECT 636.400 63.600 637.200 64.400 ;
        RECT 636.400 61.600 637.200 62.400 ;
        RECT 636.500 54.400 637.100 61.600 ;
        RECT 634.800 53.600 635.600 54.400 ;
        RECT 636.400 53.600 637.200 54.400 ;
        RECT 634.900 52.400 635.500 53.600 ;
        RECT 636.500 52.400 637.100 53.600 ;
        RECT 625.200 51.600 626.000 52.400 ;
        RECT 633.200 51.600 634.000 52.400 ;
        RECT 634.800 51.600 635.600 52.400 ;
        RECT 636.400 51.600 637.200 52.400 ;
        RECT 625.300 38.400 625.900 51.600 ;
        RECT 630.000 43.600 630.800 44.400 ;
        RECT 633.200 43.600 634.000 44.400 ;
        RECT 636.400 43.600 637.200 44.400 ;
        RECT 628.400 41.600 629.200 42.400 ;
        RECT 625.200 37.600 626.000 38.400 ;
        RECT 622.100 33.700 624.300 34.300 ;
        RECT 618.800 32.300 619.600 32.400 ;
        RECT 614.000 27.600 614.800 28.400 ;
        RECT 614.100 22.400 614.700 27.600 ;
        RECT 615.600 26.200 616.400 31.800 ;
        RECT 618.800 31.700 621.100 32.300 ;
        RECT 618.800 31.600 619.600 31.700 ;
        RECT 618.900 30.400 619.500 31.600 ;
        RECT 618.800 29.600 619.600 30.400 ;
        RECT 617.200 27.600 618.000 28.400 ;
        RECT 618.800 27.600 619.600 28.400 ;
        RECT 614.000 21.600 614.800 22.400 ;
        RECT 614.000 17.600 614.800 18.400 ;
        RECT 609.200 11.600 610.000 12.400 ;
        RECT 614.100 10.400 614.700 17.600 ;
        RECT 618.900 14.400 619.500 27.600 ;
        RECT 618.800 13.600 619.600 14.400 ;
        RECT 620.500 12.400 621.100 31.700 ;
        RECT 622.000 31.600 622.800 32.400 ;
        RECT 620.400 11.600 621.200 12.400 ;
        RECT 609.200 9.600 610.000 10.400 ;
        RECT 614.000 9.600 614.800 10.400 ;
        RECT 623.700 8.400 624.300 33.700 ;
        RECT 626.800 33.600 627.600 34.400 ;
        RECT 628.500 28.400 629.100 41.600 ;
        RECT 630.100 30.400 630.700 43.600 ;
        RECT 631.600 31.600 632.400 32.400 ;
        RECT 631.700 30.400 632.300 31.600 ;
        RECT 630.000 29.600 630.800 30.400 ;
        RECT 631.600 29.600 632.400 30.400 ;
        RECT 630.100 28.400 630.700 29.600 ;
        RECT 628.400 27.600 629.200 28.400 ;
        RECT 630.000 27.600 630.800 28.400 ;
        RECT 625.200 19.600 626.000 20.400 ;
        RECT 625.300 10.400 625.900 19.600 ;
        RECT 628.500 16.400 629.100 27.600 ;
        RECT 633.300 18.400 633.900 43.600 ;
        RECT 636.500 38.400 637.100 43.600 ;
        RECT 638.100 42.400 638.700 67.600 ;
        RECT 639.600 63.600 640.400 64.400 ;
        RECT 639.700 46.300 640.300 63.600 ;
        RECT 642.800 53.600 643.600 54.400 ;
        RECT 646.000 53.600 646.800 54.400 ;
        RECT 641.200 51.600 642.000 52.400 ;
        RECT 639.700 45.700 641.900 46.300 ;
        RECT 639.600 43.600 640.400 44.400 ;
        RECT 638.000 41.600 638.800 42.400 ;
        RECT 636.400 37.600 637.200 38.400 ;
        RECT 638.000 37.600 638.800 38.400 ;
        RECT 634.800 33.600 635.600 34.400 ;
        RECT 633.200 17.600 634.000 18.400 ;
        RECT 634.900 16.400 635.500 33.600 ;
        RECT 636.500 30.400 637.100 37.600 ;
        RECT 638.100 36.400 638.700 37.600 ;
        RECT 638.000 35.600 638.800 36.400 ;
        RECT 638.100 30.400 638.700 35.600 ;
        RECT 636.400 29.600 637.200 30.400 ;
        RECT 638.000 29.600 638.800 30.400 ;
        RECT 636.400 25.600 637.200 26.400 ;
        RECT 636.500 18.400 637.100 25.600 ;
        RECT 636.400 17.600 637.200 18.400 ;
        RECT 639.700 16.400 640.300 43.600 ;
        RECT 641.300 30.400 641.900 45.700 ;
        RECT 641.200 29.600 642.000 30.400 ;
        RECT 642.900 20.400 643.500 53.600 ;
        RECT 644.400 49.600 645.200 50.400 ;
        RECT 646.100 48.400 646.700 53.600 ;
        RECT 647.700 52.400 648.300 91.700 ;
        RECT 649.200 64.200 650.000 75.800 ;
        RECT 652.400 69.600 653.200 70.400 ;
        RECT 654.100 66.400 654.700 103.600 ;
        RECT 655.600 86.200 656.400 97.800 ;
        RECT 658.900 96.400 659.500 175.600 ;
        RECT 660.500 150.400 661.100 181.600 ;
        RECT 660.400 149.600 661.200 150.400 ;
        RECT 662.100 150.300 662.700 181.600 ;
        RECT 663.700 152.400 664.300 195.600 ;
        RECT 665.300 190.400 665.900 213.600 ;
        RECT 671.700 212.400 672.300 213.600 ;
        RECT 671.600 211.600 672.400 212.400 ;
        RECT 671.600 193.600 672.400 194.400 ;
        RECT 671.700 192.400 672.300 193.600 ;
        RECT 671.600 191.600 672.400 192.400 ;
        RECT 665.200 190.300 666.000 190.400 ;
        RECT 666.800 190.300 667.600 190.400 ;
        RECT 665.200 189.700 667.600 190.300 ;
        RECT 665.200 189.600 666.000 189.700 ;
        RECT 666.800 189.600 667.600 189.700 ;
        RECT 671.600 189.600 672.400 190.400 ;
        RECT 665.300 182.400 665.900 189.600 ;
        RECT 666.800 185.600 667.600 186.400 ;
        RECT 670.000 185.600 670.800 186.400 ;
        RECT 671.600 183.600 672.400 184.400 ;
        RECT 665.200 181.600 666.000 182.400 ;
        RECT 671.700 178.400 672.300 183.600 ;
        RECT 673.300 182.400 673.900 243.600 ;
        RECT 674.800 229.600 675.600 230.400 ;
        RECT 674.800 227.600 675.600 228.400 ;
        RECT 673.200 181.600 674.000 182.400 ;
        RECT 674.900 180.400 675.500 227.600 ;
        RECT 678.100 194.400 678.700 345.600 ;
        RECT 679.600 343.600 680.400 344.400 ;
        RECT 679.700 200.400 680.300 343.600 ;
        RECT 681.200 331.600 682.000 332.400 ;
        RECT 681.300 320.400 681.900 331.600 ;
        RECT 682.800 326.200 683.600 337.800 ;
        RECT 687.600 337.600 688.400 338.400 ;
        RECT 687.700 330.400 688.300 337.600 ;
        RECT 687.600 329.600 688.400 330.400 ;
        RECT 681.200 319.600 682.000 320.400 ;
        RECT 681.200 304.200 682.000 315.800 ;
        RECT 686.000 313.600 686.800 314.400 ;
        RECT 686.100 312.400 686.700 313.600 ;
        RECT 686.000 311.600 686.800 312.400 ;
        RECT 681.200 301.600 682.000 302.400 ;
        RECT 681.300 298.400 681.900 301.600 ;
        RECT 681.200 297.600 682.000 298.400 ;
        RECT 681.200 264.200 682.000 275.800 ;
        RECT 684.400 266.200 685.200 271.800 ;
        RECT 682.800 246.200 683.600 257.800 ;
        RECT 687.600 257.600 688.400 258.400 ;
        RECT 681.200 224.200 682.000 235.800 ;
        RECT 686.000 223.600 686.800 224.400 ;
        RECT 686.100 206.400 686.700 223.600 ;
        RECT 686.000 205.600 686.800 206.400 ;
        RECT 682.800 203.600 683.600 204.400 ;
        RECT 679.600 199.600 680.400 200.400 ;
        RECT 682.900 198.400 683.500 203.600 ;
        RECT 682.800 197.600 683.600 198.400 ;
        RECT 678.000 193.600 678.800 194.400 ;
        RECT 676.400 191.600 677.200 192.400 ;
        RECT 679.600 191.800 680.400 192.600 ;
        RECT 686.200 191.800 687.000 192.600 ;
        RECT 676.500 190.400 677.100 191.600 ;
        RECT 676.400 189.600 677.200 190.400 ;
        RECT 679.600 188.400 680.200 191.800 ;
        RECT 683.600 188.400 684.400 188.600 ;
        RECT 676.400 187.600 677.200 188.400 ;
        RECT 678.000 187.600 678.800 188.400 ;
        RECT 679.600 187.800 684.400 188.400 ;
        RECT 678.100 184.400 678.700 187.600 ;
        RECT 679.600 187.000 680.200 187.800 ;
        RECT 681.000 187.000 681.800 187.200 ;
        RECT 684.400 187.000 685.200 187.200 ;
        RECT 686.400 187.000 687.000 191.800 ;
        RECT 687.600 189.600 688.400 190.400 ;
        RECT 687.700 188.400 688.300 189.600 ;
        RECT 687.600 187.600 688.400 188.400 ;
        RECT 679.600 186.200 680.400 187.000 ;
        RECT 681.000 186.400 685.200 187.000 ;
        RECT 686.200 186.200 687.000 187.000 ;
        RECT 678.000 183.600 678.800 184.400 ;
        RECT 681.200 183.600 682.000 184.400 ;
        RECT 674.800 179.600 675.600 180.400 ;
        RECT 665.200 164.200 666.000 177.800 ;
        RECT 666.800 164.200 667.600 177.800 ;
        RECT 668.400 164.200 669.200 177.800 ;
        RECT 670.000 166.200 670.800 177.800 ;
        RECT 671.600 177.600 672.400 178.400 ;
        RECT 671.600 175.600 672.400 176.400 ;
        RECT 671.700 174.400 672.300 175.600 ;
        RECT 671.600 173.600 672.400 174.400 ;
        RECT 668.400 155.600 669.200 156.400 ;
        RECT 668.500 152.400 669.100 155.600 ;
        RECT 670.000 153.600 670.800 154.400 ;
        RECT 671.700 152.400 672.300 173.600 ;
        RECT 673.200 166.200 674.000 177.800 ;
        RECT 674.800 173.600 675.600 174.400 ;
        RECT 674.800 171.600 675.600 172.400 ;
        RECT 676.400 166.200 677.200 177.800 ;
        RECT 676.400 163.600 677.200 164.400 ;
        RECT 678.000 164.200 678.800 177.800 ;
        RECT 679.600 164.200 680.400 177.800 ;
        RECT 681.300 174.400 681.900 183.600 ;
        RECT 682.800 181.600 683.600 182.400 ;
        RECT 681.200 173.600 682.000 174.400 ;
        RECT 682.900 168.400 683.500 181.600 ;
        RECT 684.400 179.600 685.200 180.400 ;
        RECT 682.800 167.600 683.600 168.400 ;
        RECT 663.600 151.600 664.400 152.400 ;
        RECT 668.400 151.600 669.200 152.400 ;
        RECT 671.600 151.600 672.400 152.400 ;
        RECT 662.100 149.700 664.300 150.300 ;
        RECT 663.700 148.400 664.300 149.700 ;
        RECT 668.400 149.600 669.200 150.400 ;
        RECT 663.600 147.600 664.400 148.400 ;
        RECT 663.700 134.400 664.300 147.600 ;
        RECT 670.000 145.600 670.800 146.400 ;
        RECT 670.100 138.400 670.700 145.600 ;
        RECT 674.800 144.200 675.600 155.800 ;
        RECT 670.000 137.600 670.800 138.400 ;
        RECT 671.600 137.600 672.400 138.400 ;
        RECT 663.600 133.600 664.400 134.400 ;
        RECT 665.200 131.600 666.000 132.400 ;
        RECT 668.400 131.600 669.200 132.400 ;
        RECT 660.400 129.600 661.200 130.400 ;
        RECT 668.400 129.600 669.200 130.400 ;
        RECT 660.500 118.400 661.100 129.600 ;
        RECT 660.400 117.600 661.200 118.400 ;
        RECT 666.800 111.600 667.600 112.400 ;
        RECT 660.400 109.600 661.200 110.400 ;
        RECT 658.800 95.600 659.600 96.400 ;
        RECT 657.200 93.600 658.000 94.400 ;
        RECT 657.300 92.400 657.900 93.600 ;
        RECT 657.200 91.600 658.000 92.400 ;
        RECT 657.300 68.400 657.900 91.600 ;
        RECT 657.200 67.600 658.000 68.400 ;
        RECT 654.000 65.600 654.800 66.400 ;
        RECT 654.100 58.300 654.700 65.600 ;
        RECT 658.800 64.200 659.600 75.800 ;
        RECT 654.100 57.700 656.300 58.300 ;
        RECT 654.000 55.600 654.800 56.400 ;
        RECT 649.200 53.600 650.000 54.400 ;
        RECT 650.800 53.600 651.600 54.400 ;
        RECT 647.600 51.600 648.400 52.400 ;
        RECT 646.000 47.600 646.800 48.400 ;
        RECT 647.600 47.600 648.400 48.400 ;
        RECT 647.600 33.600 648.400 34.400 ;
        RECT 647.700 30.400 648.300 33.600 ;
        RECT 649.300 30.400 649.900 53.600 ;
        RECT 654.100 52.400 654.700 55.600 ;
        RECT 655.700 54.400 656.300 57.700 ;
        RECT 660.500 54.400 661.100 109.600 ;
        RECT 663.600 91.800 664.400 92.600 ;
        RECT 663.700 78.400 664.300 91.800 ;
        RECT 665.200 86.200 666.000 97.800 ;
        RECT 666.900 80.300 667.500 111.600 ;
        RECT 671.700 108.400 672.300 137.600 ;
        RECT 674.800 126.200 675.600 137.800 ;
        RECT 674.800 119.600 675.600 120.400 ;
        RECT 674.900 110.400 675.500 119.600 ;
        RECT 674.800 109.600 675.600 110.400 ;
        RECT 671.600 107.600 672.400 108.400 ;
        RECT 673.200 107.600 674.000 108.400 ;
        RECT 668.400 90.200 669.200 95.800 ;
        RECT 670.000 90.200 670.800 95.800 ;
        RECT 670.000 87.600 670.800 88.400 ;
        RECT 665.300 79.700 667.500 80.300 ;
        RECT 663.600 77.600 664.400 78.400 ;
        RECT 662.000 66.200 662.800 71.800 ;
        RECT 663.600 71.600 664.400 72.400 ;
        RECT 655.600 53.600 656.400 54.400 ;
        RECT 660.400 53.600 661.200 54.400 ;
        RECT 665.300 52.400 665.900 79.700 ;
        RECT 670.100 78.400 670.700 87.600 ;
        RECT 666.800 77.600 667.600 78.400 ;
        RECT 670.000 77.600 670.800 78.400 ;
        RECT 670.000 75.600 670.800 76.400 ;
        RECT 666.800 69.600 667.600 70.400 ;
        RECT 668.400 67.600 669.200 68.400 ;
        RECT 668.500 66.400 669.100 67.600 ;
        RECT 668.400 65.600 669.200 66.400 ;
        RECT 668.500 54.400 669.100 65.600 ;
        RECT 666.800 53.600 667.600 54.400 ;
        RECT 668.400 53.600 669.200 54.400 ;
        RECT 666.900 52.400 667.500 53.600 ;
        RECT 650.800 51.600 651.600 52.400 ;
        RECT 654.000 51.600 654.800 52.400 ;
        RECT 658.800 51.600 659.600 52.400 ;
        RECT 660.400 51.600 661.200 52.400 ;
        RECT 663.600 51.600 664.400 52.400 ;
        RECT 665.200 51.600 666.000 52.400 ;
        RECT 666.800 51.600 667.600 52.400 ;
        RECT 668.400 51.600 669.200 52.400 ;
        RECT 650.800 49.600 651.600 50.400 ;
        RECT 650.900 48.400 651.500 49.600 ;
        RECT 650.800 47.600 651.600 48.400 ;
        RECT 658.900 44.400 659.500 51.600 ;
        RECT 658.800 43.600 659.600 44.400 ;
        RECT 654.000 33.600 654.800 34.400 ;
        RECT 654.100 32.400 654.700 33.600 ;
        RECT 660.500 32.400 661.100 51.600 ;
        RECT 663.700 46.400 664.300 51.600 ;
        RECT 663.600 45.600 664.400 46.400 ;
        RECT 662.000 43.600 662.800 44.400 ;
        RECT 662.100 32.400 662.700 43.600 ;
        RECT 663.700 36.400 664.300 45.600 ;
        RECT 666.900 38.400 667.500 51.600 ;
        RECT 668.500 50.400 669.100 51.600 ;
        RECT 668.400 49.600 669.200 50.400 ;
        RECT 666.800 37.600 667.600 38.400 ;
        RECT 663.600 35.600 664.400 36.400 ;
        RECT 666.800 35.600 667.600 36.400 ;
        RECT 666.900 32.400 667.500 35.600 ;
        RECT 650.800 31.600 651.600 32.400 ;
        RECT 654.000 31.600 654.800 32.400 ;
        RECT 660.400 31.600 661.200 32.400 ;
        RECT 662.000 31.600 662.800 32.400 ;
        RECT 666.800 31.600 667.600 32.400 ;
        RECT 650.900 30.400 651.500 31.600 ;
        RECT 647.600 29.600 648.400 30.400 ;
        RECT 649.200 29.600 650.000 30.400 ;
        RECT 650.800 29.600 651.600 30.400 ;
        RECT 649.300 28.400 649.900 29.600 ;
        RECT 647.600 27.600 648.400 28.400 ;
        RECT 649.200 27.600 650.000 28.400 ;
        RECT 649.200 21.600 650.000 22.400 ;
        RECT 642.800 19.600 643.600 20.400 ;
        RECT 642.900 18.400 643.500 19.600 ;
        RECT 641.200 17.600 642.000 18.400 ;
        RECT 642.800 17.600 643.600 18.400 ;
        RECT 628.400 15.600 629.200 16.400 ;
        RECT 630.000 15.600 630.800 16.400 ;
        RECT 634.800 15.600 635.600 16.400 ;
        RECT 639.600 15.600 640.400 16.400 ;
        RECT 628.500 14.400 629.100 15.600 ;
        RECT 628.400 13.600 629.200 14.400 ;
        RECT 630.100 12.400 630.700 15.600 ;
        RECT 641.300 14.400 641.900 17.600 ;
        RECT 631.600 13.600 632.400 14.400 ;
        RECT 641.200 13.600 642.000 14.400 ;
        RECT 630.000 11.600 630.800 12.400 ;
        RECT 639.600 11.600 640.400 12.400 ;
        RECT 625.200 9.600 626.000 10.400 ;
        RECT 630.000 9.600 630.800 10.400 ;
        RECT 636.400 9.600 637.200 10.400 ;
        RECT 636.500 8.400 637.100 9.600 ;
        RECT 623.600 7.600 624.400 8.400 ;
        RECT 636.400 7.600 637.200 8.400 ;
        RECT 647.600 6.200 648.400 17.800 ;
        RECT 649.300 14.400 649.900 21.600 ;
        RECT 654.100 18.400 654.700 31.600 ;
        RECT 660.500 30.400 661.100 31.600 ;
        RECT 658.800 29.600 659.600 30.400 ;
        RECT 660.400 29.600 661.200 30.400 ;
        RECT 662.000 29.600 662.800 30.400 ;
        RECT 658.900 28.400 659.500 29.600 ;
        RECT 662.100 28.400 662.700 29.600 ;
        RECT 658.800 27.600 659.600 28.400 ;
        RECT 660.400 27.600 661.200 28.400 ;
        RECT 662.000 27.600 662.800 28.400 ;
        RECT 655.600 23.600 656.400 24.400 ;
        RECT 654.000 17.600 654.800 18.400 ;
        RECT 649.200 13.600 650.000 14.400 ;
        RECT 655.700 12.400 656.300 23.600 ;
        RECT 654.000 11.600 654.800 12.400 ;
        RECT 655.600 11.600 656.400 12.400 ;
        RECT 654.100 10.400 654.700 11.600 ;
        RECT 654.000 9.600 654.800 10.400 ;
        RECT 657.200 6.200 658.000 17.800 ;
        RECT 662.000 17.600 662.800 18.400 ;
        RECT 658.800 13.600 659.600 14.400 ;
        RECT 660.400 10.200 661.200 15.800 ;
        RECT 666.800 6.200 667.600 17.800 ;
        RECT 670.100 14.400 670.700 75.600 ;
        RECT 671.700 68.400 672.300 107.600 ;
        RECT 673.200 86.200 674.000 97.800 ;
        RECT 676.500 84.400 677.100 163.600 ;
        RECT 684.500 162.400 685.100 179.600 ;
        RECT 681.200 161.600 682.000 162.400 ;
        RECT 684.400 161.600 685.200 162.400 ;
        RECT 678.000 151.600 678.800 152.400 ;
        RECT 678.100 150.400 678.700 151.600 ;
        RECT 678.000 149.600 678.800 150.400 ;
        RECT 679.600 149.600 680.400 150.400 ;
        RECT 679.600 131.600 680.400 132.400 ;
        RECT 681.300 124.400 681.900 161.600 ;
        RECT 682.800 145.600 683.600 146.400 ;
        RECT 682.900 136.400 683.500 145.600 ;
        RECT 684.400 144.200 685.200 155.800 ;
        RECT 687.600 146.200 688.400 151.800 ;
        RECT 682.800 135.600 683.600 136.400 ;
        RECT 684.400 126.200 685.200 137.800 ;
        RECT 687.600 130.200 688.400 135.800 ;
        RECT 681.200 123.600 682.000 124.400 ;
        RECT 684.400 123.600 685.200 124.400 ;
        RECT 678.000 111.600 678.800 112.400 ;
        RECT 679.600 111.600 680.400 112.400 ;
        RECT 678.100 110.400 678.700 111.600 ;
        RECT 679.700 110.400 680.300 111.600 ;
        RECT 678.000 109.600 678.800 110.400 ;
        RECT 679.600 109.600 680.400 110.400 ;
        RECT 681.200 109.600 682.000 110.400 ;
        RECT 681.300 104.400 681.900 109.600 ;
        RECT 678.000 103.600 678.800 104.400 ;
        RECT 681.200 103.600 682.000 104.400 ;
        RECT 682.800 103.600 683.600 104.400 ;
        RECT 676.400 83.600 677.200 84.400 ;
        RECT 671.600 67.600 672.400 68.400 ;
        RECT 673.200 67.600 674.000 68.400 ;
        RECT 671.600 65.600 672.400 66.400 ;
        RECT 671.700 50.400 672.300 65.600 ;
        RECT 678.100 58.400 678.700 103.600 ;
        RECT 682.900 100.400 683.500 103.600 ;
        RECT 682.800 99.600 683.600 100.400 ;
        RECT 679.600 91.600 680.400 92.400 ;
        RECT 678.000 57.600 678.800 58.400 ;
        RECT 673.200 55.600 674.000 56.400 ;
        RECT 673.300 54.400 673.900 55.600 ;
        RECT 673.200 53.600 674.000 54.400 ;
        RECT 674.800 53.600 675.600 54.400 ;
        RECT 671.600 49.600 672.400 50.400 ;
        RECT 671.600 47.600 672.400 48.400 ;
        RECT 671.700 38.400 672.300 47.600 ;
        RECT 671.600 37.600 672.400 38.400 ;
        RECT 671.600 31.600 672.400 32.400 ;
        RECT 671.700 30.400 672.300 31.600 ;
        RECT 674.900 30.400 675.500 53.600 ;
        RECT 676.400 51.600 677.200 52.400 ;
        RECT 678.000 51.600 678.800 52.400 ;
        RECT 676.500 50.400 677.100 51.600 ;
        RECT 676.400 49.600 677.200 50.400 ;
        RECT 679.700 44.400 680.300 91.600 ;
        RECT 682.800 86.200 683.600 97.800 ;
        RECT 682.800 83.600 683.600 84.400 ;
        RECT 682.900 58.400 683.500 83.600 ;
        RECT 684.500 76.400 685.100 123.600 ;
        RECT 686.000 109.600 686.800 110.400 ;
        RECT 687.600 109.600 688.400 110.400 ;
        RECT 686.100 98.400 686.700 109.600 ;
        RECT 687.700 98.400 688.300 109.600 ;
        RECT 686.000 97.600 686.800 98.400 ;
        RECT 687.600 97.600 688.400 98.400 ;
        RECT 684.400 75.600 685.200 76.400 ;
        RECT 684.400 73.600 685.200 74.400 ;
        RECT 682.800 57.600 683.600 58.400 ;
        RECT 681.200 49.600 682.000 50.400 ;
        RECT 684.500 46.400 685.100 73.600 ;
        RECT 686.000 55.600 686.800 56.400 ;
        RECT 686.100 52.400 686.700 55.600 ;
        RECT 687.600 53.600 688.400 54.400 ;
        RECT 686.000 51.600 686.800 52.400 ;
        RECT 681.200 45.600 682.000 46.400 ;
        RECT 684.400 45.600 685.200 46.400 ;
        RECT 679.600 43.600 680.400 44.400 ;
        RECT 681.300 38.400 681.900 45.600 ;
        RECT 681.200 37.600 682.000 38.400 ;
        RECT 684.400 33.600 685.200 34.400 ;
        RECT 676.400 31.800 677.200 32.600 ;
        RECT 683.000 31.800 683.800 32.600 ;
        RECT 671.600 29.600 672.400 30.400 ;
        RECT 674.800 29.600 675.600 30.400 ;
        RECT 676.400 28.400 677.000 31.800 ;
        RECT 680.400 28.400 681.200 28.600 ;
        RECT 673.200 27.600 674.000 28.400 ;
        RECT 674.800 27.600 675.600 28.400 ;
        RECT 676.400 27.800 681.200 28.400 ;
        RECT 673.300 26.400 673.900 27.600 ;
        RECT 676.400 27.000 677.000 27.800 ;
        RECT 677.800 27.000 678.600 27.200 ;
        RECT 681.200 27.000 682.000 27.200 ;
        RECT 683.200 27.000 683.800 31.800 ;
        RECT 684.500 28.400 685.100 33.600 ;
        RECT 684.400 27.600 685.200 28.400 ;
        RECT 673.200 25.600 674.000 26.400 ;
        RECT 676.400 26.200 677.200 27.000 ;
        RECT 677.800 26.400 682.000 27.000 ;
        RECT 683.000 26.200 683.800 27.000 ;
        RECT 687.700 26.400 688.300 53.600 ;
        RECT 687.600 25.600 688.400 26.400 ;
        RECT 681.200 23.600 682.000 24.400 ;
        RECT 681.300 18.400 681.900 23.600 ;
        RECT 670.000 13.600 670.800 14.400 ;
        RECT 670.100 12.400 670.700 13.600 ;
        RECT 670.000 11.600 670.800 12.400 ;
        RECT 673.200 11.600 674.000 12.400 ;
        RECT 676.400 6.200 677.200 17.800 ;
        RECT 681.200 17.600 682.000 18.400 ;
        RECT 679.600 10.200 680.400 15.800 ;
        RECT 687.700 14.400 688.300 25.600 ;
        RECT 687.600 13.600 688.400 14.400 ;
        RECT 684.400 11.600 685.200 12.400 ;
        RECT 681.200 9.600 682.000 10.400 ;
      LAYER via2 ;
        RECT 14.000 429.600 14.800 430.400 ;
        RECT 90.800 189.600 91.600 190.400 ;
        RECT 167.600 149.600 168.400 150.400 ;
        RECT 156.400 109.600 157.200 110.400 ;
        RECT 84.400 13.600 85.200 14.400 ;
        RECT 270.000 229.600 270.800 230.400 ;
        RECT 446.000 469.600 446.800 470.400 ;
        RECT 492.400 491.600 493.200 492.400 ;
        RECT 230.000 187.600 230.800 188.400 ;
        RECT 159.600 29.600 160.400 30.400 ;
        RECT 303.600 147.600 304.400 148.400 ;
        RECT 326.000 267.600 326.800 268.400 ;
        RECT 338.800 187.600 339.600 188.400 ;
        RECT 591.600 389.600 592.400 390.400 ;
        RECT 545.200 269.600 546.000 270.400 ;
        RECT 450.800 211.600 451.600 212.400 ;
        RECT 412.400 13.600 413.200 14.400 ;
        RECT 612.400 211.600 613.200 212.400 ;
        RECT 538.800 69.600 539.600 70.400 ;
        RECT 673.200 309.600 674.000 310.400 ;
      LAYER metal3 ;
        RECT 631.600 498.300 632.400 498.400 ;
        RECT 671.600 498.300 672.400 498.400 ;
        RECT 631.600 497.700 672.400 498.300 ;
        RECT 631.600 497.600 632.400 497.700 ;
        RECT 671.600 497.600 672.400 497.700 ;
        RECT 86.000 496.300 86.800 496.400 ;
        RECT 161.200 496.300 162.000 496.400 ;
        RECT 86.000 495.700 162.000 496.300 ;
        RECT 86.000 495.600 86.800 495.700 ;
        RECT 161.200 495.600 162.000 495.700 ;
        RECT 183.600 496.300 184.400 496.400 ;
        RECT 222.000 496.300 222.800 496.400 ;
        RECT 239.600 496.300 240.400 496.400 ;
        RECT 314.800 496.300 315.600 496.400 ;
        RECT 362.800 496.300 363.600 496.400 ;
        RECT 183.600 495.700 240.400 496.300 ;
        RECT 183.600 495.600 184.400 495.700 ;
        RECT 222.000 495.600 222.800 495.700 ;
        RECT 239.600 495.600 240.400 495.700 ;
        RECT 292.500 495.700 363.600 496.300 ;
        RECT 292.500 494.400 293.100 495.700 ;
        RECT 314.800 495.600 315.600 495.700 ;
        RECT 362.800 495.600 363.600 495.700 ;
        RECT 386.800 496.300 387.600 496.400 ;
        RECT 430.000 496.300 430.800 496.400 ;
        RECT 386.800 495.700 430.800 496.300 ;
        RECT 386.800 495.600 387.600 495.700 ;
        RECT 430.000 495.600 430.800 495.700 ;
        RECT 462.000 496.300 462.800 496.400 ;
        RECT 508.400 496.300 509.200 496.400 ;
        RECT 462.000 495.700 509.200 496.300 ;
        RECT 462.000 495.600 462.800 495.700 ;
        RECT 508.400 495.600 509.200 495.700 ;
        RECT 511.600 496.300 512.400 496.400 ;
        RECT 532.400 496.300 533.200 496.400 ;
        RECT 511.600 495.700 533.200 496.300 ;
        RECT 511.600 495.600 512.400 495.700 ;
        RECT 532.400 495.600 533.200 495.700 ;
        RECT 567.600 496.300 568.400 496.400 ;
        RECT 578.800 496.300 579.600 496.400 ;
        RECT 606.000 496.300 606.800 496.400 ;
        RECT 668.400 496.300 669.200 496.400 ;
        RECT 567.600 495.700 669.200 496.300 ;
        RECT 567.600 495.600 568.400 495.700 ;
        RECT 578.800 495.600 579.600 495.700 ;
        RECT 606.000 495.600 606.800 495.700 ;
        RECT 668.400 495.600 669.200 495.700 ;
        RECT 14.000 494.300 14.800 494.400 ;
        RECT 34.800 494.300 35.600 494.400 ;
        RECT 14.000 493.700 35.600 494.300 ;
        RECT 14.000 493.600 14.800 493.700 ;
        RECT 34.800 493.600 35.600 493.700 ;
        RECT 58.800 494.300 59.600 494.400 ;
        RECT 87.600 494.300 88.400 494.400 ;
        RECT 58.800 493.700 88.400 494.300 ;
        RECT 58.800 493.600 59.600 493.700 ;
        RECT 87.600 493.600 88.400 493.700 ;
        RECT 110.000 494.300 110.800 494.400 ;
        RECT 148.400 494.300 149.200 494.400 ;
        RECT 110.000 493.700 149.200 494.300 ;
        RECT 110.000 493.600 110.800 493.700 ;
        RECT 148.400 493.600 149.200 493.700 ;
        RECT 161.200 494.300 162.000 494.400 ;
        RECT 201.200 494.300 202.000 494.400 ;
        RECT 161.200 493.700 202.000 494.300 ;
        RECT 161.200 493.600 162.000 493.700 ;
        RECT 201.200 493.600 202.000 493.700 ;
        RECT 204.400 494.300 205.200 494.400 ;
        RECT 225.200 494.300 226.000 494.400 ;
        RECT 204.400 493.700 226.000 494.300 ;
        RECT 204.400 493.600 205.200 493.700 ;
        RECT 225.200 493.600 226.000 493.700 ;
        RECT 249.200 494.300 250.000 494.400 ;
        RECT 274.800 494.300 275.600 494.400 ;
        RECT 292.400 494.300 293.200 494.400 ;
        RECT 249.200 493.700 293.200 494.300 ;
        RECT 249.200 493.600 250.000 493.700 ;
        RECT 274.800 493.600 275.600 493.700 ;
        RECT 292.400 493.600 293.200 493.700 ;
        RECT 303.600 494.300 304.400 494.400 ;
        RECT 334.000 494.300 334.800 494.400 ;
        RECT 303.600 493.700 334.800 494.300 ;
        RECT 303.600 493.600 304.400 493.700 ;
        RECT 334.000 493.600 334.800 493.700 ;
        RECT 345.200 494.300 346.000 494.400 ;
        RECT 366.000 494.300 366.800 494.400 ;
        RECT 345.200 493.700 366.800 494.300 ;
        RECT 345.200 493.600 346.000 493.700 ;
        RECT 366.000 493.600 366.800 493.700 ;
        RECT 406.000 493.600 406.800 494.400 ;
        RECT 433.200 494.300 434.000 494.400 ;
        RECT 439.600 494.300 440.400 494.400 ;
        RECT 433.200 493.700 440.400 494.300 ;
        RECT 433.200 493.600 434.000 493.700 ;
        RECT 439.600 493.600 440.400 493.700 ;
        RECT 465.200 494.300 466.000 494.400 ;
        RECT 476.400 494.300 477.200 494.400 ;
        RECT 465.200 493.700 477.200 494.300 ;
        RECT 465.200 493.600 466.000 493.700 ;
        RECT 476.400 493.600 477.200 493.700 ;
        RECT 529.200 494.300 530.000 494.400 ;
        RECT 538.800 494.300 539.600 494.400 ;
        RECT 545.200 494.300 546.000 494.400 ;
        RECT 529.200 493.700 546.000 494.300 ;
        RECT 529.200 493.600 530.000 493.700 ;
        RECT 538.800 493.600 539.600 493.700 ;
        RECT 545.200 493.600 546.000 493.700 ;
        RECT 585.200 494.300 586.000 494.400 ;
        RECT 625.200 494.300 626.000 494.400 ;
        RECT 585.200 493.700 626.000 494.300 ;
        RECT 585.200 493.600 586.000 493.700 ;
        RECT 625.200 493.600 626.000 493.700 ;
        RECT 25.200 492.300 26.000 492.400 ;
        RECT 49.200 492.300 50.000 492.400 ;
        RECT 25.200 491.700 50.000 492.300 ;
        RECT 25.200 491.600 26.000 491.700 ;
        RECT 49.200 491.600 50.000 491.700 ;
        RECT 127.600 492.300 128.400 492.400 ;
        RECT 135.600 492.300 136.400 492.400 ;
        RECT 127.600 491.700 136.400 492.300 ;
        RECT 127.600 491.600 128.400 491.700 ;
        RECT 135.600 491.600 136.400 491.700 ;
        RECT 166.000 492.300 166.800 492.400 ;
        RECT 186.800 492.300 187.600 492.400 ;
        RECT 166.000 491.700 187.600 492.300 ;
        RECT 166.000 491.600 166.800 491.700 ;
        RECT 186.800 491.600 187.600 491.700 ;
        RECT 198.000 492.300 198.800 492.400 ;
        RECT 214.000 492.300 214.800 492.400 ;
        RECT 198.000 491.700 214.800 492.300 ;
        RECT 198.000 491.600 198.800 491.700 ;
        RECT 214.000 491.600 214.800 491.700 ;
        RECT 236.400 492.300 237.200 492.400 ;
        RECT 262.000 492.300 262.800 492.400 ;
        RECT 236.400 491.700 262.800 492.300 ;
        RECT 236.400 491.600 237.200 491.700 ;
        RECT 262.000 491.600 262.800 491.700 ;
        RECT 290.800 492.300 291.600 492.400 ;
        RECT 302.000 492.300 302.800 492.400 ;
        RECT 290.800 491.700 302.800 492.300 ;
        RECT 290.800 491.600 291.600 491.700 ;
        RECT 302.000 491.600 302.800 491.700 ;
        RECT 322.800 492.300 323.600 492.400 ;
        RECT 354.800 492.300 355.600 492.400 ;
        RECT 322.800 491.700 355.600 492.300 ;
        RECT 322.800 491.600 323.600 491.700 ;
        RECT 354.800 491.600 355.600 491.700 ;
        RECT 362.800 492.300 363.600 492.400 ;
        RECT 402.800 492.300 403.600 492.400 ;
        RECT 362.800 491.700 403.600 492.300 ;
        RECT 406.100 492.300 406.700 493.600 ;
        RECT 436.400 492.300 437.200 492.400 ;
        RECT 406.100 491.700 437.200 492.300 ;
        RECT 362.800 491.600 363.600 491.700 ;
        RECT 402.800 491.600 403.600 491.700 ;
        RECT 436.400 491.600 437.200 491.700 ;
        RECT 486.000 492.300 486.800 492.400 ;
        RECT 492.400 492.300 493.200 492.400 ;
        RECT 526.000 492.300 526.800 492.400 ;
        RECT 486.000 491.700 526.800 492.300 ;
        RECT 486.000 491.600 486.800 491.700 ;
        RECT 492.400 491.600 493.200 491.700 ;
        RECT 526.000 491.600 526.800 491.700 ;
        RECT 542.000 492.300 542.800 492.400 ;
        RECT 570.800 492.300 571.600 492.400 ;
        RECT 542.000 491.700 571.600 492.300 ;
        RECT 542.000 491.600 542.800 491.700 ;
        RECT 570.800 491.600 571.600 491.700 ;
        RECT 586.800 492.300 587.600 492.400 ;
        RECT 602.800 492.300 603.600 492.400 ;
        RECT 586.800 491.700 603.600 492.300 ;
        RECT 586.800 491.600 587.600 491.700 ;
        RECT 602.800 491.600 603.600 491.700 ;
        RECT 36.400 490.300 37.200 490.400 ;
        RECT 39.600 490.300 40.400 490.400 ;
        RECT 36.400 489.700 40.400 490.300 ;
        RECT 36.400 489.600 37.200 489.700 ;
        RECT 39.600 489.600 40.400 489.700 ;
        RECT 41.200 490.300 42.000 490.400 ;
        RECT 46.000 490.300 46.800 490.400 ;
        RECT 86.000 490.300 86.800 490.400 ;
        RECT 41.200 489.700 86.800 490.300 ;
        RECT 41.200 489.600 42.000 489.700 ;
        RECT 46.000 489.600 46.800 489.700 ;
        RECT 86.000 489.600 86.800 489.700 ;
        RECT 94.000 490.300 94.800 490.400 ;
        RECT 151.600 490.300 152.400 490.400 ;
        RECT 94.000 489.700 152.400 490.300 ;
        RECT 94.000 489.600 94.800 489.700 ;
        RECT 151.600 489.600 152.400 489.700 ;
        RECT 156.400 490.300 157.200 490.400 ;
        RECT 164.400 490.300 165.200 490.400 ;
        RECT 156.400 489.700 165.200 490.300 ;
        RECT 156.400 489.600 157.200 489.700 ;
        RECT 164.400 489.600 165.200 489.700 ;
        RECT 529.200 490.300 530.000 490.400 ;
        RECT 538.800 490.300 539.600 490.400 ;
        RECT 529.200 489.700 539.600 490.300 ;
        RECT 529.200 489.600 530.000 489.700 ;
        RECT 538.800 489.600 539.600 489.700 ;
        RECT 87.600 488.300 88.400 488.400 ;
        RECT 95.600 488.300 96.400 488.400 ;
        RECT 87.600 487.700 96.400 488.300 ;
        RECT 87.600 487.600 88.400 487.700 ;
        RECT 95.600 487.600 96.400 487.700 ;
        RECT 154.800 488.300 155.600 488.400 ;
        RECT 167.600 488.300 168.400 488.400 ;
        RECT 154.800 487.700 168.400 488.300 ;
        RECT 154.800 487.600 155.600 487.700 ;
        RECT 167.600 487.600 168.400 487.700 ;
        RECT 522.800 488.300 523.600 488.400 ;
        RECT 559.600 488.300 560.400 488.400 ;
        RECT 522.800 487.700 560.400 488.300 ;
        RECT 522.800 487.600 523.600 487.700 ;
        RECT 559.600 487.600 560.400 487.700 ;
        RECT 70.000 486.300 70.800 486.400 ;
        RECT 175.600 486.300 176.400 486.400 ;
        RECT 70.000 485.700 176.400 486.300 ;
        RECT 70.000 485.600 70.800 485.700 ;
        RECT 175.600 485.600 176.400 485.700 ;
        RECT 511.600 486.300 512.400 486.400 ;
        RECT 535.600 486.300 536.400 486.400 ;
        RECT 511.600 485.700 536.400 486.300 ;
        RECT 511.600 485.600 512.400 485.700 ;
        RECT 535.600 485.600 536.400 485.700 ;
        RECT 78.000 484.300 78.800 484.400 ;
        RECT 89.200 484.300 90.000 484.400 ;
        RECT 78.000 483.700 90.000 484.300 ;
        RECT 78.000 483.600 78.800 483.700 ;
        RECT 89.200 483.600 90.000 483.700 ;
        RECT 122.800 484.300 123.600 484.400 ;
        RECT 134.000 484.300 134.800 484.400 ;
        RECT 137.200 484.300 138.000 484.400 ;
        RECT 122.800 483.700 138.000 484.300 ;
        RECT 122.800 483.600 123.600 483.700 ;
        RECT 134.000 483.600 134.800 483.700 ;
        RECT 137.200 483.600 138.000 483.700 ;
        RECT 159.600 484.300 160.400 484.400 ;
        RECT 206.000 484.300 206.800 484.400 ;
        RECT 159.600 483.700 206.800 484.300 ;
        RECT 159.600 483.600 160.400 483.700 ;
        RECT 206.000 483.600 206.800 483.700 ;
        RECT 330.800 484.300 331.600 484.400 ;
        RECT 334.000 484.300 334.800 484.400 ;
        RECT 330.800 483.700 334.800 484.300 ;
        RECT 330.800 483.600 331.600 483.700 ;
        RECT 334.000 483.600 334.800 483.700 ;
        RECT 401.200 484.300 402.000 484.400 ;
        RECT 406.000 484.300 406.800 484.400 ;
        RECT 401.200 483.700 406.800 484.300 ;
        RECT 401.200 483.600 402.000 483.700 ;
        RECT 406.000 483.600 406.800 483.700 ;
        RECT 548.400 484.300 549.200 484.400 ;
        RECT 551.600 484.300 552.400 484.400 ;
        RECT 548.400 483.700 552.400 484.300 ;
        RECT 548.400 483.600 549.200 483.700 ;
        RECT 551.600 483.600 552.400 483.700 ;
        RECT 634.800 484.300 635.600 484.400 ;
        RECT 652.400 484.300 653.200 484.400 ;
        RECT 634.800 483.700 653.200 484.300 ;
        RECT 634.800 483.600 635.600 483.700 ;
        RECT 652.400 483.600 653.200 483.700 ;
        RECT 10.800 482.300 11.600 482.400 ;
        RECT 14.000 482.300 14.800 482.400 ;
        RECT 10.800 481.700 14.800 482.300 ;
        RECT 10.800 481.600 11.600 481.700 ;
        RECT 14.000 481.600 14.800 481.700 ;
        RECT 148.400 482.300 149.200 482.400 ;
        RECT 252.400 482.300 253.200 482.400 ;
        RECT 281.200 482.300 282.000 482.400 ;
        RECT 148.400 481.700 282.000 482.300 ;
        RECT 148.400 481.600 149.200 481.700 ;
        RECT 252.400 481.600 253.200 481.700 ;
        RECT 281.200 481.600 282.000 481.700 ;
        RECT 332.400 482.300 333.200 482.400 ;
        RECT 346.800 482.300 347.600 482.400 ;
        RECT 359.600 482.300 360.400 482.400 ;
        RECT 332.400 481.700 360.400 482.300 ;
        RECT 332.400 481.600 333.200 481.700 ;
        RECT 346.800 481.600 347.600 481.700 ;
        RECT 359.600 481.600 360.400 481.700 ;
        RECT 500.400 482.300 501.200 482.400 ;
        RECT 503.600 482.300 504.400 482.400 ;
        RECT 500.400 481.700 504.400 482.300 ;
        RECT 500.400 481.600 501.200 481.700 ;
        RECT 503.600 481.600 504.400 481.700 ;
        RECT 409.200 478.300 410.000 478.400 ;
        RECT 422.000 478.300 422.800 478.400 ;
        RECT 409.200 477.700 422.800 478.300 ;
        RECT 409.200 477.600 410.000 477.700 ;
        RECT 422.000 477.600 422.800 477.700 ;
        RECT 426.800 478.300 427.600 478.400 ;
        RECT 433.200 478.300 434.000 478.400 ;
        RECT 527.600 478.300 528.400 478.400 ;
        RECT 426.800 477.700 528.400 478.300 ;
        RECT 426.800 477.600 427.600 477.700 ;
        RECT 433.200 477.600 434.000 477.700 ;
        RECT 527.600 477.600 528.400 477.700 ;
        RECT 39.600 476.300 40.400 476.400 ;
        RECT 94.000 476.300 94.800 476.400 ;
        RECT 39.600 475.700 94.800 476.300 ;
        RECT 39.600 475.600 40.400 475.700 ;
        RECT 94.000 475.600 94.800 475.700 ;
        RECT 71.600 474.300 72.400 474.400 ;
        RECT 78.000 474.300 78.800 474.400 ;
        RECT 71.600 473.700 78.800 474.300 ;
        RECT 71.600 473.600 72.400 473.700 ;
        RECT 78.000 473.600 78.800 473.700 ;
        RECT 84.400 474.300 85.200 474.400 ;
        RECT 98.800 474.300 99.600 474.400 ;
        RECT 84.400 473.700 99.600 474.300 ;
        RECT 84.400 473.600 85.200 473.700 ;
        RECT 98.800 473.600 99.600 473.700 ;
        RECT 164.400 474.300 165.200 474.400 ;
        RECT 167.600 474.300 168.400 474.400 ;
        RECT 164.400 473.700 168.400 474.300 ;
        RECT 164.400 473.600 165.200 473.700 ;
        RECT 167.600 473.600 168.400 473.700 ;
        RECT 326.000 474.300 326.800 474.400 ;
        RECT 377.200 474.300 378.000 474.400 ;
        RECT 326.000 473.700 378.000 474.300 ;
        RECT 326.000 473.600 326.800 473.700 ;
        RECT 377.200 473.600 378.000 473.700 ;
        RECT 647.600 474.300 648.400 474.400 ;
        RECT 666.800 474.300 667.600 474.400 ;
        RECT 647.600 473.700 667.600 474.300 ;
        RECT 647.600 473.600 648.400 473.700 ;
        RECT 666.800 473.600 667.600 473.700 ;
        RECT 33.200 472.300 34.000 472.400 ;
        RECT 36.400 472.300 37.200 472.400 ;
        RECT 42.800 472.300 43.600 472.400 ;
        RECT 33.200 471.700 43.600 472.300 ;
        RECT 33.200 471.600 34.000 471.700 ;
        RECT 36.400 471.600 37.200 471.700 ;
        RECT 42.800 471.600 43.600 471.700 ;
        RECT 68.400 472.300 69.200 472.400 ;
        RECT 132.400 472.300 133.200 472.400 ;
        RECT 68.400 471.700 133.200 472.300 ;
        RECT 68.400 471.600 69.200 471.700 ;
        RECT 132.400 471.600 133.200 471.700 ;
        RECT 172.400 472.300 173.200 472.400 ;
        RECT 180.400 472.300 181.200 472.400 ;
        RECT 172.400 471.700 181.200 472.300 ;
        RECT 172.400 471.600 173.200 471.700 ;
        RECT 180.400 471.600 181.200 471.700 ;
        RECT 276.400 471.600 277.200 472.400 ;
        RECT 316.400 472.300 317.200 472.400 ;
        RECT 319.600 472.300 320.400 472.400 ;
        RECT 316.400 471.700 320.400 472.300 ;
        RECT 316.400 471.600 317.200 471.700 ;
        RECT 319.600 471.600 320.400 471.700 ;
        RECT 330.800 472.300 331.600 472.400 ;
        RECT 358.000 472.300 358.800 472.400 ;
        RECT 330.800 471.700 358.800 472.300 ;
        RECT 330.800 471.600 331.600 471.700 ;
        RECT 358.000 471.600 358.800 471.700 ;
        RECT 366.000 472.300 366.800 472.400 ;
        RECT 372.400 472.300 373.200 472.400 ;
        RECT 366.000 471.700 373.200 472.300 ;
        RECT 366.000 471.600 366.800 471.700 ;
        RECT 372.400 471.600 373.200 471.700 ;
        RECT 375.600 472.300 376.400 472.400 ;
        RECT 398.000 472.300 398.800 472.400 ;
        RECT 375.600 471.700 398.800 472.300 ;
        RECT 375.600 471.600 376.400 471.700 ;
        RECT 398.000 471.600 398.800 471.700 ;
        RECT 420.400 472.300 421.200 472.400 ;
        RECT 428.400 472.300 429.200 472.400 ;
        RECT 420.400 471.700 429.200 472.300 ;
        RECT 420.400 471.600 421.200 471.700 ;
        RECT 428.400 471.600 429.200 471.700 ;
        RECT 526.000 472.300 526.800 472.400 ;
        RECT 530.800 472.300 531.600 472.400 ;
        RECT 526.000 471.700 531.600 472.300 ;
        RECT 526.000 471.600 526.800 471.700 ;
        RECT 530.800 471.600 531.600 471.700 ;
        RECT 583.600 472.300 584.400 472.400 ;
        RECT 601.200 472.300 602.000 472.400 ;
        RECT 583.600 471.700 602.000 472.300 ;
        RECT 583.600 471.600 584.400 471.700 ;
        RECT 601.200 471.600 602.000 471.700 ;
        RECT 609.200 472.300 610.000 472.400 ;
        RECT 617.200 472.300 618.000 472.400 ;
        RECT 634.800 472.300 635.600 472.400 ;
        RECT 609.200 471.700 635.600 472.300 ;
        RECT 609.200 471.600 610.000 471.700 ;
        RECT 617.200 471.600 618.000 471.700 ;
        RECT 634.800 471.600 635.600 471.700 ;
        RECT 652.400 472.300 653.200 472.400 ;
        RECT 654.000 472.300 654.800 472.400 ;
        RECT 652.400 471.700 654.800 472.300 ;
        RECT 652.400 471.600 653.200 471.700 ;
        RECT 654.000 471.600 654.800 471.700 ;
        RECT 73.200 470.300 74.000 470.400 ;
        RECT 82.800 470.300 83.600 470.400 ;
        RECT 73.200 469.700 83.600 470.300 ;
        RECT 73.200 469.600 74.000 469.700 ;
        RECT 82.800 469.600 83.600 469.700 ;
        RECT 105.200 470.300 106.000 470.400 ;
        RECT 126.000 470.300 126.800 470.400 ;
        RECT 105.200 469.700 126.800 470.300 ;
        RECT 105.200 469.600 106.000 469.700 ;
        RECT 126.000 469.600 126.800 469.700 ;
        RECT 130.800 470.300 131.600 470.400 ;
        RECT 138.800 470.300 139.600 470.400 ;
        RECT 162.800 470.300 163.600 470.400 ;
        RECT 130.800 469.700 163.600 470.300 ;
        RECT 130.800 469.600 131.600 469.700 ;
        RECT 138.800 469.600 139.600 469.700 ;
        RECT 162.800 469.600 163.600 469.700 ;
        RECT 169.200 470.300 170.000 470.400 ;
        RECT 178.800 470.300 179.600 470.400 ;
        RECT 194.800 470.300 195.600 470.400 ;
        RECT 169.200 469.700 195.600 470.300 ;
        RECT 169.200 469.600 170.000 469.700 ;
        RECT 178.800 469.600 179.600 469.700 ;
        RECT 194.800 469.600 195.600 469.700 ;
        RECT 215.600 470.300 216.400 470.400 ;
        RECT 241.200 470.300 242.000 470.400 ;
        RECT 215.600 469.700 242.000 470.300 ;
        RECT 215.600 469.600 216.400 469.700 ;
        RECT 241.200 469.600 242.000 469.700 ;
        RECT 273.200 470.300 274.000 470.400 ;
        RECT 276.400 470.300 277.200 470.400 ;
        RECT 273.200 469.700 277.200 470.300 ;
        RECT 273.200 469.600 274.000 469.700 ;
        RECT 276.400 469.600 277.200 469.700 ;
        RECT 300.400 470.300 301.200 470.400 ;
        RECT 327.600 470.300 328.400 470.400 ;
        RECT 335.600 470.300 336.400 470.400 ;
        RECT 346.800 470.300 347.600 470.400 ;
        RECT 300.400 469.700 347.600 470.300 ;
        RECT 300.400 469.600 301.200 469.700 ;
        RECT 327.600 469.600 328.400 469.700 ;
        RECT 335.600 469.600 336.400 469.700 ;
        RECT 346.800 469.600 347.600 469.700 ;
        RECT 348.400 470.300 349.200 470.400 ;
        RECT 353.200 470.300 354.000 470.400 ;
        RECT 348.400 469.700 354.000 470.300 ;
        RECT 348.400 469.600 349.200 469.700 ;
        RECT 353.200 469.600 354.000 469.700 ;
        RECT 420.400 470.300 421.200 470.400 ;
        RECT 423.600 470.300 424.400 470.400 ;
        RECT 420.400 469.700 424.400 470.300 ;
        RECT 420.400 469.600 421.200 469.700 ;
        RECT 423.600 469.600 424.400 469.700 ;
        RECT 430.000 470.300 430.800 470.400 ;
        RECT 446.000 470.300 446.800 470.400 ;
        RECT 430.000 469.700 446.800 470.300 ;
        RECT 430.000 469.600 430.800 469.700 ;
        RECT 446.000 469.600 446.800 469.700 ;
        RECT 550.000 470.300 550.800 470.400 ;
        RECT 578.800 470.300 579.600 470.400 ;
        RECT 550.000 469.700 579.600 470.300 ;
        RECT 550.000 469.600 550.800 469.700 ;
        RECT 578.800 469.600 579.600 469.700 ;
        RECT 599.600 470.300 600.400 470.400 ;
        RECT 606.000 470.300 606.800 470.400 ;
        RECT 612.400 470.300 613.200 470.400 ;
        RECT 622.000 470.300 622.800 470.400 ;
        RECT 599.600 469.700 622.800 470.300 ;
        RECT 599.600 469.600 600.400 469.700 ;
        RECT 606.000 469.600 606.800 469.700 ;
        RECT 612.400 469.600 613.200 469.700 ;
        RECT 622.000 469.600 622.800 469.700 ;
        RECT 626.800 470.300 627.600 470.400 ;
        RECT 634.800 470.300 635.600 470.400 ;
        RECT 626.800 469.700 635.600 470.300 ;
        RECT 626.800 469.600 627.600 469.700 ;
        RECT 634.800 469.600 635.600 469.700 ;
        RECT 644.400 470.300 645.200 470.400 ;
        RECT 655.600 470.300 656.400 470.400 ;
        RECT 644.400 469.700 656.400 470.300 ;
        RECT 644.400 469.600 645.200 469.700 ;
        RECT 655.600 469.600 656.400 469.700 ;
        RECT 670.000 469.600 670.800 470.400 ;
        RECT 22.000 468.300 22.800 468.400 ;
        RECT 38.000 468.300 38.800 468.400 ;
        RECT 22.000 467.700 38.800 468.300 ;
        RECT 22.000 467.600 22.800 467.700 ;
        RECT 38.000 467.600 38.800 467.700 ;
        RECT 46.000 468.300 46.800 468.400 ;
        RECT 92.400 468.300 93.200 468.400 ;
        RECT 94.000 468.300 94.800 468.400 ;
        RECT 159.600 468.300 160.400 468.400 ;
        RECT 46.000 467.700 160.400 468.300 ;
        RECT 46.000 467.600 46.800 467.700 ;
        RECT 92.400 467.600 93.200 467.700 ;
        RECT 94.000 467.600 94.800 467.700 ;
        RECT 159.600 467.600 160.400 467.700 ;
        RECT 177.200 468.300 178.000 468.400 ;
        RECT 180.400 468.300 181.200 468.400 ;
        RECT 230.000 468.300 230.800 468.400 ;
        RECT 177.200 467.700 230.800 468.300 ;
        RECT 177.200 467.600 178.000 467.700 ;
        RECT 180.400 467.600 181.200 467.700 ;
        RECT 230.000 467.600 230.800 467.700 ;
        RECT 231.600 468.300 232.400 468.400 ;
        RECT 252.400 468.300 253.200 468.400 ;
        RECT 231.600 467.700 253.200 468.300 ;
        RECT 231.600 467.600 232.400 467.700 ;
        RECT 252.400 467.600 253.200 467.700 ;
        RECT 310.000 468.300 310.800 468.400 ;
        RECT 324.400 468.300 325.200 468.400 ;
        RECT 332.400 468.300 333.200 468.400 ;
        RECT 310.000 467.700 321.900 468.300 ;
        RECT 310.000 467.600 310.800 467.700 ;
        RECT 321.300 466.400 321.900 467.700 ;
        RECT 324.400 467.700 333.200 468.300 ;
        RECT 324.400 467.600 325.200 467.700 ;
        RECT 332.400 467.600 333.200 467.700 ;
        RECT 343.600 468.300 344.400 468.400 ;
        RECT 361.200 468.300 362.000 468.400 ;
        RECT 343.600 467.700 362.000 468.300 ;
        RECT 343.600 467.600 344.400 467.700 ;
        RECT 361.200 467.600 362.000 467.700 ;
        RECT 390.000 468.300 390.800 468.400 ;
        RECT 415.600 468.300 416.400 468.400 ;
        RECT 390.000 467.700 416.400 468.300 ;
        RECT 390.000 467.600 390.800 467.700 ;
        RECT 415.600 467.600 416.400 467.700 ;
        RECT 436.400 468.300 437.200 468.400 ;
        RECT 465.200 468.300 466.000 468.400 ;
        RECT 436.400 467.700 466.000 468.300 ;
        RECT 436.400 467.600 437.200 467.700 ;
        RECT 465.200 467.600 466.000 467.700 ;
        RECT 492.400 468.300 493.200 468.400 ;
        RECT 542.000 468.300 542.800 468.400 ;
        RECT 492.400 467.700 542.800 468.300 ;
        RECT 492.400 467.600 493.200 467.700 ;
        RECT 542.000 467.600 542.800 467.700 ;
        RECT 569.200 468.300 570.000 468.400 ;
        RECT 577.200 468.300 578.000 468.400 ;
        RECT 569.200 467.700 578.000 468.300 ;
        RECT 569.200 467.600 570.000 467.700 ;
        RECT 577.200 467.600 578.000 467.700 ;
        RECT 585.200 468.300 586.000 468.400 ;
        RECT 596.400 468.300 597.200 468.400 ;
        RECT 585.200 467.700 597.200 468.300 ;
        RECT 585.200 467.600 586.000 467.700 ;
        RECT 596.400 467.600 597.200 467.700 ;
        RECT 601.200 468.300 602.000 468.400 ;
        RECT 609.200 468.300 610.000 468.400 ;
        RECT 601.200 467.700 610.000 468.300 ;
        RECT 634.900 468.300 635.500 469.600 ;
        RECT 644.400 468.300 645.200 468.400 ;
        RECT 634.900 467.700 645.200 468.300 ;
        RECT 601.200 467.600 602.000 467.700 ;
        RECT 609.200 467.600 610.000 467.700 ;
        RECT 644.400 467.600 645.200 467.700 ;
        RECT 650.800 468.300 651.600 468.400 ;
        RECT 657.200 468.300 658.000 468.400 ;
        RECT 650.800 467.700 658.000 468.300 ;
        RECT 650.800 467.600 651.600 467.700 ;
        RECT 657.200 467.600 658.000 467.700 ;
        RECT 674.800 468.300 675.600 468.400 ;
        RECT 681.200 468.300 682.000 468.400 ;
        RECT 674.800 467.700 682.000 468.300 ;
        RECT 674.800 467.600 675.600 467.700 ;
        RECT 681.200 467.600 682.000 467.700 ;
        RECT 71.600 466.300 72.400 466.400 ;
        RECT 76.400 466.300 77.200 466.400 ;
        RECT 71.600 465.700 77.200 466.300 ;
        RECT 71.600 465.600 72.400 465.700 ;
        RECT 76.400 465.600 77.200 465.700 ;
        RECT 82.800 466.300 83.600 466.400 ;
        RECT 111.600 466.300 112.400 466.400 ;
        RECT 82.800 465.700 112.400 466.300 ;
        RECT 82.800 465.600 83.600 465.700 ;
        RECT 111.600 465.600 112.400 465.700 ;
        RECT 124.400 466.300 125.200 466.400 ;
        RECT 129.200 466.300 130.000 466.400 ;
        RECT 124.400 465.700 130.000 466.300 ;
        RECT 124.400 465.600 125.200 465.700 ;
        RECT 129.200 465.600 130.000 465.700 ;
        RECT 164.400 466.300 165.200 466.400 ;
        RECT 174.000 466.300 174.800 466.400 ;
        RECT 183.600 466.300 184.400 466.400 ;
        RECT 164.400 465.700 184.400 466.300 ;
        RECT 164.400 465.600 165.200 465.700 ;
        RECT 174.000 465.600 174.800 465.700 ;
        RECT 183.600 465.600 184.400 465.700 ;
        RECT 279.600 466.300 280.400 466.400 ;
        RECT 294.000 466.300 294.800 466.400 ;
        RECT 279.600 465.700 294.800 466.300 ;
        RECT 279.600 465.600 280.400 465.700 ;
        RECT 294.000 465.600 294.800 465.700 ;
        RECT 298.800 466.300 299.600 466.400 ;
        RECT 310.000 466.300 310.800 466.400 ;
        RECT 298.800 465.700 310.800 466.300 ;
        RECT 298.800 465.600 299.600 465.700 ;
        RECT 310.000 465.600 310.800 465.700 ;
        RECT 321.200 466.300 322.000 466.400 ;
        RECT 340.400 466.300 341.200 466.400 ;
        RECT 343.600 466.300 344.400 466.400 ;
        RECT 321.200 465.700 344.400 466.300 ;
        RECT 321.200 465.600 322.000 465.700 ;
        RECT 340.400 465.600 341.200 465.700 ;
        RECT 343.600 465.600 344.400 465.700 ;
        RECT 346.800 466.300 347.600 466.400 ;
        RECT 353.200 466.300 354.000 466.400 ;
        RECT 370.800 466.300 371.600 466.400 ;
        RECT 382.000 466.300 382.800 466.400 ;
        RECT 346.800 465.700 382.800 466.300 ;
        RECT 346.800 465.600 347.600 465.700 ;
        RECT 353.200 465.600 354.000 465.700 ;
        RECT 370.800 465.600 371.600 465.700 ;
        RECT 382.000 465.600 382.800 465.700 ;
        RECT 423.600 466.300 424.400 466.400 ;
        RECT 454.000 466.300 454.800 466.400 ;
        RECT 423.600 465.700 454.800 466.300 ;
        RECT 423.600 465.600 424.400 465.700 ;
        RECT 454.000 465.600 454.800 465.700 ;
        RECT 474.800 466.300 475.600 466.400 ;
        RECT 484.400 466.300 485.200 466.400 ;
        RECT 492.400 466.300 493.200 466.400 ;
        RECT 474.800 465.700 493.200 466.300 ;
        RECT 474.800 465.600 475.600 465.700 ;
        RECT 484.400 465.600 485.200 465.700 ;
        RECT 492.400 465.600 493.200 465.700 ;
        RECT 495.600 466.300 496.400 466.400 ;
        RECT 508.400 466.300 509.200 466.400 ;
        RECT 513.200 466.300 514.000 466.400 ;
        RECT 495.600 465.700 514.000 466.300 ;
        RECT 495.600 465.600 496.400 465.700 ;
        RECT 508.400 465.600 509.200 465.700 ;
        RECT 513.200 465.600 514.000 465.700 ;
        RECT 518.000 466.300 518.800 466.400 ;
        RECT 559.600 466.300 560.400 466.400 ;
        RECT 567.600 466.300 568.400 466.400 ;
        RECT 575.600 466.300 576.400 466.400 ;
        RECT 518.000 465.700 576.400 466.300 ;
        RECT 518.000 465.600 518.800 465.700 ;
        RECT 559.600 465.600 560.400 465.700 ;
        RECT 567.600 465.600 568.400 465.700 ;
        RECT 575.600 465.600 576.400 465.700 ;
        RECT 577.200 466.300 578.000 466.400 ;
        RECT 590.000 466.300 590.800 466.400 ;
        RECT 577.200 465.700 590.800 466.300 ;
        RECT 577.200 465.600 578.000 465.700 ;
        RECT 590.000 465.600 590.800 465.700 ;
        RECT 610.800 466.300 611.600 466.400 ;
        RECT 620.400 466.300 621.200 466.400 ;
        RECT 631.600 466.300 632.400 466.400 ;
        RECT 636.400 466.300 637.200 466.400 ;
        RECT 639.600 466.300 640.400 466.400 ;
        RECT 610.800 465.700 640.400 466.300 ;
        RECT 610.800 465.600 611.600 465.700 ;
        RECT 620.400 465.600 621.200 465.700 ;
        RECT 631.600 465.600 632.400 465.700 ;
        RECT 636.400 465.600 637.200 465.700 ;
        RECT 639.600 465.600 640.400 465.700 ;
        RECT 641.200 466.300 642.000 466.400 ;
        RECT 649.200 466.300 650.000 466.400 ;
        RECT 641.200 465.700 650.000 466.300 ;
        RECT 641.200 465.600 642.000 465.700 ;
        RECT 649.200 465.600 650.000 465.700 ;
        RECT 58.800 464.300 59.600 464.400 ;
        RECT 68.400 464.300 69.200 464.400 ;
        RECT 58.800 463.700 69.200 464.300 ;
        RECT 58.800 463.600 59.600 463.700 ;
        RECT 68.400 463.600 69.200 463.700 ;
        RECT 81.200 464.300 82.000 464.400 ;
        RECT 98.800 464.300 99.600 464.400 ;
        RECT 81.200 463.700 99.600 464.300 ;
        RECT 81.200 463.600 82.000 463.700 ;
        RECT 98.800 463.600 99.600 463.700 ;
        RECT 127.600 464.300 128.400 464.400 ;
        RECT 134.000 464.300 134.800 464.400 ;
        RECT 127.600 463.700 134.800 464.300 ;
        RECT 127.600 463.600 128.400 463.700 ;
        RECT 134.000 463.600 134.800 463.700 ;
        RECT 140.400 464.300 141.200 464.400 ;
        RECT 146.800 464.300 147.600 464.400 ;
        RECT 140.400 463.700 147.600 464.300 ;
        RECT 140.400 463.600 141.200 463.700 ;
        RECT 146.800 463.600 147.600 463.700 ;
        RECT 156.400 464.300 157.200 464.400 ;
        RECT 161.200 464.300 162.000 464.400 ;
        RECT 182.000 464.300 182.800 464.400 ;
        RECT 156.400 463.700 182.800 464.300 ;
        RECT 156.400 463.600 157.200 463.700 ;
        RECT 161.200 463.600 162.000 463.700 ;
        RECT 182.000 463.600 182.800 463.700 ;
        RECT 338.800 464.300 339.600 464.400 ;
        RECT 343.600 464.300 344.400 464.400 ;
        RECT 338.800 463.700 344.400 464.300 ;
        RECT 338.800 463.600 339.600 463.700 ;
        RECT 343.600 463.600 344.400 463.700 ;
        RECT 434.800 464.300 435.600 464.400 ;
        RECT 518.000 464.300 518.800 464.400 ;
        RECT 434.800 463.700 518.800 464.300 ;
        RECT 434.800 463.600 435.600 463.700 ;
        RECT 518.000 463.600 518.800 463.700 ;
        RECT 550.000 464.300 550.800 464.400 ;
        RECT 553.200 464.300 554.000 464.400 ;
        RECT 550.000 463.700 554.000 464.300 ;
        RECT 590.100 464.300 590.700 465.600 ;
        RECT 634.800 464.300 635.600 464.400 ;
        RECT 642.800 464.300 643.600 464.400 ;
        RECT 590.100 463.700 643.600 464.300 ;
        RECT 550.000 463.600 550.800 463.700 ;
        RECT 553.200 463.600 554.000 463.700 ;
        RECT 634.800 463.600 635.600 463.700 ;
        RECT 642.800 463.600 643.600 463.700 ;
        RECT 658.800 464.300 659.600 464.400 ;
        RECT 673.200 464.300 674.000 464.400 ;
        RECT 658.800 463.700 674.000 464.300 ;
        RECT 658.800 463.600 659.600 463.700 ;
        RECT 673.200 463.600 674.000 463.700 ;
        RECT 86.000 462.300 86.800 462.400 ;
        RECT 100.400 462.300 101.200 462.400 ;
        RECT 119.600 462.300 120.400 462.400 ;
        RECT 86.000 461.700 120.400 462.300 ;
        RECT 86.000 461.600 86.800 461.700 ;
        RECT 100.400 461.600 101.200 461.700 ;
        RECT 119.600 461.600 120.400 461.700 ;
        RECT 129.200 462.300 130.000 462.400 ;
        RECT 150.000 462.300 150.800 462.400 ;
        RECT 129.200 461.700 150.800 462.300 ;
        RECT 129.200 461.600 130.000 461.700 ;
        RECT 150.000 461.600 150.800 461.700 ;
        RECT 198.000 462.300 198.800 462.400 ;
        RECT 220.400 462.300 221.200 462.400 ;
        RECT 198.000 461.700 221.200 462.300 ;
        RECT 198.000 461.600 198.800 461.700 ;
        RECT 220.400 461.600 221.200 461.700 ;
        RECT 319.600 462.300 320.400 462.400 ;
        RECT 350.000 462.300 350.800 462.400 ;
        RECT 319.600 461.700 350.800 462.300 ;
        RECT 319.600 461.600 320.400 461.700 ;
        RECT 350.000 461.600 350.800 461.700 ;
        RECT 359.600 462.300 360.400 462.400 ;
        RECT 386.800 462.300 387.600 462.400 ;
        RECT 359.600 461.700 387.600 462.300 ;
        RECT 359.600 461.600 360.400 461.700 ;
        RECT 386.800 461.600 387.600 461.700 ;
        RECT 393.200 462.300 394.000 462.400 ;
        RECT 454.000 462.300 454.800 462.400 ;
        RECT 462.000 462.300 462.800 462.400 ;
        RECT 393.200 461.700 462.800 462.300 ;
        RECT 393.200 461.600 394.000 461.700 ;
        RECT 454.000 461.600 454.800 461.700 ;
        RECT 462.000 461.600 462.800 461.700 ;
        RECT 593.200 462.300 594.000 462.400 ;
        RECT 610.800 462.300 611.600 462.400 ;
        RECT 593.200 461.700 611.600 462.300 ;
        RECT 593.200 461.600 594.000 461.700 ;
        RECT 610.800 461.600 611.600 461.700 ;
        RECT 617.200 462.300 618.000 462.400 ;
        RECT 622.000 462.300 622.800 462.400 ;
        RECT 631.600 462.300 632.400 462.400 ;
        RECT 617.200 461.700 632.400 462.300 ;
        RECT 617.200 461.600 618.000 461.700 ;
        RECT 622.000 461.600 622.800 461.700 ;
        RECT 631.600 461.600 632.400 461.700 ;
        RECT 18.800 460.300 19.600 460.400 ;
        RECT 55.600 460.300 56.400 460.400 ;
        RECT 84.400 460.300 85.200 460.400 ;
        RECT 18.800 459.700 85.200 460.300 ;
        RECT 18.800 459.600 19.600 459.700 ;
        RECT 55.600 459.600 56.400 459.700 ;
        RECT 84.400 459.600 85.200 459.700 ;
        RECT 281.200 460.300 282.000 460.400 ;
        RECT 295.600 460.300 296.400 460.400 ;
        RECT 281.200 459.700 296.400 460.300 ;
        RECT 281.200 459.600 282.000 459.700 ;
        RECT 295.600 459.600 296.400 459.700 ;
        RECT 350.000 460.300 350.800 460.400 ;
        RECT 370.800 460.300 371.600 460.400 ;
        RECT 390.000 460.300 390.800 460.400 ;
        RECT 350.000 459.700 390.800 460.300 ;
        RECT 350.000 459.600 350.800 459.700 ;
        RECT 370.800 459.600 371.600 459.700 ;
        RECT 390.000 459.600 390.800 459.700 ;
        RECT 393.200 460.300 394.000 460.400 ;
        RECT 434.800 460.300 435.600 460.400 ;
        RECT 393.200 459.700 435.600 460.300 ;
        RECT 393.200 459.600 394.000 459.700 ;
        RECT 434.800 459.600 435.600 459.700 ;
        RECT 514.800 460.300 515.600 460.400 ;
        RECT 542.000 460.300 542.800 460.400 ;
        RECT 514.800 459.700 542.800 460.300 ;
        RECT 514.800 459.600 515.600 459.700 ;
        RECT 542.000 459.600 542.800 459.700 ;
        RECT 551.600 460.300 552.400 460.400 ;
        RECT 569.200 460.300 570.000 460.400 ;
        RECT 551.600 459.700 570.000 460.300 ;
        RECT 551.600 459.600 552.400 459.700 ;
        RECT 569.200 459.600 570.000 459.700 ;
        RECT 647.600 460.300 648.400 460.400 ;
        RECT 655.600 460.300 656.400 460.400 ;
        RECT 647.600 459.700 656.400 460.300 ;
        RECT 647.600 459.600 648.400 459.700 ;
        RECT 655.600 459.600 656.400 459.700 ;
        RECT 172.400 458.300 173.200 458.400 ;
        RECT 175.600 458.300 176.400 458.400 ;
        RECT 172.400 457.700 176.400 458.300 ;
        RECT 172.400 457.600 173.200 457.700 ;
        RECT 175.600 457.600 176.400 457.700 ;
        RECT 202.800 458.300 203.600 458.400 ;
        RECT 244.400 458.300 245.200 458.400 ;
        RECT 202.800 457.700 245.200 458.300 ;
        RECT 202.800 457.600 203.600 457.700 ;
        RECT 244.400 457.600 245.200 457.700 ;
        RECT 330.800 458.300 331.600 458.400 ;
        RECT 348.400 458.300 349.200 458.400 ;
        RECT 330.800 457.700 349.200 458.300 ;
        RECT 330.800 457.600 331.600 457.700 ;
        RECT 348.400 457.600 349.200 457.700 ;
        RECT 606.000 458.300 606.800 458.400 ;
        RECT 644.400 458.300 645.200 458.400 ;
        RECT 606.000 457.700 645.200 458.300 ;
        RECT 606.000 457.600 606.800 457.700 ;
        RECT 644.400 457.600 645.200 457.700 ;
        RECT 652.400 458.300 653.200 458.400 ;
        RECT 657.200 458.300 658.000 458.400 ;
        RECT 652.400 457.700 658.000 458.300 ;
        RECT 652.400 457.600 653.200 457.700 ;
        RECT 657.200 457.600 658.000 457.700 ;
        RECT 42.800 455.600 43.600 456.400 ;
        RECT 78.000 456.300 78.800 456.400 ;
        RECT 87.600 456.300 88.400 456.400 ;
        RECT 98.800 456.300 99.600 456.400 ;
        RECT 118.000 456.300 118.800 456.400 ;
        RECT 129.200 456.300 130.000 456.400 ;
        RECT 78.000 455.700 130.000 456.300 ;
        RECT 78.000 455.600 78.800 455.700 ;
        RECT 87.600 455.600 88.400 455.700 ;
        RECT 98.800 455.600 99.600 455.700 ;
        RECT 118.000 455.600 118.800 455.700 ;
        RECT 129.200 455.600 130.000 455.700 ;
        RECT 282.800 456.300 283.600 456.400 ;
        RECT 292.400 456.300 293.200 456.400 ;
        RECT 282.800 455.700 293.200 456.300 ;
        RECT 282.800 455.600 283.600 455.700 ;
        RECT 292.400 455.600 293.200 455.700 ;
        RECT 305.200 456.300 306.000 456.400 ;
        RECT 308.400 456.300 309.200 456.400 ;
        RECT 305.200 455.700 309.200 456.300 ;
        RECT 305.200 455.600 306.000 455.700 ;
        RECT 308.400 455.600 309.200 455.700 ;
        RECT 335.600 456.300 336.400 456.400 ;
        RECT 345.200 456.300 346.000 456.400 ;
        RECT 351.600 456.300 352.400 456.400 ;
        RECT 335.600 455.700 352.400 456.300 ;
        RECT 335.600 455.600 336.400 455.700 ;
        RECT 345.200 455.600 346.000 455.700 ;
        RECT 351.600 455.600 352.400 455.700 ;
        RECT 356.400 456.300 357.200 456.400 ;
        RECT 375.600 456.300 376.400 456.400 ;
        RECT 356.400 455.700 376.400 456.300 ;
        RECT 356.400 455.600 357.200 455.700 ;
        RECT 375.600 455.600 376.400 455.700 ;
        RECT 402.800 456.300 403.600 456.400 ;
        RECT 410.800 456.300 411.600 456.400 ;
        RECT 402.800 455.700 411.600 456.300 ;
        RECT 402.800 455.600 403.600 455.700 ;
        RECT 410.800 455.600 411.600 455.700 ;
        RECT 450.800 456.300 451.600 456.400 ;
        RECT 478.000 456.300 478.800 456.400 ;
        RECT 450.800 455.700 478.800 456.300 ;
        RECT 450.800 455.600 451.600 455.700 ;
        RECT 478.000 455.600 478.800 455.700 ;
        RECT 481.200 456.300 482.000 456.400 ;
        RECT 497.200 456.300 498.000 456.400 ;
        RECT 481.200 455.700 498.000 456.300 ;
        RECT 481.200 455.600 482.000 455.700 ;
        RECT 497.200 455.600 498.000 455.700 ;
        RECT 510.000 456.300 510.800 456.400 ;
        RECT 530.800 456.300 531.600 456.400 ;
        RECT 510.000 455.700 531.600 456.300 ;
        RECT 510.000 455.600 510.800 455.700 ;
        RECT 530.800 455.600 531.600 455.700 ;
        RECT 612.400 456.300 613.200 456.400 ;
        RECT 615.600 456.300 616.400 456.400 ;
        RECT 625.200 456.300 626.000 456.400 ;
        RECT 612.400 455.700 626.000 456.300 ;
        RECT 612.400 455.600 613.200 455.700 ;
        RECT 615.600 455.600 616.400 455.700 ;
        RECT 625.200 455.600 626.000 455.700 ;
        RECT 34.800 454.300 35.600 454.400 ;
        RECT 46.000 454.300 46.800 454.400 ;
        RECT 34.800 453.700 46.800 454.300 ;
        RECT 34.800 453.600 35.600 453.700 ;
        RECT 46.000 453.600 46.800 453.700 ;
        RECT 86.000 454.300 86.800 454.400 ;
        RECT 110.000 454.300 110.800 454.400 ;
        RECT 124.400 454.300 125.200 454.400 ;
        RECT 86.000 453.700 125.200 454.300 ;
        RECT 86.000 453.600 86.800 453.700 ;
        RECT 110.000 453.600 110.800 453.700 ;
        RECT 124.400 453.600 125.200 453.700 ;
        RECT 162.800 454.300 163.600 454.400 ;
        RECT 164.400 454.300 165.200 454.400 ;
        RECT 162.800 453.700 165.200 454.300 ;
        RECT 162.800 453.600 163.600 453.700 ;
        RECT 164.400 453.600 165.200 453.700 ;
        RECT 170.800 453.600 171.600 454.400 ;
        RECT 185.200 454.300 186.000 454.400 ;
        RECT 199.600 454.300 200.400 454.400 ;
        RECT 185.200 453.700 200.400 454.300 ;
        RECT 185.200 453.600 186.000 453.700 ;
        RECT 199.600 453.600 200.400 453.700 ;
        RECT 279.600 454.300 280.400 454.400 ;
        RECT 300.400 454.300 301.200 454.400 ;
        RECT 279.600 453.700 301.200 454.300 ;
        RECT 279.600 453.600 280.400 453.700 ;
        RECT 300.400 453.600 301.200 453.700 ;
        RECT 311.600 454.300 312.400 454.400 ;
        RECT 319.600 454.300 320.400 454.400 ;
        RECT 311.600 453.700 320.400 454.300 ;
        RECT 311.600 453.600 312.400 453.700 ;
        RECT 319.600 453.600 320.400 453.700 ;
        RECT 330.800 454.300 331.600 454.400 ;
        RECT 338.800 454.300 339.600 454.400 ;
        RECT 346.800 454.300 347.600 454.400 ;
        RECT 330.800 453.700 347.600 454.300 ;
        RECT 330.800 453.600 331.600 453.700 ;
        RECT 338.800 453.600 339.600 453.700 ;
        RECT 346.800 453.600 347.600 453.700 ;
        RECT 354.800 454.300 355.600 454.400 ;
        RECT 366.000 454.300 366.800 454.400 ;
        RECT 354.800 453.700 366.800 454.300 ;
        RECT 354.800 453.600 355.600 453.700 ;
        RECT 366.000 453.600 366.800 453.700 ;
        RECT 378.800 454.300 379.600 454.400 ;
        RECT 382.000 454.300 382.800 454.400 ;
        RECT 378.800 453.700 382.800 454.300 ;
        RECT 378.800 453.600 379.600 453.700 ;
        RECT 382.000 453.600 382.800 453.700 ;
        RECT 398.000 454.300 398.800 454.400 ;
        RECT 414.000 454.300 414.800 454.400 ;
        RECT 398.000 453.700 414.800 454.300 ;
        RECT 398.000 453.600 398.800 453.700 ;
        RECT 414.000 453.600 414.800 453.700 ;
        RECT 442.800 454.300 443.600 454.400 ;
        RECT 473.200 454.300 474.000 454.400 ;
        RECT 442.800 453.700 474.000 454.300 ;
        RECT 442.800 453.600 443.600 453.700 ;
        RECT 473.200 453.600 474.000 453.700 ;
        RECT 526.000 454.300 526.800 454.400 ;
        RECT 546.800 454.300 547.600 454.400 ;
        RECT 526.000 453.700 547.600 454.300 ;
        RECT 526.000 453.600 526.800 453.700 ;
        RECT 546.800 453.600 547.600 453.700 ;
        RECT 591.600 454.300 592.400 454.400 ;
        RECT 594.800 454.300 595.600 454.400 ;
        RECT 606.000 454.300 606.800 454.400 ;
        RECT 591.600 453.700 606.800 454.300 ;
        RECT 591.600 453.600 592.400 453.700 ;
        RECT 594.800 453.600 595.600 453.700 ;
        RECT 606.000 453.600 606.800 453.700 ;
        RECT 609.200 454.300 610.000 454.400 ;
        RECT 633.200 454.300 634.000 454.400 ;
        RECT 641.200 454.300 642.000 454.400 ;
        RECT 609.200 453.700 642.000 454.300 ;
        RECT 609.200 453.600 610.000 453.700 ;
        RECT 633.200 453.600 634.000 453.700 ;
        RECT 641.200 453.600 642.000 453.700 ;
        RECT 30.000 452.300 30.800 452.400 ;
        RECT 44.400 452.300 45.200 452.400 ;
        RECT 30.000 451.700 45.200 452.300 ;
        RECT 30.000 451.600 30.800 451.700 ;
        RECT 44.400 451.600 45.200 451.700 ;
        RECT 66.800 452.300 67.600 452.400 ;
        RECT 73.200 452.300 74.000 452.400 ;
        RECT 66.800 451.700 74.000 452.300 ;
        RECT 66.800 451.600 67.600 451.700 ;
        RECT 73.200 451.600 74.000 451.700 ;
        RECT 106.800 452.300 107.600 452.400 ;
        RECT 127.600 452.300 128.400 452.400 ;
        RECT 106.800 451.700 128.400 452.300 ;
        RECT 106.800 451.600 107.600 451.700 ;
        RECT 127.600 451.600 128.400 451.700 ;
        RECT 145.200 452.300 146.000 452.400 ;
        RECT 150.000 452.300 150.800 452.400 ;
        RECT 145.200 451.700 150.800 452.300 ;
        RECT 145.200 451.600 146.000 451.700 ;
        RECT 150.000 451.600 150.800 451.700 ;
        RECT 154.800 452.300 155.600 452.400 ;
        RECT 162.800 452.300 163.600 452.400 ;
        RECT 154.800 451.700 163.600 452.300 ;
        RECT 154.800 451.600 155.600 451.700 ;
        RECT 162.800 451.600 163.600 451.700 ;
        RECT 164.400 452.300 165.200 452.400 ;
        RECT 170.800 452.300 171.600 452.400 ;
        RECT 164.400 451.700 171.600 452.300 ;
        RECT 164.400 451.600 165.200 451.700 ;
        RECT 170.800 451.600 171.600 451.700 ;
        RECT 174.000 452.300 174.800 452.400 ;
        RECT 180.400 452.300 181.200 452.400 ;
        RECT 174.000 451.700 181.200 452.300 ;
        RECT 174.000 451.600 174.800 451.700 ;
        RECT 180.400 451.600 181.200 451.700 ;
        RECT 196.400 452.300 197.200 452.400 ;
        RECT 209.200 452.300 210.000 452.400 ;
        RECT 196.400 451.700 210.000 452.300 ;
        RECT 196.400 451.600 197.200 451.700 ;
        RECT 209.200 451.600 210.000 451.700 ;
        RECT 214.000 452.300 214.800 452.400 ;
        RECT 218.800 452.300 219.600 452.400 ;
        RECT 214.000 451.700 219.600 452.300 ;
        RECT 214.000 451.600 214.800 451.700 ;
        RECT 218.800 451.600 219.600 451.700 ;
        RECT 257.200 452.300 258.000 452.400 ;
        RECT 260.400 452.300 261.200 452.400 ;
        RECT 257.200 451.700 261.200 452.300 ;
        RECT 257.200 451.600 258.000 451.700 ;
        RECT 260.400 451.600 261.200 451.700 ;
        RECT 271.600 452.300 272.400 452.400 ;
        RECT 279.600 452.300 280.400 452.400 ;
        RECT 271.600 451.700 280.400 452.300 ;
        RECT 271.600 451.600 272.400 451.700 ;
        RECT 279.600 451.600 280.400 451.700 ;
        RECT 322.800 452.300 323.600 452.400 ;
        RECT 332.400 452.300 333.200 452.400 ;
        RECT 322.800 451.700 333.200 452.300 ;
        RECT 322.800 451.600 323.600 451.700 ;
        RECT 332.400 451.600 333.200 451.700 ;
        RECT 348.400 452.300 349.200 452.400 ;
        RECT 356.400 452.300 357.200 452.400 ;
        RECT 348.400 451.700 357.200 452.300 ;
        RECT 348.400 451.600 349.200 451.700 ;
        RECT 356.400 451.600 357.200 451.700 ;
        RECT 358.000 452.300 358.800 452.400 ;
        RECT 369.200 452.300 370.000 452.400 ;
        RECT 372.400 452.300 373.200 452.400 ;
        RECT 358.000 451.700 373.200 452.300 ;
        RECT 358.000 451.600 358.800 451.700 ;
        RECT 369.200 451.600 370.000 451.700 ;
        RECT 372.400 451.600 373.200 451.700 ;
        RECT 374.000 452.300 374.800 452.400 ;
        RECT 388.400 452.300 389.200 452.400 ;
        RECT 374.000 451.700 389.200 452.300 ;
        RECT 374.000 451.600 374.800 451.700 ;
        RECT 388.400 451.600 389.200 451.700 ;
        RECT 562.800 452.300 563.600 452.400 ;
        RECT 570.800 452.300 571.600 452.400 ;
        RECT 562.800 451.700 571.600 452.300 ;
        RECT 562.800 451.600 563.600 451.700 ;
        RECT 570.800 451.600 571.600 451.700 ;
        RECT 582.000 452.300 582.800 452.400 ;
        RECT 622.000 452.300 622.800 452.400 ;
        RECT 582.000 451.700 622.800 452.300 ;
        RECT 582.000 451.600 582.800 451.700 ;
        RECT 622.000 451.600 622.800 451.700 ;
        RECT 14.000 450.300 14.800 450.400 ;
        RECT 22.000 450.300 22.800 450.400 ;
        RECT 14.000 449.700 22.800 450.300 ;
        RECT 14.000 449.600 14.800 449.700 ;
        RECT 22.000 449.600 22.800 449.700 ;
        RECT 31.600 450.300 32.400 450.400 ;
        RECT 41.200 450.300 42.000 450.400 ;
        RECT 42.800 450.300 43.600 450.400 ;
        RECT 31.600 449.700 43.600 450.300 ;
        RECT 31.600 449.600 32.400 449.700 ;
        RECT 41.200 449.600 42.000 449.700 ;
        RECT 42.800 449.600 43.600 449.700 ;
        RECT 49.200 450.300 50.000 450.400 ;
        RECT 63.600 450.300 64.400 450.400 ;
        RECT 65.200 450.300 66.000 450.400 ;
        RECT 49.200 449.700 66.000 450.300 ;
        RECT 49.200 449.600 50.000 449.700 ;
        RECT 63.600 449.600 64.400 449.700 ;
        RECT 65.200 449.600 66.000 449.700 ;
        RECT 70.000 450.300 70.800 450.400 ;
        RECT 84.400 450.300 85.200 450.400 ;
        RECT 70.000 449.700 85.200 450.300 ;
        RECT 70.000 449.600 70.800 449.700 ;
        RECT 84.400 449.600 85.200 449.700 ;
        RECT 142.000 450.300 142.800 450.400 ;
        RECT 161.200 450.300 162.000 450.400 ;
        RECT 142.000 449.700 162.000 450.300 ;
        RECT 142.000 449.600 142.800 449.700 ;
        RECT 161.200 449.600 162.000 449.700 ;
        RECT 174.000 450.300 174.800 450.400 ;
        RECT 185.200 450.300 186.000 450.400 ;
        RECT 174.000 449.700 186.000 450.300 ;
        RECT 174.000 449.600 174.800 449.700 ;
        RECT 185.200 449.600 186.000 449.700 ;
        RECT 367.600 450.300 368.400 450.400 ;
        RECT 377.200 450.300 378.000 450.400 ;
        RECT 380.400 450.300 381.200 450.400 ;
        RECT 367.600 449.700 381.200 450.300 ;
        RECT 367.600 449.600 368.400 449.700 ;
        RECT 377.200 449.600 378.000 449.700 ;
        RECT 380.400 449.600 381.200 449.700 ;
        RECT 476.400 450.300 477.200 450.400 ;
        RECT 478.000 450.300 478.800 450.400 ;
        RECT 476.400 449.700 478.800 450.300 ;
        RECT 476.400 449.600 477.200 449.700 ;
        RECT 478.000 449.600 478.800 449.700 ;
        RECT 542.000 450.300 542.800 450.400 ;
        RECT 550.000 450.300 550.800 450.400 ;
        RECT 542.000 449.700 550.800 450.300 ;
        RECT 542.000 449.600 542.800 449.700 ;
        RECT 550.000 449.600 550.800 449.700 ;
        RECT 554.800 450.300 555.600 450.400 ;
        RECT 596.400 450.300 597.200 450.400 ;
        RECT 554.800 449.700 597.200 450.300 ;
        RECT 554.800 449.600 555.600 449.700 ;
        RECT 596.400 449.600 597.200 449.700 ;
        RECT 599.600 450.300 600.400 450.400 ;
        RECT 617.200 450.300 618.000 450.400 ;
        RECT 599.600 449.700 618.000 450.300 ;
        RECT 599.600 449.600 600.400 449.700 ;
        RECT 617.200 449.600 618.000 449.700 ;
        RECT 620.400 450.300 621.200 450.400 ;
        RECT 628.400 450.300 629.200 450.400 ;
        RECT 620.400 449.700 629.200 450.300 ;
        RECT 620.400 449.600 621.200 449.700 ;
        RECT 628.400 449.600 629.200 449.700 ;
        RECT 663.600 450.300 664.400 450.400 ;
        RECT 670.000 450.300 670.800 450.400 ;
        RECT 663.600 449.700 670.800 450.300 ;
        RECT 663.600 449.600 664.400 449.700 ;
        RECT 670.000 449.600 670.800 449.700 ;
        RECT 2.800 448.300 3.600 448.400 ;
        RECT 39.600 448.300 40.400 448.400 ;
        RECT 2.800 447.700 40.400 448.300 ;
        RECT 2.800 447.600 3.600 447.700 ;
        RECT 39.600 447.600 40.400 447.700 ;
        RECT 156.400 448.300 157.200 448.400 ;
        RECT 182.000 448.300 182.800 448.400 ;
        RECT 193.200 448.300 194.000 448.400 ;
        RECT 156.400 447.700 194.000 448.300 ;
        RECT 156.400 447.600 157.200 447.700 ;
        RECT 182.000 447.600 182.800 447.700 ;
        RECT 193.200 447.600 194.000 447.700 ;
        RECT 222.000 448.300 222.800 448.400 ;
        RECT 226.800 448.300 227.600 448.400 ;
        RECT 222.000 447.700 227.600 448.300 ;
        RECT 222.000 447.600 222.800 447.700 ;
        RECT 226.800 447.600 227.600 447.700 ;
        RECT 314.800 448.300 315.600 448.400 ;
        RECT 321.200 448.300 322.000 448.400 ;
        RECT 327.600 448.300 328.400 448.400 ;
        RECT 314.800 447.700 328.400 448.300 ;
        RECT 314.800 447.600 315.600 447.700 ;
        RECT 321.200 447.600 322.000 447.700 ;
        RECT 327.600 447.600 328.400 447.700 ;
        RECT 382.000 448.300 382.800 448.400 ;
        RECT 388.400 448.300 389.200 448.400 ;
        RECT 382.000 447.700 389.200 448.300 ;
        RECT 382.000 447.600 382.800 447.700 ;
        RECT 388.400 447.600 389.200 447.700 ;
        RECT 495.600 448.300 496.400 448.400 ;
        RECT 593.200 448.300 594.000 448.400 ;
        RECT 602.800 448.300 603.600 448.400 ;
        RECT 495.600 447.700 603.600 448.300 ;
        RECT 495.600 447.600 496.400 447.700 ;
        RECT 593.200 447.600 594.000 447.700 ;
        RECT 602.800 447.600 603.600 447.700 ;
        RECT 626.800 448.300 627.600 448.400 ;
        RECT 630.000 448.300 630.800 448.400 ;
        RECT 626.800 447.700 630.800 448.300 ;
        RECT 626.800 447.600 627.600 447.700 ;
        RECT 630.000 447.600 630.800 447.700 ;
        RECT 631.600 447.600 632.400 448.400 ;
        RECT 636.400 448.300 637.200 448.400 ;
        RECT 652.400 448.300 653.200 448.400 ;
        RECT 668.400 448.300 669.200 448.400 ;
        RECT 636.400 447.700 669.200 448.300 ;
        RECT 636.400 447.600 637.200 447.700 ;
        RECT 652.400 447.600 653.200 447.700 ;
        RECT 668.400 447.600 669.200 447.700 ;
        RECT 20.400 446.300 21.200 446.400 ;
        RECT 55.600 446.300 56.400 446.400 ;
        RECT 20.400 445.700 56.400 446.300 ;
        RECT 20.400 445.600 21.200 445.700 ;
        RECT 55.600 445.600 56.400 445.700 ;
        RECT 71.600 446.300 72.400 446.400 ;
        RECT 86.000 446.300 86.800 446.400 ;
        RECT 71.600 445.700 86.800 446.300 ;
        RECT 71.600 445.600 72.400 445.700 ;
        RECT 86.000 445.600 86.800 445.700 ;
        RECT 111.600 446.300 112.400 446.400 ;
        RECT 127.600 446.300 128.400 446.400 ;
        RECT 111.600 445.700 128.400 446.300 ;
        RECT 111.600 445.600 112.400 445.700 ;
        RECT 127.600 445.600 128.400 445.700 ;
        RECT 306.800 446.300 307.600 446.400 ;
        RECT 326.000 446.300 326.800 446.400 ;
        RECT 362.800 446.300 363.600 446.400 ;
        RECT 306.800 445.700 363.600 446.300 ;
        RECT 306.800 445.600 307.600 445.700 ;
        RECT 326.000 445.600 326.800 445.700 ;
        RECT 362.800 445.600 363.600 445.700 ;
        RECT 399.600 446.300 400.400 446.400 ;
        RECT 436.400 446.300 437.200 446.400 ;
        RECT 550.000 446.300 550.800 446.400 ;
        RECT 399.600 445.700 550.800 446.300 ;
        RECT 399.600 445.600 400.400 445.700 ;
        RECT 436.400 445.600 437.200 445.700 ;
        RECT 550.000 445.600 550.800 445.700 ;
        RECT 612.400 446.300 613.200 446.400 ;
        RECT 628.400 446.300 629.200 446.400 ;
        RECT 612.400 445.700 629.200 446.300 ;
        RECT 612.400 445.600 613.200 445.700 ;
        RECT 628.400 445.600 629.200 445.700 ;
        RECT 1.200 444.300 2.000 444.400 ;
        RECT 26.800 444.300 27.600 444.400 ;
        RECT 39.600 444.300 40.400 444.400 ;
        RECT 1.200 443.700 40.400 444.300 ;
        RECT 1.200 443.600 2.000 443.700 ;
        RECT 26.800 443.600 27.600 443.700 ;
        RECT 39.600 443.600 40.400 443.700 ;
        RECT 73.200 444.300 74.000 444.400 ;
        RECT 97.200 444.300 98.000 444.400 ;
        RECT 73.200 443.700 98.000 444.300 ;
        RECT 73.200 443.600 74.000 443.700 ;
        RECT 97.200 443.600 98.000 443.700 ;
        RECT 103.600 444.300 104.400 444.400 ;
        RECT 116.400 444.300 117.200 444.400 ;
        RECT 103.600 443.700 117.200 444.300 ;
        RECT 103.600 443.600 104.400 443.700 ;
        RECT 116.400 443.600 117.200 443.700 ;
        RECT 276.400 444.300 277.200 444.400 ;
        RECT 281.200 444.300 282.000 444.400 ;
        RECT 276.400 443.700 282.000 444.300 ;
        RECT 276.400 443.600 277.200 443.700 ;
        RECT 281.200 443.600 282.000 443.700 ;
        RECT 329.200 444.300 330.000 444.400 ;
        RECT 335.600 444.300 336.400 444.400 ;
        RECT 342.000 444.300 342.800 444.400 ;
        RECT 372.400 444.300 373.200 444.400 ;
        RECT 329.200 443.700 373.200 444.300 ;
        RECT 329.200 443.600 330.000 443.700 ;
        RECT 335.600 443.600 336.400 443.700 ;
        RECT 342.000 443.600 342.800 443.700 ;
        RECT 372.400 443.600 373.200 443.700 ;
        RECT 390.000 444.300 390.800 444.400 ;
        RECT 394.800 444.300 395.600 444.400 ;
        RECT 390.000 443.700 395.600 444.300 ;
        RECT 390.000 443.600 390.800 443.700 ;
        RECT 394.800 443.600 395.600 443.700 ;
        RECT 486.000 444.300 486.800 444.400 ;
        RECT 498.800 444.300 499.600 444.400 ;
        RECT 486.000 443.700 499.600 444.300 ;
        RECT 486.000 443.600 486.800 443.700 ;
        RECT 498.800 443.600 499.600 443.700 ;
        RECT 514.800 444.300 515.600 444.400 ;
        RECT 546.800 444.300 547.600 444.400 ;
        RECT 514.800 443.700 547.600 444.300 ;
        RECT 514.800 443.600 515.600 443.700 ;
        RECT 546.800 443.600 547.600 443.700 ;
        RECT 23.600 442.300 24.400 442.400 ;
        RECT 36.400 442.300 37.200 442.400 ;
        RECT 23.600 441.700 37.200 442.300 ;
        RECT 23.600 441.600 24.400 441.700 ;
        RECT 36.400 441.600 37.200 441.700 ;
        RECT 318.000 442.300 318.800 442.400 ;
        RECT 340.400 442.300 341.200 442.400 ;
        RECT 318.000 441.700 341.200 442.300 ;
        RECT 318.000 441.600 318.800 441.700 ;
        RECT 340.400 441.600 341.200 441.700 ;
        RECT 350.000 442.300 350.800 442.400 ;
        RECT 354.800 442.300 355.600 442.400 ;
        RECT 369.200 442.300 370.000 442.400 ;
        RECT 350.000 441.700 370.000 442.300 ;
        RECT 350.000 441.600 350.800 441.700 ;
        RECT 354.800 441.600 355.600 441.700 ;
        RECT 369.200 441.600 370.000 441.700 ;
        RECT 401.200 442.300 402.000 442.400 ;
        RECT 407.600 442.300 408.400 442.400 ;
        RECT 401.200 441.700 408.400 442.300 ;
        RECT 401.200 441.600 402.000 441.700 ;
        RECT 407.600 441.600 408.400 441.700 ;
        RECT 438.000 442.300 438.800 442.400 ;
        RECT 446.000 442.300 446.800 442.400 ;
        RECT 438.000 441.700 446.800 442.300 ;
        RECT 438.000 441.600 438.800 441.700 ;
        RECT 446.000 441.600 446.800 441.700 ;
        RECT 649.200 442.300 650.000 442.400 ;
        RECT 650.800 442.300 651.600 442.400 ;
        RECT 649.200 441.700 651.600 442.300 ;
        RECT 649.200 441.600 650.000 441.700 ;
        RECT 650.800 441.600 651.600 441.700 ;
        RECT 137.200 440.300 138.000 440.400 ;
        RECT 148.400 440.300 149.200 440.400 ;
        RECT 169.200 440.300 170.000 440.400 ;
        RECT 198.000 440.300 198.800 440.400 ;
        RECT 137.200 439.700 198.800 440.300 ;
        RECT 137.200 439.600 138.000 439.700 ;
        RECT 148.400 439.600 149.200 439.700 ;
        RECT 169.200 439.600 170.000 439.700 ;
        RECT 198.000 439.600 198.800 439.700 ;
        RECT 362.800 440.300 363.600 440.400 ;
        RECT 383.600 440.300 384.400 440.400 ;
        RECT 362.800 439.700 384.400 440.300 ;
        RECT 362.800 439.600 363.600 439.700 ;
        RECT 383.600 439.600 384.400 439.700 ;
        RECT 426.800 440.300 427.600 440.400 ;
        RECT 438.000 440.300 438.800 440.400 ;
        RECT 426.800 439.700 438.800 440.300 ;
        RECT 426.800 439.600 427.600 439.700 ;
        RECT 438.000 439.600 438.800 439.700 ;
        RECT 478.000 440.300 478.800 440.400 ;
        RECT 484.400 440.300 485.200 440.400 ;
        RECT 478.000 439.700 485.200 440.300 ;
        RECT 478.000 439.600 478.800 439.700 ;
        RECT 484.400 439.600 485.200 439.700 ;
        RECT 41.200 438.300 42.000 438.400 ;
        RECT 65.200 438.300 66.000 438.400 ;
        RECT 70.000 438.300 70.800 438.400 ;
        RECT 154.800 438.300 155.600 438.400 ;
        RECT 41.200 437.700 155.600 438.300 ;
        RECT 41.200 437.600 42.000 437.700 ;
        RECT 65.200 437.600 66.000 437.700 ;
        RECT 70.000 437.600 70.800 437.700 ;
        RECT 154.800 437.600 155.600 437.700 ;
        RECT 218.800 438.300 219.600 438.400 ;
        RECT 231.600 438.300 232.400 438.400 ;
        RECT 218.800 437.700 232.400 438.300 ;
        RECT 218.800 437.600 219.600 437.700 ;
        RECT 231.600 437.600 232.400 437.700 ;
        RECT 342.000 438.300 342.800 438.400 ;
        RECT 346.800 438.300 347.600 438.400 ;
        RECT 342.000 437.700 347.600 438.300 ;
        RECT 342.000 437.600 342.800 437.700 ;
        RECT 346.800 437.600 347.600 437.700 ;
        RECT 366.000 437.600 366.800 438.400 ;
        RECT 482.800 438.300 483.600 438.400 ;
        RECT 495.600 438.300 496.400 438.400 ;
        RECT 482.800 437.700 496.400 438.300 ;
        RECT 482.800 437.600 483.600 437.700 ;
        RECT 495.600 437.600 496.400 437.700 ;
        RECT 513.200 438.300 514.000 438.400 ;
        RECT 518.000 438.300 518.800 438.400 ;
        RECT 513.200 437.700 518.800 438.300 ;
        RECT 513.200 437.600 514.000 437.700 ;
        RECT 518.000 437.600 518.800 437.700 ;
        RECT 521.200 438.300 522.000 438.400 ;
        RECT 543.600 438.300 544.400 438.400 ;
        RECT 551.600 438.300 552.400 438.400 ;
        RECT 521.200 437.700 552.400 438.300 ;
        RECT 521.200 437.600 522.000 437.700 ;
        RECT 543.600 437.600 544.400 437.700 ;
        RECT 551.600 437.600 552.400 437.700 ;
        RECT 42.800 435.600 43.600 436.400 ;
        RECT 55.600 436.300 56.400 436.400 ;
        RECT 138.800 436.300 139.600 436.400 ;
        RECT 55.600 435.700 139.600 436.300 ;
        RECT 55.600 435.600 56.400 435.700 ;
        RECT 138.800 435.600 139.600 435.700 ;
        RECT 161.200 436.300 162.000 436.400 ;
        RECT 178.800 436.300 179.600 436.400 ;
        RECT 161.200 435.700 179.600 436.300 ;
        RECT 161.200 435.600 162.000 435.700 ;
        RECT 178.800 435.600 179.600 435.700 ;
        RECT 322.800 436.300 323.600 436.400 ;
        RECT 330.800 436.300 331.600 436.400 ;
        RECT 322.800 435.700 331.600 436.300 ;
        RECT 322.800 435.600 323.600 435.700 ;
        RECT 330.800 435.600 331.600 435.700 ;
        RECT 345.200 436.300 346.000 436.400 ;
        RECT 348.400 436.300 349.200 436.400 ;
        RECT 345.200 435.700 349.200 436.300 ;
        RECT 345.200 435.600 346.000 435.700 ;
        RECT 348.400 435.600 349.200 435.700 ;
        RECT 366.000 436.300 366.800 436.400 ;
        RECT 369.200 436.300 370.000 436.400 ;
        RECT 366.000 435.700 370.000 436.300 ;
        RECT 366.000 435.600 366.800 435.700 ;
        RECT 369.200 435.600 370.000 435.700 ;
        RECT 382.000 436.300 382.800 436.400 ;
        RECT 406.000 436.300 406.800 436.400 ;
        RECT 382.000 435.700 406.800 436.300 ;
        RECT 382.000 435.600 382.800 435.700 ;
        RECT 406.000 435.600 406.800 435.700 ;
        RECT 44.400 434.300 45.200 434.400 ;
        RECT 76.400 434.300 77.200 434.400 ;
        RECT 44.400 433.700 77.200 434.300 ;
        RECT 44.400 433.600 45.200 433.700 ;
        RECT 76.400 433.600 77.200 433.700 ;
        RECT 151.600 434.300 152.400 434.400 ;
        RECT 169.200 434.300 170.000 434.400 ;
        RECT 151.600 433.700 170.000 434.300 ;
        RECT 151.600 433.600 152.400 433.700 ;
        RECT 169.200 433.600 170.000 433.700 ;
        RECT 225.200 434.300 226.000 434.400 ;
        RECT 247.600 434.300 248.400 434.400 ;
        RECT 225.200 433.700 248.400 434.300 ;
        RECT 225.200 433.600 226.000 433.700 ;
        RECT 247.600 433.600 248.400 433.700 ;
        RECT 319.600 434.300 320.400 434.400 ;
        RECT 327.600 434.300 328.400 434.400 ;
        RECT 364.400 434.300 365.200 434.400 ;
        RECT 370.800 434.300 371.600 434.400 ;
        RECT 372.400 434.300 373.200 434.400 ;
        RECT 319.600 433.700 373.200 434.300 ;
        RECT 319.600 433.600 320.400 433.700 ;
        RECT 327.600 433.600 328.400 433.700 ;
        RECT 364.400 433.600 365.200 433.700 ;
        RECT 370.800 433.600 371.600 433.700 ;
        RECT 372.400 433.600 373.200 433.700 ;
        RECT 506.800 434.300 507.600 434.400 ;
        RECT 638.000 434.300 638.800 434.400 ;
        RECT 647.600 434.300 648.400 434.400 ;
        RECT 655.600 434.300 656.400 434.400 ;
        RECT 506.800 433.700 656.400 434.300 ;
        RECT 506.800 433.600 507.600 433.700 ;
        RECT 638.000 433.600 638.800 433.700 ;
        RECT 647.600 433.600 648.400 433.700 ;
        RECT 655.600 433.600 656.400 433.700 ;
        RECT 1.200 432.300 2.000 432.400 ;
        RECT 26.800 432.300 27.600 432.400 ;
        RECT 33.200 432.300 34.000 432.400 ;
        RECT 66.800 432.300 67.600 432.400 ;
        RECT 1.200 431.700 34.000 432.300 ;
        RECT 1.200 431.600 2.000 431.700 ;
        RECT 26.800 431.600 27.600 431.700 ;
        RECT 33.200 431.600 34.000 431.700 ;
        RECT 57.300 431.700 67.600 432.300 ;
        RECT 57.300 430.400 57.900 431.700 ;
        RECT 66.800 431.600 67.600 431.700 ;
        RECT 84.400 432.300 85.200 432.400 ;
        RECT 98.800 432.300 99.600 432.400 ;
        RECT 84.400 431.700 99.600 432.300 ;
        RECT 84.400 431.600 85.200 431.700 ;
        RECT 98.800 431.600 99.600 431.700 ;
        RECT 146.800 432.300 147.600 432.400 ;
        RECT 159.600 432.300 160.400 432.400 ;
        RECT 146.800 431.700 160.400 432.300 ;
        RECT 146.800 431.600 147.600 431.700 ;
        RECT 159.600 431.600 160.400 431.700 ;
        RECT 169.200 432.300 170.000 432.400 ;
        RECT 177.200 432.300 178.000 432.400 ;
        RECT 169.200 431.700 178.000 432.300 ;
        RECT 169.200 431.600 170.000 431.700 ;
        RECT 177.200 431.600 178.000 431.700 ;
        RECT 217.200 432.300 218.000 432.400 ;
        RECT 228.400 432.300 229.200 432.400 ;
        RECT 234.800 432.300 235.600 432.400 ;
        RECT 217.200 431.700 235.600 432.300 ;
        RECT 217.200 431.600 218.000 431.700 ;
        RECT 228.400 431.600 229.200 431.700 ;
        RECT 234.800 431.600 235.600 431.700 ;
        RECT 298.800 432.300 299.600 432.400 ;
        RECT 303.600 432.300 304.400 432.400 ;
        RECT 298.800 431.700 304.400 432.300 ;
        RECT 298.800 431.600 299.600 431.700 ;
        RECT 303.600 431.600 304.400 431.700 ;
        RECT 332.400 432.300 333.200 432.400 ;
        RECT 345.200 432.300 346.000 432.400 ;
        RECT 356.400 432.300 357.200 432.400 ;
        RECT 367.600 432.300 368.400 432.400 ;
        RECT 374.000 432.300 374.800 432.400 ;
        RECT 332.400 431.700 357.200 432.300 ;
        RECT 332.400 431.600 333.200 431.700 ;
        RECT 345.200 431.600 346.000 431.700 ;
        RECT 356.400 431.600 357.200 431.700 ;
        RECT 366.100 431.700 374.800 432.300 ;
        RECT 14.000 430.300 14.800 430.400 ;
        RECT 23.600 430.300 24.400 430.400 ;
        RECT 14.000 429.700 24.400 430.300 ;
        RECT 14.000 429.600 14.800 429.700 ;
        RECT 23.600 429.600 24.400 429.700 ;
        RECT 34.800 430.300 35.600 430.400 ;
        RECT 36.400 430.300 37.200 430.400 ;
        RECT 42.800 430.300 43.600 430.400 ;
        RECT 57.200 430.300 58.000 430.400 ;
        RECT 34.800 429.700 58.000 430.300 ;
        RECT 34.800 429.600 35.600 429.700 ;
        RECT 36.400 429.600 37.200 429.700 ;
        RECT 42.800 429.600 43.600 429.700 ;
        RECT 57.200 429.600 58.000 429.700 ;
        RECT 65.200 430.300 66.000 430.400 ;
        RECT 84.400 430.300 85.200 430.400 ;
        RECT 65.200 429.700 85.200 430.300 ;
        RECT 65.200 429.600 66.000 429.700 ;
        RECT 84.400 429.600 85.200 429.700 ;
        RECT 121.200 430.300 122.000 430.400 ;
        RECT 122.800 430.300 123.600 430.400 ;
        RECT 134.000 430.300 134.800 430.400 ;
        RECT 121.200 429.700 134.800 430.300 ;
        RECT 121.200 429.600 122.000 429.700 ;
        RECT 122.800 429.600 123.600 429.700 ;
        RECT 134.000 429.600 134.800 429.700 ;
        RECT 153.200 430.300 154.000 430.400 ;
        RECT 159.600 430.300 160.400 430.400 ;
        RECT 153.200 429.700 160.400 430.300 ;
        RECT 153.200 429.600 154.000 429.700 ;
        RECT 159.600 429.600 160.400 429.700 ;
        RECT 162.800 430.300 163.600 430.400 ;
        RECT 180.400 430.300 181.200 430.400 ;
        RECT 162.800 429.700 181.200 430.300 ;
        RECT 162.800 429.600 163.600 429.700 ;
        RECT 180.400 429.600 181.200 429.700 ;
        RECT 190.000 430.300 190.800 430.400 ;
        RECT 201.200 430.300 202.000 430.400 ;
        RECT 190.000 429.700 202.000 430.300 ;
        RECT 190.000 429.600 190.800 429.700 ;
        RECT 201.200 429.600 202.000 429.700 ;
        RECT 210.800 430.300 211.600 430.400 ;
        RECT 225.200 430.300 226.000 430.400 ;
        RECT 210.800 429.700 226.000 430.300 ;
        RECT 210.800 429.600 211.600 429.700 ;
        RECT 225.200 429.600 226.000 429.700 ;
        RECT 295.600 430.300 296.400 430.400 ;
        RECT 300.400 430.300 301.200 430.400 ;
        RECT 305.200 430.300 306.000 430.400 ;
        RECT 313.200 430.300 314.000 430.400 ;
        RECT 295.600 429.700 314.000 430.300 ;
        RECT 295.600 429.600 296.400 429.700 ;
        RECT 300.400 429.600 301.200 429.700 ;
        RECT 305.200 429.600 306.000 429.700 ;
        RECT 313.200 429.600 314.000 429.700 ;
        RECT 318.000 430.300 318.800 430.400 ;
        RECT 334.000 430.300 334.800 430.400 ;
        RECT 340.400 430.300 341.200 430.400 ;
        RECT 366.100 430.300 366.700 431.700 ;
        RECT 367.600 431.600 368.400 431.700 ;
        RECT 374.000 431.600 374.800 431.700 ;
        RECT 380.400 432.300 381.200 432.400 ;
        RECT 383.600 432.300 384.400 432.400 ;
        RECT 386.800 432.300 387.600 432.400 ;
        RECT 380.400 431.700 387.600 432.300 ;
        RECT 380.400 431.600 381.200 431.700 ;
        RECT 383.600 431.600 384.400 431.700 ;
        RECT 386.800 431.600 387.600 431.700 ;
        RECT 388.400 432.300 389.200 432.400 ;
        RECT 449.200 432.300 450.000 432.400 ;
        RECT 388.400 431.700 450.000 432.300 ;
        RECT 388.400 431.600 389.200 431.700 ;
        RECT 449.200 431.600 450.000 431.700 ;
        RECT 532.400 431.600 533.200 432.400 ;
        RECT 546.800 432.300 547.600 432.400 ;
        RECT 554.800 432.300 555.600 432.400 ;
        RECT 558.000 432.300 558.800 432.400 ;
        RECT 546.800 431.700 558.800 432.300 ;
        RECT 546.800 431.600 547.600 431.700 ;
        RECT 554.800 431.600 555.600 431.700 ;
        RECT 558.000 431.600 558.800 431.700 ;
        RECT 583.600 432.300 584.400 432.400 ;
        RECT 596.400 432.300 597.200 432.400 ;
        RECT 609.200 432.300 610.000 432.400 ;
        RECT 583.600 431.700 610.000 432.300 ;
        RECT 583.600 431.600 584.400 431.700 ;
        RECT 596.400 431.600 597.200 431.700 ;
        RECT 609.200 431.600 610.000 431.700 ;
        RECT 318.000 429.700 341.200 430.300 ;
        RECT 318.000 429.600 318.800 429.700 ;
        RECT 334.000 429.600 334.800 429.700 ;
        RECT 340.400 429.600 341.200 429.700 ;
        RECT 346.900 429.700 366.700 430.300 ;
        RECT 367.600 430.300 368.400 430.400 ;
        RECT 390.000 430.300 390.800 430.400 ;
        RECT 367.600 429.700 390.800 430.300 ;
        RECT 74.800 428.300 75.600 428.400 ;
        RECT 78.000 428.300 78.800 428.400 ;
        RECT 74.800 427.700 78.800 428.300 ;
        RECT 74.800 427.600 75.600 427.700 ;
        RECT 78.000 427.600 78.800 427.700 ;
        RECT 153.200 428.300 154.000 428.400 ;
        RECT 161.200 428.300 162.000 428.400 ;
        RECT 153.200 427.700 162.000 428.300 ;
        RECT 153.200 427.600 154.000 427.700 ;
        RECT 161.200 427.600 162.000 427.700 ;
        RECT 164.400 428.300 165.200 428.400 ;
        RECT 178.800 428.300 179.600 428.400 ;
        RECT 186.800 428.300 187.600 428.400 ;
        RECT 191.600 428.300 192.400 428.400 ;
        RECT 164.400 427.700 192.400 428.300 ;
        RECT 164.400 427.600 165.200 427.700 ;
        RECT 178.800 427.600 179.600 427.700 ;
        RECT 186.800 427.600 187.600 427.700 ;
        RECT 191.600 427.600 192.400 427.700 ;
        RECT 215.600 428.300 216.400 428.400 ;
        RECT 246.000 428.300 246.800 428.400 ;
        RECT 260.400 428.300 261.200 428.400 ;
        RECT 215.600 427.700 235.500 428.300 ;
        RECT 215.600 427.600 216.400 427.700 ;
        RECT 234.900 426.400 235.500 427.700 ;
        RECT 246.000 427.700 261.200 428.300 ;
        RECT 246.000 427.600 246.800 427.700 ;
        RECT 260.400 427.600 261.200 427.700 ;
        RECT 273.200 428.300 274.000 428.400 ;
        RECT 282.800 428.300 283.600 428.400 ;
        RECT 273.200 427.700 283.600 428.300 ;
        RECT 273.200 427.600 274.000 427.700 ;
        RECT 282.800 427.600 283.600 427.700 ;
        RECT 295.600 428.300 296.400 428.400 ;
        RECT 297.200 428.300 298.000 428.400 ;
        RECT 295.600 427.700 298.000 428.300 ;
        RECT 295.600 427.600 296.400 427.700 ;
        RECT 297.200 427.600 298.000 427.700 ;
        RECT 305.200 428.300 306.000 428.400 ;
        RECT 313.200 428.300 314.000 428.400 ;
        RECT 305.200 427.700 314.000 428.300 ;
        RECT 305.200 427.600 306.000 427.700 ;
        RECT 313.200 427.600 314.000 427.700 ;
        RECT 332.400 428.300 333.200 428.400 ;
        RECT 346.900 428.300 347.500 429.700 ;
        RECT 367.600 429.600 368.400 429.700 ;
        RECT 390.000 429.600 390.800 429.700 ;
        RECT 450.800 430.300 451.600 430.400 ;
        RECT 468.400 430.300 469.200 430.400 ;
        RECT 502.000 430.300 502.800 430.400 ;
        RECT 450.800 429.700 502.800 430.300 ;
        RECT 450.800 429.600 451.600 429.700 ;
        RECT 468.400 429.600 469.200 429.700 ;
        RECT 502.000 429.600 502.800 429.700 ;
        RECT 503.600 430.300 504.400 430.400 ;
        RECT 508.400 430.300 509.200 430.400 ;
        RECT 529.200 430.300 530.000 430.400 ;
        RECT 503.600 429.700 530.000 430.300 ;
        RECT 503.600 429.600 504.400 429.700 ;
        RECT 508.400 429.600 509.200 429.700 ;
        RECT 529.200 429.600 530.000 429.700 ;
        RECT 550.000 430.300 550.800 430.400 ;
        RECT 583.600 430.300 584.400 430.400 ;
        RECT 550.000 429.700 584.400 430.300 ;
        RECT 550.000 429.600 550.800 429.700 ;
        RECT 583.600 429.600 584.400 429.700 ;
        RECT 630.000 430.300 630.800 430.400 ;
        RECT 631.600 430.300 632.400 430.400 ;
        RECT 630.000 429.700 632.400 430.300 ;
        RECT 630.000 429.600 630.800 429.700 ;
        RECT 631.600 429.600 632.400 429.700 ;
        RECT 332.400 427.700 347.500 428.300 ;
        RECT 348.400 428.300 349.200 428.400 ;
        RECT 359.600 428.300 360.400 428.400 ;
        RECT 348.400 427.700 360.400 428.300 ;
        RECT 332.400 427.600 333.200 427.700 ;
        RECT 348.400 427.600 349.200 427.700 ;
        RECT 359.600 427.600 360.400 427.700 ;
        RECT 375.600 428.300 376.400 428.400 ;
        RECT 385.200 428.300 386.000 428.400 ;
        RECT 375.600 427.700 386.000 428.300 ;
        RECT 375.600 427.600 376.400 427.700 ;
        RECT 385.200 427.600 386.000 427.700 ;
        RECT 391.600 428.300 392.400 428.400 ;
        RECT 396.400 428.300 397.200 428.400 ;
        RECT 391.600 427.700 397.200 428.300 ;
        RECT 391.600 427.600 392.400 427.700 ;
        RECT 396.400 427.600 397.200 427.700 ;
        RECT 463.600 428.300 464.400 428.400 ;
        RECT 506.800 428.300 507.600 428.400 ;
        RECT 463.600 427.700 507.600 428.300 ;
        RECT 463.600 427.600 464.400 427.700 ;
        RECT 506.800 427.600 507.600 427.700 ;
        RECT 522.800 428.300 523.600 428.400 ;
        RECT 534.000 428.300 534.800 428.400 ;
        RECT 535.600 428.300 536.400 428.400 ;
        RECT 561.200 428.300 562.000 428.400 ;
        RECT 522.800 427.700 562.000 428.300 ;
        RECT 522.800 427.600 523.600 427.700 ;
        RECT 534.000 427.600 534.800 427.700 ;
        RECT 535.600 427.600 536.400 427.700 ;
        RECT 561.200 427.600 562.000 427.700 ;
        RECT 574.000 428.300 574.800 428.400 ;
        RECT 599.600 428.300 600.400 428.400 ;
        RECT 574.000 427.700 600.400 428.300 ;
        RECT 574.000 427.600 574.800 427.700 ;
        RECT 599.600 427.600 600.400 427.700 ;
        RECT 631.600 428.300 632.400 428.400 ;
        RECT 658.800 428.300 659.600 428.400 ;
        RECT 631.600 427.700 659.600 428.300 ;
        RECT 631.600 427.600 632.400 427.700 ;
        RECT 658.800 427.600 659.600 427.700 ;
        RECT 63.600 426.300 64.400 426.400 ;
        RECT 79.600 426.300 80.400 426.400 ;
        RECT 87.600 426.300 88.400 426.400 ;
        RECT 63.600 425.700 88.400 426.300 ;
        RECT 63.600 425.600 64.400 425.700 ;
        RECT 79.600 425.600 80.400 425.700 ;
        RECT 87.600 425.600 88.400 425.700 ;
        RECT 180.400 426.300 181.200 426.400 ;
        RECT 185.200 426.300 186.000 426.400 ;
        RECT 180.400 425.700 186.000 426.300 ;
        RECT 180.400 425.600 181.200 425.700 ;
        RECT 185.200 425.600 186.000 425.700 ;
        RECT 188.400 426.300 189.200 426.400 ;
        RECT 193.200 426.300 194.000 426.400 ;
        RECT 188.400 425.700 194.000 426.300 ;
        RECT 188.400 425.600 189.200 425.700 ;
        RECT 193.200 425.600 194.000 425.700 ;
        RECT 214.000 426.300 214.800 426.400 ;
        RECT 217.200 426.300 218.000 426.400 ;
        RECT 214.000 425.700 218.000 426.300 ;
        RECT 214.000 425.600 214.800 425.700 ;
        RECT 217.200 425.600 218.000 425.700 ;
        RECT 234.800 426.300 235.600 426.400 ;
        RECT 241.200 426.300 242.000 426.400 ;
        RECT 234.800 425.700 242.000 426.300 ;
        RECT 234.800 425.600 235.600 425.700 ;
        RECT 241.200 425.600 242.000 425.700 ;
        RECT 244.400 426.300 245.200 426.400 ;
        RECT 257.200 426.300 258.000 426.400 ;
        RECT 281.200 426.300 282.000 426.400 ;
        RECT 244.400 425.700 282.000 426.300 ;
        RECT 244.400 425.600 245.200 425.700 ;
        RECT 257.200 425.600 258.000 425.700 ;
        RECT 281.200 425.600 282.000 425.700 ;
        RECT 292.400 426.300 293.200 426.400 ;
        RECT 298.800 426.300 299.600 426.400 ;
        RECT 292.400 425.700 299.600 426.300 ;
        RECT 292.400 425.600 293.200 425.700 ;
        RECT 298.800 425.600 299.600 425.700 ;
        RECT 306.800 426.300 307.600 426.400 ;
        RECT 319.600 426.300 320.400 426.400 ;
        RECT 306.800 425.700 320.400 426.300 ;
        RECT 306.800 425.600 307.600 425.700 ;
        RECT 319.600 425.600 320.400 425.700 ;
        RECT 321.200 426.300 322.000 426.400 ;
        RECT 326.000 426.300 326.800 426.400 ;
        RECT 321.200 425.700 326.800 426.300 ;
        RECT 321.200 425.600 322.000 425.700 ;
        RECT 326.000 425.600 326.800 425.700 ;
        RECT 329.200 426.300 330.000 426.400 ;
        RECT 335.600 426.300 336.400 426.400 ;
        RECT 329.200 425.700 336.400 426.300 ;
        RECT 329.200 425.600 330.000 425.700 ;
        RECT 335.600 425.600 336.400 425.700 ;
        RECT 337.200 426.300 338.000 426.400 ;
        RECT 343.600 426.300 344.400 426.400 ;
        RECT 337.200 425.700 344.400 426.300 ;
        RECT 337.200 425.600 338.000 425.700 ;
        RECT 343.600 425.600 344.400 425.700 ;
        RECT 346.800 426.300 347.600 426.400 ;
        RECT 354.800 426.300 355.600 426.400 ;
        RECT 346.800 425.700 355.600 426.300 ;
        RECT 346.800 425.600 347.600 425.700 ;
        RECT 354.800 425.600 355.600 425.700 ;
        RECT 361.200 426.300 362.000 426.400 ;
        RECT 378.800 426.300 379.600 426.400 ;
        RECT 361.200 425.700 379.600 426.300 ;
        RECT 361.200 425.600 362.000 425.700 ;
        RECT 378.800 425.600 379.600 425.700 ;
        RECT 394.800 426.300 395.600 426.400 ;
        RECT 398.000 426.300 398.800 426.400 ;
        RECT 442.800 426.300 443.600 426.400 ;
        RECT 394.800 425.700 443.600 426.300 ;
        RECT 394.800 425.600 395.600 425.700 ;
        RECT 398.000 425.600 398.800 425.700 ;
        RECT 442.800 425.600 443.600 425.700 ;
        RECT 481.200 426.300 482.000 426.400 ;
        RECT 519.600 426.300 520.400 426.400 ;
        RECT 481.200 425.700 520.400 426.300 ;
        RECT 481.200 425.600 482.000 425.700 ;
        RECT 519.600 425.600 520.400 425.700 ;
        RECT 526.000 426.300 526.800 426.400 ;
        RECT 542.000 426.300 542.800 426.400 ;
        RECT 561.200 426.300 562.000 426.400 ;
        RECT 526.000 425.700 562.000 426.300 ;
        RECT 526.000 425.600 526.800 425.700 ;
        RECT 542.000 425.600 542.800 425.700 ;
        RECT 561.200 425.600 562.000 425.700 ;
        RECT 570.800 426.300 571.600 426.400 ;
        RECT 594.800 426.300 595.600 426.400 ;
        RECT 617.200 426.300 618.000 426.400 ;
        RECT 666.800 426.300 667.600 426.400 ;
        RECT 570.800 425.700 667.600 426.300 ;
        RECT 570.800 425.600 571.600 425.700 ;
        RECT 594.800 425.600 595.600 425.700 ;
        RECT 617.200 425.600 618.000 425.700 ;
        RECT 666.800 425.600 667.600 425.700 ;
        RECT 46.000 424.300 46.800 424.400 ;
        RECT 87.600 424.300 88.400 424.400 ;
        RECT 46.000 423.700 88.400 424.300 ;
        RECT 46.000 423.600 46.800 423.700 ;
        RECT 87.600 423.600 88.400 423.700 ;
        RECT 159.600 424.300 160.400 424.400 ;
        RECT 164.400 424.300 165.200 424.400 ;
        RECT 159.600 423.700 165.200 424.300 ;
        RECT 159.600 423.600 160.400 423.700 ;
        RECT 164.400 423.600 165.200 423.700 ;
        RECT 185.200 424.300 186.000 424.400 ;
        RECT 206.000 424.300 206.800 424.400 ;
        RECT 185.200 423.700 206.800 424.300 ;
        RECT 185.200 423.600 186.000 423.700 ;
        RECT 206.000 423.600 206.800 423.700 ;
        RECT 308.400 424.300 309.200 424.400 ;
        RECT 322.800 424.300 323.600 424.400 ;
        RECT 308.400 423.700 323.600 424.300 ;
        RECT 308.400 423.600 309.200 423.700 ;
        RECT 322.800 423.600 323.600 423.700 ;
        RECT 346.800 424.300 347.600 424.400 ;
        RECT 348.400 424.300 349.200 424.400 ;
        RECT 346.800 423.700 349.200 424.300 ;
        RECT 346.800 423.600 347.600 423.700 ;
        RECT 348.400 423.600 349.200 423.700 ;
        RECT 356.400 424.300 357.200 424.400 ;
        RECT 366.000 424.300 366.800 424.400 ;
        RECT 356.400 423.700 366.800 424.300 ;
        RECT 356.400 423.600 357.200 423.700 ;
        RECT 366.000 423.600 366.800 423.700 ;
        RECT 370.800 424.300 371.600 424.400 ;
        RECT 388.400 424.300 389.200 424.400 ;
        RECT 370.800 423.700 389.200 424.300 ;
        RECT 370.800 423.600 371.600 423.700 ;
        RECT 388.400 423.600 389.200 423.700 ;
        RECT 502.000 424.300 502.800 424.400 ;
        RECT 518.000 424.300 518.800 424.400 ;
        RECT 502.000 423.700 518.800 424.300 ;
        RECT 502.000 423.600 502.800 423.700 ;
        RECT 518.000 423.600 518.800 423.700 ;
        RECT 519.600 424.300 520.400 424.400 ;
        RECT 526.000 424.300 526.800 424.400 ;
        RECT 519.600 423.700 526.800 424.300 ;
        RECT 519.600 423.600 520.400 423.700 ;
        RECT 526.000 423.600 526.800 423.700 ;
        RECT 529.200 424.300 530.000 424.400 ;
        RECT 535.600 424.300 536.400 424.400 ;
        RECT 562.800 424.300 563.600 424.400 ;
        RECT 529.200 423.700 563.600 424.300 ;
        RECT 529.200 423.600 530.000 423.700 ;
        RECT 535.600 423.600 536.400 423.700 ;
        RECT 562.800 423.600 563.600 423.700 ;
        RECT 601.200 424.300 602.000 424.400 ;
        RECT 607.600 424.300 608.400 424.400 ;
        RECT 601.200 423.700 608.400 424.300 ;
        RECT 601.200 423.600 602.000 423.700 ;
        RECT 607.600 423.600 608.400 423.700 ;
        RECT 615.600 424.300 616.400 424.400 ;
        RECT 633.200 424.300 634.000 424.400 ;
        RECT 615.600 423.700 634.000 424.300 ;
        RECT 615.600 423.600 616.400 423.700 ;
        RECT 633.200 423.600 634.000 423.700 ;
        RECT 647.600 424.300 648.400 424.400 ;
        RECT 650.800 424.300 651.600 424.400 ;
        RECT 647.600 423.700 651.600 424.300 ;
        RECT 647.600 423.600 648.400 423.700 ;
        RECT 650.800 423.600 651.600 423.700 ;
        RECT 73.200 422.300 74.000 422.400 ;
        RECT 78.000 422.300 78.800 422.400 ;
        RECT 119.600 422.300 120.400 422.400 ;
        RECT 134.000 422.300 134.800 422.400 ;
        RECT 170.800 422.300 171.600 422.400 ;
        RECT 73.200 421.700 171.600 422.300 ;
        RECT 73.200 421.600 74.000 421.700 ;
        RECT 78.000 421.600 78.800 421.700 ;
        RECT 119.600 421.600 120.400 421.700 ;
        RECT 134.000 421.600 134.800 421.700 ;
        RECT 170.800 421.600 171.600 421.700 ;
        RECT 209.200 422.300 210.000 422.400 ;
        RECT 244.400 422.300 245.200 422.400 ;
        RECT 209.200 421.700 245.200 422.300 ;
        RECT 209.200 421.600 210.000 421.700 ;
        RECT 244.400 421.600 245.200 421.700 ;
        RECT 321.200 422.300 322.000 422.400 ;
        RECT 340.400 422.300 341.200 422.400 ;
        RECT 321.200 421.700 341.200 422.300 ;
        RECT 321.200 421.600 322.000 421.700 ;
        RECT 340.400 421.600 341.200 421.700 ;
        RECT 343.600 422.300 344.400 422.400 ;
        RECT 345.200 422.300 346.000 422.400 ;
        RECT 343.600 421.700 346.000 422.300 ;
        RECT 343.600 421.600 344.400 421.700 ;
        RECT 345.200 421.600 346.000 421.700 ;
        RECT 346.800 422.300 347.600 422.400 ;
        RECT 383.600 422.300 384.400 422.400 ;
        RECT 346.800 421.700 384.400 422.300 ;
        RECT 346.800 421.600 347.600 421.700 ;
        RECT 383.600 421.600 384.400 421.700 ;
        RECT 425.200 422.300 426.000 422.400 ;
        RECT 430.000 422.300 430.800 422.400 ;
        RECT 425.200 421.700 430.800 422.300 ;
        RECT 425.200 421.600 426.000 421.700 ;
        RECT 430.000 421.600 430.800 421.700 ;
        RECT 470.000 422.300 470.800 422.400 ;
        RECT 484.400 422.300 485.200 422.400 ;
        RECT 470.000 421.700 485.200 422.300 ;
        RECT 470.000 421.600 470.800 421.700 ;
        RECT 484.400 421.600 485.200 421.700 ;
        RECT 505.200 422.300 506.000 422.400 ;
        RECT 527.600 422.300 528.400 422.400 ;
        RECT 505.200 421.700 528.400 422.300 ;
        RECT 505.200 421.600 506.000 421.700 ;
        RECT 527.600 421.600 528.400 421.700 ;
        RECT 551.600 422.300 552.400 422.400 ;
        RECT 569.200 422.300 570.000 422.400 ;
        RECT 551.600 421.700 570.000 422.300 ;
        RECT 551.600 421.600 552.400 421.700 ;
        RECT 569.200 421.600 570.000 421.700 ;
        RECT 644.400 422.300 645.200 422.400 ;
        RECT 670.000 422.300 670.800 422.400 ;
        RECT 644.400 421.700 670.800 422.300 ;
        RECT 644.400 421.600 645.200 421.700 ;
        RECT 670.000 421.600 670.800 421.700 ;
        RECT 65.200 419.600 66.000 420.400 ;
        RECT 90.800 419.600 91.600 420.400 ;
        RECT 100.400 420.300 101.200 420.400 ;
        RECT 103.600 420.300 104.400 420.400 ;
        RECT 100.400 419.700 104.400 420.300 ;
        RECT 100.400 419.600 101.200 419.700 ;
        RECT 103.600 419.600 104.400 419.700 ;
        RECT 140.400 420.300 141.200 420.400 ;
        RECT 167.600 420.300 168.400 420.400 ;
        RECT 174.000 420.300 174.800 420.400 ;
        RECT 140.400 419.700 174.800 420.300 ;
        RECT 140.400 419.600 141.200 419.700 ;
        RECT 167.600 419.600 168.400 419.700 ;
        RECT 174.000 419.600 174.800 419.700 ;
        RECT 212.400 420.300 213.200 420.400 ;
        RECT 215.600 420.300 216.400 420.400 ;
        RECT 212.400 419.700 216.400 420.300 ;
        RECT 212.400 419.600 213.200 419.700 ;
        RECT 215.600 419.600 216.400 419.700 ;
        RECT 270.000 420.300 270.800 420.400 ;
        RECT 279.600 420.300 280.400 420.400 ;
        RECT 270.000 419.700 280.400 420.300 ;
        RECT 270.000 419.600 270.800 419.700 ;
        RECT 279.600 419.600 280.400 419.700 ;
        RECT 281.200 420.300 282.000 420.400 ;
        RECT 286.000 420.300 286.800 420.400 ;
        RECT 281.200 419.700 286.800 420.300 ;
        RECT 281.200 419.600 282.000 419.700 ;
        RECT 286.000 419.600 286.800 419.700 ;
        RECT 334.000 420.300 334.800 420.400 ;
        RECT 343.600 420.300 344.400 420.400 ;
        RECT 334.000 419.700 344.400 420.300 ;
        RECT 334.000 419.600 334.800 419.700 ;
        RECT 343.600 419.600 344.400 419.700 ;
        RECT 350.000 420.300 350.800 420.400 ;
        RECT 353.200 420.300 354.000 420.400 ;
        RECT 370.800 420.300 371.600 420.400 ;
        RECT 385.200 420.300 386.000 420.400 ;
        RECT 350.000 419.700 386.000 420.300 ;
        RECT 350.000 419.600 350.800 419.700 ;
        RECT 353.200 419.600 354.000 419.700 ;
        RECT 370.800 419.600 371.600 419.700 ;
        RECT 385.200 419.600 386.000 419.700 ;
        RECT 436.400 420.300 437.200 420.400 ;
        RECT 441.200 420.300 442.000 420.400 ;
        RECT 436.400 419.700 442.000 420.300 ;
        RECT 436.400 419.600 437.200 419.700 ;
        RECT 441.200 419.600 442.000 419.700 ;
        RECT 449.200 420.300 450.000 420.400 ;
        RECT 540.400 420.300 541.200 420.400 ;
        RECT 554.800 420.300 555.600 420.400 ;
        RECT 449.200 419.700 555.600 420.300 ;
        RECT 449.200 419.600 450.000 419.700 ;
        RECT 540.400 419.600 541.200 419.700 ;
        RECT 554.800 419.600 555.600 419.700 ;
        RECT 34.800 418.300 35.600 418.400 ;
        RECT 55.600 418.300 56.400 418.400 ;
        RECT 58.800 418.300 59.600 418.400 ;
        RECT 34.800 417.700 59.600 418.300 ;
        RECT 34.800 417.600 35.600 417.700 ;
        RECT 55.600 417.600 56.400 417.700 ;
        RECT 58.800 417.600 59.600 417.700 ;
        RECT 90.800 418.300 91.600 418.400 ;
        RECT 97.200 418.300 98.000 418.400 ;
        RECT 90.800 417.700 98.000 418.300 ;
        RECT 90.800 417.600 91.600 417.700 ;
        RECT 97.200 417.600 98.000 417.700 ;
        RECT 154.800 418.300 155.600 418.400 ;
        RECT 182.000 418.300 182.800 418.400 ;
        RECT 154.800 417.700 182.800 418.300 ;
        RECT 154.800 417.600 155.600 417.700 ;
        RECT 182.000 417.600 182.800 417.700 ;
        RECT 292.400 418.300 293.200 418.400 ;
        RECT 358.000 418.300 358.800 418.400 ;
        RECT 362.800 418.300 363.600 418.400 ;
        RECT 378.800 418.300 379.600 418.400 ;
        RECT 292.400 417.700 379.600 418.300 ;
        RECT 292.400 417.600 293.200 417.700 ;
        RECT 358.000 417.600 358.800 417.700 ;
        RECT 362.800 417.600 363.600 417.700 ;
        RECT 378.800 417.600 379.600 417.700 ;
        RECT 383.600 418.300 384.400 418.400 ;
        RECT 399.600 418.300 400.400 418.400 ;
        RECT 383.600 417.700 400.400 418.300 ;
        RECT 383.600 417.600 384.400 417.700 ;
        RECT 399.600 417.600 400.400 417.700 ;
        RECT 463.600 418.300 464.400 418.400 ;
        RECT 492.400 418.300 493.200 418.400 ;
        RECT 463.600 417.700 493.200 418.300 ;
        RECT 463.600 417.600 464.400 417.700 ;
        RECT 492.400 417.600 493.200 417.700 ;
        RECT 554.800 418.300 555.600 418.400 ;
        RECT 598.000 418.300 598.800 418.400 ;
        RECT 554.800 417.700 598.800 418.300 ;
        RECT 554.800 417.600 555.600 417.700 ;
        RECT 598.000 417.600 598.800 417.700 ;
        RECT 22.000 416.300 22.800 416.400 ;
        RECT 30.000 416.300 30.800 416.400 ;
        RECT 22.000 415.700 30.800 416.300 ;
        RECT 22.000 415.600 22.800 415.700 ;
        RECT 30.000 415.600 30.800 415.700 ;
        RECT 31.600 416.300 32.400 416.400 ;
        RECT 42.800 416.300 43.600 416.400 ;
        RECT 50.800 416.300 51.600 416.400 ;
        RECT 31.600 415.700 51.600 416.300 ;
        RECT 31.600 415.600 32.400 415.700 ;
        RECT 42.800 415.600 43.600 415.700 ;
        RECT 50.800 415.600 51.600 415.700 ;
        RECT 130.800 416.300 131.600 416.400 ;
        RECT 135.600 416.300 136.400 416.400 ;
        RECT 130.800 415.700 136.400 416.300 ;
        RECT 130.800 415.600 131.600 415.700 ;
        RECT 135.600 415.600 136.400 415.700 ;
        RECT 169.200 416.300 170.000 416.400 ;
        RECT 170.800 416.300 171.600 416.400 ;
        RECT 169.200 415.700 171.600 416.300 ;
        RECT 169.200 415.600 170.000 415.700 ;
        RECT 170.800 415.600 171.600 415.700 ;
        RECT 236.400 416.300 237.200 416.400 ;
        RECT 257.200 416.300 258.000 416.400 ;
        RECT 278.000 416.300 278.800 416.400 ;
        RECT 236.400 415.700 278.800 416.300 ;
        RECT 236.400 415.600 237.200 415.700 ;
        RECT 257.200 415.600 258.000 415.700 ;
        RECT 278.000 415.600 278.800 415.700 ;
        RECT 303.600 416.300 304.400 416.400 ;
        RECT 316.400 416.300 317.200 416.400 ;
        RECT 303.600 415.700 317.200 416.300 ;
        RECT 303.600 415.600 304.400 415.700 ;
        RECT 316.400 415.600 317.200 415.700 ;
        RECT 324.400 416.300 325.200 416.400 ;
        RECT 334.000 416.300 334.800 416.400 ;
        RECT 346.800 416.300 347.600 416.400 ;
        RECT 324.400 415.700 347.600 416.300 ;
        RECT 324.400 415.600 325.200 415.700 ;
        RECT 334.000 415.600 334.800 415.700 ;
        RECT 346.800 415.600 347.600 415.700 ;
        RECT 348.400 416.300 349.200 416.400 ;
        RECT 361.200 416.300 362.000 416.400 ;
        RECT 348.400 415.700 362.000 416.300 ;
        RECT 348.400 415.600 349.200 415.700 ;
        RECT 361.200 415.600 362.000 415.700 ;
        RECT 377.200 416.300 378.000 416.400 ;
        RECT 390.000 416.300 390.800 416.400 ;
        RECT 391.600 416.300 392.400 416.400 ;
        RECT 377.200 415.700 392.400 416.300 ;
        RECT 377.200 415.600 378.000 415.700 ;
        RECT 390.000 415.600 390.800 415.700 ;
        RECT 391.600 415.600 392.400 415.700 ;
        RECT 394.800 416.300 395.600 416.400 ;
        RECT 401.200 416.300 402.000 416.400 ;
        RECT 394.800 415.700 402.000 416.300 ;
        RECT 394.800 415.600 395.600 415.700 ;
        RECT 401.200 415.600 402.000 415.700 ;
        RECT 422.000 416.300 422.800 416.400 ;
        RECT 433.200 416.300 434.000 416.400 ;
        RECT 452.400 416.300 453.200 416.400 ;
        RECT 466.800 416.300 467.600 416.400 ;
        RECT 422.000 415.700 467.600 416.300 ;
        RECT 422.000 415.600 422.800 415.700 ;
        RECT 433.200 415.600 434.000 415.700 ;
        RECT 452.400 415.600 453.200 415.700 ;
        RECT 466.800 415.600 467.600 415.700 ;
        RECT 540.400 416.300 541.200 416.400 ;
        RECT 586.800 416.300 587.600 416.400 ;
        RECT 540.400 415.700 587.600 416.300 ;
        RECT 540.400 415.600 541.200 415.700 ;
        RECT 586.800 415.600 587.600 415.700 ;
        RECT 596.400 416.300 597.200 416.400 ;
        RECT 612.400 416.300 613.200 416.400 ;
        RECT 596.400 415.700 613.200 416.300 ;
        RECT 596.400 415.600 597.200 415.700 ;
        RECT 612.400 415.600 613.200 415.700 ;
        RECT 670.000 416.300 670.800 416.400 ;
        RECT 676.400 416.300 677.200 416.400 ;
        RECT 670.000 415.700 677.200 416.300 ;
        RECT 670.000 415.600 670.800 415.700 ;
        RECT 676.400 415.600 677.200 415.700 ;
        RECT 22.000 414.300 22.800 414.400 ;
        RECT 26.800 414.300 27.600 414.400 ;
        RECT 22.000 413.700 27.600 414.300 ;
        RECT 22.000 413.600 22.800 413.700 ;
        RECT 26.800 413.600 27.600 413.700 ;
        RECT 50.800 414.300 51.600 414.400 ;
        RECT 79.600 414.300 80.400 414.400 ;
        RECT 50.800 413.700 80.400 414.300 ;
        RECT 50.800 413.600 51.600 413.700 ;
        RECT 79.600 413.600 80.400 413.700 ;
        RECT 84.400 414.300 85.200 414.400 ;
        RECT 98.800 414.300 99.600 414.400 ;
        RECT 84.400 413.700 99.600 414.300 ;
        RECT 84.400 413.600 85.200 413.700 ;
        RECT 98.800 413.600 99.600 413.700 ;
        RECT 103.600 414.300 104.400 414.400 ;
        RECT 116.400 414.300 117.200 414.400 ;
        RECT 103.600 413.700 117.200 414.300 ;
        RECT 103.600 413.600 104.400 413.700 ;
        RECT 116.400 413.600 117.200 413.700 ;
        RECT 124.400 414.300 125.200 414.400 ;
        RECT 137.200 414.300 138.000 414.400 ;
        RECT 124.400 413.700 138.000 414.300 ;
        RECT 124.400 413.600 125.200 413.700 ;
        RECT 137.200 413.600 138.000 413.700 ;
        RECT 151.600 414.300 152.400 414.400 ;
        RECT 170.800 414.300 171.600 414.400 ;
        RECT 183.600 414.300 184.400 414.400 ;
        RECT 194.800 414.300 195.600 414.400 ;
        RECT 151.600 413.700 195.600 414.300 ;
        RECT 151.600 413.600 152.400 413.700 ;
        RECT 170.800 413.600 171.600 413.700 ;
        RECT 183.600 413.600 184.400 413.700 ;
        RECT 194.800 413.600 195.600 413.700 ;
        RECT 220.400 414.300 221.200 414.400 ;
        RECT 226.800 414.300 227.600 414.400 ;
        RECT 238.000 414.300 238.800 414.400 ;
        RECT 220.400 413.700 238.800 414.300 ;
        RECT 220.400 413.600 221.200 413.700 ;
        RECT 226.800 413.600 227.600 413.700 ;
        RECT 238.000 413.600 238.800 413.700 ;
        RECT 247.600 414.300 248.400 414.400 ;
        RECT 258.800 414.300 259.600 414.400 ;
        RECT 247.600 413.700 259.600 414.300 ;
        RECT 247.600 413.600 248.400 413.700 ;
        RECT 258.800 413.600 259.600 413.700 ;
        RECT 326.000 414.300 326.800 414.400 ;
        RECT 362.800 414.300 363.600 414.400 ;
        RECT 386.800 414.300 387.600 414.400 ;
        RECT 326.000 413.700 387.600 414.300 ;
        RECT 326.000 413.600 326.800 413.700 ;
        RECT 362.800 413.600 363.600 413.700 ;
        RECT 386.800 413.600 387.600 413.700 ;
        RECT 393.200 414.300 394.000 414.400 ;
        RECT 398.000 414.300 398.800 414.400 ;
        RECT 393.200 413.700 398.800 414.300 ;
        RECT 393.200 413.600 394.000 413.700 ;
        RECT 398.000 413.600 398.800 413.700 ;
        RECT 486.000 414.300 486.800 414.400 ;
        RECT 489.200 414.300 490.000 414.400 ;
        RECT 486.000 413.700 490.000 414.300 ;
        RECT 486.000 413.600 486.800 413.700 ;
        RECT 489.200 413.600 490.000 413.700 ;
        RECT 497.200 414.300 498.000 414.400 ;
        RECT 502.000 414.300 502.800 414.400 ;
        RECT 497.200 413.700 502.800 414.300 ;
        RECT 497.200 413.600 498.000 413.700 ;
        RECT 502.000 413.600 502.800 413.700 ;
        RECT 506.800 414.300 507.600 414.400 ;
        RECT 529.200 414.300 530.000 414.400 ;
        RECT 506.800 413.700 530.000 414.300 ;
        RECT 506.800 413.600 507.600 413.700 ;
        RECT 529.200 413.600 530.000 413.700 ;
        RECT 561.200 414.300 562.000 414.400 ;
        RECT 564.400 414.300 565.200 414.400 ;
        RECT 561.200 413.700 565.200 414.300 ;
        RECT 561.200 413.600 562.000 413.700 ;
        RECT 564.400 413.600 565.200 413.700 ;
        RECT 566.000 414.300 566.800 414.400 ;
        RECT 567.600 414.300 568.400 414.400 ;
        RECT 566.000 413.700 568.400 414.300 ;
        RECT 566.000 413.600 566.800 413.700 ;
        RECT 567.600 413.600 568.400 413.700 ;
        RECT 622.000 414.300 622.800 414.400 ;
        RECT 623.600 414.300 624.400 414.400 ;
        RECT 631.600 414.300 632.400 414.400 ;
        RECT 622.000 413.700 632.400 414.300 ;
        RECT 622.000 413.600 622.800 413.700 ;
        RECT 623.600 413.600 624.400 413.700 ;
        RECT 631.600 413.600 632.400 413.700 ;
        RECT 670.000 414.300 670.800 414.400 ;
        RECT 682.800 414.300 683.600 414.400 ;
        RECT 670.000 413.700 683.600 414.300 ;
        RECT 670.000 413.600 670.800 413.700 ;
        RECT 682.800 413.600 683.600 413.700 ;
        RECT 7.600 412.300 8.400 412.400 ;
        RECT 23.600 412.300 24.400 412.400 ;
        RECT 7.600 411.700 24.400 412.300 ;
        RECT 7.600 411.600 8.400 411.700 ;
        RECT 23.600 411.600 24.400 411.700 ;
        RECT 52.400 412.300 53.200 412.400 ;
        RECT 58.800 412.300 59.600 412.400 ;
        RECT 52.400 411.700 59.600 412.300 ;
        RECT 52.400 411.600 53.200 411.700 ;
        RECT 58.800 411.600 59.600 411.700 ;
        RECT 62.000 412.300 62.800 412.400 ;
        RECT 68.400 412.300 69.200 412.400 ;
        RECT 62.000 411.700 69.200 412.300 ;
        RECT 62.000 411.600 62.800 411.700 ;
        RECT 68.400 411.600 69.200 411.700 ;
        RECT 92.400 412.300 93.200 412.400 ;
        RECT 129.200 412.300 130.000 412.400 ;
        RECT 150.000 412.300 150.800 412.400 ;
        RECT 92.400 411.700 150.800 412.300 ;
        RECT 92.400 411.600 93.200 411.700 ;
        RECT 129.200 411.600 130.000 411.700 ;
        RECT 150.000 411.600 150.800 411.700 ;
        RECT 164.400 412.300 165.200 412.400 ;
        RECT 177.200 412.300 178.000 412.400 ;
        RECT 180.400 412.300 181.200 412.400 ;
        RECT 164.400 411.700 181.200 412.300 ;
        RECT 164.400 411.600 165.200 411.700 ;
        RECT 177.200 411.600 178.000 411.700 ;
        RECT 180.400 411.600 181.200 411.700 ;
        RECT 223.600 412.300 224.400 412.400 ;
        RECT 244.400 412.300 245.200 412.400 ;
        RECT 223.600 411.700 245.200 412.300 ;
        RECT 223.600 411.600 224.400 411.700 ;
        RECT 244.400 411.600 245.200 411.700 ;
        RECT 327.600 412.300 328.400 412.400 ;
        RECT 353.200 412.300 354.000 412.400 ;
        RECT 327.600 411.700 354.000 412.300 ;
        RECT 327.600 411.600 328.400 411.700 ;
        RECT 353.200 411.600 354.000 411.700 ;
        RECT 356.400 412.300 357.200 412.400 ;
        RECT 359.600 412.300 360.400 412.400 ;
        RECT 356.400 411.700 360.400 412.300 ;
        RECT 356.400 411.600 357.200 411.700 ;
        RECT 359.600 411.600 360.400 411.700 ;
        RECT 372.400 412.300 373.200 412.400 ;
        RECT 375.600 412.300 376.400 412.400 ;
        RECT 382.000 412.300 382.800 412.400 ;
        RECT 372.400 411.700 382.800 412.300 ;
        RECT 372.400 411.600 373.200 411.700 ;
        RECT 375.600 411.600 376.400 411.700 ;
        RECT 382.000 411.600 382.800 411.700 ;
        RECT 388.400 412.300 389.200 412.400 ;
        RECT 402.800 412.300 403.600 412.400 ;
        RECT 388.400 411.700 403.600 412.300 ;
        RECT 388.400 411.600 389.200 411.700 ;
        RECT 402.800 411.600 403.600 411.700 ;
        RECT 447.600 412.300 448.400 412.400 ;
        RECT 450.800 412.300 451.600 412.400 ;
        RECT 454.000 412.300 454.800 412.400 ;
        RECT 447.600 411.700 454.800 412.300 ;
        RECT 447.600 411.600 448.400 411.700 ;
        RECT 450.800 411.600 451.600 411.700 ;
        RECT 454.000 411.600 454.800 411.700 ;
        RECT 487.600 412.300 488.400 412.400 ;
        RECT 495.600 412.300 496.400 412.400 ;
        RECT 503.600 412.300 504.400 412.400 ;
        RECT 538.800 412.300 539.600 412.400 ;
        RECT 551.600 412.300 552.400 412.400 ;
        RECT 487.600 411.700 552.400 412.300 ;
        RECT 487.600 411.600 488.400 411.700 ;
        RECT 495.600 411.600 496.400 411.700 ;
        RECT 503.600 411.600 504.400 411.700 ;
        RECT 538.800 411.600 539.600 411.700 ;
        RECT 551.600 411.600 552.400 411.700 ;
        RECT 554.800 412.300 555.600 412.400 ;
        RECT 559.600 412.300 560.400 412.400 ;
        RECT 554.800 411.700 560.400 412.300 ;
        RECT 554.800 411.600 555.600 411.700 ;
        RECT 559.600 411.600 560.400 411.700 ;
        RECT 567.600 412.300 568.400 412.400 ;
        RECT 622.000 412.300 622.800 412.400 ;
        RECT 567.600 411.700 622.800 412.300 ;
        RECT 567.600 411.600 568.400 411.700 ;
        RECT 622.000 411.600 622.800 411.700 ;
        RECT 18.800 410.300 19.600 410.400 ;
        RECT 26.800 410.300 27.600 410.400 ;
        RECT 18.800 409.700 27.600 410.300 ;
        RECT 18.800 409.600 19.600 409.700 ;
        RECT 26.800 409.600 27.600 409.700 ;
        RECT 57.200 410.300 58.000 410.400 ;
        RECT 62.000 410.300 62.800 410.400 ;
        RECT 57.200 409.700 62.800 410.300 ;
        RECT 57.200 409.600 58.000 409.700 ;
        RECT 62.000 409.600 62.800 409.700 ;
        RECT 63.600 410.300 64.400 410.400 ;
        RECT 65.200 410.300 66.000 410.400 ;
        RECT 114.800 410.300 115.600 410.400 ;
        RECT 63.600 409.700 115.600 410.300 ;
        RECT 63.600 409.600 64.400 409.700 ;
        RECT 65.200 409.600 66.000 409.700 ;
        RECT 114.800 409.600 115.600 409.700 ;
        RECT 137.200 410.300 138.000 410.400 ;
        RECT 154.800 410.300 155.600 410.400 ;
        RECT 137.200 409.700 155.600 410.300 ;
        RECT 137.200 409.600 138.000 409.700 ;
        RECT 154.800 409.600 155.600 409.700 ;
        RECT 174.000 410.300 174.800 410.400 ;
        RECT 188.400 410.300 189.200 410.400 ;
        RECT 174.000 409.700 189.200 410.300 ;
        RECT 174.000 409.600 174.800 409.700 ;
        RECT 188.400 409.600 189.200 409.700 ;
        RECT 241.200 410.300 242.000 410.400 ;
        RECT 247.600 410.300 248.400 410.400 ;
        RECT 241.200 409.700 248.400 410.300 ;
        RECT 241.200 409.600 242.000 409.700 ;
        RECT 247.600 409.600 248.400 409.700 ;
        RECT 303.600 410.300 304.400 410.400 ;
        RECT 332.400 410.300 333.200 410.400 ;
        RECT 335.600 410.300 336.400 410.400 ;
        RECT 303.600 409.700 336.400 410.300 ;
        RECT 303.600 409.600 304.400 409.700 ;
        RECT 332.400 409.600 333.200 409.700 ;
        RECT 335.600 409.600 336.400 409.700 ;
        RECT 351.600 410.300 352.400 410.400 ;
        RECT 361.200 410.300 362.000 410.400 ;
        RECT 351.600 409.700 362.000 410.300 ;
        RECT 351.600 409.600 352.400 409.700 ;
        RECT 361.200 409.600 362.000 409.700 ;
        RECT 369.200 410.300 370.000 410.400 ;
        RECT 380.400 410.300 381.200 410.400 ;
        RECT 409.200 410.300 410.000 410.400 ;
        RECT 369.200 409.700 410.000 410.300 ;
        RECT 369.200 409.600 370.000 409.700 ;
        RECT 380.400 409.600 381.200 409.700 ;
        RECT 409.200 409.600 410.000 409.700 ;
        RECT 500.400 410.300 501.200 410.400 ;
        RECT 503.600 410.300 504.400 410.400 ;
        RECT 500.400 409.700 504.400 410.300 ;
        RECT 500.400 409.600 501.200 409.700 ;
        RECT 503.600 409.600 504.400 409.700 ;
        RECT 542.000 410.300 542.800 410.400 ;
        RECT 548.400 410.300 549.200 410.400 ;
        RECT 542.000 409.700 549.200 410.300 ;
        RECT 542.000 409.600 542.800 409.700 ;
        RECT 548.400 409.600 549.200 409.700 ;
        RECT 550.000 410.300 550.800 410.400 ;
        RECT 556.400 410.300 557.200 410.400 ;
        RECT 550.000 409.700 557.200 410.300 ;
        RECT 550.000 409.600 550.800 409.700 ;
        RECT 556.400 409.600 557.200 409.700 ;
        RECT 559.600 410.300 560.400 410.400 ;
        RECT 575.600 410.300 576.400 410.400 ;
        RECT 559.600 409.700 576.400 410.300 ;
        RECT 559.600 409.600 560.400 409.700 ;
        RECT 575.600 409.600 576.400 409.700 ;
        RECT 626.800 410.300 627.600 410.400 ;
        RECT 636.400 410.300 637.200 410.400 ;
        RECT 650.800 410.300 651.600 410.400 ;
        RECT 626.800 409.700 651.600 410.300 ;
        RECT 626.800 409.600 627.600 409.700 ;
        RECT 636.400 409.600 637.200 409.700 ;
        RECT 650.800 409.600 651.600 409.700 ;
        RECT 25.200 408.300 26.000 408.400 ;
        RECT 28.400 408.300 29.200 408.400 ;
        RECT 25.200 407.700 29.200 408.300 ;
        RECT 25.200 407.600 26.000 407.700 ;
        RECT 28.400 407.600 29.200 407.700 ;
        RECT 39.600 408.300 40.400 408.400 ;
        RECT 65.200 408.300 66.000 408.400 ;
        RECT 39.600 407.700 66.000 408.300 ;
        RECT 39.600 407.600 40.400 407.700 ;
        RECT 65.200 407.600 66.000 407.700 ;
        RECT 94.000 408.300 94.800 408.400 ;
        RECT 127.600 408.300 128.400 408.400 ;
        RECT 148.400 408.300 149.200 408.400 ;
        RECT 94.000 407.700 149.200 408.300 ;
        RECT 94.000 407.600 94.800 407.700 ;
        RECT 127.600 407.600 128.400 407.700 ;
        RECT 148.400 407.600 149.200 407.700 ;
        RECT 311.600 408.300 312.400 408.400 ;
        RECT 322.800 408.300 323.600 408.400 ;
        RECT 337.200 408.300 338.000 408.400 ;
        RECT 311.600 407.700 338.000 408.300 ;
        RECT 311.600 407.600 312.400 407.700 ;
        RECT 322.800 407.600 323.600 407.700 ;
        RECT 337.200 407.600 338.000 407.700 ;
        RECT 343.600 408.300 344.400 408.400 ;
        RECT 351.600 408.300 352.400 408.400 ;
        RECT 343.600 407.700 352.400 408.300 ;
        RECT 343.600 407.600 344.400 407.700 ;
        RECT 351.600 407.600 352.400 407.700 ;
        RECT 359.600 408.300 360.400 408.400 ;
        RECT 364.400 408.300 365.200 408.400 ;
        RECT 359.600 407.700 365.200 408.300 ;
        RECT 359.600 407.600 360.400 407.700 ;
        RECT 364.400 407.600 365.200 407.700 ;
        RECT 366.000 408.300 366.800 408.400 ;
        RECT 369.200 408.300 370.000 408.400 ;
        RECT 366.000 407.700 370.000 408.300 ;
        RECT 366.000 407.600 366.800 407.700 ;
        RECT 369.200 407.600 370.000 407.700 ;
        RECT 372.400 408.300 373.200 408.400 ;
        RECT 377.200 408.300 378.000 408.400 ;
        RECT 372.400 407.700 378.000 408.300 ;
        RECT 372.400 407.600 373.200 407.700 ;
        RECT 377.200 407.600 378.000 407.700 ;
        RECT 378.800 408.300 379.600 408.400 ;
        RECT 385.200 408.300 386.000 408.400 ;
        RECT 393.200 408.300 394.000 408.400 ;
        RECT 378.800 407.700 394.000 408.300 ;
        RECT 378.800 407.600 379.600 407.700 ;
        RECT 385.200 407.600 386.000 407.700 ;
        RECT 393.200 407.600 394.000 407.700 ;
        RECT 474.800 408.300 475.600 408.400 ;
        RECT 510.000 408.300 510.800 408.400 ;
        RECT 518.000 408.300 518.800 408.400 ;
        RECT 474.800 407.700 518.800 408.300 ;
        RECT 474.800 407.600 475.600 407.700 ;
        RECT 510.000 407.600 510.800 407.700 ;
        RECT 518.000 407.600 518.800 407.700 ;
        RECT 548.400 408.300 549.200 408.400 ;
        RECT 551.600 408.300 552.400 408.400 ;
        RECT 548.400 407.700 552.400 408.300 ;
        RECT 548.400 407.600 549.200 407.700 ;
        RECT 551.600 407.600 552.400 407.700 ;
        RECT 567.600 407.600 568.400 408.400 ;
        RECT 570.800 408.300 571.600 408.400 ;
        RECT 606.000 408.300 606.800 408.400 ;
        RECT 570.800 407.700 606.800 408.300 ;
        RECT 570.800 407.600 571.600 407.700 ;
        RECT 606.000 407.600 606.800 407.700 ;
        RECT 647.600 408.300 648.400 408.400 ;
        RECT 650.800 408.300 651.600 408.400 ;
        RECT 647.600 407.700 651.600 408.300 ;
        RECT 647.600 407.600 648.400 407.700 ;
        RECT 650.800 407.600 651.600 407.700 ;
        RECT 47.600 406.300 48.400 406.400 ;
        RECT 62.000 406.300 62.800 406.400 ;
        RECT 79.600 406.300 80.400 406.400 ;
        RECT 47.600 405.700 80.400 406.300 ;
        RECT 47.600 405.600 48.400 405.700 ;
        RECT 62.000 405.600 62.800 405.700 ;
        RECT 79.600 405.600 80.400 405.700 ;
        RECT 114.800 406.300 115.600 406.400 ;
        RECT 126.000 406.300 126.800 406.400 ;
        RECT 172.400 406.300 173.200 406.400 ;
        RECT 114.800 405.700 173.200 406.300 ;
        RECT 114.800 405.600 115.600 405.700 ;
        RECT 126.000 405.600 126.800 405.700 ;
        RECT 172.400 405.600 173.200 405.700 ;
        RECT 254.000 406.300 254.800 406.400 ;
        RECT 268.400 406.300 269.200 406.400 ;
        RECT 254.000 405.700 269.200 406.300 ;
        RECT 254.000 405.600 254.800 405.700 ;
        RECT 268.400 405.600 269.200 405.700 ;
        RECT 313.200 406.300 314.000 406.400 ;
        RECT 314.800 406.300 315.600 406.400 ;
        RECT 313.200 405.700 315.600 406.300 ;
        RECT 313.200 405.600 314.000 405.700 ;
        RECT 314.800 405.600 315.600 405.700 ;
        RECT 334.000 406.300 334.800 406.400 ;
        RECT 340.400 406.300 341.200 406.400 ;
        RECT 382.000 406.300 382.800 406.400 ;
        RECT 334.000 405.700 382.800 406.300 ;
        RECT 334.000 405.600 334.800 405.700 ;
        RECT 340.400 405.600 341.200 405.700 ;
        RECT 382.000 405.600 382.800 405.700 ;
        RECT 386.800 406.300 387.600 406.400 ;
        RECT 396.400 406.300 397.200 406.400 ;
        RECT 386.800 405.700 397.200 406.300 ;
        RECT 386.800 405.600 387.600 405.700 ;
        RECT 396.400 405.600 397.200 405.700 ;
        RECT 54.000 404.300 54.800 404.400 ;
        RECT 78.000 404.300 78.800 404.400 ;
        RECT 132.400 404.300 133.200 404.400 ;
        RECT 193.200 404.300 194.000 404.400 ;
        RECT 54.000 403.700 194.000 404.300 ;
        RECT 54.000 403.600 54.800 403.700 ;
        RECT 78.000 403.600 78.800 403.700 ;
        RECT 132.400 403.600 133.200 403.700 ;
        RECT 193.200 403.600 194.000 403.700 ;
        RECT 286.000 404.300 286.800 404.400 ;
        RECT 297.200 404.300 298.000 404.400 ;
        RECT 286.000 403.700 298.000 404.300 ;
        RECT 286.000 403.600 286.800 403.700 ;
        RECT 297.200 403.600 298.000 403.700 ;
        RECT 340.400 404.300 341.200 404.400 ;
        RECT 366.000 404.300 366.800 404.400 ;
        RECT 340.400 403.700 366.800 404.300 ;
        RECT 340.400 403.600 341.200 403.700 ;
        RECT 366.000 403.600 366.800 403.700 ;
        RECT 374.000 404.300 374.800 404.400 ;
        RECT 391.600 404.300 392.400 404.400 ;
        RECT 374.000 403.700 392.400 404.300 ;
        RECT 374.000 403.600 374.800 403.700 ;
        RECT 391.600 403.600 392.400 403.700 ;
        RECT 482.800 404.300 483.600 404.400 ;
        RECT 487.600 404.300 488.400 404.400 ;
        RECT 482.800 403.700 488.400 404.300 ;
        RECT 482.800 403.600 483.600 403.700 ;
        RECT 487.600 403.600 488.400 403.700 ;
        RECT 494.000 404.300 494.800 404.400 ;
        RECT 529.200 404.300 530.000 404.400 ;
        RECT 494.000 403.700 530.000 404.300 ;
        RECT 494.000 403.600 494.800 403.700 ;
        RECT 529.200 403.600 530.000 403.700 ;
        RECT 530.800 404.300 531.600 404.400 ;
        RECT 532.400 404.300 533.200 404.400 ;
        RECT 530.800 403.700 533.200 404.300 ;
        RECT 530.800 403.600 531.600 403.700 ;
        RECT 532.400 403.600 533.200 403.700 ;
        RECT 20.400 402.300 21.200 402.400 ;
        RECT 50.800 402.300 51.600 402.400 ;
        RECT 55.600 402.300 56.400 402.400 ;
        RECT 98.800 402.300 99.600 402.400 ;
        RECT 20.400 401.700 99.600 402.300 ;
        RECT 20.400 401.600 21.200 401.700 ;
        RECT 50.800 401.600 51.600 401.700 ;
        RECT 55.600 401.600 56.400 401.700 ;
        RECT 98.800 401.600 99.600 401.700 ;
        RECT 201.200 402.300 202.000 402.400 ;
        RECT 204.400 402.300 205.200 402.400 ;
        RECT 201.200 401.700 205.200 402.300 ;
        RECT 201.200 401.600 202.000 401.700 ;
        RECT 204.400 401.600 205.200 401.700 ;
        RECT 284.400 402.300 285.200 402.400 ;
        RECT 290.800 402.300 291.600 402.400 ;
        RECT 284.400 401.700 291.600 402.300 ;
        RECT 284.400 401.600 285.200 401.700 ;
        RECT 290.800 401.600 291.600 401.700 ;
        RECT 346.800 402.300 347.600 402.400 ;
        RECT 350.000 402.300 350.800 402.400 ;
        RECT 358.000 402.300 358.800 402.400 ;
        RECT 346.800 401.700 358.800 402.300 ;
        RECT 346.800 401.600 347.600 401.700 ;
        RECT 350.000 401.600 350.800 401.700 ;
        RECT 358.000 401.600 358.800 401.700 ;
        RECT 361.200 402.300 362.000 402.400 ;
        RECT 390.000 402.300 390.800 402.400 ;
        RECT 406.000 402.300 406.800 402.400 ;
        RECT 361.200 401.700 406.800 402.300 ;
        RECT 361.200 401.600 362.000 401.700 ;
        RECT 390.000 401.600 390.800 401.700 ;
        RECT 406.000 401.600 406.800 401.700 ;
        RECT 506.800 402.300 507.600 402.400 ;
        RECT 521.200 402.300 522.000 402.400 ;
        RECT 506.800 401.700 522.000 402.300 ;
        RECT 506.800 401.600 507.600 401.700 ;
        RECT 521.200 401.600 522.000 401.700 ;
        RECT 638.000 401.600 638.800 402.400 ;
        RECT 30.000 400.300 30.800 400.400 ;
        RECT 63.600 400.300 64.400 400.400 ;
        RECT 30.000 399.700 64.400 400.300 ;
        RECT 30.000 399.600 30.800 399.700 ;
        RECT 63.600 399.600 64.400 399.700 ;
        RECT 66.800 400.300 67.600 400.400 ;
        RECT 102.000 400.300 102.800 400.400 ;
        RECT 66.800 399.700 102.800 400.300 ;
        RECT 66.800 399.600 67.600 399.700 ;
        RECT 102.000 399.600 102.800 399.700 ;
        RECT 138.800 400.300 139.600 400.400 ;
        RECT 178.800 400.300 179.600 400.400 ;
        RECT 138.800 399.700 179.600 400.300 ;
        RECT 138.800 399.600 139.600 399.700 ;
        RECT 178.800 399.600 179.600 399.700 ;
        RECT 274.800 400.300 275.600 400.400 ;
        RECT 300.400 400.300 301.200 400.400 ;
        RECT 274.800 399.700 301.200 400.300 ;
        RECT 274.800 399.600 275.600 399.700 ;
        RECT 300.400 399.600 301.200 399.700 ;
        RECT 318.000 400.300 318.800 400.400 ;
        RECT 321.200 400.300 322.000 400.400 ;
        RECT 318.000 399.700 322.000 400.300 ;
        RECT 318.000 399.600 318.800 399.700 ;
        RECT 321.200 399.600 322.000 399.700 ;
        RECT 334.000 400.300 334.800 400.400 ;
        RECT 340.400 400.300 341.200 400.400 ;
        RECT 334.000 399.700 341.200 400.300 ;
        RECT 334.000 399.600 334.800 399.700 ;
        RECT 340.400 399.600 341.200 399.700 ;
        RECT 354.800 400.300 355.600 400.400 ;
        RECT 375.600 400.300 376.400 400.400 ;
        RECT 354.800 399.700 376.400 400.300 ;
        RECT 354.800 399.600 355.600 399.700 ;
        RECT 375.600 399.600 376.400 399.700 ;
        RECT 377.200 400.300 378.000 400.400 ;
        RECT 391.600 400.300 392.400 400.400 ;
        RECT 394.800 400.300 395.600 400.400 ;
        RECT 377.200 399.700 395.600 400.300 ;
        RECT 377.200 399.600 378.000 399.700 ;
        RECT 391.600 399.600 392.400 399.700 ;
        RECT 394.800 399.600 395.600 399.700 ;
        RECT 431.600 400.300 432.400 400.400 ;
        RECT 505.200 400.300 506.000 400.400 ;
        RECT 431.600 399.700 506.000 400.300 ;
        RECT 431.600 399.600 432.400 399.700 ;
        RECT 505.200 399.600 506.000 399.700 ;
        RECT 607.600 400.300 608.400 400.400 ;
        RECT 628.400 400.300 629.200 400.400 ;
        RECT 607.600 399.700 629.200 400.300 ;
        RECT 607.600 399.600 608.400 399.700 ;
        RECT 628.400 399.600 629.200 399.700 ;
        RECT 650.800 400.300 651.600 400.400 ;
        RECT 681.200 400.300 682.000 400.400 ;
        RECT 650.800 399.700 682.000 400.300 ;
        RECT 650.800 399.600 651.600 399.700 ;
        RECT 681.200 399.600 682.000 399.700 ;
        RECT 23.600 398.300 24.400 398.400 ;
        RECT 42.800 398.300 43.600 398.400 ;
        RECT 23.600 397.700 43.600 398.300 ;
        RECT 23.600 397.600 24.400 397.700 ;
        RECT 42.800 397.600 43.600 397.700 ;
        RECT 68.400 398.300 69.200 398.400 ;
        RECT 140.400 398.300 141.200 398.400 ;
        RECT 68.400 397.700 141.200 398.300 ;
        RECT 68.400 397.600 69.200 397.700 ;
        RECT 140.400 397.600 141.200 397.700 ;
        RECT 278.000 398.300 278.800 398.400 ;
        RECT 318.000 398.300 318.800 398.400 ;
        RECT 374.000 398.300 374.800 398.400 ;
        RECT 278.000 397.700 374.800 398.300 ;
        RECT 278.000 397.600 278.800 397.700 ;
        RECT 318.000 397.600 318.800 397.700 ;
        RECT 374.000 397.600 374.800 397.700 ;
        RECT 490.800 398.300 491.600 398.400 ;
        RECT 510.000 398.300 510.800 398.400 ;
        RECT 490.800 397.700 510.800 398.300 ;
        RECT 490.800 397.600 491.600 397.700 ;
        RECT 510.000 397.600 510.800 397.700 ;
        RECT 678.000 398.300 678.800 398.400 ;
        RECT 681.200 398.300 682.000 398.400 ;
        RECT 678.000 397.700 682.000 398.300 ;
        RECT 678.000 397.600 678.800 397.700 ;
        RECT 681.200 397.600 682.000 397.700 ;
        RECT 36.400 396.300 37.200 396.400 ;
        RECT 71.600 396.300 72.400 396.400 ;
        RECT 36.400 395.700 72.400 396.300 ;
        RECT 36.400 395.600 37.200 395.700 ;
        RECT 71.600 395.600 72.400 395.700 ;
        RECT 89.200 396.300 90.000 396.400 ;
        RECT 95.600 396.300 96.400 396.400 ;
        RECT 89.200 395.700 96.400 396.300 ;
        RECT 89.200 395.600 90.000 395.700 ;
        RECT 95.600 395.600 96.400 395.700 ;
        RECT 103.600 396.300 104.400 396.400 ;
        RECT 122.800 396.300 123.600 396.400 ;
        RECT 103.600 395.700 123.600 396.300 ;
        RECT 103.600 395.600 104.400 395.700 ;
        RECT 122.800 395.600 123.600 395.700 ;
        RECT 126.000 396.300 126.800 396.400 ;
        RECT 129.200 396.300 130.000 396.400 ;
        RECT 126.000 395.700 130.000 396.300 ;
        RECT 126.000 395.600 126.800 395.700 ;
        RECT 129.200 395.600 130.000 395.700 ;
        RECT 132.400 396.300 133.200 396.400 ;
        RECT 138.800 396.300 139.600 396.400 ;
        RECT 132.400 395.700 139.600 396.300 ;
        RECT 132.400 395.600 133.200 395.700 ;
        RECT 138.800 395.600 139.600 395.700 ;
        RECT 177.200 396.300 178.000 396.400 ;
        RECT 271.600 396.300 272.400 396.400 ;
        RECT 177.200 395.700 272.400 396.300 ;
        RECT 177.200 395.600 178.000 395.700 ;
        RECT 271.600 395.600 272.400 395.700 ;
        RECT 314.800 396.300 315.600 396.400 ;
        RECT 319.600 396.300 320.400 396.400 ;
        RECT 350.000 396.300 350.800 396.400 ;
        RECT 314.800 395.700 350.800 396.300 ;
        RECT 314.800 395.600 315.600 395.700 ;
        RECT 319.600 395.600 320.400 395.700 ;
        RECT 350.000 395.600 350.800 395.700 ;
        RECT 358.000 396.300 358.800 396.400 ;
        RECT 361.200 396.300 362.000 396.400 ;
        RECT 358.000 395.700 362.000 396.300 ;
        RECT 358.000 395.600 358.800 395.700 ;
        RECT 361.200 395.600 362.000 395.700 ;
        RECT 478.000 396.300 478.800 396.400 ;
        RECT 481.200 396.300 482.000 396.400 ;
        RECT 478.000 395.700 482.000 396.300 ;
        RECT 478.000 395.600 478.800 395.700 ;
        RECT 481.200 395.600 482.000 395.700 ;
        RECT 487.600 396.300 488.400 396.400 ;
        RECT 503.600 396.300 504.400 396.400 ;
        RECT 487.600 395.700 504.400 396.300 ;
        RECT 487.600 395.600 488.400 395.700 ;
        RECT 503.600 395.600 504.400 395.700 ;
        RECT 522.800 396.300 523.600 396.400 ;
        RECT 535.600 396.300 536.400 396.400 ;
        RECT 545.200 396.300 546.000 396.400 ;
        RECT 522.800 395.700 546.000 396.300 ;
        RECT 522.800 395.600 523.600 395.700 ;
        RECT 535.600 395.600 536.400 395.700 ;
        RECT 545.200 395.600 546.000 395.700 ;
        RECT 564.400 396.300 565.200 396.400 ;
        RECT 590.000 396.300 590.800 396.400 ;
        RECT 612.400 396.300 613.200 396.400 ;
        RECT 620.400 396.300 621.200 396.400 ;
        RECT 622.000 396.300 622.800 396.400 ;
        RECT 564.400 395.700 622.800 396.300 ;
        RECT 564.400 395.600 565.200 395.700 ;
        RECT 590.000 395.600 590.800 395.700 ;
        RECT 612.400 395.600 613.200 395.700 ;
        RECT 620.400 395.600 621.200 395.700 ;
        RECT 622.000 395.600 622.800 395.700 ;
        RECT 14.000 394.300 14.800 394.400 ;
        RECT 47.600 394.300 48.400 394.400 ;
        RECT 14.000 393.700 48.400 394.300 ;
        RECT 14.000 393.600 14.800 393.700 ;
        RECT 47.600 393.600 48.400 393.700 ;
        RECT 81.200 394.300 82.000 394.400 ;
        RECT 108.400 394.300 109.200 394.400 ;
        RECT 81.200 393.700 109.200 394.300 ;
        RECT 81.200 393.600 82.000 393.700 ;
        RECT 108.400 393.600 109.200 393.700 ;
        RECT 113.200 394.300 114.000 394.400 ;
        RECT 118.000 394.300 118.800 394.400 ;
        RECT 113.200 393.700 118.800 394.300 ;
        RECT 113.200 393.600 114.000 393.700 ;
        RECT 118.000 393.600 118.800 393.700 ;
        RECT 119.600 394.300 120.400 394.400 ;
        RECT 124.400 394.300 125.200 394.400 ;
        RECT 135.600 394.300 136.400 394.400 ;
        RECT 119.600 393.700 136.400 394.300 ;
        RECT 119.600 393.600 120.400 393.700 ;
        RECT 124.400 393.600 125.200 393.700 ;
        RECT 135.600 393.600 136.400 393.700 ;
        RECT 142.000 394.300 142.800 394.400 ;
        RECT 143.600 394.300 144.400 394.400 ;
        RECT 188.400 394.300 189.200 394.400 ;
        RECT 142.000 393.700 144.400 394.300 ;
        RECT 142.000 393.600 142.800 393.700 ;
        RECT 143.600 393.600 144.400 393.700 ;
        RECT 177.300 393.700 189.200 394.300 ;
        RECT 177.300 392.400 177.900 393.700 ;
        RECT 188.400 393.600 189.200 393.700 ;
        RECT 226.800 394.300 227.600 394.400 ;
        RECT 233.200 394.300 234.000 394.400 ;
        RECT 242.800 394.300 243.600 394.400 ;
        RECT 226.800 393.700 243.600 394.300 ;
        RECT 226.800 393.600 227.600 393.700 ;
        RECT 233.200 393.600 234.000 393.700 ;
        RECT 242.800 393.600 243.600 393.700 ;
        RECT 250.800 394.300 251.600 394.400 ;
        RECT 258.800 394.300 259.600 394.400 ;
        RECT 250.800 393.700 259.600 394.300 ;
        RECT 250.800 393.600 251.600 393.700 ;
        RECT 258.800 393.600 259.600 393.700 ;
        RECT 305.200 394.300 306.000 394.400 ;
        RECT 326.000 394.300 326.800 394.400 ;
        RECT 305.200 393.700 326.800 394.300 ;
        RECT 305.200 393.600 306.000 393.700 ;
        RECT 326.000 393.600 326.800 393.700 ;
        RECT 334.000 394.300 334.800 394.400 ;
        RECT 343.600 394.300 344.400 394.400 ;
        RECT 334.000 393.700 344.400 394.300 ;
        RECT 334.000 393.600 334.800 393.700 ;
        RECT 343.600 393.600 344.400 393.700 ;
        RECT 345.200 394.300 346.000 394.400 ;
        RECT 362.800 394.300 363.600 394.400 ;
        RECT 369.200 394.300 370.000 394.400 ;
        RECT 345.200 393.700 370.000 394.300 ;
        RECT 345.200 393.600 346.000 393.700 ;
        RECT 362.800 393.600 363.600 393.700 ;
        RECT 369.200 393.600 370.000 393.700 ;
        RECT 374.000 394.300 374.800 394.400 ;
        RECT 417.200 394.300 418.000 394.400 ;
        RECT 374.000 393.700 418.000 394.300 ;
        RECT 374.000 393.600 374.800 393.700 ;
        RECT 417.200 393.600 418.000 393.700 ;
        RECT 486.000 394.300 486.800 394.400 ;
        RECT 498.800 394.300 499.600 394.400 ;
        RECT 514.800 394.300 515.600 394.400 ;
        RECT 486.000 393.700 515.600 394.300 ;
        RECT 486.000 393.600 486.800 393.700 ;
        RECT 498.800 393.600 499.600 393.700 ;
        RECT 514.800 393.600 515.600 393.700 ;
        RECT 519.600 394.300 520.400 394.400 ;
        RECT 546.800 394.300 547.600 394.400 ;
        RECT 519.600 393.700 547.600 394.300 ;
        RECT 519.600 393.600 520.400 393.700 ;
        RECT 546.800 393.600 547.600 393.700 ;
        RECT 569.200 394.300 570.000 394.400 ;
        RECT 604.400 394.300 605.200 394.400 ;
        RECT 569.200 393.700 605.200 394.300 ;
        RECT 569.200 393.600 570.000 393.700 ;
        RECT 604.400 393.600 605.200 393.700 ;
        RECT 609.200 394.300 610.000 394.400 ;
        RECT 654.000 394.300 654.800 394.400 ;
        RECT 609.200 393.700 654.800 394.300 ;
        RECT 609.200 393.600 610.000 393.700 ;
        RECT 654.000 393.600 654.800 393.700 ;
        RECT 20.400 392.300 21.200 392.400 ;
        RECT 25.200 392.300 26.000 392.400 ;
        RECT 20.400 391.700 26.000 392.300 ;
        RECT 20.400 391.600 21.200 391.700 ;
        RECT 25.200 391.600 26.000 391.700 ;
        RECT 42.800 392.300 43.600 392.400 ;
        RECT 49.200 392.300 50.000 392.400 ;
        RECT 42.800 391.700 50.000 392.300 ;
        RECT 42.800 391.600 43.600 391.700 ;
        RECT 49.200 391.600 50.000 391.700 ;
        RECT 78.000 392.300 78.800 392.400 ;
        RECT 84.400 392.300 85.200 392.400 ;
        RECT 78.000 391.700 85.200 392.300 ;
        RECT 78.000 391.600 78.800 391.700 ;
        RECT 84.400 391.600 85.200 391.700 ;
        RECT 103.600 392.300 104.400 392.400 ;
        RECT 121.200 392.300 122.000 392.400 ;
        RECT 103.600 391.700 122.000 392.300 ;
        RECT 103.600 391.600 104.400 391.700 ;
        RECT 121.200 391.600 122.000 391.700 ;
        RECT 129.200 392.300 130.000 392.400 ;
        RECT 143.600 392.300 144.400 392.400 ;
        RECT 129.200 391.700 144.400 392.300 ;
        RECT 129.200 391.600 130.000 391.700 ;
        RECT 143.600 391.600 144.400 391.700 ;
        RECT 158.000 392.300 158.800 392.400 ;
        RECT 172.400 392.300 173.200 392.400 ;
        RECT 158.000 391.700 173.200 392.300 ;
        RECT 158.000 391.600 158.800 391.700 ;
        RECT 172.400 391.600 173.200 391.700 ;
        RECT 175.600 392.300 176.400 392.400 ;
        RECT 177.200 392.300 178.000 392.400 ;
        RECT 175.600 391.700 178.000 392.300 ;
        RECT 175.600 391.600 176.400 391.700 ;
        RECT 177.200 391.600 178.000 391.700 ;
        RECT 186.800 392.300 187.600 392.400 ;
        RECT 193.200 392.300 194.000 392.400 ;
        RECT 201.200 392.300 202.000 392.400 ;
        RECT 186.800 391.700 202.000 392.300 ;
        RECT 186.800 391.600 187.600 391.700 ;
        RECT 193.200 391.600 194.000 391.700 ;
        RECT 201.200 391.600 202.000 391.700 ;
        RECT 220.400 392.300 221.200 392.400 ;
        RECT 234.800 392.300 235.600 392.400 ;
        RECT 238.000 392.300 238.800 392.400 ;
        RECT 220.400 391.700 238.800 392.300 ;
        RECT 220.400 391.600 221.200 391.700 ;
        RECT 234.800 391.600 235.600 391.700 ;
        RECT 238.000 391.600 238.800 391.700 ;
        RECT 314.800 392.300 315.600 392.400 ;
        RECT 337.200 392.300 338.000 392.400 ;
        RECT 314.800 391.700 338.000 392.300 ;
        RECT 314.800 391.600 315.600 391.700 ;
        RECT 337.200 391.600 338.000 391.700 ;
        RECT 343.600 392.300 344.400 392.400 ;
        RECT 362.800 392.300 363.600 392.400 ;
        RECT 343.600 391.700 363.600 392.300 ;
        RECT 343.600 391.600 344.400 391.700 ;
        RECT 362.800 391.600 363.600 391.700 ;
        RECT 366.000 392.300 366.800 392.400 ;
        RECT 375.600 392.300 376.400 392.400 ;
        RECT 386.800 392.300 387.600 392.400 ;
        RECT 366.000 391.700 387.600 392.300 ;
        RECT 366.000 391.600 366.800 391.700 ;
        RECT 375.600 391.600 376.400 391.700 ;
        RECT 386.800 391.600 387.600 391.700 ;
        RECT 492.400 392.300 493.200 392.400 ;
        RECT 506.800 392.300 507.600 392.400 ;
        RECT 492.400 391.700 507.600 392.300 ;
        RECT 492.400 391.600 493.200 391.700 ;
        RECT 506.800 391.600 507.600 391.700 ;
        RECT 545.200 392.300 546.000 392.400 ;
        RECT 554.800 392.300 555.600 392.400 ;
        RECT 545.200 391.700 555.600 392.300 ;
        RECT 545.200 391.600 546.000 391.700 ;
        RECT 554.800 391.600 555.600 391.700 ;
        RECT 562.800 392.300 563.600 392.400 ;
        RECT 618.800 392.300 619.600 392.400 ;
        RECT 678.000 392.300 678.800 392.400 ;
        RECT 562.800 391.700 678.800 392.300 ;
        RECT 562.800 391.600 563.600 391.700 ;
        RECT 618.800 391.600 619.600 391.700 ;
        RECT 678.000 391.600 678.800 391.700 ;
        RECT 25.200 390.300 26.000 390.400 ;
        RECT 33.200 390.300 34.000 390.400 ;
        RECT 39.600 390.300 40.400 390.400 ;
        RECT 25.200 389.700 40.400 390.300 ;
        RECT 25.200 389.600 26.000 389.700 ;
        RECT 33.200 389.600 34.000 389.700 ;
        RECT 39.600 389.600 40.400 389.700 ;
        RECT 47.600 390.300 48.400 390.400 ;
        RECT 52.400 390.300 53.200 390.400 ;
        RECT 47.600 389.700 53.200 390.300 ;
        RECT 47.600 389.600 48.400 389.700 ;
        RECT 52.400 389.600 53.200 389.700 ;
        RECT 58.800 389.600 59.600 390.400 ;
        RECT 82.800 390.300 83.600 390.400 ;
        RECT 108.400 390.300 109.200 390.400 ;
        RECT 82.800 389.700 109.200 390.300 ;
        RECT 82.800 389.600 83.600 389.700 ;
        RECT 108.400 389.600 109.200 389.700 ;
        RECT 118.000 390.300 118.800 390.400 ;
        RECT 127.600 390.300 128.400 390.400 ;
        RECT 134.000 390.300 134.800 390.400 ;
        RECT 118.000 389.700 134.800 390.300 ;
        RECT 118.000 389.600 118.800 389.700 ;
        RECT 127.600 389.600 128.400 389.700 ;
        RECT 134.000 389.600 134.800 389.700 ;
        RECT 140.400 390.300 141.200 390.400 ;
        RECT 148.400 390.300 149.200 390.400 ;
        RECT 140.400 389.700 149.200 390.300 ;
        RECT 140.400 389.600 141.200 389.700 ;
        RECT 148.400 389.600 149.200 389.700 ;
        RECT 194.800 390.300 195.600 390.400 ;
        RECT 199.600 390.300 200.400 390.400 ;
        RECT 194.800 389.700 200.400 390.300 ;
        RECT 194.800 389.600 195.600 389.700 ;
        RECT 199.600 389.600 200.400 389.700 ;
        RECT 202.800 390.300 203.600 390.400 ;
        RECT 276.400 390.300 277.200 390.400 ;
        RECT 202.800 389.700 277.200 390.300 ;
        RECT 202.800 389.600 203.600 389.700 ;
        RECT 276.400 389.600 277.200 389.700 ;
        RECT 303.600 390.300 304.400 390.400 ;
        RECT 388.400 390.300 389.200 390.400 ;
        RECT 303.600 389.700 389.200 390.300 ;
        RECT 303.600 389.600 304.400 389.700 ;
        RECT 388.400 389.600 389.200 389.700 ;
        RECT 439.600 390.300 440.400 390.400 ;
        RECT 449.200 390.300 450.000 390.400 ;
        RECT 439.600 389.700 450.000 390.300 ;
        RECT 439.600 389.600 440.400 389.700 ;
        RECT 449.200 389.600 450.000 389.700 ;
        RECT 486.000 390.300 486.800 390.400 ;
        RECT 506.800 390.300 507.600 390.400 ;
        RECT 486.000 389.700 507.600 390.300 ;
        RECT 486.000 389.600 486.800 389.700 ;
        RECT 506.800 389.600 507.600 389.700 ;
        RECT 508.400 390.300 509.200 390.400 ;
        RECT 514.800 390.300 515.600 390.400 ;
        RECT 521.200 390.300 522.000 390.400 ;
        RECT 508.400 389.700 522.000 390.300 ;
        RECT 508.400 389.600 509.200 389.700 ;
        RECT 514.800 389.600 515.600 389.700 ;
        RECT 521.200 389.600 522.000 389.700 ;
        RECT 527.600 390.300 528.400 390.400 ;
        RECT 591.600 390.300 592.400 390.400 ;
        RECT 527.600 389.700 592.400 390.300 ;
        RECT 527.600 389.600 528.400 389.700 ;
        RECT 591.600 389.600 592.400 389.700 ;
        RECT 610.800 390.300 611.600 390.400 ;
        RECT 623.600 390.300 624.400 390.400 ;
        RECT 610.800 389.700 624.400 390.300 ;
        RECT 610.800 389.600 611.600 389.700 ;
        RECT 623.600 389.600 624.400 389.700 ;
        RECT 641.200 390.300 642.000 390.400 ;
        RECT 646.000 390.300 646.800 390.400 ;
        RECT 641.200 389.700 646.800 390.300 ;
        RECT 641.200 389.600 642.000 389.700 ;
        RECT 646.000 389.600 646.800 389.700 ;
        RECT 30.000 388.300 30.800 388.400 ;
        RECT 38.000 388.300 38.800 388.400 ;
        RECT 30.000 387.700 38.800 388.300 ;
        RECT 30.000 387.600 30.800 387.700 ;
        RECT 38.000 387.600 38.800 387.700 ;
        RECT 57.200 388.300 58.000 388.400 ;
        RECT 60.400 388.300 61.200 388.400 ;
        RECT 57.200 387.700 61.200 388.300 ;
        RECT 57.200 387.600 58.000 387.700 ;
        RECT 60.400 387.600 61.200 387.700 ;
        RECT 65.200 388.300 66.000 388.400 ;
        RECT 70.000 388.300 70.800 388.400 ;
        RECT 65.200 387.700 70.800 388.300 ;
        RECT 65.200 387.600 66.000 387.700 ;
        RECT 70.000 387.600 70.800 387.700 ;
        RECT 87.600 388.300 88.400 388.400 ;
        RECT 119.600 388.300 120.400 388.400 ;
        RECT 87.600 387.700 120.400 388.300 ;
        RECT 87.600 387.600 88.400 387.700 ;
        RECT 119.600 387.600 120.400 387.700 ;
        RECT 127.600 388.300 128.400 388.400 ;
        RECT 138.800 388.300 139.600 388.400 ;
        RECT 145.200 388.300 146.000 388.400 ;
        RECT 127.600 387.700 146.000 388.300 ;
        RECT 127.600 387.600 128.400 387.700 ;
        RECT 138.800 387.600 139.600 387.700 ;
        RECT 145.200 387.600 146.000 387.700 ;
        RECT 148.400 388.300 149.200 388.400 ;
        RECT 167.600 388.300 168.400 388.400 ;
        RECT 148.400 387.700 168.400 388.300 ;
        RECT 148.400 387.600 149.200 387.700 ;
        RECT 167.600 387.600 168.400 387.700 ;
        RECT 177.200 388.300 178.000 388.400 ;
        RECT 188.400 388.300 189.200 388.400 ;
        RECT 177.200 387.700 189.200 388.300 ;
        RECT 177.200 387.600 178.000 387.700 ;
        RECT 188.400 387.600 189.200 387.700 ;
        RECT 199.600 388.300 200.400 388.400 ;
        RECT 210.800 388.300 211.600 388.400 ;
        RECT 199.600 387.700 211.600 388.300 ;
        RECT 199.600 387.600 200.400 387.700 ;
        RECT 210.800 387.600 211.600 387.700 ;
        RECT 239.600 388.300 240.400 388.400 ;
        RECT 247.600 388.300 248.400 388.400 ;
        RECT 239.600 387.700 248.400 388.300 ;
        RECT 239.600 387.600 240.400 387.700 ;
        RECT 247.600 387.600 248.400 387.700 ;
        RECT 292.400 388.300 293.200 388.400 ;
        RECT 302.000 388.300 302.800 388.400 ;
        RECT 313.200 388.300 314.000 388.400 ;
        RECT 292.400 387.700 314.000 388.300 ;
        RECT 292.400 387.600 293.200 387.700 ;
        RECT 302.000 387.600 302.800 387.700 ;
        RECT 313.200 387.600 314.000 387.700 ;
        RECT 329.200 388.300 330.000 388.400 ;
        RECT 359.600 388.300 360.400 388.400 ;
        RECT 372.400 388.300 373.200 388.400 ;
        RECT 329.200 387.700 373.200 388.300 ;
        RECT 329.200 387.600 330.000 387.700 ;
        RECT 359.600 387.600 360.400 387.700 ;
        RECT 372.400 387.600 373.200 387.700 ;
        RECT 383.600 388.300 384.400 388.400 ;
        RECT 428.400 388.300 429.200 388.400 ;
        RECT 383.600 387.700 429.200 388.300 ;
        RECT 383.600 387.600 384.400 387.700 ;
        RECT 428.400 387.600 429.200 387.700 ;
        RECT 430.000 388.300 430.800 388.400 ;
        RECT 436.400 388.300 437.200 388.400 ;
        RECT 441.200 388.300 442.000 388.400 ;
        RECT 430.000 387.700 442.000 388.300 ;
        RECT 430.000 387.600 430.800 387.700 ;
        RECT 436.400 387.600 437.200 387.700 ;
        RECT 441.200 387.600 442.000 387.700 ;
        RECT 447.600 388.300 448.400 388.400 ;
        RECT 482.800 388.300 483.600 388.400 ;
        RECT 447.600 387.700 483.600 388.300 ;
        RECT 447.600 387.600 448.400 387.700 ;
        RECT 482.800 387.600 483.600 387.700 ;
        RECT 484.400 388.300 485.200 388.400 ;
        RECT 490.800 388.300 491.600 388.400 ;
        RECT 503.600 388.300 504.400 388.400 ;
        RECT 484.400 387.700 504.400 388.300 ;
        RECT 484.400 387.600 485.200 387.700 ;
        RECT 490.800 387.600 491.600 387.700 ;
        RECT 503.600 387.600 504.400 387.700 ;
        RECT 505.200 388.300 506.000 388.400 ;
        RECT 510.000 388.300 510.800 388.400 ;
        RECT 516.400 388.300 517.200 388.400 ;
        RECT 522.800 388.300 523.600 388.400 ;
        RECT 505.200 387.700 523.600 388.300 ;
        RECT 505.200 387.600 506.000 387.700 ;
        RECT 510.000 387.600 510.800 387.700 ;
        RECT 516.400 387.600 517.200 387.700 ;
        RECT 522.800 387.600 523.600 387.700 ;
        RECT 534.000 388.300 534.800 388.400 ;
        RECT 578.800 388.300 579.600 388.400 ;
        RECT 614.000 388.300 614.800 388.400 ;
        RECT 534.000 387.700 614.800 388.300 ;
        RECT 534.000 387.600 534.800 387.700 ;
        RECT 578.800 387.600 579.600 387.700 ;
        RECT 614.000 387.600 614.800 387.700 ;
        RECT 618.800 388.300 619.600 388.400 ;
        RECT 662.000 388.300 662.800 388.400 ;
        RECT 618.800 387.700 662.800 388.300 ;
        RECT 618.800 387.600 619.600 387.700 ;
        RECT 662.000 387.600 662.800 387.700 ;
        RECT 33.200 386.300 34.000 386.400 ;
        RECT 66.800 386.300 67.600 386.400 ;
        RECT 33.200 385.700 67.600 386.300 ;
        RECT 33.200 385.600 34.000 385.700 ;
        RECT 66.800 385.600 67.600 385.700 ;
        RECT 97.200 386.300 98.000 386.400 ;
        RECT 129.200 386.300 130.000 386.400 ;
        RECT 97.200 385.700 130.000 386.300 ;
        RECT 97.200 385.600 98.000 385.700 ;
        RECT 129.200 385.600 130.000 385.700 ;
        RECT 142.000 386.300 142.800 386.400 ;
        RECT 143.600 386.300 144.400 386.400 ;
        RECT 142.000 385.700 144.400 386.300 ;
        RECT 142.000 385.600 142.800 385.700 ;
        RECT 143.600 385.600 144.400 385.700 ;
        RECT 150.000 386.300 150.800 386.400 ;
        RECT 151.600 386.300 152.400 386.400 ;
        RECT 150.000 385.700 152.400 386.300 ;
        RECT 150.000 385.600 150.800 385.700 ;
        RECT 151.600 385.600 152.400 385.700 ;
        RECT 186.800 386.300 187.600 386.400 ;
        RECT 196.400 386.300 197.200 386.400 ;
        RECT 186.800 385.700 197.200 386.300 ;
        RECT 186.800 385.600 187.600 385.700 ;
        RECT 196.400 385.600 197.200 385.700 ;
        RECT 241.200 386.300 242.000 386.400 ;
        RECT 252.400 386.300 253.200 386.400 ;
        RECT 241.200 385.700 253.200 386.300 ;
        RECT 241.200 385.600 242.000 385.700 ;
        RECT 252.400 385.600 253.200 385.700 ;
        RECT 324.400 386.300 325.200 386.400 ;
        RECT 335.600 386.300 336.400 386.400 ;
        RECT 324.400 385.700 336.400 386.300 ;
        RECT 324.400 385.600 325.200 385.700 ;
        RECT 335.600 385.600 336.400 385.700 ;
        RECT 343.600 386.300 344.400 386.400 ;
        RECT 346.800 386.300 347.600 386.400 ;
        RECT 359.600 386.300 360.400 386.400 ;
        RECT 343.600 385.700 360.400 386.300 ;
        RECT 343.600 385.600 344.400 385.700 ;
        RECT 346.800 385.600 347.600 385.700 ;
        RECT 359.600 385.600 360.400 385.700 ;
        RECT 478.000 386.300 478.800 386.400 ;
        RECT 494.000 386.300 494.800 386.400 ;
        RECT 478.000 385.700 494.800 386.300 ;
        RECT 478.000 385.600 478.800 385.700 ;
        RECT 494.000 385.600 494.800 385.700 ;
        RECT 516.400 386.300 517.200 386.400 ;
        RECT 519.600 386.300 520.400 386.400 ;
        RECT 516.400 385.700 520.400 386.300 ;
        RECT 516.400 385.600 517.200 385.700 ;
        RECT 519.600 385.600 520.400 385.700 ;
        RECT 521.200 386.300 522.000 386.400 ;
        RECT 535.600 386.300 536.400 386.400 ;
        RECT 521.200 385.700 536.400 386.300 ;
        RECT 521.200 385.600 522.000 385.700 ;
        RECT 535.600 385.600 536.400 385.700 ;
        RECT 556.400 386.300 557.200 386.400 ;
        RECT 588.400 386.300 589.200 386.400 ;
        RECT 556.400 385.700 589.200 386.300 ;
        RECT 556.400 385.600 557.200 385.700 ;
        RECT 588.400 385.600 589.200 385.700 ;
        RECT 609.200 386.300 610.000 386.400 ;
        RECT 610.800 386.300 611.600 386.400 ;
        RECT 626.800 386.300 627.600 386.400 ;
        RECT 609.200 385.700 627.600 386.300 ;
        RECT 609.200 385.600 610.000 385.700 ;
        RECT 610.800 385.600 611.600 385.700 ;
        RECT 626.800 385.600 627.600 385.700 ;
        RECT 634.800 386.300 635.600 386.400 ;
        RECT 647.600 386.300 648.400 386.400 ;
        RECT 634.800 385.700 648.400 386.300 ;
        RECT 634.800 385.600 635.600 385.700 ;
        RECT 647.600 385.600 648.400 385.700 ;
        RECT 49.200 384.300 50.000 384.400 ;
        RECT 79.600 384.300 80.400 384.400 ;
        RECT 49.200 383.700 80.400 384.300 ;
        RECT 49.200 383.600 50.000 383.700 ;
        RECT 79.600 383.600 80.400 383.700 ;
        RECT 116.400 384.300 117.200 384.400 ;
        RECT 127.600 384.300 128.400 384.400 ;
        RECT 116.400 383.700 128.400 384.300 ;
        RECT 116.400 383.600 117.200 383.700 ;
        RECT 127.600 383.600 128.400 383.700 ;
        RECT 129.200 384.300 130.000 384.400 ;
        RECT 166.000 384.300 166.800 384.400 ;
        RECT 190.000 384.300 190.800 384.400 ;
        RECT 194.800 384.300 195.600 384.400 ;
        RECT 217.200 384.300 218.000 384.400 ;
        RECT 231.600 384.300 232.400 384.400 ;
        RECT 236.400 384.300 237.200 384.400 ;
        RECT 129.200 383.700 237.200 384.300 ;
        RECT 129.200 383.600 130.000 383.700 ;
        RECT 166.000 383.600 166.800 383.700 ;
        RECT 190.000 383.600 190.800 383.700 ;
        RECT 194.800 383.600 195.600 383.700 ;
        RECT 217.200 383.600 218.000 383.700 ;
        RECT 231.600 383.600 232.400 383.700 ;
        RECT 236.400 383.600 237.200 383.700 ;
        RECT 254.000 384.300 254.800 384.400 ;
        RECT 292.400 384.300 293.200 384.400 ;
        RECT 295.600 384.300 296.400 384.400 ;
        RECT 254.000 383.700 296.400 384.300 ;
        RECT 254.000 383.600 254.800 383.700 ;
        RECT 292.400 383.600 293.200 383.700 ;
        RECT 295.600 383.600 296.400 383.700 ;
        RECT 303.600 384.300 304.400 384.400 ;
        RECT 308.400 384.300 309.200 384.400 ;
        RECT 311.600 384.300 312.400 384.400 ;
        RECT 303.600 383.700 312.400 384.300 ;
        RECT 303.600 383.600 304.400 383.700 ;
        RECT 308.400 383.600 309.200 383.700 ;
        RECT 311.600 383.600 312.400 383.700 ;
        RECT 313.200 384.300 314.000 384.400 ;
        RECT 398.000 384.300 398.800 384.400 ;
        RECT 313.200 383.700 398.800 384.300 ;
        RECT 313.200 383.600 314.000 383.700 ;
        RECT 398.000 383.600 398.800 383.700 ;
        RECT 468.400 384.300 469.200 384.400 ;
        RECT 484.400 384.300 485.200 384.400 ;
        RECT 468.400 383.700 485.200 384.300 ;
        RECT 468.400 383.600 469.200 383.700 ;
        RECT 484.400 383.600 485.200 383.700 ;
        RECT 494.000 384.300 494.800 384.400 ;
        RECT 530.800 384.300 531.600 384.400 ;
        RECT 494.000 383.700 531.600 384.300 ;
        RECT 494.000 383.600 494.800 383.700 ;
        RECT 530.800 383.600 531.600 383.700 ;
        RECT 561.200 384.300 562.000 384.400 ;
        RECT 570.800 384.300 571.600 384.400 ;
        RECT 561.200 383.700 571.600 384.300 ;
        RECT 561.200 383.600 562.000 383.700 ;
        RECT 570.800 383.600 571.600 383.700 ;
        RECT 583.600 384.300 584.400 384.400 ;
        RECT 586.800 384.300 587.600 384.400 ;
        RECT 615.600 384.300 616.400 384.400 ;
        RECT 583.600 383.700 616.400 384.300 ;
        RECT 583.600 383.600 584.400 383.700 ;
        RECT 586.800 383.600 587.600 383.700 ;
        RECT 615.600 383.600 616.400 383.700 ;
        RECT 23.600 382.300 24.400 382.400 ;
        RECT 30.000 382.300 30.800 382.400 ;
        RECT 74.800 382.300 75.600 382.400 ;
        RECT 23.600 381.700 75.600 382.300 ;
        RECT 23.600 381.600 24.400 381.700 ;
        RECT 30.000 381.600 30.800 381.700 ;
        RECT 74.800 381.600 75.600 381.700 ;
        RECT 114.800 382.300 115.600 382.400 ;
        RECT 135.600 382.300 136.400 382.400 ;
        RECT 151.600 382.300 152.400 382.400 ;
        RECT 114.800 381.700 152.400 382.300 ;
        RECT 114.800 381.600 115.600 381.700 ;
        RECT 135.600 381.600 136.400 381.700 ;
        RECT 151.600 381.600 152.400 381.700 ;
        RECT 162.800 382.300 163.600 382.400 ;
        RECT 166.000 382.300 166.800 382.400 ;
        RECT 180.400 382.300 181.200 382.400 ;
        RECT 162.800 381.700 181.200 382.300 ;
        RECT 162.800 381.600 163.600 381.700 ;
        RECT 166.000 381.600 166.800 381.700 ;
        RECT 180.400 381.600 181.200 381.700 ;
        RECT 228.400 382.300 229.200 382.400 ;
        RECT 241.200 382.300 242.000 382.400 ;
        RECT 228.400 381.700 242.000 382.300 ;
        RECT 228.400 381.600 229.200 381.700 ;
        RECT 241.200 381.600 242.000 381.700 ;
        RECT 290.800 382.300 291.600 382.400 ;
        RECT 295.600 382.300 296.400 382.400 ;
        RECT 290.800 381.700 296.400 382.300 ;
        RECT 290.800 381.600 291.600 381.700 ;
        RECT 295.600 381.600 296.400 381.700 ;
        RECT 318.000 382.300 318.800 382.400 ;
        RECT 337.200 382.300 338.000 382.400 ;
        RECT 318.000 381.700 338.000 382.300 ;
        RECT 318.000 381.600 318.800 381.700 ;
        RECT 337.200 381.600 338.000 381.700 ;
        RECT 342.000 382.300 342.800 382.400 ;
        RECT 351.600 382.300 352.400 382.400 ;
        RECT 362.800 382.300 363.600 382.400 ;
        RECT 342.000 381.700 363.600 382.300 ;
        RECT 342.000 381.600 342.800 381.700 ;
        RECT 351.600 381.600 352.400 381.700 ;
        RECT 362.800 381.600 363.600 381.700 ;
        RECT 398.000 382.300 398.800 382.400 ;
        RECT 399.600 382.300 400.400 382.400 ;
        RECT 398.000 381.700 400.400 382.300 ;
        RECT 398.000 381.600 398.800 381.700 ;
        RECT 399.600 381.600 400.400 381.700 ;
        RECT 407.600 382.300 408.400 382.400 ;
        RECT 425.200 382.300 426.000 382.400 ;
        RECT 407.600 381.700 426.000 382.300 ;
        RECT 407.600 381.600 408.400 381.700 ;
        RECT 425.200 381.600 426.000 381.700 ;
        RECT 463.600 382.300 464.400 382.400 ;
        RECT 489.200 382.300 490.000 382.400 ;
        RECT 463.600 381.700 490.000 382.300 ;
        RECT 463.600 381.600 464.400 381.700 ;
        RECT 489.200 381.600 490.000 381.700 ;
        RECT 503.600 382.300 504.400 382.400 ;
        RECT 511.600 382.300 512.400 382.400 ;
        RECT 503.600 381.700 512.400 382.300 ;
        RECT 503.600 381.600 504.400 381.700 ;
        RECT 511.600 381.600 512.400 381.700 ;
        RECT 518.000 382.300 518.800 382.400 ;
        RECT 540.400 382.300 541.200 382.400 ;
        RECT 564.400 382.300 565.200 382.400 ;
        RECT 567.600 382.300 568.400 382.400 ;
        RECT 518.000 381.700 568.400 382.300 ;
        RECT 518.000 381.600 518.800 381.700 ;
        RECT 540.400 381.600 541.200 381.700 ;
        RECT 564.400 381.600 565.200 381.700 ;
        RECT 567.600 381.600 568.400 381.700 ;
        RECT 585.200 382.300 586.000 382.400 ;
        RECT 604.400 382.300 605.200 382.400 ;
        RECT 585.200 381.700 605.200 382.300 ;
        RECT 585.200 381.600 586.000 381.700 ;
        RECT 604.400 381.600 605.200 381.700 ;
        RECT 22.000 380.300 22.800 380.400 ;
        RECT 95.600 380.300 96.400 380.400 ;
        RECT 22.000 379.700 96.400 380.300 ;
        RECT 22.000 379.600 22.800 379.700 ;
        RECT 95.600 379.600 96.400 379.700 ;
        RECT 145.200 380.300 146.000 380.400 ;
        RECT 150.000 380.300 150.800 380.400 ;
        RECT 158.000 380.300 158.800 380.400 ;
        RECT 145.200 379.700 158.800 380.300 ;
        RECT 145.200 379.600 146.000 379.700 ;
        RECT 150.000 379.600 150.800 379.700 ;
        RECT 158.000 379.600 158.800 379.700 ;
        RECT 169.200 380.300 170.000 380.400 ;
        RECT 212.400 380.300 213.200 380.400 ;
        RECT 250.800 380.300 251.600 380.400 ;
        RECT 169.200 379.700 251.600 380.300 ;
        RECT 169.200 379.600 170.000 379.700 ;
        RECT 212.400 379.600 213.200 379.700 ;
        RECT 250.800 379.600 251.600 379.700 ;
        RECT 319.600 380.300 320.400 380.400 ;
        RECT 324.400 380.300 325.200 380.400 ;
        RECT 319.600 379.700 325.200 380.300 ;
        RECT 319.600 379.600 320.400 379.700 ;
        RECT 324.400 379.600 325.200 379.700 ;
        RECT 358.000 380.300 358.800 380.400 ;
        RECT 362.800 380.300 363.600 380.400 ;
        RECT 358.000 379.700 363.600 380.300 ;
        RECT 358.000 379.600 358.800 379.700 ;
        RECT 362.800 379.600 363.600 379.700 ;
        RECT 366.000 380.300 366.800 380.400 ;
        RECT 367.600 380.300 368.400 380.400 ;
        RECT 366.000 379.700 368.400 380.300 ;
        RECT 366.000 379.600 366.800 379.700 ;
        RECT 367.600 379.600 368.400 379.700 ;
        RECT 426.800 380.300 427.600 380.400 ;
        RECT 490.800 380.300 491.600 380.400 ;
        RECT 426.800 379.700 491.600 380.300 ;
        RECT 426.800 379.600 427.600 379.700 ;
        RECT 490.800 379.600 491.600 379.700 ;
        RECT 522.800 380.300 523.600 380.400 ;
        RECT 537.200 380.300 538.000 380.400 ;
        RECT 522.800 379.700 538.000 380.300 ;
        RECT 522.800 379.600 523.600 379.700 ;
        RECT 537.200 379.600 538.000 379.700 ;
        RECT 639.600 380.300 640.400 380.400 ;
        RECT 670.000 380.300 670.800 380.400 ;
        RECT 639.600 379.700 670.800 380.300 ;
        RECT 639.600 379.600 640.400 379.700 ;
        RECT 670.000 379.600 670.800 379.700 ;
        RECT 36.400 378.300 37.200 378.400 ;
        RECT 47.600 378.300 48.400 378.400 ;
        RECT 36.400 377.700 48.400 378.300 ;
        RECT 36.400 377.600 37.200 377.700 ;
        RECT 47.600 377.600 48.400 377.700 ;
        RECT 54.000 378.300 54.800 378.400 ;
        RECT 65.200 378.300 66.000 378.400 ;
        RECT 54.000 377.700 66.000 378.300 ;
        RECT 54.000 377.600 54.800 377.700 ;
        RECT 65.200 377.600 66.000 377.700 ;
        RECT 148.400 378.300 149.200 378.400 ;
        RECT 185.200 378.300 186.000 378.400 ;
        RECT 148.400 377.700 186.000 378.300 ;
        RECT 148.400 377.600 149.200 377.700 ;
        RECT 185.200 377.600 186.000 377.700 ;
        RECT 186.800 378.300 187.600 378.400 ;
        RECT 196.400 378.300 197.200 378.400 ;
        RECT 254.000 378.300 254.800 378.400 ;
        RECT 186.800 377.700 254.800 378.300 ;
        RECT 186.800 377.600 187.600 377.700 ;
        RECT 196.400 377.600 197.200 377.700 ;
        RECT 254.000 377.600 254.800 377.700 ;
        RECT 321.200 378.300 322.000 378.400 ;
        RECT 332.400 378.300 333.200 378.400 ;
        RECT 321.200 377.700 333.200 378.300 ;
        RECT 321.200 377.600 322.000 377.700 ;
        RECT 332.400 377.600 333.200 377.700 ;
        RECT 338.800 378.300 339.600 378.400 ;
        RECT 346.800 378.300 347.600 378.400 ;
        RECT 377.200 378.300 378.000 378.400 ;
        RECT 338.800 377.700 378.000 378.300 ;
        RECT 338.800 377.600 339.600 377.700 ;
        RECT 346.800 377.600 347.600 377.700 ;
        RECT 377.200 377.600 378.000 377.700 ;
        RECT 494.000 378.300 494.800 378.400 ;
        RECT 526.000 378.300 526.800 378.400 ;
        RECT 494.000 377.700 526.800 378.300 ;
        RECT 494.000 377.600 494.800 377.700 ;
        RECT 526.000 377.600 526.800 377.700 ;
        RECT 530.800 378.300 531.600 378.400 ;
        RECT 543.600 378.300 544.400 378.400 ;
        RECT 530.800 377.700 544.400 378.300 ;
        RECT 530.800 377.600 531.600 377.700 ;
        RECT 543.600 377.600 544.400 377.700 ;
        RECT 567.600 378.300 568.400 378.400 ;
        RECT 570.800 378.300 571.600 378.400 ;
        RECT 567.600 377.700 571.600 378.300 ;
        RECT 567.600 377.600 568.400 377.700 ;
        RECT 570.800 377.600 571.600 377.700 ;
        RECT 577.200 378.300 578.000 378.400 ;
        RECT 580.400 378.300 581.200 378.400 ;
        RECT 577.200 377.700 581.200 378.300 ;
        RECT 577.200 377.600 578.000 377.700 ;
        RECT 580.400 377.600 581.200 377.700 ;
        RECT 618.800 378.300 619.600 378.400 ;
        RECT 634.800 378.300 635.600 378.400 ;
        RECT 618.800 377.700 635.600 378.300 ;
        RECT 618.800 377.600 619.600 377.700 ;
        RECT 634.800 377.600 635.600 377.700 ;
        RECT 638.000 378.300 638.800 378.400 ;
        RECT 642.800 378.300 643.600 378.400 ;
        RECT 638.000 377.700 643.600 378.300 ;
        RECT 638.000 377.600 638.800 377.700 ;
        RECT 642.800 377.600 643.600 377.700 ;
        RECT 33.200 376.300 34.000 376.400 ;
        RECT 46.000 376.300 46.800 376.400 ;
        RECT 33.200 375.700 46.800 376.300 ;
        RECT 33.200 375.600 34.000 375.700 ;
        RECT 46.000 375.600 46.800 375.700 ;
        RECT 57.200 376.300 58.000 376.400 ;
        RECT 63.600 376.300 64.400 376.400 ;
        RECT 57.200 375.700 64.400 376.300 ;
        RECT 57.200 375.600 58.000 375.700 ;
        RECT 63.600 375.600 64.400 375.700 ;
        RECT 66.800 376.300 67.600 376.400 ;
        RECT 70.000 376.300 70.800 376.400 ;
        RECT 66.800 375.700 70.800 376.300 ;
        RECT 66.800 375.600 67.600 375.700 ;
        RECT 70.000 375.600 70.800 375.700 ;
        RECT 71.600 376.300 72.400 376.400 ;
        RECT 82.800 376.300 83.600 376.400 ;
        RECT 134.000 376.300 134.800 376.400 ;
        RECT 137.200 376.300 138.000 376.400 ;
        RECT 71.600 375.700 138.000 376.300 ;
        RECT 71.600 375.600 72.400 375.700 ;
        RECT 82.800 375.600 83.600 375.700 ;
        RECT 134.000 375.600 134.800 375.700 ;
        RECT 137.200 375.600 138.000 375.700 ;
        RECT 177.200 376.300 178.000 376.400 ;
        RECT 193.200 376.300 194.000 376.400 ;
        RECT 177.200 375.700 194.000 376.300 ;
        RECT 177.200 375.600 178.000 375.700 ;
        RECT 193.200 375.600 194.000 375.700 ;
        RECT 206.000 376.300 206.800 376.400 ;
        RECT 230.000 376.300 230.800 376.400 ;
        RECT 206.000 375.700 230.800 376.300 ;
        RECT 206.000 375.600 206.800 375.700 ;
        RECT 230.000 375.600 230.800 375.700 ;
        RECT 234.800 376.300 235.600 376.400 ;
        RECT 250.800 376.300 251.600 376.400 ;
        RECT 234.800 375.700 251.600 376.300 ;
        RECT 234.800 375.600 235.600 375.700 ;
        RECT 250.800 375.600 251.600 375.700 ;
        RECT 282.800 376.300 283.600 376.400 ;
        RECT 287.600 376.300 288.400 376.400 ;
        RECT 292.400 376.300 293.200 376.400 ;
        RECT 282.800 375.700 293.200 376.300 ;
        RECT 282.800 375.600 283.600 375.700 ;
        RECT 287.600 375.600 288.400 375.700 ;
        RECT 292.400 375.600 293.200 375.700 ;
        RECT 298.800 376.300 299.600 376.400 ;
        RECT 306.800 376.300 307.600 376.400 ;
        RECT 298.800 375.700 307.600 376.300 ;
        RECT 298.800 375.600 299.600 375.700 ;
        RECT 306.800 375.600 307.600 375.700 ;
        RECT 310.000 376.300 310.800 376.400 ;
        RECT 316.400 376.300 317.200 376.400 ;
        RECT 310.000 375.700 317.200 376.300 ;
        RECT 310.000 375.600 310.800 375.700 ;
        RECT 316.400 375.600 317.200 375.700 ;
        RECT 321.200 376.300 322.000 376.400 ;
        RECT 326.000 376.300 326.800 376.400 ;
        RECT 321.200 375.700 326.800 376.300 ;
        RECT 321.200 375.600 322.000 375.700 ;
        RECT 326.000 375.600 326.800 375.700 ;
        RECT 342.000 376.300 342.800 376.400 ;
        RECT 353.200 376.300 354.000 376.400 ;
        RECT 342.000 375.700 354.000 376.300 ;
        RECT 342.000 375.600 342.800 375.700 ;
        RECT 353.200 375.600 354.000 375.700 ;
        RECT 361.200 376.300 362.000 376.400 ;
        RECT 367.600 376.300 368.400 376.400 ;
        RECT 361.200 375.700 368.400 376.300 ;
        RECT 361.200 375.600 362.000 375.700 ;
        RECT 367.600 375.600 368.400 375.700 ;
        RECT 433.200 376.300 434.000 376.400 ;
        RECT 452.400 376.300 453.200 376.400 ;
        RECT 466.800 376.300 467.600 376.400 ;
        RECT 433.200 375.700 467.600 376.300 ;
        RECT 433.200 375.600 434.000 375.700 ;
        RECT 452.400 375.600 453.200 375.700 ;
        RECT 466.800 375.600 467.600 375.700 ;
        RECT 489.200 376.300 490.000 376.400 ;
        RECT 500.400 376.300 501.200 376.400 ;
        RECT 489.200 375.700 501.200 376.300 ;
        RECT 489.200 375.600 490.000 375.700 ;
        RECT 500.400 375.600 501.200 375.700 ;
        RECT 526.000 376.300 526.800 376.400 ;
        RECT 540.400 376.300 541.200 376.400 ;
        RECT 569.200 376.300 570.000 376.400 ;
        RECT 526.000 375.700 570.000 376.300 ;
        RECT 526.000 375.600 526.800 375.700 ;
        RECT 540.400 375.600 541.200 375.700 ;
        RECT 569.200 375.600 570.000 375.700 ;
        RECT 572.400 376.300 573.200 376.400 ;
        RECT 582.000 376.300 582.800 376.400 ;
        RECT 572.400 375.700 582.800 376.300 ;
        RECT 572.400 375.600 573.200 375.700 ;
        RECT 582.000 375.600 582.800 375.700 ;
        RECT 590.000 375.600 590.800 376.400 ;
        RECT 599.600 376.300 600.400 376.400 ;
        RECT 638.000 376.300 638.800 376.400 ;
        RECT 641.200 376.300 642.000 376.400 ;
        RECT 599.600 375.700 642.000 376.300 ;
        RECT 599.600 375.600 600.400 375.700 ;
        RECT 638.000 375.600 638.800 375.700 ;
        RECT 641.200 375.600 642.000 375.700 ;
        RECT 18.800 374.300 19.600 374.400 ;
        RECT 28.400 374.300 29.200 374.400 ;
        RECT 52.400 374.300 53.200 374.400 ;
        RECT 65.200 374.300 66.000 374.400 ;
        RECT 18.800 373.700 66.000 374.300 ;
        RECT 18.800 373.600 19.600 373.700 ;
        RECT 28.400 373.600 29.200 373.700 ;
        RECT 52.400 373.600 53.200 373.700 ;
        RECT 65.200 373.600 66.000 373.700 ;
        RECT 70.000 374.300 70.800 374.400 ;
        RECT 81.200 374.300 82.000 374.400 ;
        RECT 70.000 373.700 82.000 374.300 ;
        RECT 70.000 373.600 70.800 373.700 ;
        RECT 81.200 373.600 82.000 373.700 ;
        RECT 122.800 374.300 123.600 374.400 ;
        RECT 126.000 374.300 126.800 374.400 ;
        RECT 122.800 373.700 126.800 374.300 ;
        RECT 122.800 373.600 123.600 373.700 ;
        RECT 126.000 373.600 126.800 373.700 ;
        RECT 138.800 374.300 139.600 374.400 ;
        RECT 174.000 374.300 174.800 374.400 ;
        RECT 138.800 373.700 174.800 374.300 ;
        RECT 138.800 373.600 139.600 373.700 ;
        RECT 174.000 373.600 174.800 373.700 ;
        RECT 178.800 374.300 179.600 374.400 ;
        RECT 214.000 374.300 214.800 374.400 ;
        RECT 178.800 373.700 214.800 374.300 ;
        RECT 178.800 373.600 179.600 373.700 ;
        RECT 214.000 373.600 214.800 373.700 ;
        RECT 220.400 374.300 221.200 374.400 ;
        RECT 230.000 374.300 230.800 374.400 ;
        RECT 220.400 373.700 230.800 374.300 ;
        RECT 220.400 373.600 221.200 373.700 ;
        RECT 230.000 373.600 230.800 373.700 ;
        RECT 236.400 374.300 237.200 374.400 ;
        RECT 271.600 374.300 272.400 374.400 ;
        RECT 236.400 373.700 272.400 374.300 ;
        RECT 236.400 373.600 237.200 373.700 ;
        RECT 271.600 373.600 272.400 373.700 ;
        RECT 284.400 374.300 285.200 374.400 ;
        RECT 294.000 374.300 294.800 374.400 ;
        RECT 284.400 373.700 294.800 374.300 ;
        RECT 284.400 373.600 285.200 373.700 ;
        RECT 294.000 373.600 294.800 373.700 ;
        RECT 319.600 374.300 320.400 374.400 ;
        RECT 324.400 374.300 325.200 374.400 ;
        RECT 319.600 373.700 325.200 374.300 ;
        RECT 319.600 373.600 320.400 373.700 ;
        RECT 324.400 373.600 325.200 373.700 ;
        RECT 511.600 374.300 512.400 374.400 ;
        RECT 534.000 374.300 534.800 374.400 ;
        RECT 511.600 373.700 534.800 374.300 ;
        RECT 511.600 373.600 512.400 373.700 ;
        RECT 534.000 373.600 534.800 373.700 ;
        RECT 537.200 374.300 538.000 374.400 ;
        RECT 607.600 374.300 608.400 374.400 ;
        RECT 618.800 374.300 619.600 374.400 ;
        RECT 537.200 373.700 619.600 374.300 ;
        RECT 537.200 373.600 538.000 373.700 ;
        RECT 607.600 373.600 608.400 373.700 ;
        RECT 618.800 373.600 619.600 373.700 ;
        RECT 628.400 374.300 629.200 374.400 ;
        RECT 631.600 374.300 632.400 374.400 ;
        RECT 628.400 373.700 632.400 374.300 ;
        RECT 628.400 373.600 629.200 373.700 ;
        RECT 631.600 373.600 632.400 373.700 ;
        RECT 642.800 374.300 643.600 374.400 ;
        RECT 647.600 374.300 648.400 374.400 ;
        RECT 642.800 373.700 648.400 374.300 ;
        RECT 642.800 373.600 643.600 373.700 ;
        RECT 647.600 373.600 648.400 373.700 ;
        RECT 657.200 374.300 658.000 374.400 ;
        RECT 658.800 374.300 659.600 374.400 ;
        RECT 657.200 373.700 659.600 374.300 ;
        RECT 657.200 373.600 658.000 373.700 ;
        RECT 658.800 373.600 659.600 373.700 ;
        RECT 673.200 374.300 674.000 374.400 ;
        RECT 679.600 374.300 680.400 374.400 ;
        RECT 673.200 373.700 680.400 374.300 ;
        RECT 673.200 373.600 674.000 373.700 ;
        RECT 679.600 373.600 680.400 373.700 ;
        RECT 7.600 372.300 8.400 372.400 ;
        RECT 30.000 372.300 30.800 372.400 ;
        RECT 7.600 371.700 30.800 372.300 ;
        RECT 7.600 371.600 8.400 371.700 ;
        RECT 30.000 371.600 30.800 371.700 ;
        RECT 44.400 372.300 45.200 372.400 ;
        RECT 68.400 372.300 69.200 372.400 ;
        RECT 44.400 371.700 69.200 372.300 ;
        RECT 44.400 371.600 45.200 371.700 ;
        RECT 68.400 371.600 69.200 371.700 ;
        RECT 79.600 372.300 80.400 372.400 ;
        RECT 90.800 372.300 91.600 372.400 ;
        RECT 79.600 371.700 91.600 372.300 ;
        RECT 79.600 371.600 80.400 371.700 ;
        RECT 90.800 371.600 91.600 371.700 ;
        RECT 94.000 372.300 94.800 372.400 ;
        RECT 95.600 372.300 96.400 372.400 ;
        RECT 94.000 371.700 96.400 372.300 ;
        RECT 94.000 371.600 94.800 371.700 ;
        RECT 95.600 371.600 96.400 371.700 ;
        RECT 108.400 372.300 109.200 372.400 ;
        RECT 119.600 372.300 120.400 372.400 ;
        RECT 137.200 372.300 138.000 372.400 ;
        RECT 108.400 371.700 138.000 372.300 ;
        RECT 108.400 371.600 109.200 371.700 ;
        RECT 119.600 371.600 120.400 371.700 ;
        RECT 137.200 371.600 138.000 371.700 ;
        RECT 161.200 372.300 162.000 372.400 ;
        RECT 170.800 372.300 171.600 372.400 ;
        RECT 161.200 371.700 171.600 372.300 ;
        RECT 161.200 371.600 162.000 371.700 ;
        RECT 170.800 371.600 171.600 371.700 ;
        RECT 175.600 372.300 176.400 372.400 ;
        RECT 183.600 372.300 184.400 372.400 ;
        RECT 175.600 371.700 184.400 372.300 ;
        RECT 175.600 371.600 176.400 371.700 ;
        RECT 183.600 371.600 184.400 371.700 ;
        RECT 226.800 372.300 227.600 372.400 ;
        RECT 284.400 372.300 285.200 372.400 ;
        RECT 286.000 372.300 286.800 372.400 ;
        RECT 226.800 371.700 286.800 372.300 ;
        RECT 226.800 371.600 227.600 371.700 ;
        RECT 284.400 371.600 285.200 371.700 ;
        RECT 286.000 371.600 286.800 371.700 ;
        RECT 326.000 372.300 326.800 372.400 ;
        RECT 329.200 372.300 330.000 372.400 ;
        RECT 326.000 371.700 330.000 372.300 ;
        RECT 326.000 371.600 326.800 371.700 ;
        RECT 329.200 371.600 330.000 371.700 ;
        RECT 340.400 372.300 341.200 372.400 ;
        RECT 346.800 372.300 347.600 372.400 ;
        RECT 340.400 371.700 347.600 372.300 ;
        RECT 340.400 371.600 341.200 371.700 ;
        RECT 346.800 371.600 347.600 371.700 ;
        RECT 361.200 372.300 362.000 372.400 ;
        RECT 362.800 372.300 363.600 372.400 ;
        RECT 375.600 372.300 376.400 372.400 ;
        RECT 361.200 371.700 376.400 372.300 ;
        RECT 361.200 371.600 362.000 371.700 ;
        RECT 362.800 371.600 363.600 371.700 ;
        RECT 375.600 371.600 376.400 371.700 ;
        RECT 402.800 372.300 403.600 372.400 ;
        RECT 412.400 372.300 413.200 372.400 ;
        RECT 402.800 371.700 413.200 372.300 ;
        RECT 402.800 371.600 403.600 371.700 ;
        RECT 412.400 371.600 413.200 371.700 ;
        RECT 446.000 372.300 446.800 372.400 ;
        RECT 457.200 372.300 458.000 372.400 ;
        RECT 446.000 371.700 458.000 372.300 ;
        RECT 446.000 371.600 446.800 371.700 ;
        RECT 457.200 371.600 458.000 371.700 ;
        RECT 490.800 372.300 491.600 372.400 ;
        RECT 500.400 372.300 501.200 372.400 ;
        RECT 511.600 372.300 512.400 372.400 ;
        RECT 490.800 371.700 512.400 372.300 ;
        RECT 490.800 371.600 491.600 371.700 ;
        RECT 500.400 371.600 501.200 371.700 ;
        RECT 511.600 371.600 512.400 371.700 ;
        RECT 516.400 372.300 517.200 372.400 ;
        RECT 556.400 372.300 557.200 372.400 ;
        RECT 569.200 372.300 570.000 372.400 ;
        RECT 516.400 371.700 570.000 372.300 ;
        RECT 516.400 371.600 517.200 371.700 ;
        RECT 556.400 371.600 557.200 371.700 ;
        RECT 569.200 371.600 570.000 371.700 ;
        RECT 578.800 372.300 579.600 372.400 ;
        RECT 582.000 372.300 582.800 372.400 ;
        RECT 591.600 372.300 592.400 372.400 ;
        RECT 578.800 371.700 592.400 372.300 ;
        RECT 578.800 371.600 579.600 371.700 ;
        RECT 582.000 371.600 582.800 371.700 ;
        RECT 591.600 371.600 592.400 371.700 ;
        RECT 598.000 372.300 598.800 372.400 ;
        RECT 602.800 372.300 603.600 372.400 ;
        RECT 598.000 371.700 603.600 372.300 ;
        RECT 598.000 371.600 598.800 371.700 ;
        RECT 602.800 371.600 603.600 371.700 ;
        RECT 634.800 372.300 635.600 372.400 ;
        RECT 639.600 372.300 640.400 372.400 ;
        RECT 634.800 371.700 640.400 372.300 ;
        RECT 634.800 371.600 635.600 371.700 ;
        RECT 639.600 371.600 640.400 371.700 ;
        RECT 42.800 370.300 43.600 370.400 ;
        RECT 55.600 370.300 56.400 370.400 ;
        RECT 42.800 369.700 56.400 370.300 ;
        RECT 42.800 369.600 43.600 369.700 ;
        RECT 55.600 369.600 56.400 369.700 ;
        RECT 62.000 370.300 62.800 370.400 ;
        RECT 73.200 370.300 74.000 370.400 ;
        RECT 103.600 370.300 104.400 370.400 ;
        RECT 62.000 369.700 74.000 370.300 ;
        RECT 62.000 369.600 62.800 369.700 ;
        RECT 73.200 369.600 74.000 369.700 ;
        RECT 98.900 369.700 104.400 370.300 ;
        RECT 62.000 368.300 62.800 368.400 ;
        RECT 98.900 368.300 99.500 369.700 ;
        RECT 103.600 369.600 104.400 369.700 ;
        RECT 111.600 370.300 112.400 370.400 ;
        RECT 122.800 370.300 123.600 370.400 ;
        RECT 111.600 369.700 123.600 370.300 ;
        RECT 111.600 369.600 112.400 369.700 ;
        RECT 122.800 369.600 123.600 369.700 ;
        RECT 162.800 370.300 163.600 370.400 ;
        RECT 186.800 370.300 187.600 370.400 ;
        RECT 162.800 369.700 187.600 370.300 ;
        RECT 162.800 369.600 163.600 369.700 ;
        RECT 186.800 369.600 187.600 369.700 ;
        RECT 204.400 370.300 205.200 370.400 ;
        RECT 241.200 370.300 242.000 370.400 ;
        RECT 204.400 369.700 242.000 370.300 ;
        RECT 204.400 369.600 205.200 369.700 ;
        RECT 241.200 369.600 242.000 369.700 ;
        RECT 319.600 370.300 320.400 370.400 ;
        RECT 337.200 370.300 338.000 370.400 ;
        RECT 350.000 370.300 350.800 370.400 ;
        RECT 319.600 369.700 338.000 370.300 ;
        RECT 319.600 369.600 320.400 369.700 ;
        RECT 337.200 369.600 338.000 369.700 ;
        RECT 338.900 369.700 350.800 370.300 ;
        RECT 62.000 367.700 99.500 368.300 ;
        RECT 100.400 368.300 101.200 368.400 ;
        RECT 114.800 368.300 115.600 368.400 ;
        RECT 100.400 367.700 115.600 368.300 ;
        RECT 62.000 367.600 62.800 367.700 ;
        RECT 100.400 367.600 101.200 367.700 ;
        RECT 114.800 367.600 115.600 367.700 ;
        RECT 116.400 368.300 117.200 368.400 ;
        RECT 118.000 368.300 118.800 368.400 ;
        RECT 134.000 368.300 134.800 368.400 ;
        RECT 233.200 368.300 234.000 368.400 ;
        RECT 116.400 367.700 134.800 368.300 ;
        RECT 116.400 367.600 117.200 367.700 ;
        RECT 118.000 367.600 118.800 367.700 ;
        RECT 134.000 367.600 134.800 367.700 ;
        RECT 218.900 367.700 234.000 368.300 ;
        RECT 66.800 366.300 67.600 366.400 ;
        RECT 78.000 366.300 78.800 366.400 ;
        RECT 66.800 365.700 78.800 366.300 ;
        RECT 66.800 365.600 67.600 365.700 ;
        RECT 78.000 365.600 78.800 365.700 ;
        RECT 94.000 366.300 94.800 366.400 ;
        RECT 108.400 366.300 109.200 366.400 ;
        RECT 94.000 365.700 109.200 366.300 ;
        RECT 94.000 365.600 94.800 365.700 ;
        RECT 108.400 365.600 109.200 365.700 ;
        RECT 122.800 366.300 123.600 366.400 ;
        RECT 218.900 366.300 219.500 367.700 ;
        RECT 233.200 367.600 234.000 367.700 ;
        RECT 316.400 368.300 317.200 368.400 ;
        RECT 338.900 368.300 339.500 369.700 ;
        RECT 350.000 369.600 350.800 369.700 ;
        RECT 358.000 370.300 358.800 370.400 ;
        RECT 366.000 370.300 366.800 370.400 ;
        RECT 370.800 370.300 371.600 370.400 ;
        RECT 358.000 369.700 371.600 370.300 ;
        RECT 358.000 369.600 358.800 369.700 ;
        RECT 366.000 369.600 366.800 369.700 ;
        RECT 370.800 369.600 371.600 369.700 ;
        RECT 372.400 370.300 373.200 370.400 ;
        RECT 378.800 370.300 379.600 370.400 ;
        RECT 372.400 369.700 379.600 370.300 ;
        RECT 372.400 369.600 373.200 369.700 ;
        RECT 378.800 369.600 379.600 369.700 ;
        RECT 380.400 370.300 381.200 370.400 ;
        RECT 385.200 370.300 386.000 370.400 ;
        RECT 380.400 369.700 386.000 370.300 ;
        RECT 380.400 369.600 381.200 369.700 ;
        RECT 385.200 369.600 386.000 369.700 ;
        RECT 388.400 370.300 389.200 370.400 ;
        RECT 393.200 370.300 394.000 370.400 ;
        RECT 388.400 369.700 394.000 370.300 ;
        RECT 388.400 369.600 389.200 369.700 ;
        RECT 393.200 369.600 394.000 369.700 ;
        RECT 482.800 370.300 483.600 370.400 ;
        RECT 503.600 370.300 504.400 370.400 ;
        RECT 482.800 369.700 504.400 370.300 ;
        RECT 482.800 369.600 483.600 369.700 ;
        RECT 503.600 369.600 504.400 369.700 ;
        RECT 529.200 370.300 530.000 370.400 ;
        RECT 532.400 370.300 533.200 370.400 ;
        RECT 545.200 370.300 546.000 370.400 ;
        RECT 578.900 370.300 579.500 371.600 ;
        RECT 609.200 370.300 610.000 370.400 ;
        RECT 618.800 370.300 619.600 370.400 ;
        RECT 529.200 369.700 579.500 370.300 ;
        RECT 580.500 369.700 619.600 370.300 ;
        RECT 529.200 369.600 530.000 369.700 ;
        RECT 532.400 369.600 533.200 369.700 ;
        RECT 545.200 369.600 546.000 369.700 ;
        RECT 316.400 367.700 339.500 368.300 ;
        RECT 340.400 368.300 341.200 368.400 ;
        RECT 348.400 368.300 349.200 368.400 ;
        RECT 394.800 368.300 395.600 368.400 ;
        RECT 340.400 367.700 395.600 368.300 ;
        RECT 316.400 367.600 317.200 367.700 ;
        RECT 340.400 367.600 341.200 367.700 ;
        RECT 348.400 367.600 349.200 367.700 ;
        RECT 394.800 367.600 395.600 367.700 ;
        RECT 410.800 368.300 411.600 368.400 ;
        RECT 449.200 368.300 450.000 368.400 ;
        RECT 410.800 367.700 450.000 368.300 ;
        RECT 410.800 367.600 411.600 367.700 ;
        RECT 449.200 367.600 450.000 367.700 ;
        RECT 510.000 368.300 510.800 368.400 ;
        RECT 546.800 368.300 547.600 368.400 ;
        RECT 510.000 367.700 547.600 368.300 ;
        RECT 510.000 367.600 510.800 367.700 ;
        RECT 546.800 367.600 547.600 367.700 ;
        RECT 562.800 368.300 563.600 368.400 ;
        RECT 570.800 368.300 571.600 368.400 ;
        RECT 562.800 367.700 571.600 368.300 ;
        RECT 562.800 367.600 563.600 367.700 ;
        RECT 570.800 367.600 571.600 367.700 ;
        RECT 572.400 368.300 573.200 368.400 ;
        RECT 580.500 368.300 581.100 369.700 ;
        RECT 609.200 369.600 610.000 369.700 ;
        RECT 618.800 369.600 619.600 369.700 ;
        RECT 625.200 370.300 626.000 370.400 ;
        RECT 628.400 370.300 629.200 370.400 ;
        RECT 625.200 369.700 629.200 370.300 ;
        RECT 625.200 369.600 626.000 369.700 ;
        RECT 628.400 369.600 629.200 369.700 ;
        RECT 639.600 370.300 640.400 370.400 ;
        RECT 644.400 370.300 645.200 370.400 ;
        RECT 639.600 369.700 645.200 370.300 ;
        RECT 639.600 369.600 640.400 369.700 ;
        RECT 644.400 369.600 645.200 369.700 ;
        RECT 572.400 367.700 581.100 368.300 ;
        RECT 588.400 368.300 589.200 368.400 ;
        RECT 593.200 368.300 594.000 368.400 ;
        RECT 588.400 367.700 594.000 368.300 ;
        RECT 572.400 367.600 573.200 367.700 ;
        RECT 588.400 367.600 589.200 367.700 ;
        RECT 593.200 367.600 594.000 367.700 ;
        RECT 622.000 368.300 622.800 368.400 ;
        RECT 636.400 368.300 637.200 368.400 ;
        RECT 622.000 367.700 637.200 368.300 ;
        RECT 622.000 367.600 622.800 367.700 ;
        RECT 636.400 367.600 637.200 367.700 ;
        RECT 647.600 368.300 648.400 368.400 ;
        RECT 649.200 368.300 650.000 368.400 ;
        RECT 647.600 367.700 650.000 368.300 ;
        RECT 647.600 367.600 648.400 367.700 ;
        RECT 649.200 367.600 650.000 367.700 ;
        RECT 650.800 368.300 651.600 368.400 ;
        RECT 657.200 368.300 658.000 368.400 ;
        RECT 650.800 367.700 658.000 368.300 ;
        RECT 650.800 367.600 651.600 367.700 ;
        RECT 657.200 367.600 658.000 367.700 ;
        RECT 122.800 365.700 219.500 366.300 ;
        RECT 220.400 366.300 221.200 366.400 ;
        RECT 281.200 366.300 282.000 366.400 ;
        RECT 220.400 365.700 282.000 366.300 ;
        RECT 122.800 365.600 123.600 365.700 ;
        RECT 220.400 365.600 221.200 365.700 ;
        RECT 281.200 365.600 282.000 365.700 ;
        RECT 300.400 366.300 301.200 366.400 ;
        RECT 324.400 366.300 325.200 366.400 ;
        RECT 300.400 365.700 325.200 366.300 ;
        RECT 300.400 365.600 301.200 365.700 ;
        RECT 324.400 365.600 325.200 365.700 ;
        RECT 327.600 366.300 328.400 366.400 ;
        RECT 343.600 366.300 344.400 366.400 ;
        RECT 327.600 365.700 344.400 366.300 ;
        RECT 327.600 365.600 328.400 365.700 ;
        RECT 343.600 365.600 344.400 365.700 ;
        RECT 348.400 366.300 349.200 366.400 ;
        RECT 369.200 366.300 370.000 366.400 ;
        RECT 348.400 365.700 370.000 366.300 ;
        RECT 348.400 365.600 349.200 365.700 ;
        RECT 369.200 365.600 370.000 365.700 ;
        RECT 375.600 366.300 376.400 366.400 ;
        RECT 380.400 366.300 381.200 366.400 ;
        RECT 375.600 365.700 381.200 366.300 ;
        RECT 375.600 365.600 376.400 365.700 ;
        RECT 380.400 365.600 381.200 365.700 ;
        RECT 382.000 366.300 382.800 366.400 ;
        RECT 393.200 366.300 394.000 366.400 ;
        RECT 382.000 365.700 394.000 366.300 ;
        RECT 382.000 365.600 382.800 365.700 ;
        RECT 393.200 365.600 394.000 365.700 ;
        RECT 417.200 366.300 418.000 366.400 ;
        RECT 422.000 366.300 422.800 366.400 ;
        RECT 417.200 365.700 422.800 366.300 ;
        RECT 417.200 365.600 418.000 365.700 ;
        RECT 422.000 365.600 422.800 365.700 ;
        RECT 535.600 366.300 536.400 366.400 ;
        RECT 598.000 366.300 598.800 366.400 ;
        RECT 612.400 366.300 613.200 366.400 ;
        RECT 535.600 365.700 613.200 366.300 ;
        RECT 535.600 365.600 536.400 365.700 ;
        RECT 598.000 365.600 598.800 365.700 ;
        RECT 612.400 365.600 613.200 365.700 ;
        RECT 94.000 364.300 94.800 364.400 ;
        RECT 97.200 364.300 98.000 364.400 ;
        RECT 94.000 363.700 98.000 364.300 ;
        RECT 94.000 363.600 94.800 363.700 ;
        RECT 97.200 363.600 98.000 363.700 ;
        RECT 103.600 364.300 104.400 364.400 ;
        RECT 239.600 364.300 240.400 364.400 ;
        RECT 103.600 363.700 240.400 364.300 ;
        RECT 103.600 363.600 104.400 363.700 ;
        RECT 239.600 363.600 240.400 363.700 ;
        RECT 302.000 364.300 302.800 364.400 ;
        RECT 402.800 364.300 403.600 364.400 ;
        RECT 433.200 364.300 434.000 364.400 ;
        RECT 302.000 363.700 434.000 364.300 ;
        RECT 302.000 363.600 302.800 363.700 ;
        RECT 402.800 363.600 403.600 363.700 ;
        RECT 433.200 363.600 434.000 363.700 ;
        RECT 530.800 364.300 531.600 364.400 ;
        RECT 626.800 364.300 627.600 364.400 ;
        RECT 530.800 363.700 627.600 364.300 ;
        RECT 530.800 363.600 531.600 363.700 ;
        RECT 626.800 363.600 627.600 363.700 ;
        RECT 127.600 362.300 128.400 362.400 ;
        RECT 166.000 362.300 166.800 362.400 ;
        RECT 127.600 361.700 166.800 362.300 ;
        RECT 127.600 361.600 128.400 361.700 ;
        RECT 166.000 361.600 166.800 361.700 ;
        RECT 278.000 362.300 278.800 362.400 ;
        RECT 326.000 362.300 326.800 362.400 ;
        RECT 278.000 361.700 326.800 362.300 ;
        RECT 278.000 361.600 278.800 361.700 ;
        RECT 326.000 361.600 326.800 361.700 ;
        RECT 334.000 362.300 334.800 362.400 ;
        RECT 372.400 362.300 373.200 362.400 ;
        RECT 334.000 361.700 373.200 362.300 ;
        RECT 334.000 361.600 334.800 361.700 ;
        RECT 372.400 361.600 373.200 361.700 ;
        RECT 375.600 362.300 376.400 362.400 ;
        RECT 398.000 362.300 398.800 362.400 ;
        RECT 375.600 361.700 398.800 362.300 ;
        RECT 375.600 361.600 376.400 361.700 ;
        RECT 398.000 361.600 398.800 361.700 ;
        RECT 433.200 362.300 434.000 362.400 ;
        RECT 436.400 362.300 437.200 362.400 ;
        RECT 433.200 361.700 437.200 362.300 ;
        RECT 433.200 361.600 434.000 361.700 ;
        RECT 436.400 361.600 437.200 361.700 ;
        RECT 519.600 362.300 520.400 362.400 ;
        RECT 543.600 362.300 544.400 362.400 ;
        RECT 519.600 361.700 544.400 362.300 ;
        RECT 519.600 361.600 520.400 361.700 ;
        RECT 543.600 361.600 544.400 361.700 ;
        RECT 647.600 362.300 648.400 362.400 ;
        RECT 649.200 362.300 650.000 362.400 ;
        RECT 654.000 362.300 654.800 362.400 ;
        RECT 679.600 362.300 680.400 362.400 ;
        RECT 647.600 361.700 680.400 362.300 ;
        RECT 647.600 361.600 648.400 361.700 ;
        RECT 649.200 361.600 650.000 361.700 ;
        RECT 654.000 361.600 654.800 361.700 ;
        RECT 679.600 361.600 680.400 361.700 ;
        RECT 18.800 360.300 19.600 360.400 ;
        RECT 42.800 360.300 43.600 360.400 ;
        RECT 18.800 359.700 43.600 360.300 ;
        RECT 18.800 359.600 19.600 359.700 ;
        RECT 42.800 359.600 43.600 359.700 ;
        RECT 212.400 360.300 213.200 360.400 ;
        RECT 310.000 360.300 310.800 360.400 ;
        RECT 332.400 360.300 333.200 360.400 ;
        RECT 212.400 359.700 333.200 360.300 ;
        RECT 212.400 359.600 213.200 359.700 ;
        RECT 310.000 359.600 310.800 359.700 ;
        RECT 332.400 359.600 333.200 359.700 ;
        RECT 335.600 360.300 336.400 360.400 ;
        RECT 342.000 360.300 342.800 360.400 ;
        RECT 335.600 359.700 342.800 360.300 ;
        RECT 335.600 359.600 336.400 359.700 ;
        RECT 342.000 359.600 342.800 359.700 ;
        RECT 377.200 360.300 378.000 360.400 ;
        RECT 380.400 360.300 381.200 360.400 ;
        RECT 377.200 359.700 381.200 360.300 ;
        RECT 377.200 359.600 378.000 359.700 ;
        RECT 380.400 359.600 381.200 359.700 ;
        RECT 538.800 360.300 539.600 360.400 ;
        RECT 542.000 360.300 542.800 360.400 ;
        RECT 538.800 359.700 542.800 360.300 ;
        RECT 538.800 359.600 539.600 359.700 ;
        RECT 542.000 359.600 542.800 359.700 ;
        RECT 548.400 360.300 549.200 360.400 ;
        RECT 564.400 360.300 565.200 360.400 ;
        RECT 548.400 359.700 565.200 360.300 ;
        RECT 548.400 359.600 549.200 359.700 ;
        RECT 564.400 359.600 565.200 359.700 ;
        RECT 590.000 360.300 590.800 360.400 ;
        RECT 650.800 360.300 651.600 360.400 ;
        RECT 590.000 359.700 651.600 360.300 ;
        RECT 590.000 359.600 590.800 359.700 ;
        RECT 650.800 359.600 651.600 359.700 ;
        RECT 666.800 360.300 667.600 360.400 ;
        RECT 670.000 360.300 670.800 360.400 ;
        RECT 666.800 359.700 670.800 360.300 ;
        RECT 666.800 359.600 667.600 359.700 ;
        RECT 670.000 359.600 670.800 359.700 ;
        RECT 38.000 358.300 38.800 358.400 ;
        RECT 46.000 358.300 46.800 358.400 ;
        RECT 92.400 358.300 93.200 358.400 ;
        RECT 106.800 358.300 107.600 358.400 ;
        RECT 38.000 357.700 107.600 358.300 ;
        RECT 38.000 357.600 38.800 357.700 ;
        RECT 46.000 357.600 46.800 357.700 ;
        RECT 92.400 357.600 93.200 357.700 ;
        RECT 106.800 357.600 107.600 357.700 ;
        RECT 116.400 358.300 117.200 358.400 ;
        RECT 121.200 358.300 122.000 358.400 ;
        RECT 116.400 357.700 122.000 358.300 ;
        RECT 116.400 357.600 117.200 357.700 ;
        RECT 121.200 357.600 122.000 357.700 ;
        RECT 150.000 358.300 150.800 358.400 ;
        RECT 151.600 358.300 152.400 358.400 ;
        RECT 150.000 357.700 152.400 358.300 ;
        RECT 150.000 357.600 150.800 357.700 ;
        RECT 151.600 357.600 152.400 357.700 ;
        RECT 314.800 358.300 315.600 358.400 ;
        RECT 329.200 358.300 330.000 358.400 ;
        RECT 314.800 357.700 330.000 358.300 ;
        RECT 314.800 357.600 315.600 357.700 ;
        RECT 329.200 357.600 330.000 357.700 ;
        RECT 330.800 358.300 331.600 358.400 ;
        RECT 334.000 358.300 334.800 358.400 ;
        RECT 330.800 357.700 334.800 358.300 ;
        RECT 330.800 357.600 331.600 357.700 ;
        RECT 334.000 357.600 334.800 357.700 ;
        RECT 350.000 358.300 350.800 358.400 ;
        RECT 366.000 358.300 366.800 358.400 ;
        RECT 350.000 357.700 366.800 358.300 ;
        RECT 350.000 357.600 350.800 357.700 ;
        RECT 366.000 357.600 366.800 357.700 ;
        RECT 401.200 358.300 402.000 358.400 ;
        RECT 423.600 358.300 424.400 358.400 ;
        RECT 428.400 358.300 429.200 358.400 ;
        RECT 442.800 358.300 443.600 358.400 ;
        RECT 401.200 357.700 443.600 358.300 ;
        RECT 401.200 357.600 402.000 357.700 ;
        RECT 423.600 357.600 424.400 357.700 ;
        RECT 428.400 357.600 429.200 357.700 ;
        RECT 442.800 357.600 443.600 357.700 ;
        RECT 481.200 358.300 482.000 358.400 ;
        RECT 487.600 358.300 488.400 358.400 ;
        RECT 481.200 357.700 488.400 358.300 ;
        RECT 481.200 357.600 482.000 357.700 ;
        RECT 487.600 357.600 488.400 357.700 ;
        RECT 546.800 358.300 547.600 358.400 ;
        RECT 633.200 358.300 634.000 358.400 ;
        RECT 546.800 357.700 634.000 358.300 ;
        RECT 546.800 357.600 547.600 357.700 ;
        RECT 633.200 357.600 634.000 357.700 ;
        RECT 655.600 358.300 656.400 358.400 ;
        RECT 670.000 358.300 670.800 358.400 ;
        RECT 655.600 357.700 670.800 358.300 ;
        RECT 655.600 357.600 656.400 357.700 ;
        RECT 670.000 357.600 670.800 357.700 ;
        RECT 25.200 356.300 26.000 356.400 ;
        RECT 34.800 356.300 35.600 356.400 ;
        RECT 25.200 355.700 35.600 356.300 ;
        RECT 25.200 355.600 26.000 355.700 ;
        RECT 34.800 355.600 35.600 355.700 ;
        RECT 58.800 356.300 59.600 356.400 ;
        RECT 70.000 356.300 70.800 356.400 ;
        RECT 58.800 355.700 70.800 356.300 ;
        RECT 58.800 355.600 59.600 355.700 ;
        RECT 70.000 355.600 70.800 355.700 ;
        RECT 95.600 356.300 96.400 356.400 ;
        RECT 132.400 356.300 133.200 356.400 ;
        RECT 135.600 356.300 136.400 356.400 ;
        RECT 169.200 356.300 170.000 356.400 ;
        RECT 95.600 355.700 170.000 356.300 ;
        RECT 95.600 355.600 96.400 355.700 ;
        RECT 132.400 355.600 133.200 355.700 ;
        RECT 135.600 355.600 136.400 355.700 ;
        RECT 169.200 355.600 170.000 355.700 ;
        RECT 204.400 356.300 205.200 356.400 ;
        RECT 281.200 356.300 282.000 356.400 ;
        RECT 290.800 356.300 291.600 356.400 ;
        RECT 204.400 355.700 291.600 356.300 ;
        RECT 204.400 355.600 205.200 355.700 ;
        RECT 281.200 355.600 282.000 355.700 ;
        RECT 290.800 355.600 291.600 355.700 ;
        RECT 311.600 356.300 312.400 356.400 ;
        RECT 314.800 356.300 315.600 356.400 ;
        RECT 343.600 356.300 344.400 356.400 ;
        RECT 346.800 356.300 347.600 356.400 ;
        RECT 311.600 355.700 347.600 356.300 ;
        RECT 311.600 355.600 312.400 355.700 ;
        RECT 314.800 355.600 315.600 355.700 ;
        RECT 343.600 355.600 344.400 355.700 ;
        RECT 346.800 355.600 347.600 355.700 ;
        RECT 348.400 356.300 349.200 356.400 ;
        RECT 356.400 356.300 357.200 356.400 ;
        RECT 348.400 355.700 357.200 356.300 ;
        RECT 348.400 355.600 349.200 355.700 ;
        RECT 356.400 355.600 357.200 355.700 ;
        RECT 519.600 356.300 520.400 356.400 ;
        RECT 532.400 356.300 533.200 356.400 ;
        RECT 519.600 355.700 533.200 356.300 ;
        RECT 519.600 355.600 520.400 355.700 ;
        RECT 532.400 355.600 533.200 355.700 ;
        RECT 550.000 356.300 550.800 356.400 ;
        RECT 561.200 356.300 562.000 356.400 ;
        RECT 578.800 356.300 579.600 356.400 ;
        RECT 550.000 355.700 579.600 356.300 ;
        RECT 550.000 355.600 550.800 355.700 ;
        RECT 561.200 355.600 562.000 355.700 ;
        RECT 578.800 355.600 579.600 355.700 ;
        RECT 606.000 356.300 606.800 356.400 ;
        RECT 631.600 356.300 632.400 356.400 ;
        RECT 606.000 355.700 632.400 356.300 ;
        RECT 606.000 355.600 606.800 355.700 ;
        RECT 631.600 355.600 632.400 355.700 ;
        RECT 30.000 354.300 30.800 354.400 ;
        RECT 39.600 354.300 40.400 354.400 ;
        RECT 30.000 353.700 40.400 354.300 ;
        RECT 30.000 353.600 30.800 353.700 ;
        RECT 39.600 353.600 40.400 353.700 ;
        RECT 68.400 354.300 69.200 354.400 ;
        RECT 78.000 354.300 78.800 354.400 ;
        RECT 68.400 353.700 78.800 354.300 ;
        RECT 68.400 353.600 69.200 353.700 ;
        RECT 78.000 353.600 78.800 353.700 ;
        RECT 106.800 354.300 107.600 354.400 ;
        RECT 114.800 354.300 115.600 354.400 ;
        RECT 106.800 353.700 115.600 354.300 ;
        RECT 106.800 353.600 107.600 353.700 ;
        RECT 114.800 353.600 115.600 353.700 ;
        RECT 119.600 354.300 120.400 354.400 ;
        RECT 126.000 354.300 126.800 354.400 ;
        RECT 119.600 353.700 126.800 354.300 ;
        RECT 119.600 353.600 120.400 353.700 ;
        RECT 126.000 353.600 126.800 353.700 ;
        RECT 156.400 354.300 157.200 354.400 ;
        RECT 162.800 354.300 163.600 354.400 ;
        RECT 228.400 354.300 229.200 354.400 ;
        RECT 156.400 353.700 229.200 354.300 ;
        RECT 156.400 353.600 157.200 353.700 ;
        RECT 162.800 353.600 163.600 353.700 ;
        RECT 228.400 353.600 229.200 353.700 ;
        RECT 236.400 354.300 237.200 354.400 ;
        RECT 273.200 354.300 274.000 354.400 ;
        RECT 236.400 353.700 274.000 354.300 ;
        RECT 236.400 353.600 237.200 353.700 ;
        RECT 273.200 353.600 274.000 353.700 ;
        RECT 311.600 354.300 312.400 354.400 ;
        RECT 316.400 354.300 317.200 354.400 ;
        RECT 327.600 354.300 328.400 354.400 ;
        RECT 330.800 354.300 331.600 354.400 ;
        RECT 311.600 353.700 331.600 354.300 ;
        RECT 311.600 353.600 312.400 353.700 ;
        RECT 316.400 353.600 317.200 353.700 ;
        RECT 327.600 353.600 328.400 353.700 ;
        RECT 330.800 353.600 331.600 353.700 ;
        RECT 332.400 354.300 333.200 354.400 ;
        RECT 374.000 354.300 374.800 354.400 ;
        RECT 332.400 353.700 374.800 354.300 ;
        RECT 332.400 353.600 333.200 353.700 ;
        RECT 374.000 353.600 374.800 353.700 ;
        RECT 375.600 354.300 376.400 354.400 ;
        RECT 382.000 354.300 382.800 354.400 ;
        RECT 375.600 353.700 382.800 354.300 ;
        RECT 375.600 353.600 376.400 353.700 ;
        RECT 382.000 353.600 382.800 353.700 ;
        RECT 522.800 354.300 523.600 354.400 ;
        RECT 530.800 354.300 531.600 354.400 ;
        RECT 522.800 353.700 531.600 354.300 ;
        RECT 522.800 353.600 523.600 353.700 ;
        RECT 530.800 353.600 531.600 353.700 ;
        RECT 542.000 354.300 542.800 354.400 ;
        RECT 566.000 354.300 566.800 354.400 ;
        RECT 542.000 353.700 566.800 354.300 ;
        RECT 542.000 353.600 542.800 353.700 ;
        RECT 566.000 353.600 566.800 353.700 ;
        RECT 580.400 354.300 581.200 354.400 ;
        RECT 623.600 354.300 624.400 354.400 ;
        RECT 580.400 353.700 624.400 354.300 ;
        RECT 580.400 353.600 581.200 353.700 ;
        RECT 623.600 353.600 624.400 353.700 ;
        RECT 626.800 354.300 627.600 354.400 ;
        RECT 636.400 354.300 637.200 354.400 ;
        RECT 626.800 353.700 637.200 354.300 ;
        RECT 626.800 353.600 627.600 353.700 ;
        RECT 636.400 353.600 637.200 353.700 ;
        RECT 638.000 353.600 638.800 354.400 ;
        RECT 23.600 352.300 24.400 352.400 ;
        RECT 26.800 352.300 27.600 352.400 ;
        RECT 23.600 351.700 27.600 352.300 ;
        RECT 23.600 351.600 24.400 351.700 ;
        RECT 26.800 351.600 27.600 351.700 ;
        RECT 38.000 352.300 38.800 352.400 ;
        RECT 65.200 352.300 66.000 352.400 ;
        RECT 70.000 352.300 70.800 352.400 ;
        RECT 38.000 351.700 53.100 352.300 ;
        RECT 38.000 351.600 38.800 351.700 ;
        RECT 52.500 350.400 53.100 351.700 ;
        RECT 65.200 351.700 70.800 352.300 ;
        RECT 65.200 351.600 66.000 351.700 ;
        RECT 70.000 351.600 70.800 351.700 ;
        RECT 71.600 352.300 72.400 352.400 ;
        RECT 74.800 352.300 75.600 352.400 ;
        RECT 71.600 351.700 75.600 352.300 ;
        RECT 71.600 351.600 72.400 351.700 ;
        RECT 74.800 351.600 75.600 351.700 ;
        RECT 89.200 352.300 90.000 352.400 ;
        RECT 90.800 352.300 91.600 352.400 ;
        RECT 89.200 351.700 91.600 352.300 ;
        RECT 89.200 351.600 90.000 351.700 ;
        RECT 90.800 351.600 91.600 351.700 ;
        RECT 100.400 352.300 101.200 352.400 ;
        RECT 126.000 352.300 126.800 352.400 ;
        RECT 100.400 351.700 126.800 352.300 ;
        RECT 100.400 351.600 101.200 351.700 ;
        RECT 126.000 351.600 126.800 351.700 ;
        RECT 130.800 352.300 131.600 352.400 ;
        RECT 138.800 352.300 139.600 352.400 ;
        RECT 130.800 351.700 139.600 352.300 ;
        RECT 130.800 351.600 131.600 351.700 ;
        RECT 138.800 351.600 139.600 351.700 ;
        RECT 154.800 352.300 155.600 352.400 ;
        RECT 158.000 352.300 158.800 352.400 ;
        RECT 154.800 351.700 158.800 352.300 ;
        RECT 154.800 351.600 155.600 351.700 ;
        RECT 158.000 351.600 158.800 351.700 ;
        RECT 159.600 352.300 160.400 352.400 ;
        RECT 164.400 352.300 165.200 352.400 ;
        RECT 159.600 351.700 165.200 352.300 ;
        RECT 159.600 351.600 160.400 351.700 ;
        RECT 164.400 351.600 165.200 351.700 ;
        RECT 222.000 352.300 222.800 352.400 ;
        RECT 228.400 352.300 229.200 352.400 ;
        RECT 222.000 351.700 229.200 352.300 ;
        RECT 222.000 351.600 222.800 351.700 ;
        RECT 228.400 351.600 229.200 351.700 ;
        RECT 297.200 352.300 298.000 352.400 ;
        RECT 302.000 352.300 302.800 352.400 ;
        RECT 297.200 351.700 302.800 352.300 ;
        RECT 297.200 351.600 298.000 351.700 ;
        RECT 302.000 351.600 302.800 351.700 ;
        RECT 305.200 352.300 306.000 352.400 ;
        RECT 318.000 352.300 318.800 352.400 ;
        RECT 305.200 351.700 318.800 352.300 ;
        RECT 305.200 351.600 306.000 351.700 ;
        RECT 318.000 351.600 318.800 351.700 ;
        RECT 322.800 352.300 323.600 352.400 ;
        RECT 338.800 352.300 339.600 352.400 ;
        RECT 434.800 352.300 435.600 352.400 ;
        RECT 538.800 352.300 539.600 352.400 ;
        RECT 545.200 352.300 546.000 352.400 ;
        RECT 548.400 352.300 549.200 352.400 ;
        RECT 322.800 351.700 336.300 352.300 ;
        RECT 322.800 351.600 323.600 351.700 ;
        RECT 23.600 350.300 24.400 350.400 ;
        RECT 34.800 350.300 35.600 350.400 ;
        RECT 23.600 349.700 35.600 350.300 ;
        RECT 23.600 349.600 24.400 349.700 ;
        RECT 34.800 349.600 35.600 349.700 ;
        RECT 42.800 350.300 43.600 350.400 ;
        RECT 47.600 350.300 48.400 350.400 ;
        RECT 42.800 349.700 48.400 350.300 ;
        RECT 42.800 349.600 43.600 349.700 ;
        RECT 47.600 349.600 48.400 349.700 ;
        RECT 52.400 350.300 53.200 350.400 ;
        RECT 55.600 350.300 56.400 350.400 ;
        RECT 52.400 349.700 56.400 350.300 ;
        RECT 52.400 349.600 53.200 349.700 ;
        RECT 55.600 349.600 56.400 349.700 ;
        RECT 63.600 350.300 64.400 350.400 ;
        RECT 78.000 350.300 78.800 350.400 ;
        RECT 63.600 349.700 78.800 350.300 ;
        RECT 63.600 349.600 64.400 349.700 ;
        RECT 78.000 349.600 78.800 349.700 ;
        RECT 86.000 350.300 86.800 350.400 ;
        RECT 114.800 350.300 115.600 350.400 ;
        RECT 86.000 349.700 115.600 350.300 ;
        RECT 86.000 349.600 86.800 349.700 ;
        RECT 114.800 349.600 115.600 349.700 ;
        RECT 118.000 350.300 118.800 350.400 ;
        RECT 121.200 350.300 122.000 350.400 ;
        RECT 118.000 349.700 122.000 350.300 ;
        RECT 118.000 349.600 118.800 349.700 ;
        RECT 121.200 349.600 122.000 349.700 ;
        RECT 126.000 350.300 126.800 350.400 ;
        RECT 132.400 350.300 133.200 350.400 ;
        RECT 126.000 349.700 133.200 350.300 ;
        RECT 126.000 349.600 126.800 349.700 ;
        RECT 132.400 349.600 133.200 349.700 ;
        RECT 167.600 349.600 168.400 350.400 ;
        RECT 223.600 350.300 224.400 350.400 ;
        RECT 231.600 350.300 232.400 350.400 ;
        RECT 223.600 349.700 232.400 350.300 ;
        RECT 223.600 349.600 224.400 349.700 ;
        RECT 231.600 349.600 232.400 349.700 ;
        RECT 241.200 350.300 242.000 350.400 ;
        RECT 244.400 350.300 245.200 350.400 ;
        RECT 241.200 349.700 245.200 350.300 ;
        RECT 241.200 349.600 242.000 349.700 ;
        RECT 244.400 349.600 245.200 349.700 ;
        RECT 254.000 350.300 254.800 350.400 ;
        RECT 257.200 350.300 258.000 350.400 ;
        RECT 254.000 349.700 258.000 350.300 ;
        RECT 254.000 349.600 254.800 349.700 ;
        RECT 257.200 349.600 258.000 349.700 ;
        RECT 313.200 350.300 314.000 350.400 ;
        RECT 321.200 350.300 322.000 350.400 ;
        RECT 313.200 349.700 322.000 350.300 ;
        RECT 313.200 349.600 314.000 349.700 ;
        RECT 321.200 349.600 322.000 349.700 ;
        RECT 324.400 350.300 325.200 350.400 ;
        RECT 334.000 350.300 334.800 350.400 ;
        RECT 324.400 349.700 334.800 350.300 ;
        RECT 335.700 350.300 336.300 351.700 ;
        RECT 338.800 351.700 357.100 352.300 ;
        RECT 338.800 351.600 339.600 351.700 ;
        RECT 356.500 350.400 357.100 351.700 ;
        RECT 434.800 351.700 528.300 352.300 ;
        RECT 434.800 351.600 435.600 351.700 ;
        RECT 343.600 350.300 344.400 350.400 ;
        RECT 353.200 350.300 354.000 350.400 ;
        RECT 335.700 349.700 354.000 350.300 ;
        RECT 324.400 349.600 325.200 349.700 ;
        RECT 334.000 349.600 334.800 349.700 ;
        RECT 343.600 349.600 344.400 349.700 ;
        RECT 353.200 349.600 354.000 349.700 ;
        RECT 356.400 350.300 357.200 350.400 ;
        RECT 370.800 350.300 371.600 350.400 ;
        RECT 382.000 350.300 382.800 350.400 ;
        RECT 356.400 349.700 382.800 350.300 ;
        RECT 356.400 349.600 357.200 349.700 ;
        RECT 370.800 349.600 371.600 349.700 ;
        RECT 382.000 349.600 382.800 349.700 ;
        RECT 415.600 350.300 416.400 350.400 ;
        RECT 425.200 350.300 426.000 350.400 ;
        RECT 415.600 349.700 426.000 350.300 ;
        RECT 415.600 349.600 416.400 349.700 ;
        RECT 425.200 349.600 426.000 349.700 ;
        RECT 466.800 350.300 467.600 350.400 ;
        RECT 478.000 350.300 478.800 350.400 ;
        RECT 466.800 349.700 478.800 350.300 ;
        RECT 466.800 349.600 467.600 349.700 ;
        RECT 478.000 349.600 478.800 349.700 ;
        RECT 510.000 350.300 510.800 350.400 ;
        RECT 526.000 350.300 526.800 350.400 ;
        RECT 510.000 349.700 526.800 350.300 ;
        RECT 527.700 350.300 528.300 351.700 ;
        RECT 538.800 351.700 546.000 352.300 ;
        RECT 538.800 351.600 539.600 351.700 ;
        RECT 545.200 351.600 546.000 351.700 ;
        RECT 546.900 351.700 549.200 352.300 ;
        RECT 546.900 350.300 547.500 351.700 ;
        RECT 548.400 351.600 549.200 351.700 ;
        RECT 551.600 352.300 552.400 352.400 ;
        RECT 558.000 352.300 558.800 352.400 ;
        RECT 551.600 351.700 558.800 352.300 ;
        RECT 551.600 351.600 552.400 351.700 ;
        RECT 558.000 351.600 558.800 351.700 ;
        RECT 562.800 352.300 563.600 352.400 ;
        RECT 572.400 352.300 573.200 352.400 ;
        RECT 562.800 351.700 573.200 352.300 ;
        RECT 562.800 351.600 563.600 351.700 ;
        RECT 572.400 351.600 573.200 351.700 ;
        RECT 578.800 352.300 579.600 352.400 ;
        RECT 585.200 352.300 586.000 352.400 ;
        RECT 578.800 351.700 586.000 352.300 ;
        RECT 578.800 351.600 579.600 351.700 ;
        RECT 585.200 351.600 586.000 351.700 ;
        RECT 620.400 352.300 621.200 352.400 ;
        RECT 634.800 352.300 635.600 352.400 ;
        RECT 620.400 351.700 635.600 352.300 ;
        RECT 620.400 351.600 621.200 351.700 ;
        RECT 634.800 351.600 635.600 351.700 ;
        RECT 646.000 352.300 646.800 352.400 ;
        RECT 660.400 352.300 661.200 352.400 ;
        RECT 646.000 351.700 661.200 352.300 ;
        RECT 646.000 351.600 646.800 351.700 ;
        RECT 660.400 351.600 661.200 351.700 ;
        RECT 527.700 349.700 547.500 350.300 ;
        RECT 548.400 350.300 549.200 350.400 ;
        RECT 551.600 350.300 552.400 350.400 ;
        RECT 548.400 349.700 552.400 350.300 ;
        RECT 510.000 349.600 510.800 349.700 ;
        RECT 526.000 349.600 526.800 349.700 ;
        RECT 548.400 349.600 549.200 349.700 ;
        RECT 551.600 349.600 552.400 349.700 ;
        RECT 556.400 350.300 557.200 350.400 ;
        RECT 586.800 350.300 587.600 350.400 ;
        RECT 556.400 349.700 587.600 350.300 ;
        RECT 556.400 349.600 557.200 349.700 ;
        RECT 586.800 349.600 587.600 349.700 ;
        RECT 599.600 350.300 600.400 350.400 ;
        RECT 614.000 350.300 614.800 350.400 ;
        RECT 599.600 349.700 614.800 350.300 ;
        RECT 599.600 349.600 600.400 349.700 ;
        RECT 614.000 349.600 614.800 349.700 ;
        RECT 623.600 350.300 624.400 350.400 ;
        RECT 647.600 350.300 648.400 350.400 ;
        RECT 660.400 350.300 661.200 350.400 ;
        RECT 623.600 349.700 661.200 350.300 ;
        RECT 623.600 349.600 624.400 349.700 ;
        RECT 647.600 349.600 648.400 349.700 ;
        RECT 660.400 349.600 661.200 349.700 ;
        RECT 7.600 348.300 8.400 348.400 ;
        RECT 26.800 348.300 27.600 348.400 ;
        RECT 7.600 347.700 27.600 348.300 ;
        RECT 7.600 347.600 8.400 347.700 ;
        RECT 26.800 347.600 27.600 347.700 ;
        RECT 34.800 348.300 35.600 348.400 ;
        RECT 62.000 348.300 62.800 348.400 ;
        RECT 34.800 347.700 62.800 348.300 ;
        RECT 34.800 347.600 35.600 347.700 ;
        RECT 62.000 347.600 62.800 347.700 ;
        RECT 73.200 348.300 74.000 348.400 ;
        RECT 105.200 348.300 106.000 348.400 ;
        RECT 142.000 348.300 142.800 348.400 ;
        RECT 153.200 348.300 154.000 348.400 ;
        RECT 161.200 348.300 162.000 348.400 ;
        RECT 73.200 347.700 162.000 348.300 ;
        RECT 73.200 347.600 74.000 347.700 ;
        RECT 105.200 347.600 106.000 347.700 ;
        RECT 142.000 347.600 142.800 347.700 ;
        RECT 153.200 347.600 154.000 347.700 ;
        RECT 161.200 347.600 162.000 347.700 ;
        RECT 225.200 348.300 226.000 348.400 ;
        RECT 230.000 348.300 230.800 348.400 ;
        RECT 225.200 347.700 230.800 348.300 ;
        RECT 225.200 347.600 226.000 347.700 ;
        RECT 230.000 347.600 230.800 347.700 ;
        RECT 238.000 348.300 238.800 348.400 ;
        RECT 254.000 348.300 254.800 348.400 ;
        RECT 238.000 347.700 254.800 348.300 ;
        RECT 238.000 347.600 238.800 347.700 ;
        RECT 254.000 347.600 254.800 347.700 ;
        RECT 297.200 348.300 298.000 348.400 ;
        RECT 303.600 348.300 304.400 348.400 ;
        RECT 311.600 348.300 312.400 348.400 ;
        RECT 297.200 347.700 312.400 348.300 ;
        RECT 297.200 347.600 298.000 347.700 ;
        RECT 303.600 347.600 304.400 347.700 ;
        RECT 311.600 347.600 312.400 347.700 ;
        RECT 313.200 348.300 314.000 348.400 ;
        RECT 319.600 348.300 320.400 348.400 ;
        RECT 313.200 347.700 320.400 348.300 ;
        RECT 313.200 347.600 314.000 347.700 ;
        RECT 319.600 347.600 320.400 347.700 ;
        RECT 321.200 348.300 322.000 348.400 ;
        RECT 324.400 348.300 325.200 348.400 ;
        RECT 337.200 348.300 338.000 348.400 ;
        RECT 366.000 348.300 366.800 348.400 ;
        RECT 367.600 348.300 368.400 348.400 ;
        RECT 375.600 348.300 376.400 348.400 ;
        RECT 386.800 348.300 387.600 348.400 ;
        RECT 321.200 347.700 387.600 348.300 ;
        RECT 321.200 347.600 322.000 347.700 ;
        RECT 324.400 347.600 325.200 347.700 ;
        RECT 337.200 347.600 338.000 347.700 ;
        RECT 366.000 347.600 366.800 347.700 ;
        RECT 367.600 347.600 368.400 347.700 ;
        RECT 375.600 347.600 376.400 347.700 ;
        RECT 386.800 347.600 387.600 347.700 ;
        RECT 406.000 348.300 406.800 348.400 ;
        RECT 414.000 348.300 414.800 348.400 ;
        RECT 406.000 347.700 414.800 348.300 ;
        RECT 406.000 347.600 406.800 347.700 ;
        RECT 414.000 347.600 414.800 347.700 ;
        RECT 430.000 347.600 430.800 348.400 ;
        RECT 471.600 348.300 472.400 348.400 ;
        RECT 476.400 348.300 477.200 348.400 ;
        RECT 478.000 348.300 478.800 348.400 ;
        RECT 490.800 348.300 491.600 348.400 ;
        RECT 471.600 347.700 491.600 348.300 ;
        RECT 471.600 347.600 472.400 347.700 ;
        RECT 476.400 347.600 477.200 347.700 ;
        RECT 478.000 347.600 478.800 347.700 ;
        RECT 490.800 347.600 491.600 347.700 ;
        RECT 495.600 348.300 496.400 348.400 ;
        RECT 503.600 348.300 504.400 348.400 ;
        RECT 495.600 347.700 504.400 348.300 ;
        RECT 495.600 347.600 496.400 347.700 ;
        RECT 503.600 347.600 504.400 347.700 ;
        RECT 527.600 348.300 528.400 348.400 ;
        RECT 534.000 348.300 534.800 348.400 ;
        RECT 527.600 347.700 534.800 348.300 ;
        RECT 527.600 347.600 528.400 347.700 ;
        RECT 534.000 347.600 534.800 347.700 ;
        RECT 553.200 348.300 554.000 348.400 ;
        RECT 562.800 348.300 563.600 348.400 ;
        RECT 553.200 347.700 563.600 348.300 ;
        RECT 553.200 347.600 554.000 347.700 ;
        RECT 562.800 347.600 563.600 347.700 ;
        RECT 582.000 348.300 582.800 348.400 ;
        RECT 610.800 348.300 611.600 348.400 ;
        RECT 582.000 347.700 611.600 348.300 ;
        RECT 582.000 347.600 582.800 347.700 ;
        RECT 610.800 347.600 611.600 347.700 ;
        RECT 622.000 348.300 622.800 348.400 ;
        RECT 633.200 348.300 634.000 348.400 ;
        RECT 641.200 348.300 642.000 348.400 ;
        RECT 662.000 348.300 662.800 348.400 ;
        RECT 622.000 347.700 635.500 348.300 ;
        RECT 622.000 347.600 622.800 347.700 ;
        RECT 633.200 347.600 634.000 347.700 ;
        RECT 25.200 346.300 26.000 346.400 ;
        RECT 33.200 346.300 34.000 346.400 ;
        RECT 71.600 346.300 72.400 346.400 ;
        RECT 25.200 345.700 72.400 346.300 ;
        RECT 25.200 345.600 26.000 345.700 ;
        RECT 33.200 345.600 34.000 345.700 ;
        RECT 71.600 345.600 72.400 345.700 ;
        RECT 87.600 346.300 88.400 346.400 ;
        RECT 113.200 346.300 114.000 346.400 ;
        RECT 129.200 346.300 130.000 346.400 ;
        RECT 87.600 345.700 130.000 346.300 ;
        RECT 87.600 345.600 88.400 345.700 ;
        RECT 113.200 345.600 114.000 345.700 ;
        RECT 129.200 345.600 130.000 345.700 ;
        RECT 132.400 346.300 133.200 346.400 ;
        RECT 138.800 346.300 139.600 346.400 ;
        RECT 132.400 345.700 139.600 346.300 ;
        RECT 132.400 345.600 133.200 345.700 ;
        RECT 138.800 345.600 139.600 345.700 ;
        RECT 140.400 346.300 141.200 346.400 ;
        RECT 162.800 346.300 163.600 346.400 ;
        RECT 140.400 345.700 163.600 346.300 ;
        RECT 140.400 345.600 141.200 345.700 ;
        RECT 162.800 345.600 163.600 345.700 ;
        RECT 220.400 346.300 221.200 346.400 ;
        RECT 270.000 346.300 270.800 346.400 ;
        RECT 220.400 345.700 270.800 346.300 ;
        RECT 220.400 345.600 221.200 345.700 ;
        RECT 270.000 345.600 270.800 345.700 ;
        RECT 308.400 346.300 309.200 346.400 ;
        RECT 319.600 346.300 320.400 346.400 ;
        RECT 308.400 345.700 320.400 346.300 ;
        RECT 308.400 345.600 309.200 345.700 ;
        RECT 319.600 345.600 320.400 345.700 ;
        RECT 329.200 346.300 330.000 346.400 ;
        RECT 340.400 346.300 341.200 346.400 ;
        RECT 329.200 345.700 341.200 346.300 ;
        RECT 329.200 345.600 330.000 345.700 ;
        RECT 340.400 345.600 341.200 345.700 ;
        RECT 342.000 346.300 342.800 346.400 ;
        RECT 348.400 346.300 349.200 346.400 ;
        RECT 342.000 345.700 349.200 346.300 ;
        RECT 342.000 345.600 342.800 345.700 ;
        RECT 348.400 345.600 349.200 345.700 ;
        RECT 364.400 346.300 365.200 346.400 ;
        RECT 366.000 346.300 366.800 346.400 ;
        RECT 364.400 345.700 366.800 346.300 ;
        RECT 364.400 345.600 365.200 345.700 ;
        RECT 366.000 345.600 366.800 345.700 ;
        RECT 385.200 346.300 386.000 346.400 ;
        RECT 406.000 346.300 406.800 346.400 ;
        RECT 385.200 345.700 406.800 346.300 ;
        RECT 385.200 345.600 386.000 345.700 ;
        RECT 406.000 345.600 406.800 345.700 ;
        RECT 426.800 346.300 427.600 346.400 ;
        RECT 431.600 346.300 432.400 346.400 ;
        RECT 426.800 345.700 432.400 346.300 ;
        RECT 426.800 345.600 427.600 345.700 ;
        RECT 431.600 345.600 432.400 345.700 ;
        RECT 457.200 346.300 458.000 346.400 ;
        RECT 476.400 346.300 477.200 346.400 ;
        RECT 457.200 345.700 477.200 346.300 ;
        RECT 457.200 345.600 458.000 345.700 ;
        RECT 476.400 345.600 477.200 345.700 ;
        RECT 486.000 346.300 486.800 346.400 ;
        RECT 490.800 346.300 491.600 346.400 ;
        RECT 486.000 345.700 491.600 346.300 ;
        RECT 486.000 345.600 486.800 345.700 ;
        RECT 490.800 345.600 491.600 345.700 ;
        RECT 494.000 346.300 494.800 346.400 ;
        RECT 510.000 346.300 510.800 346.400 ;
        RECT 494.000 345.700 510.800 346.300 ;
        RECT 494.000 345.600 494.800 345.700 ;
        RECT 510.000 345.600 510.800 345.700 ;
        RECT 511.600 346.300 512.400 346.400 ;
        RECT 521.200 346.300 522.000 346.400 ;
        RECT 511.600 345.700 522.000 346.300 ;
        RECT 511.600 345.600 512.400 345.700 ;
        RECT 521.200 345.600 522.000 345.700 ;
        RECT 522.800 346.300 523.600 346.400 ;
        RECT 530.800 346.300 531.600 346.400 ;
        RECT 522.800 345.700 531.600 346.300 ;
        RECT 522.800 345.600 523.600 345.700 ;
        RECT 530.800 345.600 531.600 345.700 ;
        RECT 538.800 346.300 539.600 346.400 ;
        RECT 574.000 346.300 574.800 346.400 ;
        RECT 583.600 346.300 584.400 346.400 ;
        RECT 538.800 345.700 584.400 346.300 ;
        RECT 538.800 345.600 539.600 345.700 ;
        RECT 574.000 345.600 574.800 345.700 ;
        RECT 583.600 345.600 584.400 345.700 ;
        RECT 609.200 346.300 610.000 346.400 ;
        RECT 617.200 346.300 618.000 346.400 ;
        RECT 625.200 346.300 626.000 346.400 ;
        RECT 609.200 345.700 626.000 346.300 ;
        RECT 609.200 345.600 610.000 345.700 ;
        RECT 617.200 345.600 618.000 345.700 ;
        RECT 625.200 345.600 626.000 345.700 ;
        RECT 631.600 346.300 632.400 346.400 ;
        RECT 633.200 346.300 634.000 346.400 ;
        RECT 631.600 345.700 634.000 346.300 ;
        RECT 634.900 346.300 635.500 347.700 ;
        RECT 641.200 347.700 662.800 348.300 ;
        RECT 641.200 347.600 642.000 347.700 ;
        RECT 662.000 347.600 662.800 347.700 ;
        RECT 663.600 348.300 664.400 348.400 ;
        RECT 666.800 348.300 667.600 348.400 ;
        RECT 663.600 347.700 667.600 348.300 ;
        RECT 663.600 347.600 664.400 347.700 ;
        RECT 666.800 347.600 667.600 347.700 ;
        RECT 647.600 346.300 648.400 346.400 ;
        RECT 634.900 345.700 648.400 346.300 ;
        RECT 631.600 345.600 632.400 345.700 ;
        RECT 633.200 345.600 634.000 345.700 ;
        RECT 647.600 345.600 648.400 345.700 ;
        RECT 660.400 346.300 661.200 346.400 ;
        RECT 673.200 346.300 674.000 346.400 ;
        RECT 660.400 345.700 674.000 346.300 ;
        RECT 660.400 345.600 661.200 345.700 ;
        RECT 673.200 345.600 674.000 345.700 ;
        RECT 31.600 344.300 32.400 344.400 ;
        RECT 36.400 344.300 37.200 344.400 ;
        RECT 44.400 344.300 45.200 344.400 ;
        RECT 76.400 344.300 77.200 344.400 ;
        RECT 97.200 344.300 98.000 344.400 ;
        RECT 102.000 344.300 102.800 344.400 ;
        RECT 31.600 343.700 102.800 344.300 ;
        RECT 31.600 343.600 32.400 343.700 ;
        RECT 36.400 343.600 37.200 343.700 ;
        RECT 44.400 343.600 45.200 343.700 ;
        RECT 76.400 343.600 77.200 343.700 ;
        RECT 97.200 343.600 98.000 343.700 ;
        RECT 102.000 343.600 102.800 343.700 ;
        RECT 103.600 344.300 104.400 344.400 ;
        RECT 122.800 344.300 123.600 344.400 ;
        RECT 103.600 343.700 123.600 344.300 ;
        RECT 103.600 343.600 104.400 343.700 ;
        RECT 122.800 343.600 123.600 343.700 ;
        RECT 135.600 344.300 136.400 344.400 ;
        RECT 142.000 344.300 142.800 344.400 ;
        RECT 135.600 343.700 142.800 344.300 ;
        RECT 135.600 343.600 136.400 343.700 ;
        RECT 142.000 343.600 142.800 343.700 ;
        RECT 183.600 344.300 184.400 344.400 ;
        RECT 209.200 344.300 210.000 344.400 ;
        RECT 183.600 343.700 210.000 344.300 ;
        RECT 183.600 343.600 184.400 343.700 ;
        RECT 209.200 343.600 210.000 343.700 ;
        RECT 322.800 344.300 323.600 344.400 ;
        RECT 330.800 344.300 331.600 344.400 ;
        RECT 322.800 343.700 331.600 344.300 ;
        RECT 322.800 343.600 323.600 343.700 ;
        RECT 330.800 343.600 331.600 343.700 ;
        RECT 334.000 344.300 334.800 344.400 ;
        RECT 346.800 344.300 347.600 344.400 ;
        RECT 334.000 343.700 347.600 344.300 ;
        RECT 334.000 343.600 334.800 343.700 ;
        RECT 346.800 343.600 347.600 343.700 ;
        RECT 358.000 344.300 358.800 344.400 ;
        RECT 366.000 344.300 366.800 344.400 ;
        RECT 358.000 343.700 366.800 344.300 ;
        RECT 358.000 343.600 358.800 343.700 ;
        RECT 366.000 343.600 366.800 343.700 ;
        RECT 369.200 344.300 370.000 344.400 ;
        RECT 433.200 344.300 434.000 344.400 ;
        RECT 438.000 344.300 438.800 344.400 ;
        RECT 369.200 343.700 438.800 344.300 ;
        RECT 369.200 343.600 370.000 343.700 ;
        RECT 433.200 343.600 434.000 343.700 ;
        RECT 438.000 343.600 438.800 343.700 ;
        RECT 482.800 344.300 483.600 344.400 ;
        RECT 511.600 344.300 512.400 344.400 ;
        RECT 482.800 343.700 512.400 344.300 ;
        RECT 482.800 343.600 483.600 343.700 ;
        RECT 511.600 343.600 512.400 343.700 ;
        RECT 522.800 344.300 523.600 344.400 ;
        RECT 540.400 344.300 541.200 344.400 ;
        RECT 522.800 343.700 541.200 344.300 ;
        RECT 522.800 343.600 523.600 343.700 ;
        RECT 540.400 343.600 541.200 343.700 ;
        RECT 543.600 344.300 544.400 344.400 ;
        RECT 558.000 344.300 558.800 344.400 ;
        RECT 543.600 343.700 558.800 344.300 ;
        RECT 543.600 343.600 544.400 343.700 ;
        RECT 558.000 343.600 558.800 343.700 ;
        RECT 559.600 344.300 560.400 344.400 ;
        RECT 566.000 344.300 566.800 344.400 ;
        RECT 588.400 344.300 589.200 344.400 ;
        RECT 559.600 343.700 589.200 344.300 ;
        RECT 559.600 343.600 560.400 343.700 ;
        RECT 566.000 343.600 566.800 343.700 ;
        RECT 588.400 343.600 589.200 343.700 ;
        RECT 612.400 344.300 613.200 344.400 ;
        RECT 626.800 344.300 627.600 344.400 ;
        RECT 612.400 343.700 627.600 344.300 ;
        RECT 612.400 343.600 613.200 343.700 ;
        RECT 626.800 343.600 627.600 343.700 ;
        RECT 654.000 344.300 654.800 344.400 ;
        RECT 679.600 344.300 680.400 344.400 ;
        RECT 654.000 343.700 680.400 344.300 ;
        RECT 654.000 343.600 654.800 343.700 ;
        RECT 679.600 343.600 680.400 343.700 ;
        RECT 66.800 342.300 67.600 342.400 ;
        RECT 82.800 342.300 83.600 342.400 ;
        RECT 66.800 341.700 83.600 342.300 ;
        RECT 66.800 341.600 67.600 341.700 ;
        RECT 82.800 341.600 83.600 341.700 ;
        RECT 94.000 342.300 94.800 342.400 ;
        RECT 146.800 342.300 147.600 342.400 ;
        RECT 158.000 342.300 158.800 342.400 ;
        RECT 94.000 341.700 158.800 342.300 ;
        RECT 94.000 341.600 94.800 341.700 ;
        RECT 146.800 341.600 147.600 341.700 ;
        RECT 158.000 341.600 158.800 341.700 ;
        RECT 159.600 342.300 160.400 342.400 ;
        RECT 188.400 342.300 189.200 342.400 ;
        RECT 159.600 341.700 189.200 342.300 ;
        RECT 159.600 341.600 160.400 341.700 ;
        RECT 188.400 341.600 189.200 341.700 ;
        RECT 318.000 342.300 318.800 342.400 ;
        RECT 329.200 342.300 330.000 342.400 ;
        RECT 338.800 342.300 339.600 342.400 ;
        RECT 369.300 342.300 369.900 343.600 ;
        RECT 318.000 341.700 369.900 342.300 ;
        RECT 497.200 342.300 498.000 342.400 ;
        RECT 538.800 342.300 539.600 342.400 ;
        RECT 497.200 341.700 539.600 342.300 ;
        RECT 318.000 341.600 318.800 341.700 ;
        RECT 329.200 341.600 330.000 341.700 ;
        RECT 338.800 341.600 339.600 341.700 ;
        RECT 497.200 341.600 498.000 341.700 ;
        RECT 538.800 341.600 539.600 341.700 ;
        RECT 545.200 342.300 546.000 342.400 ;
        RECT 556.400 342.300 557.200 342.400 ;
        RECT 545.200 341.700 557.200 342.300 ;
        RECT 545.200 341.600 546.000 341.700 ;
        RECT 556.400 341.600 557.200 341.700 ;
        RECT 598.000 342.300 598.800 342.400 ;
        RECT 631.600 342.300 632.400 342.400 ;
        RECT 598.000 341.700 632.400 342.300 ;
        RECT 598.000 341.600 598.800 341.700 ;
        RECT 631.600 341.600 632.400 341.700 ;
        RECT 638.000 342.300 638.800 342.400 ;
        RECT 676.400 342.300 677.200 342.400 ;
        RECT 638.000 341.700 677.200 342.300 ;
        RECT 638.000 341.600 638.800 341.700 ;
        RECT 676.400 341.600 677.200 341.700 ;
        RECT 55.600 340.300 56.400 340.400 ;
        RECT 60.400 340.300 61.200 340.400 ;
        RECT 55.600 339.700 61.200 340.300 ;
        RECT 55.600 339.600 56.400 339.700 ;
        RECT 60.400 339.600 61.200 339.700 ;
        RECT 90.800 340.300 91.600 340.400 ;
        RECT 206.000 340.300 206.800 340.400 ;
        RECT 90.800 339.700 206.800 340.300 ;
        RECT 90.800 339.600 91.600 339.700 ;
        RECT 206.000 339.600 206.800 339.700 ;
        RECT 222.000 340.300 222.800 340.400 ;
        RECT 226.800 340.300 227.600 340.400 ;
        RECT 222.000 339.700 227.600 340.300 ;
        RECT 222.000 339.600 222.800 339.700 ;
        RECT 226.800 339.600 227.600 339.700 ;
        RECT 308.400 340.300 309.200 340.400 ;
        RECT 321.200 340.300 322.000 340.400 ;
        RECT 308.400 339.700 322.000 340.300 ;
        RECT 308.400 339.600 309.200 339.700 ;
        RECT 321.200 339.600 322.000 339.700 ;
        RECT 326.000 340.300 326.800 340.400 ;
        RECT 337.200 340.300 338.000 340.400 ;
        RECT 345.200 340.300 346.000 340.400 ;
        RECT 364.400 340.300 365.200 340.400 ;
        RECT 326.000 339.700 346.000 340.300 ;
        RECT 326.000 339.600 326.800 339.700 ;
        RECT 337.200 339.600 338.000 339.700 ;
        RECT 345.200 339.600 346.000 339.700 ;
        RECT 346.900 339.700 365.200 340.300 ;
        RECT 41.200 338.300 42.000 338.400 ;
        RECT 54.000 338.300 54.800 338.400 ;
        RECT 41.200 337.700 54.800 338.300 ;
        RECT 41.200 337.600 42.000 337.700 ;
        RECT 54.000 337.600 54.800 337.700 ;
        RECT 82.800 338.300 83.600 338.400 ;
        RECT 90.800 338.300 91.600 338.400 ;
        RECT 82.800 337.700 91.600 338.300 ;
        RECT 82.800 337.600 83.600 337.700 ;
        RECT 90.800 337.600 91.600 337.700 ;
        RECT 92.400 338.300 93.200 338.400 ;
        RECT 94.000 338.300 94.800 338.400 ;
        RECT 92.400 337.700 94.800 338.300 ;
        RECT 92.400 337.600 93.200 337.700 ;
        RECT 94.000 337.600 94.800 337.700 ;
        RECT 121.200 338.300 122.000 338.400 ;
        RECT 127.600 338.300 128.400 338.400 ;
        RECT 121.200 337.700 128.400 338.300 ;
        RECT 121.200 337.600 122.000 337.700 ;
        RECT 127.600 337.600 128.400 337.700 ;
        RECT 150.000 338.300 150.800 338.400 ;
        RECT 154.800 338.300 155.600 338.400 ;
        RECT 150.000 337.700 155.600 338.300 ;
        RECT 150.000 337.600 150.800 337.700 ;
        RECT 154.800 337.600 155.600 337.700 ;
        RECT 167.600 338.300 168.400 338.400 ;
        RECT 226.800 338.300 227.600 338.400 ;
        RECT 241.200 338.300 242.000 338.400 ;
        RECT 167.600 337.700 242.000 338.300 ;
        RECT 167.600 337.600 168.400 337.700 ;
        RECT 226.800 337.600 227.600 337.700 ;
        RECT 241.200 337.600 242.000 337.700 ;
        RECT 318.000 338.300 318.800 338.400 ;
        RECT 332.400 338.300 333.200 338.400 ;
        RECT 346.900 338.300 347.500 339.700 ;
        RECT 364.400 339.600 365.200 339.700 ;
        RECT 374.000 340.300 374.800 340.400 ;
        RECT 383.600 340.300 384.400 340.400 ;
        RECT 374.000 339.700 384.400 340.300 ;
        RECT 374.000 339.600 374.800 339.700 ;
        RECT 383.600 339.600 384.400 339.700 ;
        RECT 538.800 339.600 539.600 340.400 ;
        RECT 599.600 340.300 600.400 340.400 ;
        RECT 607.600 340.300 608.400 340.400 ;
        RECT 599.600 339.700 608.400 340.300 ;
        RECT 599.600 339.600 600.400 339.700 ;
        RECT 607.600 339.600 608.400 339.700 ;
        RECT 634.800 340.300 635.600 340.400 ;
        RECT 649.200 340.300 650.000 340.400 ;
        RECT 634.800 339.700 650.000 340.300 ;
        RECT 634.800 339.600 635.600 339.700 ;
        RECT 649.200 339.600 650.000 339.700 ;
        RECT 318.000 337.700 333.200 338.300 ;
        RECT 318.000 337.600 318.800 337.700 ;
        RECT 332.400 337.600 333.200 337.700 ;
        RECT 334.100 337.700 347.500 338.300 ;
        RECT 354.800 338.300 355.600 338.400 ;
        RECT 377.200 338.300 378.000 338.400 ;
        RECT 398.000 338.300 398.800 338.400 ;
        RECT 422.000 338.300 422.800 338.400 ;
        RECT 354.800 337.700 422.800 338.300 ;
        RECT 49.200 336.300 50.000 336.400 ;
        RECT 68.400 336.300 69.200 336.400 ;
        RECT 49.200 335.700 69.200 336.300 ;
        RECT 49.200 335.600 50.000 335.700 ;
        RECT 68.400 335.600 69.200 335.700 ;
        RECT 70.000 336.300 70.800 336.400 ;
        RECT 98.800 336.300 99.600 336.400 ;
        RECT 70.000 335.700 99.600 336.300 ;
        RECT 70.000 335.600 70.800 335.700 ;
        RECT 98.800 335.600 99.600 335.700 ;
        RECT 103.600 336.300 104.400 336.400 ;
        RECT 108.400 336.300 109.200 336.400 ;
        RECT 142.000 336.300 142.800 336.400 ;
        RECT 167.600 336.300 168.400 336.400 ;
        RECT 103.600 335.700 168.400 336.300 ;
        RECT 103.600 335.600 104.400 335.700 ;
        RECT 108.400 335.600 109.200 335.700 ;
        RECT 142.000 335.600 142.800 335.700 ;
        RECT 167.600 335.600 168.400 335.700 ;
        RECT 223.600 336.300 224.400 336.400 ;
        RECT 228.400 336.300 229.200 336.400 ;
        RECT 223.600 335.700 229.200 336.300 ;
        RECT 223.600 335.600 224.400 335.700 ;
        RECT 228.400 335.600 229.200 335.700 ;
        RECT 316.400 336.300 317.200 336.400 ;
        RECT 334.100 336.300 334.700 337.700 ;
        RECT 354.800 337.600 355.600 337.700 ;
        RECT 377.200 337.600 378.000 337.700 ;
        RECT 398.000 337.600 398.800 337.700 ;
        RECT 422.000 337.600 422.800 337.700 ;
        RECT 455.600 338.300 456.400 338.400 ;
        RECT 471.600 338.300 472.400 338.400 ;
        RECT 455.600 337.700 472.400 338.300 ;
        RECT 455.600 337.600 456.400 337.700 ;
        RECT 471.600 337.600 472.400 337.700 ;
        RECT 478.000 338.300 478.800 338.400 ;
        RECT 609.200 338.300 610.000 338.400 ;
        RECT 478.000 337.700 610.000 338.300 ;
        RECT 478.000 337.600 478.800 337.700 ;
        RECT 609.200 337.600 610.000 337.700 ;
        RECT 636.400 338.300 637.200 338.400 ;
        RECT 652.400 338.300 653.200 338.400 ;
        RECT 636.400 337.700 653.200 338.300 ;
        RECT 636.400 337.600 637.200 337.700 ;
        RECT 652.400 337.600 653.200 337.700 ;
        RECT 316.400 335.700 334.700 336.300 ;
        RECT 340.400 336.300 341.200 336.400 ;
        RECT 351.600 336.300 352.400 336.400 ;
        RECT 372.400 336.300 373.200 336.400 ;
        RECT 391.600 336.300 392.400 336.400 ;
        RECT 399.600 336.300 400.400 336.400 ;
        RECT 340.400 335.700 400.400 336.300 ;
        RECT 316.400 335.600 317.200 335.700 ;
        RECT 340.400 335.600 341.200 335.700 ;
        RECT 351.600 335.600 352.400 335.700 ;
        RECT 372.400 335.600 373.200 335.700 ;
        RECT 391.600 335.600 392.400 335.700 ;
        RECT 399.600 335.600 400.400 335.700 ;
        RECT 407.600 336.300 408.400 336.400 ;
        RECT 412.400 336.300 413.200 336.400 ;
        RECT 407.600 335.700 413.200 336.300 ;
        RECT 407.600 335.600 408.400 335.700 ;
        RECT 412.400 335.600 413.200 335.700 ;
        RECT 426.800 336.300 427.600 336.400 ;
        RECT 470.000 336.300 470.800 336.400 ;
        RECT 426.800 335.700 470.800 336.300 ;
        RECT 426.800 335.600 427.600 335.700 ;
        RECT 470.000 335.600 470.800 335.700 ;
        RECT 476.400 336.300 477.200 336.400 ;
        RECT 481.200 336.300 482.000 336.400 ;
        RECT 556.400 336.300 557.200 336.400 ;
        RECT 476.400 335.700 557.200 336.300 ;
        RECT 476.400 335.600 477.200 335.700 ;
        RECT 481.200 335.600 482.000 335.700 ;
        RECT 556.400 335.600 557.200 335.700 ;
        RECT 558.000 336.300 558.800 336.400 ;
        RECT 590.000 336.300 590.800 336.400 ;
        RECT 558.000 335.700 590.800 336.300 ;
        RECT 558.000 335.600 558.800 335.700 ;
        RECT 590.000 335.600 590.800 335.700 ;
        RECT 593.200 336.300 594.000 336.400 ;
        RECT 620.400 336.300 621.200 336.400 ;
        RECT 593.200 335.700 621.200 336.300 ;
        RECT 593.200 335.600 594.000 335.700 ;
        RECT 620.400 335.600 621.200 335.700 ;
        RECT 622.000 336.300 622.800 336.400 ;
        RECT 634.800 336.300 635.600 336.400 ;
        RECT 622.000 335.700 635.600 336.300 ;
        RECT 622.000 335.600 622.800 335.700 ;
        RECT 634.800 335.600 635.600 335.700 ;
        RECT 638.000 336.300 638.800 336.400 ;
        RECT 642.800 336.300 643.600 336.400 ;
        RECT 638.000 335.700 643.600 336.300 ;
        RECT 638.000 335.600 638.800 335.700 ;
        RECT 642.800 335.600 643.600 335.700 ;
        RECT 663.600 336.300 664.400 336.400 ;
        RECT 671.600 336.300 672.400 336.400 ;
        RECT 663.600 335.700 672.400 336.300 ;
        RECT 663.600 335.600 664.400 335.700 ;
        RECT 671.600 335.600 672.400 335.700 ;
        RECT 39.600 334.300 40.400 334.400 ;
        RECT 47.600 334.300 48.400 334.400 ;
        RECT 39.600 333.700 48.400 334.300 ;
        RECT 39.600 333.600 40.400 333.700 ;
        RECT 47.600 333.600 48.400 333.700 ;
        RECT 54.000 334.300 54.800 334.400 ;
        RECT 71.600 334.300 72.400 334.400 ;
        RECT 54.000 333.700 72.400 334.300 ;
        RECT 54.000 333.600 54.800 333.700 ;
        RECT 71.600 333.600 72.400 333.700 ;
        RECT 79.600 334.300 80.400 334.400 ;
        RECT 92.400 334.300 93.200 334.400 ;
        RECT 79.600 333.700 93.200 334.300 ;
        RECT 79.600 333.600 80.400 333.700 ;
        RECT 92.400 333.600 93.200 333.700 ;
        RECT 134.000 334.300 134.800 334.400 ;
        RECT 153.200 334.300 154.000 334.400 ;
        RECT 134.000 333.700 154.000 334.300 ;
        RECT 134.000 333.600 134.800 333.700 ;
        RECT 153.200 333.600 154.000 333.700 ;
        RECT 154.800 334.300 155.600 334.400 ;
        RECT 161.200 334.300 162.000 334.400 ;
        RECT 154.800 333.700 162.000 334.300 ;
        RECT 154.800 333.600 155.600 333.700 ;
        RECT 161.200 333.600 162.000 333.700 ;
        RECT 217.200 334.300 218.000 334.400 ;
        RECT 250.800 334.300 251.600 334.400 ;
        RECT 217.200 333.700 251.600 334.300 ;
        RECT 217.200 333.600 218.000 333.700 ;
        RECT 250.800 333.600 251.600 333.700 ;
        RECT 282.800 334.300 283.600 334.400 ;
        RECT 303.600 334.300 304.400 334.400 ;
        RECT 282.800 333.700 304.400 334.300 ;
        RECT 282.800 333.600 283.600 333.700 ;
        RECT 303.600 333.600 304.400 333.700 ;
        RECT 319.600 334.300 320.400 334.400 ;
        RECT 324.400 334.300 325.200 334.400 ;
        RECT 319.600 333.700 325.200 334.300 ;
        RECT 319.600 333.600 320.400 333.700 ;
        RECT 324.400 333.600 325.200 333.700 ;
        RECT 330.800 334.300 331.600 334.400 ;
        RECT 332.400 334.300 333.200 334.400 ;
        RECT 346.800 334.300 347.600 334.400 ;
        RECT 348.400 334.300 349.200 334.400 ;
        RECT 359.600 334.300 360.400 334.400 ;
        RECT 380.400 334.300 381.200 334.400 ;
        RECT 396.400 334.300 397.200 334.400 ;
        RECT 401.200 334.300 402.000 334.400 ;
        RECT 330.800 333.700 395.500 334.300 ;
        RECT 330.800 333.600 331.600 333.700 ;
        RECT 332.400 333.600 333.200 333.700 ;
        RECT 346.800 333.600 347.600 333.700 ;
        RECT 348.400 333.600 349.200 333.700 ;
        RECT 359.600 333.600 360.400 333.700 ;
        RECT 380.400 333.600 381.200 333.700 ;
        RECT 7.600 332.300 8.400 332.400 ;
        RECT 25.200 332.300 26.000 332.400 ;
        RECT 7.600 331.700 26.000 332.300 ;
        RECT 7.600 331.600 8.400 331.700 ;
        RECT 25.200 331.600 26.000 331.700 ;
        RECT 30.000 332.300 30.800 332.400 ;
        RECT 33.200 332.300 34.000 332.400 ;
        RECT 30.000 331.700 34.000 332.300 ;
        RECT 30.000 331.600 30.800 331.700 ;
        RECT 33.200 331.600 34.000 331.700 ;
        RECT 39.600 332.300 40.400 332.400 ;
        RECT 62.000 332.300 62.800 332.400 ;
        RECT 39.600 331.700 62.800 332.300 ;
        RECT 39.600 331.600 40.400 331.700 ;
        RECT 62.000 331.600 62.800 331.700 ;
        RECT 111.600 332.300 112.400 332.400 ;
        RECT 114.800 332.300 115.600 332.400 ;
        RECT 111.600 331.700 115.600 332.300 ;
        RECT 111.600 331.600 112.400 331.700 ;
        RECT 114.800 331.600 115.600 331.700 ;
        RECT 140.400 332.300 141.200 332.400 ;
        RECT 151.600 332.300 152.400 332.400 ;
        RECT 159.600 332.300 160.400 332.400 ;
        RECT 166.000 332.300 166.800 332.400 ;
        RECT 140.400 331.700 166.800 332.300 ;
        RECT 140.400 331.600 141.200 331.700 ;
        RECT 151.600 331.600 152.400 331.700 ;
        RECT 159.600 331.600 160.400 331.700 ;
        RECT 166.000 331.600 166.800 331.700 ;
        RECT 209.200 332.300 210.000 332.400 ;
        RECT 212.400 332.300 213.200 332.400 ;
        RECT 209.200 331.700 213.200 332.300 ;
        RECT 209.200 331.600 210.000 331.700 ;
        RECT 212.400 331.600 213.200 331.700 ;
        RECT 234.800 332.300 235.600 332.400 ;
        RECT 239.600 332.300 240.400 332.400 ;
        RECT 234.800 331.700 240.400 332.300 ;
        RECT 234.800 331.600 235.600 331.700 ;
        RECT 239.600 331.600 240.400 331.700 ;
        RECT 306.800 332.300 307.600 332.400 ;
        RECT 314.800 332.300 315.600 332.400 ;
        RECT 322.800 332.300 323.600 332.400 ;
        RECT 306.800 331.700 315.600 332.300 ;
        RECT 306.800 331.600 307.600 331.700 ;
        RECT 314.800 331.600 315.600 331.700 ;
        RECT 321.300 331.700 323.600 332.300 ;
        RECT 7.600 330.300 8.400 330.400 ;
        RECT 10.800 330.300 11.600 330.400 ;
        RECT 7.600 329.700 11.600 330.300 ;
        RECT 7.600 329.600 8.400 329.700 ;
        RECT 10.800 329.600 11.600 329.700 ;
        RECT 12.400 330.300 13.200 330.400 ;
        RECT 17.200 330.300 18.000 330.400 ;
        RECT 12.400 329.700 18.000 330.300 ;
        RECT 12.400 329.600 13.200 329.700 ;
        RECT 17.200 329.600 18.000 329.700 ;
        RECT 20.400 330.300 21.200 330.400 ;
        RECT 39.600 330.300 40.400 330.400 ;
        RECT 20.400 329.700 40.400 330.300 ;
        RECT 20.400 329.600 21.200 329.700 ;
        RECT 39.600 329.600 40.400 329.700 ;
        RECT 58.800 330.300 59.600 330.400 ;
        RECT 65.200 330.300 66.000 330.400 ;
        RECT 58.800 329.700 66.000 330.300 ;
        RECT 58.800 329.600 59.600 329.700 ;
        RECT 65.200 329.600 66.000 329.700 ;
        RECT 84.400 330.300 85.200 330.400 ;
        RECT 118.000 330.300 118.800 330.400 ;
        RECT 84.400 329.700 118.800 330.300 ;
        RECT 84.400 329.600 85.200 329.700 ;
        RECT 118.000 329.600 118.800 329.700 ;
        RECT 159.600 330.300 160.400 330.400 ;
        RECT 167.600 330.300 168.400 330.400 ;
        RECT 159.600 329.700 168.400 330.300 ;
        RECT 159.600 329.600 160.400 329.700 ;
        RECT 167.600 329.600 168.400 329.700 ;
        RECT 198.000 330.300 198.800 330.400 ;
        RECT 212.400 330.300 213.200 330.400 ;
        RECT 257.200 330.300 258.000 330.400 ;
        RECT 198.000 329.700 258.000 330.300 ;
        RECT 198.000 329.600 198.800 329.700 ;
        RECT 212.400 329.600 213.200 329.700 ;
        RECT 257.200 329.600 258.000 329.700 ;
        RECT 308.400 330.300 309.200 330.400 ;
        RECT 321.300 330.300 321.900 331.700 ;
        RECT 322.800 331.600 323.600 331.700 ;
        RECT 327.600 332.300 328.400 332.400 ;
        RECT 335.600 332.300 336.400 332.400 ;
        RECT 345.200 332.300 346.000 332.400 ;
        RECT 356.400 332.300 357.200 332.400 ;
        RECT 362.800 332.300 363.600 332.400 ;
        RECT 378.800 332.300 379.600 332.400 ;
        RECT 390.000 332.300 390.800 332.400 ;
        RECT 327.600 331.700 390.800 332.300 ;
        RECT 394.900 332.300 395.500 333.700 ;
        RECT 396.400 333.700 402.000 334.300 ;
        RECT 396.400 333.600 397.200 333.700 ;
        RECT 401.200 333.600 402.000 333.700 ;
        RECT 410.800 334.300 411.600 334.400 ;
        RECT 422.000 334.300 422.800 334.400 ;
        RECT 428.400 334.300 429.200 334.400 ;
        RECT 410.800 333.700 429.200 334.300 ;
        RECT 410.800 333.600 411.600 333.700 ;
        RECT 422.000 333.600 422.800 333.700 ;
        RECT 428.400 333.600 429.200 333.700 ;
        RECT 434.800 334.300 435.600 334.400 ;
        RECT 474.800 334.300 475.600 334.400 ;
        RECT 434.800 333.700 475.600 334.300 ;
        RECT 434.800 333.600 435.600 333.700 ;
        RECT 474.800 333.600 475.600 333.700 ;
        RECT 516.400 334.300 517.200 334.400 ;
        RECT 521.200 334.300 522.000 334.400 ;
        RECT 516.400 333.700 522.000 334.300 ;
        RECT 516.400 333.600 517.200 333.700 ;
        RECT 521.200 333.600 522.000 333.700 ;
        RECT 522.800 334.300 523.600 334.400 ;
        RECT 540.400 334.300 541.200 334.400 ;
        RECT 522.800 333.700 541.200 334.300 ;
        RECT 522.800 333.600 523.600 333.700 ;
        RECT 540.400 333.600 541.200 333.700 ;
        RECT 545.200 334.300 546.000 334.400 ;
        RECT 553.200 334.300 554.000 334.400 ;
        RECT 545.200 333.700 554.000 334.300 ;
        RECT 545.200 333.600 546.000 333.700 ;
        RECT 553.200 333.600 554.000 333.700 ;
        RECT 614.000 334.300 614.800 334.400 ;
        RECT 625.200 334.300 626.000 334.400 ;
        RECT 614.000 333.700 626.000 334.300 ;
        RECT 614.000 333.600 614.800 333.700 ;
        RECT 625.200 333.600 626.000 333.700 ;
        RECT 626.800 334.300 627.600 334.400 ;
        RECT 644.400 334.300 645.200 334.400 ;
        RECT 654.000 334.300 654.800 334.400 ;
        RECT 626.800 333.700 654.800 334.300 ;
        RECT 626.800 333.600 627.600 333.700 ;
        RECT 644.400 333.600 645.200 333.700 ;
        RECT 654.000 333.600 654.800 333.700 ;
        RECT 666.800 334.300 667.600 334.400 ;
        RECT 671.600 334.300 672.400 334.400 ;
        RECT 666.800 333.700 672.400 334.300 ;
        RECT 666.800 333.600 667.600 333.700 ;
        RECT 671.600 333.600 672.400 333.700 ;
        RECT 402.800 332.300 403.600 332.400 ;
        RECT 394.900 331.700 403.600 332.300 ;
        RECT 327.600 331.600 328.400 331.700 ;
        RECT 335.600 331.600 336.400 331.700 ;
        RECT 345.200 331.600 346.000 331.700 ;
        RECT 356.400 331.600 357.200 331.700 ;
        RECT 362.800 331.600 363.600 331.700 ;
        RECT 378.800 331.600 379.600 331.700 ;
        RECT 390.000 331.600 390.800 331.700 ;
        RECT 402.800 331.600 403.600 331.700 ;
        RECT 409.200 332.300 410.000 332.400 ;
        RECT 423.600 332.300 424.400 332.400 ;
        RECT 430.000 332.300 430.800 332.400 ;
        RECT 409.200 331.700 430.800 332.300 ;
        RECT 409.200 331.600 410.000 331.700 ;
        RECT 423.600 331.600 424.400 331.700 ;
        RECT 430.000 331.600 430.800 331.700 ;
        RECT 481.200 332.300 482.000 332.400 ;
        RECT 497.200 332.300 498.000 332.400 ;
        RECT 481.200 331.700 498.000 332.300 ;
        RECT 481.200 331.600 482.000 331.700 ;
        RECT 497.200 331.600 498.000 331.700 ;
        RECT 502.000 332.300 502.800 332.400 ;
        RECT 506.800 332.300 507.600 332.400 ;
        RECT 502.000 331.700 507.600 332.300 ;
        RECT 502.000 331.600 502.800 331.700 ;
        RECT 506.800 331.600 507.600 331.700 ;
        RECT 514.800 332.300 515.600 332.400 ;
        RECT 522.800 332.300 523.600 332.400 ;
        RECT 530.800 332.300 531.600 332.400 ;
        RECT 514.800 331.700 531.600 332.300 ;
        RECT 514.800 331.600 515.600 331.700 ;
        RECT 522.800 331.600 523.600 331.700 ;
        RECT 530.800 331.600 531.600 331.700 ;
        RECT 535.600 332.300 536.400 332.400 ;
        RECT 548.400 332.300 549.200 332.400 ;
        RECT 535.600 331.700 549.200 332.300 ;
        RECT 535.600 331.600 536.400 331.700 ;
        RECT 548.400 331.600 549.200 331.700 ;
        RECT 572.400 332.300 573.200 332.400 ;
        RECT 586.800 332.300 587.600 332.400 ;
        RECT 572.400 331.700 587.600 332.300 ;
        RECT 572.400 331.600 573.200 331.700 ;
        RECT 586.800 331.600 587.600 331.700 ;
        RECT 633.200 332.300 634.000 332.400 ;
        RECT 636.400 332.300 637.200 332.400 ;
        RECT 633.200 331.700 637.200 332.300 ;
        RECT 633.200 331.600 634.000 331.700 ;
        RECT 636.400 331.600 637.200 331.700 ;
        RECT 644.400 332.300 645.200 332.400 ;
        RECT 655.600 332.300 656.400 332.400 ;
        RECT 644.400 331.700 656.400 332.300 ;
        RECT 644.400 331.600 645.200 331.700 ;
        RECT 655.600 331.600 656.400 331.700 ;
        RECT 657.200 332.300 658.000 332.400 ;
        RECT 666.800 332.300 667.600 332.400 ;
        RECT 657.200 331.700 667.600 332.300 ;
        RECT 657.200 331.600 658.000 331.700 ;
        RECT 666.800 331.600 667.600 331.700 ;
        RECT 308.400 329.700 321.900 330.300 ;
        RECT 322.800 330.300 323.600 330.400 ;
        RECT 337.200 330.300 338.000 330.400 ;
        RECT 322.800 329.700 338.000 330.300 ;
        RECT 308.400 329.600 309.200 329.700 ;
        RECT 322.800 329.600 323.600 329.700 ;
        RECT 337.200 329.600 338.000 329.700 ;
        RECT 356.400 330.300 357.200 330.400 ;
        RECT 361.200 330.300 362.000 330.400 ;
        RECT 356.400 329.700 362.000 330.300 ;
        RECT 356.400 329.600 357.200 329.700 ;
        RECT 361.200 329.600 362.000 329.700 ;
        RECT 367.600 330.300 368.400 330.400 ;
        RECT 375.600 330.300 376.400 330.400 ;
        RECT 367.600 329.700 376.400 330.300 ;
        RECT 367.600 329.600 368.400 329.700 ;
        RECT 375.600 329.600 376.400 329.700 ;
        RECT 382.000 330.300 382.800 330.400 ;
        RECT 391.600 330.300 392.400 330.400 ;
        RECT 382.000 329.700 392.400 330.300 ;
        RECT 382.000 329.600 382.800 329.700 ;
        RECT 391.600 329.600 392.400 329.700 ;
        RECT 426.800 330.300 427.600 330.400 ;
        RECT 436.400 330.300 437.200 330.400 ;
        RECT 426.800 329.700 437.200 330.300 ;
        RECT 426.800 329.600 427.600 329.700 ;
        RECT 436.400 329.600 437.200 329.700 ;
        RECT 471.600 330.300 472.400 330.400 ;
        RECT 494.000 330.300 494.800 330.400 ;
        RECT 471.600 329.700 494.800 330.300 ;
        RECT 471.600 329.600 472.400 329.700 ;
        RECT 494.000 329.600 494.800 329.700 ;
        RECT 503.600 330.300 504.400 330.400 ;
        RECT 511.600 330.300 512.400 330.400 ;
        RECT 503.600 329.700 512.400 330.300 ;
        RECT 503.600 329.600 504.400 329.700 ;
        RECT 511.600 329.600 512.400 329.700 ;
        RECT 526.000 330.300 526.800 330.400 ;
        RECT 532.400 330.300 533.200 330.400 ;
        RECT 526.000 329.700 533.200 330.300 ;
        RECT 526.000 329.600 526.800 329.700 ;
        RECT 532.400 329.600 533.200 329.700 ;
        RECT 542.000 330.300 542.800 330.400 ;
        RECT 543.600 330.300 544.400 330.400 ;
        RECT 542.000 329.700 544.400 330.300 ;
        RECT 542.000 329.600 542.800 329.700 ;
        RECT 543.600 329.600 544.400 329.700 ;
        RECT 545.200 330.300 546.000 330.400 ;
        RECT 551.600 330.300 552.400 330.400 ;
        RECT 545.200 329.700 552.400 330.300 ;
        RECT 545.200 329.600 546.000 329.700 ;
        RECT 551.600 329.600 552.400 329.700 ;
        RECT 558.000 330.300 558.800 330.400 ;
        RECT 609.200 330.300 610.000 330.400 ;
        RECT 558.000 329.700 610.000 330.300 ;
        RECT 558.000 329.600 558.800 329.700 ;
        RECT 609.200 329.600 610.000 329.700 ;
        RECT 633.200 330.300 634.000 330.400 ;
        RECT 639.600 330.300 640.400 330.400 ;
        RECT 650.800 330.300 651.600 330.400 ;
        RECT 633.200 329.700 651.600 330.300 ;
        RECT 633.200 329.600 634.000 329.700 ;
        RECT 639.600 329.600 640.400 329.700 ;
        RECT 650.800 329.600 651.600 329.700 ;
        RECT 652.400 330.300 653.200 330.400 ;
        RECT 662.000 330.300 662.800 330.400 ;
        RECT 687.600 330.300 688.400 330.400 ;
        RECT 652.400 329.700 688.400 330.300 ;
        RECT 652.400 329.600 653.200 329.700 ;
        RECT 662.000 329.600 662.800 329.700 ;
        RECT 687.600 329.600 688.400 329.700 ;
        RECT 23.600 328.300 24.400 328.400 ;
        RECT 26.800 328.300 27.600 328.400 ;
        RECT 23.600 327.700 27.600 328.300 ;
        RECT 23.600 327.600 24.400 327.700 ;
        RECT 26.800 327.600 27.600 327.700 ;
        RECT 34.800 328.300 35.600 328.400 ;
        RECT 70.000 328.300 70.800 328.400 ;
        RECT 34.800 327.700 70.800 328.300 ;
        RECT 34.800 327.600 35.600 327.700 ;
        RECT 70.000 327.600 70.800 327.700 ;
        RECT 97.200 328.300 98.000 328.400 ;
        RECT 102.000 328.300 102.800 328.400 ;
        RECT 97.200 327.700 102.800 328.300 ;
        RECT 97.200 327.600 98.000 327.700 ;
        RECT 102.000 327.600 102.800 327.700 ;
        RECT 154.800 328.300 155.600 328.400 ;
        RECT 215.600 328.300 216.400 328.400 ;
        RECT 154.800 327.700 216.400 328.300 ;
        RECT 154.800 327.600 155.600 327.700 ;
        RECT 215.600 327.600 216.400 327.700 ;
        RECT 321.200 328.300 322.000 328.400 ;
        RECT 324.400 328.300 325.200 328.400 ;
        RECT 321.200 327.700 325.200 328.300 ;
        RECT 321.200 327.600 322.000 327.700 ;
        RECT 324.400 327.600 325.200 327.700 ;
        RECT 353.200 328.300 354.000 328.400 ;
        RECT 367.700 328.300 368.300 329.600 ;
        RECT 353.200 327.700 368.300 328.300 ;
        RECT 375.600 328.300 376.400 328.400 ;
        RECT 404.400 328.300 405.200 328.400 ;
        RECT 375.600 327.700 405.200 328.300 ;
        RECT 353.200 327.600 354.000 327.700 ;
        RECT 375.600 327.600 376.400 327.700 ;
        RECT 404.400 327.600 405.200 327.700 ;
        RECT 478.000 328.300 478.800 328.400 ;
        RECT 482.800 328.300 483.600 328.400 ;
        RECT 478.000 327.700 483.600 328.300 ;
        RECT 478.000 327.600 478.800 327.700 ;
        RECT 482.800 327.600 483.600 327.700 ;
        RECT 505.200 328.300 506.000 328.400 ;
        RECT 506.800 328.300 507.600 328.400 ;
        RECT 505.200 327.700 507.600 328.300 ;
        RECT 505.200 327.600 506.000 327.700 ;
        RECT 506.800 327.600 507.600 327.700 ;
        RECT 537.200 328.300 538.000 328.400 ;
        RECT 550.000 328.300 550.800 328.400 ;
        RECT 537.200 327.700 550.800 328.300 ;
        RECT 537.200 327.600 538.000 327.700 ;
        RECT 550.000 327.600 550.800 327.700 ;
        RECT 562.800 328.300 563.600 328.400 ;
        RECT 596.400 328.300 597.200 328.400 ;
        RECT 562.800 327.700 597.200 328.300 ;
        RECT 562.800 327.600 563.600 327.700 ;
        RECT 596.400 327.600 597.200 327.700 ;
        RECT 599.600 328.300 600.400 328.400 ;
        RECT 630.000 328.300 630.800 328.400 ;
        RECT 599.600 327.700 630.800 328.300 ;
        RECT 599.600 327.600 600.400 327.700 ;
        RECT 630.000 327.600 630.800 327.700 ;
        RECT 631.600 328.300 632.400 328.400 ;
        RECT 639.600 328.300 640.400 328.400 ;
        RECT 631.600 327.700 640.400 328.300 ;
        RECT 631.600 327.600 632.400 327.700 ;
        RECT 639.600 327.600 640.400 327.700 ;
        RECT 649.200 328.300 650.000 328.400 ;
        RECT 663.600 328.300 664.400 328.400 ;
        RECT 649.200 327.700 664.400 328.300 ;
        RECT 649.200 327.600 650.000 327.700 ;
        RECT 663.600 327.600 664.400 327.700 ;
        RECT 666.800 328.300 667.600 328.400 ;
        RECT 674.800 328.300 675.600 328.400 ;
        RECT 666.800 327.700 675.600 328.300 ;
        RECT 666.800 327.600 667.600 327.700 ;
        RECT 674.800 327.600 675.600 327.700 ;
        RECT 215.600 326.300 216.400 326.400 ;
        RECT 225.200 326.300 226.000 326.400 ;
        RECT 215.600 325.700 226.000 326.300 ;
        RECT 215.600 325.600 216.400 325.700 ;
        RECT 225.200 325.600 226.000 325.700 ;
        RECT 346.800 326.300 347.600 326.400 ;
        RECT 354.800 326.300 355.600 326.400 ;
        RECT 346.800 325.700 355.600 326.300 ;
        RECT 346.800 325.600 347.600 325.700 ;
        RECT 354.800 325.600 355.600 325.700 ;
        RECT 366.000 326.300 366.800 326.400 ;
        RECT 369.200 326.300 370.000 326.400 ;
        RECT 366.000 325.700 370.000 326.300 ;
        RECT 366.000 325.600 366.800 325.700 ;
        RECT 369.200 325.600 370.000 325.700 ;
        RECT 497.200 326.300 498.000 326.400 ;
        RECT 518.000 326.300 518.800 326.400 ;
        RECT 497.200 325.700 518.800 326.300 ;
        RECT 497.200 325.600 498.000 325.700 ;
        RECT 518.000 325.600 518.800 325.700 ;
        RECT 546.800 326.300 547.600 326.400 ;
        RECT 594.800 326.300 595.600 326.400 ;
        RECT 546.800 325.700 595.600 326.300 ;
        RECT 546.800 325.600 547.600 325.700 ;
        RECT 594.800 325.600 595.600 325.700 ;
        RECT 607.600 326.300 608.400 326.400 ;
        RECT 646.000 326.300 646.800 326.400 ;
        RECT 666.800 326.300 667.600 326.400 ;
        RECT 668.400 326.300 669.200 326.400 ;
        RECT 607.600 325.700 669.200 326.300 ;
        RECT 607.600 325.600 608.400 325.700 ;
        RECT 646.000 325.600 646.800 325.700 ;
        RECT 666.800 325.600 667.600 325.700 ;
        RECT 668.400 325.600 669.200 325.700 ;
        RECT 94.000 324.300 94.800 324.400 ;
        RECT 103.600 324.300 104.400 324.400 ;
        RECT 134.000 324.300 134.800 324.400 ;
        RECT 94.000 323.700 134.800 324.300 ;
        RECT 94.000 323.600 94.800 323.700 ;
        RECT 103.600 323.600 104.400 323.700 ;
        RECT 134.000 323.600 134.800 323.700 ;
        RECT 298.800 324.300 299.600 324.400 ;
        RECT 302.000 324.300 302.800 324.400 ;
        RECT 385.200 324.300 386.000 324.400 ;
        RECT 298.800 323.700 386.000 324.300 ;
        RECT 298.800 323.600 299.600 323.700 ;
        RECT 302.000 323.600 302.800 323.700 ;
        RECT 385.200 323.600 386.000 323.700 ;
        RECT 415.600 324.300 416.400 324.400 ;
        RECT 538.800 324.300 539.600 324.400 ;
        RECT 415.600 323.700 539.600 324.300 ;
        RECT 415.600 323.600 416.400 323.700 ;
        RECT 538.800 323.600 539.600 323.700 ;
        RECT 556.400 324.300 557.200 324.400 ;
        RECT 564.400 324.300 565.200 324.400 ;
        RECT 582.000 324.300 582.800 324.400 ;
        RECT 556.400 323.700 582.800 324.300 ;
        RECT 556.400 323.600 557.200 323.700 ;
        RECT 564.400 323.600 565.200 323.700 ;
        RECT 582.000 323.600 582.800 323.700 ;
        RECT 618.800 324.300 619.600 324.400 ;
        RECT 628.400 324.300 629.200 324.400 ;
        RECT 618.800 323.700 629.200 324.300 ;
        RECT 618.800 323.600 619.600 323.700 ;
        RECT 628.400 323.600 629.200 323.700 ;
        RECT 641.200 324.300 642.000 324.400 ;
        RECT 649.200 324.300 650.000 324.400 ;
        RECT 641.200 323.700 650.000 324.300 ;
        RECT 641.200 323.600 642.000 323.700 ;
        RECT 649.200 323.600 650.000 323.700 ;
        RECT 94.000 322.300 94.800 322.400 ;
        RECT 97.200 322.300 98.000 322.400 ;
        RECT 94.000 321.700 98.000 322.300 ;
        RECT 94.000 321.600 94.800 321.700 ;
        RECT 97.200 321.600 98.000 321.700 ;
        RECT 282.800 322.300 283.600 322.400 ;
        RECT 290.800 322.300 291.600 322.400 ;
        RECT 294.000 322.300 294.800 322.400 ;
        RECT 282.800 321.700 294.800 322.300 ;
        RECT 282.800 321.600 283.600 321.700 ;
        RECT 290.800 321.600 291.600 321.700 ;
        RECT 294.000 321.600 294.800 321.700 ;
        RECT 338.800 322.300 339.600 322.400 ;
        RECT 350.000 322.300 350.800 322.400 ;
        RECT 338.800 321.700 350.800 322.300 ;
        RECT 338.800 321.600 339.600 321.700 ;
        RECT 350.000 321.600 350.800 321.700 ;
        RECT 500.400 322.300 501.200 322.400 ;
        RECT 514.800 322.300 515.600 322.400 ;
        RECT 500.400 321.700 515.600 322.300 ;
        RECT 500.400 321.600 501.200 321.700 ;
        RECT 514.800 321.600 515.600 321.700 ;
        RECT 527.600 322.300 528.400 322.400 ;
        RECT 615.600 322.300 616.400 322.400 ;
        RECT 618.800 322.300 619.600 322.400 ;
        RECT 527.600 321.700 619.600 322.300 ;
        RECT 527.600 321.600 528.400 321.700 ;
        RECT 615.600 321.600 616.400 321.700 ;
        RECT 618.800 321.600 619.600 321.700 ;
        RECT 225.200 320.300 226.000 320.400 ;
        RECT 244.400 320.300 245.200 320.400 ;
        RECT 225.200 319.700 245.200 320.300 ;
        RECT 225.200 319.600 226.000 319.700 ;
        RECT 244.400 319.600 245.200 319.700 ;
        RECT 247.600 320.300 248.400 320.400 ;
        RECT 270.000 320.300 270.800 320.400 ;
        RECT 286.000 320.300 286.800 320.400 ;
        RECT 247.600 319.700 286.800 320.300 ;
        RECT 247.600 319.600 248.400 319.700 ;
        RECT 270.000 319.600 270.800 319.700 ;
        RECT 286.000 319.600 286.800 319.700 ;
        RECT 330.800 320.300 331.600 320.400 ;
        RECT 345.200 320.300 346.000 320.400 ;
        RECT 330.800 319.700 346.000 320.300 ;
        RECT 330.800 319.600 331.600 319.700 ;
        RECT 345.200 319.600 346.000 319.700 ;
        RECT 505.200 320.300 506.000 320.400 ;
        RECT 530.800 320.300 531.600 320.400 ;
        RECT 505.200 319.700 531.600 320.300 ;
        RECT 505.200 319.600 506.000 319.700 ;
        RECT 530.800 319.600 531.600 319.700 ;
        RECT 609.200 320.300 610.000 320.400 ;
        RECT 638.000 320.300 638.800 320.400 ;
        RECT 609.200 319.700 638.800 320.300 ;
        RECT 609.200 319.600 610.000 319.700 ;
        RECT 638.000 319.600 638.800 319.700 ;
        RECT 676.400 320.300 677.200 320.400 ;
        RECT 681.200 320.300 682.000 320.400 ;
        RECT 676.400 319.700 682.000 320.300 ;
        RECT 676.400 319.600 677.200 319.700 ;
        RECT 681.200 319.600 682.000 319.700 ;
        RECT 74.800 318.300 75.600 318.400 ;
        RECT 145.200 318.300 146.000 318.400 ;
        RECT 74.800 317.700 146.000 318.300 ;
        RECT 74.800 317.600 75.600 317.700 ;
        RECT 145.200 317.600 146.000 317.700 ;
        RECT 156.400 318.300 157.200 318.400 ;
        RECT 190.000 318.300 190.800 318.400 ;
        RECT 220.400 318.300 221.200 318.400 ;
        RECT 156.400 317.700 221.200 318.300 ;
        RECT 156.400 317.600 157.200 317.700 ;
        RECT 190.000 317.600 190.800 317.700 ;
        RECT 220.400 317.600 221.200 317.700 ;
        RECT 295.600 318.300 296.400 318.400 ;
        RECT 337.200 318.300 338.000 318.400 ;
        RECT 353.200 318.300 354.000 318.400 ;
        RECT 295.600 317.700 354.000 318.300 ;
        RECT 295.600 317.600 296.400 317.700 ;
        RECT 337.200 317.600 338.000 317.700 ;
        RECT 353.200 317.600 354.000 317.700 ;
        RECT 369.200 318.300 370.000 318.400 ;
        RECT 375.600 318.300 376.400 318.400 ;
        RECT 369.200 317.700 376.400 318.300 ;
        RECT 369.200 317.600 370.000 317.700 ;
        RECT 375.600 317.600 376.400 317.700 ;
        RECT 439.600 318.300 440.400 318.400 ;
        RECT 479.600 318.300 480.400 318.400 ;
        RECT 486.000 318.300 486.800 318.400 ;
        RECT 439.600 317.700 480.400 318.300 ;
        RECT 439.600 317.600 440.400 317.700 ;
        RECT 479.600 317.600 480.400 317.700 ;
        RECT 481.300 317.700 486.800 318.300 ;
        RECT 38.000 316.300 38.800 316.400 ;
        RECT 46.000 316.300 46.800 316.400 ;
        RECT 66.800 316.300 67.600 316.400 ;
        RECT 169.200 316.300 170.000 316.400 ;
        RECT 210.800 316.300 211.600 316.400 ;
        RECT 38.000 315.700 67.600 316.300 ;
        RECT 38.000 315.600 38.800 315.700 ;
        RECT 46.000 315.600 46.800 315.700 ;
        RECT 66.800 315.600 67.600 315.700 ;
        RECT 68.500 315.700 211.600 316.300 ;
        RECT 60.400 314.300 61.200 314.400 ;
        RECT 68.500 314.300 69.100 315.700 ;
        RECT 169.200 315.600 170.000 315.700 ;
        RECT 210.800 315.600 211.600 315.700 ;
        RECT 297.200 316.300 298.000 316.400 ;
        RECT 300.400 316.300 301.200 316.400 ;
        RECT 297.200 315.700 301.200 316.300 ;
        RECT 297.200 315.600 298.000 315.700 ;
        RECT 300.400 315.600 301.200 315.700 ;
        RECT 314.800 316.300 315.600 316.400 ;
        RECT 321.200 316.300 322.000 316.400 ;
        RECT 314.800 315.700 322.000 316.300 ;
        RECT 314.800 315.600 315.600 315.700 ;
        RECT 321.200 315.600 322.000 315.700 ;
        RECT 334.000 316.300 334.800 316.400 ;
        RECT 346.800 316.300 347.600 316.400 ;
        RECT 334.000 315.700 347.600 316.300 ;
        RECT 334.000 315.600 334.800 315.700 ;
        RECT 346.800 315.600 347.600 315.700 ;
        RECT 452.400 316.300 453.200 316.400 ;
        RECT 481.300 316.300 481.900 317.700 ;
        RECT 486.000 317.600 486.800 317.700 ;
        RECT 498.800 318.300 499.600 318.400 ;
        RECT 553.200 318.300 554.000 318.400 ;
        RECT 498.800 317.700 554.000 318.300 ;
        RECT 498.800 317.600 499.600 317.700 ;
        RECT 553.200 317.600 554.000 317.700 ;
        RECT 554.800 318.300 555.600 318.400 ;
        RECT 633.200 318.300 634.000 318.400 ;
        RECT 554.800 317.700 634.000 318.300 ;
        RECT 554.800 317.600 555.600 317.700 ;
        RECT 633.200 317.600 634.000 317.700 ;
        RECT 642.800 318.300 643.600 318.400 ;
        RECT 662.000 318.300 662.800 318.400 ;
        RECT 642.800 317.700 662.800 318.300 ;
        RECT 642.800 317.600 643.600 317.700 ;
        RECT 662.000 317.600 662.800 317.700 ;
        RECT 452.400 315.700 481.900 316.300 ;
        RECT 482.800 316.300 483.600 316.400 ;
        RECT 495.600 316.300 496.400 316.400 ;
        RECT 556.400 316.300 557.200 316.400 ;
        RECT 482.800 315.700 557.200 316.300 ;
        RECT 452.400 315.600 453.200 315.700 ;
        RECT 482.800 315.600 483.600 315.700 ;
        RECT 495.600 315.600 496.400 315.700 ;
        RECT 556.400 315.600 557.200 315.700 ;
        RECT 567.600 316.300 568.400 316.400 ;
        RECT 623.600 316.300 624.400 316.400 ;
        RECT 567.600 315.700 624.400 316.300 ;
        RECT 567.600 315.600 568.400 315.700 ;
        RECT 623.600 315.600 624.400 315.700 ;
        RECT 638.000 316.300 638.800 316.400 ;
        RECT 644.400 316.300 645.200 316.400 ;
        RECT 638.000 315.700 645.200 316.300 ;
        RECT 638.000 315.600 638.800 315.700 ;
        RECT 644.400 315.600 645.200 315.700 ;
        RECT 60.400 313.700 69.100 314.300 ;
        RECT 137.200 314.300 138.000 314.400 ;
        RECT 230.000 314.300 230.800 314.400 ;
        RECT 137.200 313.700 230.800 314.300 ;
        RECT 60.400 313.600 61.200 313.700 ;
        RECT 137.200 313.600 138.000 313.700 ;
        RECT 230.000 313.600 230.800 313.700 ;
        RECT 252.400 314.300 253.200 314.400 ;
        RECT 286.000 314.300 286.800 314.400 ;
        RECT 295.600 314.300 296.400 314.400 ;
        RECT 252.400 313.700 296.400 314.300 ;
        RECT 252.400 313.600 253.200 313.700 ;
        RECT 286.000 313.600 286.800 313.700 ;
        RECT 295.600 313.600 296.400 313.700 ;
        RECT 298.800 314.300 299.600 314.400 ;
        RECT 311.600 314.300 312.400 314.400 ;
        RECT 298.800 313.700 312.400 314.300 ;
        RECT 298.800 313.600 299.600 313.700 ;
        RECT 311.600 313.600 312.400 313.700 ;
        RECT 318.000 314.300 318.800 314.400 ;
        RECT 340.400 314.300 341.200 314.400 ;
        RECT 490.800 314.300 491.600 314.400 ;
        RECT 503.600 314.300 504.400 314.400 ;
        RECT 318.000 313.700 341.200 314.300 ;
        RECT 318.000 313.600 318.800 313.700 ;
        RECT 340.400 313.600 341.200 313.700 ;
        RECT 474.900 313.700 504.400 314.300 ;
        RECT 474.900 312.400 475.500 313.700 ;
        RECT 490.800 313.600 491.600 313.700 ;
        RECT 503.600 313.600 504.400 313.700 ;
        RECT 505.200 314.300 506.000 314.400 ;
        RECT 508.400 314.300 509.200 314.400 ;
        RECT 505.200 313.700 509.200 314.300 ;
        RECT 505.200 313.600 506.000 313.700 ;
        RECT 508.400 313.600 509.200 313.700 ;
        RECT 518.000 314.300 518.800 314.400 ;
        RECT 527.600 314.300 528.400 314.400 ;
        RECT 518.000 313.700 528.400 314.300 ;
        RECT 518.000 313.600 518.800 313.700 ;
        RECT 527.600 313.600 528.400 313.700 ;
        RECT 532.400 314.300 533.200 314.400 ;
        RECT 542.000 314.300 542.800 314.400 ;
        RECT 532.400 313.700 542.800 314.300 ;
        RECT 532.400 313.600 533.200 313.700 ;
        RECT 542.000 313.600 542.800 313.700 ;
        RECT 561.200 313.600 562.000 314.400 ;
        RECT 594.800 314.300 595.600 314.400 ;
        RECT 598.000 314.300 598.800 314.400 ;
        RECT 601.200 314.300 602.000 314.400 ;
        RECT 594.800 313.700 602.000 314.300 ;
        RECT 594.800 313.600 595.600 313.700 ;
        RECT 598.000 313.600 598.800 313.700 ;
        RECT 601.200 313.600 602.000 313.700 ;
        RECT 655.600 314.300 656.400 314.400 ;
        RECT 660.400 314.300 661.200 314.400 ;
        RECT 655.600 313.700 661.200 314.300 ;
        RECT 655.600 313.600 656.400 313.700 ;
        RECT 660.400 313.600 661.200 313.700 ;
        RECT 33.200 312.300 34.000 312.400 ;
        RECT 41.200 312.300 42.000 312.400 ;
        RECT 50.800 312.300 51.600 312.400 ;
        RECT 33.200 311.700 51.600 312.300 ;
        RECT 33.200 311.600 34.000 311.700 ;
        RECT 41.200 311.600 42.000 311.700 ;
        RECT 50.800 311.600 51.600 311.700 ;
        RECT 90.800 312.300 91.600 312.400 ;
        RECT 100.400 312.300 101.200 312.400 ;
        RECT 90.800 311.700 101.200 312.300 ;
        RECT 90.800 311.600 91.600 311.700 ;
        RECT 100.400 311.600 101.200 311.700 ;
        RECT 146.800 312.300 147.600 312.400 ;
        RECT 153.200 312.300 154.000 312.400 ;
        RECT 146.800 311.700 154.000 312.300 ;
        RECT 146.800 311.600 147.600 311.700 ;
        RECT 153.200 311.600 154.000 311.700 ;
        RECT 279.600 312.300 280.400 312.400 ;
        RECT 300.400 312.300 301.200 312.400 ;
        RECT 279.600 311.700 301.200 312.300 ;
        RECT 279.600 311.600 280.400 311.700 ;
        RECT 300.400 311.600 301.200 311.700 ;
        RECT 311.600 311.600 312.400 312.400 ;
        RECT 313.200 312.300 314.000 312.400 ;
        RECT 316.400 312.300 317.200 312.400 ;
        RECT 313.200 311.700 317.200 312.300 ;
        RECT 313.200 311.600 314.000 311.700 ;
        RECT 316.400 311.600 317.200 311.700 ;
        RECT 327.600 312.300 328.400 312.400 ;
        RECT 330.800 312.300 331.600 312.400 ;
        RECT 343.600 312.300 344.400 312.400 ;
        RECT 327.600 311.700 344.400 312.300 ;
        RECT 327.600 311.600 328.400 311.700 ;
        RECT 330.800 311.600 331.600 311.700 ;
        RECT 343.600 311.600 344.400 311.700 ;
        RECT 358.000 312.300 358.800 312.400 ;
        RECT 362.800 312.300 363.600 312.400 ;
        RECT 358.000 311.700 363.600 312.300 ;
        RECT 358.000 311.600 358.800 311.700 ;
        RECT 362.800 311.600 363.600 311.700 ;
        RECT 465.200 312.300 466.000 312.400 ;
        RECT 474.800 312.300 475.600 312.400 ;
        RECT 465.200 311.700 475.600 312.300 ;
        RECT 465.200 311.600 466.000 311.700 ;
        RECT 474.800 311.600 475.600 311.700 ;
        RECT 479.600 312.300 480.400 312.400 ;
        RECT 484.400 312.300 485.200 312.400 ;
        RECT 479.600 311.700 485.200 312.300 ;
        RECT 479.600 311.600 480.400 311.700 ;
        RECT 484.400 311.600 485.200 311.700 ;
        RECT 494.000 312.300 494.800 312.400 ;
        RECT 500.400 312.300 501.200 312.400 ;
        RECT 494.000 311.700 501.200 312.300 ;
        RECT 494.000 311.600 494.800 311.700 ;
        RECT 500.400 311.600 501.200 311.700 ;
        RECT 519.600 312.300 520.400 312.400 ;
        RECT 534.000 312.300 534.800 312.400 ;
        RECT 519.600 311.700 534.800 312.300 ;
        RECT 519.600 311.600 520.400 311.700 ;
        RECT 534.000 311.600 534.800 311.700 ;
        RECT 542.000 312.300 542.800 312.400 ;
        RECT 550.000 312.300 550.800 312.400 ;
        RECT 558.000 312.300 558.800 312.400 ;
        RECT 542.000 311.700 558.800 312.300 ;
        RECT 542.000 311.600 542.800 311.700 ;
        RECT 550.000 311.600 550.800 311.700 ;
        RECT 558.000 311.600 558.800 311.700 ;
        RECT 582.000 312.300 582.800 312.400 ;
        RECT 626.800 312.300 627.600 312.400 ;
        RECT 582.000 311.700 627.600 312.300 ;
        RECT 582.000 311.600 582.800 311.700 ;
        RECT 626.800 311.600 627.600 311.700 ;
        RECT 644.400 312.300 645.200 312.400 ;
        RECT 652.400 312.300 653.200 312.400 ;
        RECT 660.400 312.300 661.200 312.400 ;
        RECT 686.000 312.300 686.800 312.400 ;
        RECT 644.400 311.700 686.800 312.300 ;
        RECT 644.400 311.600 645.200 311.700 ;
        RECT 652.400 311.600 653.200 311.700 ;
        RECT 660.400 311.600 661.200 311.700 ;
        RECT 686.000 311.600 686.800 311.700 ;
        RECT 28.400 310.300 29.200 310.400 ;
        RECT 36.400 310.300 37.200 310.400 ;
        RECT 87.600 310.300 88.400 310.400 ;
        RECT 28.400 309.700 88.400 310.300 ;
        RECT 28.400 309.600 29.200 309.700 ;
        RECT 36.400 309.600 37.200 309.700 ;
        RECT 87.600 309.600 88.400 309.700 ;
        RECT 102.000 310.300 102.800 310.400 ;
        RECT 140.400 310.300 141.200 310.400 ;
        RECT 102.000 309.700 141.200 310.300 ;
        RECT 102.000 309.600 102.800 309.700 ;
        RECT 140.400 309.600 141.200 309.700 ;
        RECT 150.000 310.300 150.800 310.400 ;
        RECT 161.200 310.300 162.000 310.400 ;
        RECT 150.000 309.700 162.000 310.300 ;
        RECT 150.000 309.600 150.800 309.700 ;
        RECT 161.200 309.600 162.000 309.700 ;
        RECT 166.000 310.300 166.800 310.400 ;
        RECT 209.200 310.300 210.000 310.400 ;
        RECT 166.000 309.700 210.000 310.300 ;
        RECT 166.000 309.600 166.800 309.700 ;
        RECT 209.200 309.600 210.000 309.700 ;
        RECT 242.800 310.300 243.600 310.400 ;
        RECT 266.800 310.300 267.600 310.400 ;
        RECT 242.800 309.700 267.600 310.300 ;
        RECT 242.800 309.600 243.600 309.700 ;
        RECT 266.800 309.600 267.600 309.700 ;
        RECT 300.400 310.300 301.200 310.400 ;
        RECT 303.600 310.300 304.400 310.400 ;
        RECT 300.400 309.700 304.400 310.300 ;
        RECT 300.400 309.600 301.200 309.700 ;
        RECT 303.600 309.600 304.400 309.700 ;
        RECT 306.800 310.300 307.600 310.400 ;
        RECT 327.700 310.300 328.300 311.600 ;
        RECT 306.800 309.700 328.300 310.300 ;
        RECT 348.400 310.300 349.200 310.400 ;
        RECT 361.200 310.300 362.000 310.400 ;
        RECT 348.400 309.700 362.000 310.300 ;
        RECT 306.800 309.600 307.600 309.700 ;
        RECT 348.400 309.600 349.200 309.700 ;
        RECT 361.200 309.600 362.000 309.700 ;
        RECT 394.800 310.300 395.600 310.400 ;
        RECT 410.800 310.300 411.600 310.400 ;
        RECT 394.800 309.700 411.600 310.300 ;
        RECT 394.800 309.600 395.600 309.700 ;
        RECT 410.800 309.600 411.600 309.700 ;
        RECT 468.400 310.300 469.200 310.400 ;
        RECT 478.000 310.300 478.800 310.400 ;
        RECT 513.200 310.300 514.000 310.400 ;
        RECT 516.400 310.300 517.200 310.400 ;
        RECT 556.400 310.300 557.200 310.400 ;
        RECT 468.400 309.700 557.200 310.300 ;
        RECT 468.400 309.600 469.200 309.700 ;
        RECT 478.000 309.600 478.800 309.700 ;
        RECT 513.200 309.600 514.000 309.700 ;
        RECT 516.400 309.600 517.200 309.700 ;
        RECT 556.400 309.600 557.200 309.700 ;
        RECT 558.000 310.300 558.800 310.400 ;
        RECT 598.000 310.300 598.800 310.400 ;
        RECT 599.600 310.300 600.400 310.400 ;
        RECT 558.000 309.700 600.400 310.300 ;
        RECT 558.000 309.600 558.800 309.700 ;
        RECT 598.000 309.600 598.800 309.700 ;
        RECT 599.600 309.600 600.400 309.700 ;
        RECT 601.200 310.300 602.000 310.400 ;
        RECT 610.800 310.300 611.600 310.400 ;
        RECT 601.200 309.700 611.600 310.300 ;
        RECT 601.200 309.600 602.000 309.700 ;
        RECT 610.800 309.600 611.600 309.700 ;
        RECT 623.600 310.300 624.400 310.400 ;
        RECT 633.200 310.300 634.000 310.400 ;
        RECT 623.600 309.700 634.000 310.300 ;
        RECT 623.600 309.600 624.400 309.700 ;
        RECT 633.200 309.600 634.000 309.700 ;
        RECT 634.800 310.300 635.600 310.400 ;
        RECT 642.800 310.300 643.600 310.400 ;
        RECT 634.800 309.700 643.600 310.300 ;
        RECT 634.800 309.600 635.600 309.700 ;
        RECT 642.800 309.600 643.600 309.700 ;
        RECT 663.600 310.300 664.400 310.400 ;
        RECT 673.200 310.300 674.000 310.400 ;
        RECT 663.600 309.700 674.000 310.300 ;
        RECT 663.600 309.600 664.400 309.700 ;
        RECT 673.200 309.600 674.000 309.700 ;
        RECT 14.000 308.300 14.800 308.400 ;
        RECT 42.800 308.300 43.600 308.400 ;
        RECT 14.000 307.700 43.600 308.300 ;
        RECT 14.000 307.600 14.800 307.700 ;
        RECT 42.800 307.600 43.600 307.700 ;
        RECT 55.600 308.300 56.400 308.400 ;
        RECT 60.400 308.300 61.200 308.400 ;
        RECT 95.600 308.300 96.400 308.400 ;
        RECT 55.600 307.700 96.400 308.300 ;
        RECT 55.600 307.600 56.400 307.700 ;
        RECT 60.400 307.600 61.200 307.700 ;
        RECT 95.600 307.600 96.400 307.700 ;
        RECT 110.000 308.300 110.800 308.400 ;
        RECT 124.400 308.300 125.200 308.400 ;
        RECT 110.000 307.700 125.200 308.300 ;
        RECT 110.000 307.600 110.800 307.700 ;
        RECT 124.400 307.600 125.200 307.700 ;
        RECT 154.800 308.300 155.600 308.400 ;
        RECT 162.800 308.300 163.600 308.400 ;
        RECT 154.800 307.700 163.600 308.300 ;
        RECT 154.800 307.600 155.600 307.700 ;
        RECT 162.800 307.600 163.600 307.700 ;
        RECT 188.400 308.300 189.200 308.400 ;
        RECT 206.000 308.300 206.800 308.400 ;
        RECT 188.400 307.700 206.800 308.300 ;
        RECT 188.400 307.600 189.200 307.700 ;
        RECT 206.000 307.600 206.800 307.700 ;
        RECT 217.200 308.300 218.000 308.400 ;
        RECT 226.800 308.300 227.600 308.400 ;
        RECT 217.200 307.700 227.600 308.300 ;
        RECT 217.200 307.600 218.000 307.700 ;
        RECT 226.800 307.600 227.600 307.700 ;
        RECT 359.600 307.600 360.400 308.400 ;
        RECT 407.600 308.300 408.400 308.400 ;
        RECT 420.400 308.300 421.200 308.400 ;
        RECT 407.600 307.700 421.200 308.300 ;
        RECT 407.600 307.600 408.400 307.700 ;
        RECT 420.400 307.600 421.200 307.700 ;
        RECT 444.400 308.300 445.200 308.400 ;
        RECT 470.000 308.300 470.800 308.400 ;
        RECT 444.400 307.700 470.800 308.300 ;
        RECT 444.400 307.600 445.200 307.700 ;
        RECT 470.000 307.600 470.800 307.700 ;
        RECT 471.600 308.300 472.400 308.400 ;
        RECT 481.200 308.300 482.000 308.400 ;
        RECT 471.600 307.700 482.000 308.300 ;
        RECT 471.600 307.600 472.400 307.700 ;
        RECT 481.200 307.600 482.000 307.700 ;
        RECT 495.600 308.300 496.400 308.400 ;
        RECT 502.000 308.300 502.800 308.400 ;
        RECT 495.600 307.700 502.800 308.300 ;
        RECT 495.600 307.600 496.400 307.700 ;
        RECT 502.000 307.600 502.800 307.700 ;
        RECT 538.800 308.300 539.600 308.400 ;
        RECT 542.000 308.300 542.800 308.400 ;
        RECT 538.800 307.700 542.800 308.300 ;
        RECT 538.800 307.600 539.600 307.700 ;
        RECT 542.000 307.600 542.800 307.700 ;
        RECT 554.800 308.300 555.600 308.400 ;
        RECT 562.800 308.300 563.600 308.400 ;
        RECT 554.800 307.700 563.600 308.300 ;
        RECT 554.800 307.600 555.600 307.700 ;
        RECT 562.800 307.600 563.600 307.700 ;
        RECT 569.200 308.300 570.000 308.400 ;
        RECT 598.000 308.300 598.800 308.400 ;
        RECT 569.200 307.700 598.800 308.300 ;
        RECT 569.200 307.600 570.000 307.700 ;
        RECT 598.000 307.600 598.800 307.700 ;
        RECT 599.600 308.300 600.400 308.400 ;
        RECT 602.800 308.300 603.600 308.400 ;
        RECT 599.600 307.700 603.600 308.300 ;
        RECT 599.600 307.600 600.400 307.700 ;
        RECT 602.800 307.600 603.600 307.700 ;
        RECT 606.000 308.300 606.800 308.400 ;
        RECT 612.400 308.300 613.200 308.400 ;
        RECT 606.000 307.700 613.200 308.300 ;
        RECT 606.000 307.600 606.800 307.700 ;
        RECT 612.400 307.600 613.200 307.700 ;
        RECT 615.600 308.300 616.400 308.400 ;
        RECT 641.200 308.300 642.000 308.400 ;
        RECT 615.600 307.700 642.000 308.300 ;
        RECT 615.600 307.600 616.400 307.700 ;
        RECT 641.200 307.600 642.000 307.700 ;
        RECT 650.800 308.300 651.600 308.400 ;
        RECT 665.200 308.300 666.000 308.400 ;
        RECT 650.800 307.700 666.000 308.300 ;
        RECT 650.800 307.600 651.600 307.700 ;
        RECT 665.200 307.600 666.000 307.700 ;
        RECT 17.200 305.600 18.000 306.400 ;
        RECT 55.600 306.300 56.400 306.400 ;
        RECT 62.000 306.300 62.800 306.400 ;
        RECT 55.600 305.700 62.800 306.300 ;
        RECT 55.600 305.600 56.400 305.700 ;
        RECT 62.000 305.600 62.800 305.700 ;
        RECT 86.000 306.300 86.800 306.400 ;
        RECT 113.200 306.300 114.000 306.400 ;
        RECT 86.000 305.700 114.000 306.300 ;
        RECT 86.000 305.600 86.800 305.700 ;
        RECT 113.200 305.600 114.000 305.700 ;
        RECT 135.600 306.300 136.400 306.400 ;
        RECT 162.800 306.300 163.600 306.400 ;
        RECT 135.600 305.700 163.600 306.300 ;
        RECT 135.600 305.600 136.400 305.700 ;
        RECT 162.800 305.600 163.600 305.700 ;
        RECT 170.800 306.300 171.600 306.400 ;
        RECT 177.200 306.300 178.000 306.400 ;
        RECT 170.800 305.700 178.000 306.300 ;
        RECT 170.800 305.600 171.600 305.700 ;
        RECT 177.200 305.600 178.000 305.700 ;
        RECT 185.200 306.300 186.000 306.400 ;
        RECT 186.800 306.300 187.600 306.400 ;
        RECT 185.200 305.700 187.600 306.300 ;
        RECT 185.200 305.600 186.000 305.700 ;
        RECT 186.800 305.600 187.600 305.700 ;
        RECT 241.200 306.300 242.000 306.400 ;
        RECT 246.000 306.300 246.800 306.400 ;
        RECT 241.200 305.700 246.800 306.300 ;
        RECT 241.200 305.600 242.000 305.700 ;
        RECT 246.000 305.600 246.800 305.700 ;
        RECT 290.800 306.300 291.600 306.400 ;
        RECT 324.400 306.300 325.200 306.400 ;
        RECT 342.000 306.300 342.800 306.400 ;
        RECT 290.800 305.700 342.800 306.300 ;
        RECT 290.800 305.600 291.600 305.700 ;
        RECT 324.400 305.600 325.200 305.700 ;
        RECT 342.000 305.600 342.800 305.700 ;
        RECT 345.200 306.300 346.000 306.400 ;
        RECT 353.200 306.300 354.000 306.400 ;
        RECT 345.200 305.700 354.000 306.300 ;
        RECT 345.200 305.600 346.000 305.700 ;
        RECT 353.200 305.600 354.000 305.700 ;
        RECT 358.000 306.300 358.800 306.400 ;
        RECT 388.400 306.300 389.200 306.400 ;
        RECT 358.000 305.700 389.200 306.300 ;
        RECT 358.000 305.600 358.800 305.700 ;
        RECT 388.400 305.600 389.200 305.700 ;
        RECT 479.600 306.300 480.400 306.400 ;
        RECT 486.000 306.300 486.800 306.400 ;
        RECT 479.600 305.700 486.800 306.300 ;
        RECT 479.600 305.600 480.400 305.700 ;
        RECT 486.000 305.600 486.800 305.700 ;
        RECT 487.600 306.300 488.400 306.400 ;
        RECT 497.200 306.300 498.000 306.400 ;
        RECT 487.600 305.700 498.000 306.300 ;
        RECT 487.600 305.600 488.400 305.700 ;
        RECT 497.200 305.600 498.000 305.700 ;
        RECT 529.200 306.300 530.000 306.400 ;
        RECT 543.600 306.300 544.400 306.400 ;
        RECT 551.600 306.300 552.400 306.400 ;
        RECT 529.200 305.700 552.400 306.300 ;
        RECT 529.200 305.600 530.000 305.700 ;
        RECT 543.600 305.600 544.400 305.700 ;
        RECT 551.600 305.600 552.400 305.700 ;
        RECT 601.200 306.300 602.000 306.400 ;
        RECT 607.600 306.300 608.400 306.400 ;
        RECT 601.200 305.700 608.400 306.300 ;
        RECT 601.200 305.600 602.000 305.700 ;
        RECT 607.600 305.600 608.400 305.700 ;
        RECT 639.600 306.300 640.400 306.400 ;
        RECT 641.200 306.300 642.000 306.400 ;
        RECT 639.600 305.700 642.000 306.300 ;
        RECT 639.600 305.600 640.400 305.700 ;
        RECT 641.200 305.600 642.000 305.700 ;
        RECT 654.000 306.300 654.800 306.400 ;
        RECT 666.800 306.300 667.600 306.400 ;
        RECT 654.000 305.700 667.600 306.300 ;
        RECT 654.000 305.600 654.800 305.700 ;
        RECT 666.800 305.600 667.600 305.700 ;
        RECT 177.200 304.300 178.000 304.400 ;
        RECT 204.400 304.300 205.200 304.400 ;
        RECT 177.200 303.700 205.200 304.300 ;
        RECT 177.200 303.600 178.000 303.700 ;
        RECT 204.400 303.600 205.200 303.700 ;
        RECT 215.600 303.600 216.400 304.400 ;
        RECT 226.800 304.300 227.600 304.400 ;
        RECT 242.800 304.300 243.600 304.400 ;
        RECT 226.800 303.700 243.600 304.300 ;
        RECT 226.800 303.600 227.600 303.700 ;
        RECT 242.800 303.600 243.600 303.700 ;
        RECT 414.000 304.300 414.800 304.400 ;
        RECT 439.600 304.300 440.400 304.400 ;
        RECT 414.000 303.700 440.400 304.300 ;
        RECT 414.000 303.600 414.800 303.700 ;
        RECT 439.600 303.600 440.400 303.700 ;
        RECT 570.800 304.300 571.600 304.400 ;
        RECT 588.400 304.300 589.200 304.400 ;
        RECT 570.800 303.700 589.200 304.300 ;
        RECT 570.800 303.600 571.600 303.700 ;
        RECT 588.400 303.600 589.200 303.700 ;
        RECT 598.000 304.300 598.800 304.400 ;
        RECT 646.000 304.300 646.800 304.400 ;
        RECT 598.000 303.700 646.800 304.300 ;
        RECT 598.000 303.600 598.800 303.700 ;
        RECT 646.000 303.600 646.800 303.700 ;
        RECT 23.600 302.300 24.400 302.400 ;
        RECT 31.600 302.300 32.400 302.400 ;
        RECT 23.600 301.700 32.400 302.300 ;
        RECT 23.600 301.600 24.400 301.700 ;
        RECT 31.600 301.600 32.400 301.700 ;
        RECT 127.600 302.300 128.400 302.400 ;
        RECT 134.000 302.300 134.800 302.400 ;
        RECT 127.600 301.700 134.800 302.300 ;
        RECT 127.600 301.600 128.400 301.700 ;
        RECT 134.000 301.600 134.800 301.700 ;
        RECT 180.400 302.300 181.200 302.400 ;
        RECT 222.000 302.300 222.800 302.400 ;
        RECT 247.600 302.300 248.400 302.400 ;
        RECT 180.400 301.700 248.400 302.300 ;
        RECT 180.400 301.600 181.200 301.700 ;
        RECT 222.000 301.600 222.800 301.700 ;
        RECT 247.600 301.600 248.400 301.700 ;
        RECT 270.000 302.300 270.800 302.400 ;
        RECT 274.800 302.300 275.600 302.400 ;
        RECT 270.000 301.700 275.600 302.300 ;
        RECT 270.000 301.600 270.800 301.700 ;
        RECT 274.800 301.600 275.600 301.700 ;
        RECT 308.400 302.300 309.200 302.400 ;
        RECT 335.600 302.300 336.400 302.400 ;
        RECT 308.400 301.700 336.400 302.300 ;
        RECT 308.400 301.600 309.200 301.700 ;
        RECT 335.600 301.600 336.400 301.700 ;
        RECT 343.600 302.300 344.400 302.400 ;
        RECT 362.800 302.300 363.600 302.400 ;
        RECT 343.600 301.700 363.600 302.300 ;
        RECT 343.600 301.600 344.400 301.700 ;
        RECT 362.800 301.600 363.600 301.700 ;
        RECT 369.200 302.300 370.000 302.400 ;
        RECT 441.200 302.300 442.000 302.400 ;
        RECT 369.200 301.700 442.000 302.300 ;
        RECT 369.200 301.600 370.000 301.700 ;
        RECT 441.200 301.600 442.000 301.700 ;
        RECT 478.000 302.300 478.800 302.400 ;
        RECT 538.800 302.300 539.600 302.400 ;
        RECT 569.200 302.300 570.000 302.400 ;
        RECT 478.000 301.700 570.000 302.300 ;
        RECT 478.000 301.600 478.800 301.700 ;
        RECT 538.800 301.600 539.600 301.700 ;
        RECT 569.200 301.600 570.000 301.700 ;
        RECT 596.400 302.300 597.200 302.400 ;
        RECT 607.600 302.300 608.400 302.400 ;
        RECT 625.200 302.300 626.000 302.400 ;
        RECT 596.400 301.700 606.700 302.300 ;
        RECT 596.400 301.600 597.200 301.700 ;
        RECT 162.800 300.300 163.600 300.400 ;
        RECT 199.600 300.300 200.400 300.400 ;
        RECT 217.200 300.300 218.000 300.400 ;
        RECT 162.800 299.700 218.000 300.300 ;
        RECT 162.800 299.600 163.600 299.700 ;
        RECT 199.600 299.600 200.400 299.700 ;
        RECT 217.200 299.600 218.000 299.700 ;
        RECT 426.800 300.300 427.600 300.400 ;
        RECT 431.600 300.300 432.400 300.400 ;
        RECT 426.800 299.700 432.400 300.300 ;
        RECT 426.800 299.600 427.600 299.700 ;
        RECT 431.600 299.600 432.400 299.700 ;
        RECT 481.200 300.300 482.000 300.400 ;
        RECT 484.400 300.300 485.200 300.400 ;
        RECT 481.200 299.700 485.200 300.300 ;
        RECT 481.200 299.600 482.000 299.700 ;
        RECT 484.400 299.600 485.200 299.700 ;
        RECT 583.600 300.300 584.400 300.400 ;
        RECT 602.800 300.300 603.600 300.400 ;
        RECT 583.600 299.700 603.600 300.300 ;
        RECT 606.100 300.300 606.700 301.700 ;
        RECT 607.600 301.700 626.000 302.300 ;
        RECT 607.600 301.600 608.400 301.700 ;
        RECT 625.200 301.600 626.000 301.700 ;
        RECT 666.800 302.300 667.600 302.400 ;
        RECT 673.200 302.300 674.000 302.400 ;
        RECT 676.400 302.300 677.200 302.400 ;
        RECT 681.200 302.300 682.000 302.400 ;
        RECT 666.800 301.700 682.000 302.300 ;
        RECT 666.800 301.600 667.600 301.700 ;
        RECT 673.200 301.600 674.000 301.700 ;
        RECT 676.400 301.600 677.200 301.700 ;
        RECT 681.200 301.600 682.000 301.700 ;
        RECT 612.400 300.300 613.200 300.400 ;
        RECT 647.600 300.300 648.400 300.400 ;
        RECT 655.600 300.300 656.400 300.400 ;
        RECT 606.100 299.700 656.400 300.300 ;
        RECT 583.600 299.600 584.400 299.700 ;
        RECT 602.800 299.600 603.600 299.700 ;
        RECT 612.400 299.600 613.200 299.700 ;
        RECT 647.600 299.600 648.400 299.700 ;
        RECT 655.600 299.600 656.400 299.700 ;
        RECT 111.600 298.300 112.400 298.400 ;
        RECT 146.800 298.300 147.600 298.400 ;
        RECT 111.600 297.700 147.600 298.300 ;
        RECT 111.600 297.600 112.400 297.700 ;
        RECT 146.800 297.600 147.600 297.700 ;
        RECT 190.000 297.600 190.800 298.400 ;
        RECT 247.600 298.300 248.400 298.400 ;
        RECT 294.000 298.300 294.800 298.400 ;
        RECT 247.600 297.700 294.800 298.300 ;
        RECT 247.600 297.600 248.400 297.700 ;
        RECT 294.000 297.600 294.800 297.700 ;
        RECT 324.400 298.300 325.200 298.400 ;
        RECT 327.600 298.300 328.400 298.400 ;
        RECT 324.400 297.700 328.400 298.300 ;
        RECT 324.400 297.600 325.200 297.700 ;
        RECT 327.600 297.600 328.400 297.700 ;
        RECT 330.800 298.300 331.600 298.400 ;
        RECT 370.800 298.300 371.600 298.400 ;
        RECT 330.800 297.700 371.600 298.300 ;
        RECT 330.800 297.600 331.600 297.700 ;
        RECT 370.800 297.600 371.600 297.700 ;
        RECT 452.400 298.300 453.200 298.400 ;
        RECT 463.600 298.300 464.400 298.400 ;
        RECT 511.600 298.300 512.400 298.400 ;
        RECT 452.400 297.700 512.400 298.300 ;
        RECT 452.400 297.600 453.200 297.700 ;
        RECT 463.600 297.600 464.400 297.700 ;
        RECT 511.600 297.600 512.400 297.700 ;
        RECT 522.800 298.300 523.600 298.400 ;
        RECT 558.000 298.300 558.800 298.400 ;
        RECT 522.800 297.700 558.800 298.300 ;
        RECT 522.800 297.600 523.600 297.700 ;
        RECT 558.000 297.600 558.800 297.700 ;
        RECT 559.600 298.300 560.400 298.400 ;
        RECT 604.400 298.300 605.200 298.400 ;
        RECT 559.600 297.700 605.200 298.300 ;
        RECT 559.600 297.600 560.400 297.700 ;
        RECT 604.400 297.600 605.200 297.700 ;
        RECT 634.800 298.300 635.600 298.400 ;
        RECT 654.000 298.300 654.800 298.400 ;
        RECT 634.800 297.700 654.800 298.300 ;
        RECT 634.800 297.600 635.600 297.700 ;
        RECT 654.000 297.600 654.800 297.700 ;
        RECT 15.600 296.300 16.400 296.400 ;
        RECT 28.400 296.300 29.200 296.400 ;
        RECT 15.600 295.700 29.200 296.300 ;
        RECT 15.600 295.600 16.400 295.700 ;
        RECT 28.400 295.600 29.200 295.700 ;
        RECT 142.000 296.300 142.800 296.400 ;
        RECT 170.800 296.300 171.600 296.400 ;
        RECT 218.800 296.300 219.600 296.400 ;
        RECT 250.800 296.300 251.600 296.400 ;
        RECT 142.000 295.700 171.600 296.300 ;
        RECT 142.000 295.600 142.800 295.700 ;
        RECT 170.800 295.600 171.600 295.700 ;
        RECT 180.500 295.700 219.600 296.300 ;
        RECT 180.500 294.400 181.100 295.700 ;
        RECT 218.800 295.600 219.600 295.700 ;
        RECT 220.500 295.700 251.600 296.300 ;
        RECT 20.400 294.300 21.200 294.400 ;
        RECT 26.800 294.300 27.600 294.400 ;
        RECT 44.400 294.300 45.200 294.400 ;
        RECT 54.000 294.300 54.800 294.400 ;
        RECT 60.400 294.300 61.200 294.400 ;
        RECT 20.400 293.700 61.200 294.300 ;
        RECT 20.400 293.600 21.200 293.700 ;
        RECT 26.800 293.600 27.600 293.700 ;
        RECT 44.400 293.600 45.200 293.700 ;
        RECT 54.000 293.600 54.800 293.700 ;
        RECT 60.400 293.600 61.200 293.700 ;
        RECT 74.800 294.300 75.600 294.400 ;
        RECT 95.600 294.300 96.400 294.400 ;
        RECT 74.800 293.700 96.400 294.300 ;
        RECT 74.800 293.600 75.600 293.700 ;
        RECT 95.600 293.600 96.400 293.700 ;
        RECT 97.200 294.300 98.000 294.400 ;
        RECT 108.400 294.300 109.200 294.400 ;
        RECT 97.200 293.700 109.200 294.300 ;
        RECT 97.200 293.600 98.000 293.700 ;
        RECT 108.400 293.600 109.200 293.700 ;
        RECT 130.800 294.300 131.600 294.400 ;
        RECT 153.200 294.300 154.000 294.400 ;
        RECT 130.800 293.700 154.000 294.300 ;
        RECT 130.800 293.600 131.600 293.700 ;
        RECT 153.200 293.600 154.000 293.700 ;
        RECT 180.400 293.600 181.200 294.400 ;
        RECT 218.800 294.300 219.600 294.400 ;
        RECT 220.500 294.300 221.100 295.700 ;
        RECT 250.800 295.600 251.600 295.700 ;
        RECT 297.200 296.300 298.000 296.400 ;
        RECT 306.800 296.300 307.600 296.400 ;
        RECT 313.200 296.300 314.000 296.400 ;
        RECT 318.000 296.300 318.800 296.400 ;
        RECT 330.800 296.300 331.600 296.400 ;
        RECT 345.200 296.300 346.000 296.400 ;
        RECT 297.200 295.700 346.000 296.300 ;
        RECT 297.200 295.600 298.000 295.700 ;
        RECT 306.800 295.600 307.600 295.700 ;
        RECT 313.200 295.600 314.000 295.700 ;
        RECT 318.000 295.600 318.800 295.700 ;
        RECT 330.800 295.600 331.600 295.700 ;
        RECT 345.200 295.600 346.000 295.700 ;
        RECT 356.400 296.300 357.200 296.400 ;
        RECT 364.400 296.300 365.200 296.400 ;
        RECT 356.400 295.700 365.200 296.300 ;
        RECT 356.400 295.600 357.200 295.700 ;
        RECT 364.400 295.600 365.200 295.700 ;
        RECT 385.200 296.300 386.000 296.400 ;
        RECT 423.600 296.300 424.400 296.400 ;
        RECT 436.400 296.300 437.200 296.400 ;
        RECT 447.600 296.300 448.400 296.400 ;
        RECT 385.200 295.700 448.400 296.300 ;
        RECT 385.200 295.600 386.000 295.700 ;
        RECT 423.600 295.600 424.400 295.700 ;
        RECT 436.400 295.600 437.200 295.700 ;
        RECT 447.600 295.600 448.400 295.700 ;
        RECT 455.600 296.300 456.400 296.400 ;
        RECT 465.200 296.300 466.000 296.400 ;
        RECT 455.600 295.700 466.000 296.300 ;
        RECT 455.600 295.600 456.400 295.700 ;
        RECT 465.200 295.600 466.000 295.700 ;
        RECT 473.200 296.300 474.000 296.400 ;
        RECT 487.600 296.300 488.400 296.400 ;
        RECT 473.200 295.700 488.400 296.300 ;
        RECT 473.200 295.600 474.000 295.700 ;
        RECT 487.600 295.600 488.400 295.700 ;
        RECT 495.600 296.300 496.400 296.400 ;
        RECT 506.800 296.300 507.600 296.400 ;
        RECT 521.200 296.300 522.000 296.400 ;
        RECT 526.000 296.300 526.800 296.400 ;
        RECT 495.600 295.700 526.800 296.300 ;
        RECT 495.600 295.600 496.400 295.700 ;
        RECT 506.800 295.600 507.600 295.700 ;
        RECT 521.200 295.600 522.000 295.700 ;
        RECT 526.000 295.600 526.800 295.700 ;
        RECT 553.200 296.300 554.000 296.400 ;
        RECT 620.400 296.300 621.200 296.400 ;
        RECT 553.200 295.700 621.200 296.300 ;
        RECT 553.200 295.600 554.000 295.700 ;
        RECT 620.400 295.600 621.200 295.700 ;
        RECT 625.200 296.300 626.000 296.400 ;
        RECT 631.600 296.300 632.400 296.400 ;
        RECT 625.200 295.700 632.400 296.300 ;
        RECT 625.200 295.600 626.000 295.700 ;
        RECT 631.600 295.600 632.400 295.700 ;
        RECT 633.200 296.300 634.000 296.400 ;
        RECT 636.400 296.300 637.200 296.400 ;
        RECT 650.800 296.300 651.600 296.400 ;
        RECT 633.200 295.700 651.600 296.300 ;
        RECT 633.200 295.600 634.000 295.700 ;
        RECT 636.400 295.600 637.200 295.700 ;
        RECT 650.800 295.600 651.600 295.700 ;
        RECT 218.800 293.700 221.100 294.300 ;
        RECT 241.200 294.300 242.000 294.400 ;
        RECT 244.400 294.300 245.200 294.400 ;
        RECT 241.200 293.700 245.200 294.300 ;
        RECT 218.800 293.600 219.600 293.700 ;
        RECT 241.200 293.600 242.000 293.700 ;
        RECT 244.400 293.600 245.200 293.700 ;
        RECT 271.600 294.300 272.400 294.400 ;
        RECT 279.600 294.300 280.400 294.400 ;
        RECT 271.600 293.700 280.400 294.300 ;
        RECT 271.600 293.600 272.400 293.700 ;
        RECT 279.600 293.600 280.400 293.700 ;
        RECT 314.800 294.300 315.600 294.400 ;
        RECT 322.800 294.300 323.600 294.400 ;
        RECT 314.800 293.700 323.600 294.300 ;
        RECT 314.800 293.600 315.600 293.700 ;
        RECT 322.800 293.600 323.600 293.700 ;
        RECT 327.600 294.300 328.400 294.400 ;
        RECT 332.400 294.300 333.200 294.400 ;
        RECT 327.600 293.700 333.200 294.300 ;
        RECT 327.600 293.600 328.400 293.700 ;
        RECT 332.400 293.600 333.200 293.700 ;
        RECT 335.600 294.300 336.400 294.400 ;
        RECT 345.200 294.300 346.000 294.400 ;
        RECT 335.600 293.700 346.000 294.300 ;
        RECT 335.600 293.600 336.400 293.700 ;
        RECT 345.200 293.600 346.000 293.700 ;
        RECT 359.600 294.300 360.400 294.400 ;
        RECT 388.400 294.300 389.200 294.400 ;
        RECT 359.600 293.700 389.200 294.300 ;
        RECT 359.600 293.600 360.400 293.700 ;
        RECT 388.400 293.600 389.200 293.700 ;
        RECT 433.200 294.300 434.000 294.400 ;
        RECT 454.000 294.300 454.800 294.400 ;
        RECT 433.200 293.700 454.800 294.300 ;
        RECT 433.200 293.600 434.000 293.700 ;
        RECT 454.000 293.600 454.800 293.700 ;
        RECT 465.200 294.300 466.000 294.400 ;
        RECT 468.400 294.300 469.200 294.400 ;
        RECT 465.200 293.700 469.200 294.300 ;
        RECT 465.200 293.600 466.000 293.700 ;
        RECT 468.400 293.600 469.200 293.700 ;
        RECT 479.600 294.300 480.400 294.400 ;
        RECT 482.800 294.300 483.600 294.400 ;
        RECT 479.600 293.700 483.600 294.300 ;
        RECT 479.600 293.600 480.400 293.700 ;
        RECT 482.800 293.600 483.600 293.700 ;
        RECT 486.000 294.300 486.800 294.400 ;
        RECT 497.200 294.300 498.000 294.400 ;
        RECT 486.000 293.700 498.000 294.300 ;
        RECT 486.000 293.600 486.800 293.700 ;
        RECT 497.200 293.600 498.000 293.700 ;
        RECT 516.400 294.300 517.200 294.400 ;
        RECT 519.600 294.300 520.400 294.400 ;
        RECT 516.400 293.700 520.400 294.300 ;
        RECT 516.400 293.600 517.200 293.700 ;
        RECT 519.600 293.600 520.400 293.700 ;
        RECT 530.800 294.300 531.600 294.400 ;
        RECT 534.000 294.300 534.800 294.400 ;
        RECT 530.800 293.700 534.800 294.300 ;
        RECT 530.800 293.600 531.600 293.700 ;
        RECT 534.000 293.600 534.800 293.700 ;
        RECT 569.200 294.300 570.000 294.400 ;
        RECT 578.800 294.300 579.600 294.400 ;
        RECT 569.200 293.700 579.600 294.300 ;
        RECT 569.200 293.600 570.000 293.700 ;
        RECT 578.800 293.600 579.600 293.700 ;
        RECT 580.400 294.300 581.200 294.400 ;
        RECT 593.200 294.300 594.000 294.400 ;
        RECT 607.600 294.300 608.400 294.400 ;
        RECT 580.400 293.700 608.400 294.300 ;
        RECT 580.400 293.600 581.200 293.700 ;
        RECT 593.200 293.600 594.000 293.700 ;
        RECT 607.600 293.600 608.400 293.700 ;
        RECT 610.800 294.300 611.600 294.400 ;
        RECT 622.000 294.300 622.800 294.400 ;
        RECT 639.600 294.300 640.400 294.400 ;
        RECT 646.000 294.300 646.800 294.400 ;
        RECT 657.200 294.300 658.000 294.400 ;
        RECT 610.800 293.700 658.000 294.300 ;
        RECT 610.800 293.600 611.600 293.700 ;
        RECT 622.000 293.600 622.800 293.700 ;
        RECT 639.600 293.600 640.400 293.700 ;
        RECT 646.000 293.600 646.800 293.700 ;
        RECT 657.200 293.600 658.000 293.700 ;
        RECT 670.000 293.600 670.800 294.400 ;
        RECT 2.800 292.300 3.600 292.400 ;
        RECT 14.000 292.300 14.800 292.400 ;
        RECT 30.000 292.300 30.800 292.400 ;
        RECT 34.800 292.300 35.600 292.400 ;
        RECT 2.800 291.700 35.600 292.300 ;
        RECT 2.800 291.600 3.600 291.700 ;
        RECT 14.000 291.600 14.800 291.700 ;
        RECT 30.000 291.600 30.800 291.700 ;
        RECT 34.800 291.600 35.600 291.700 ;
        RECT 42.800 292.300 43.600 292.400 ;
        RECT 47.600 292.300 48.400 292.400 ;
        RECT 42.800 291.700 48.400 292.300 ;
        RECT 42.800 291.600 43.600 291.700 ;
        RECT 47.600 291.600 48.400 291.700 ;
        RECT 60.400 292.300 61.200 292.400 ;
        RECT 102.000 292.300 102.800 292.400 ;
        RECT 60.400 291.700 102.800 292.300 ;
        RECT 60.400 291.600 61.200 291.700 ;
        RECT 102.000 291.600 102.800 291.700 ;
        RECT 105.200 292.300 106.000 292.400 ;
        RECT 161.200 292.300 162.000 292.400 ;
        RECT 105.200 291.700 162.000 292.300 ;
        RECT 105.200 291.600 106.000 291.700 ;
        RECT 161.200 291.600 162.000 291.700 ;
        RECT 321.200 292.300 322.000 292.400 ;
        RECT 375.600 292.300 376.400 292.400 ;
        RECT 378.800 292.300 379.600 292.400 ;
        RECT 321.200 291.700 379.600 292.300 ;
        RECT 321.200 291.600 322.000 291.700 ;
        RECT 375.600 291.600 376.400 291.700 ;
        RECT 378.800 291.600 379.600 291.700 ;
        RECT 404.400 291.600 405.200 292.400 ;
        RECT 476.400 292.300 477.200 292.400 ;
        RECT 482.800 292.300 483.600 292.400 ;
        RECT 476.400 291.700 483.600 292.300 ;
        RECT 476.400 291.600 477.200 291.700 ;
        RECT 482.800 291.600 483.600 291.700 ;
        RECT 486.000 292.300 486.800 292.400 ;
        RECT 498.800 292.300 499.600 292.400 ;
        RECT 486.000 291.700 499.600 292.300 ;
        RECT 486.000 291.600 486.800 291.700 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 518.000 292.300 518.800 292.400 ;
        RECT 522.800 292.300 523.600 292.400 ;
        RECT 532.400 292.300 533.200 292.400 ;
        RECT 518.000 291.700 533.200 292.300 ;
        RECT 518.000 291.600 518.800 291.700 ;
        RECT 522.800 291.600 523.600 291.700 ;
        RECT 532.400 291.600 533.200 291.700 ;
        RECT 545.200 292.300 546.000 292.400 ;
        RECT 602.800 292.300 603.600 292.400 ;
        RECT 617.200 292.300 618.000 292.400 ;
        RECT 623.600 292.300 624.400 292.400 ;
        RECT 545.200 291.700 624.400 292.300 ;
        RECT 545.200 291.600 546.000 291.700 ;
        RECT 602.800 291.600 603.600 291.700 ;
        RECT 617.200 291.600 618.000 291.700 ;
        RECT 623.600 291.600 624.400 291.700 ;
        RECT 6.000 290.300 6.800 290.400 ;
        RECT 38.000 290.300 38.800 290.400 ;
        RECT 6.000 289.700 38.800 290.300 ;
        RECT 6.000 289.600 6.800 289.700 ;
        RECT 38.000 289.600 38.800 289.700 ;
        RECT 94.000 290.300 94.800 290.400 ;
        RECT 100.400 290.300 101.200 290.400 ;
        RECT 94.000 289.700 101.200 290.300 ;
        RECT 94.000 289.600 94.800 289.700 ;
        RECT 100.400 289.600 101.200 289.700 ;
        RECT 106.800 290.300 107.600 290.400 ;
        RECT 151.600 290.300 152.400 290.400 ;
        RECT 180.400 290.300 181.200 290.400 ;
        RECT 106.800 289.700 181.200 290.300 ;
        RECT 106.800 289.600 107.600 289.700 ;
        RECT 151.600 289.600 152.400 289.700 ;
        RECT 180.400 289.600 181.200 289.700 ;
        RECT 196.400 290.300 197.200 290.400 ;
        RECT 204.400 290.300 205.200 290.400 ;
        RECT 196.400 289.700 205.200 290.300 ;
        RECT 196.400 289.600 197.200 289.700 ;
        RECT 204.400 289.600 205.200 289.700 ;
        RECT 218.800 290.300 219.600 290.400 ;
        RECT 238.000 290.300 238.800 290.400 ;
        RECT 218.800 289.700 238.800 290.300 ;
        RECT 218.800 289.600 219.600 289.700 ;
        RECT 238.000 289.600 238.800 289.700 ;
        RECT 252.400 290.300 253.200 290.400 ;
        RECT 289.200 290.300 290.000 290.400 ;
        RECT 252.400 289.700 290.000 290.300 ;
        RECT 252.400 289.600 253.200 289.700 ;
        RECT 289.200 289.600 290.000 289.700 ;
        RECT 321.200 290.300 322.000 290.400 ;
        RECT 324.400 290.300 325.200 290.400 ;
        RECT 321.200 289.700 325.200 290.300 ;
        RECT 321.200 289.600 322.000 289.700 ;
        RECT 324.400 289.600 325.200 289.700 ;
        RECT 329.200 290.300 330.000 290.400 ;
        RECT 332.400 290.300 333.200 290.400 ;
        RECT 329.200 289.700 333.200 290.300 ;
        RECT 329.200 289.600 330.000 289.700 ;
        RECT 332.400 289.600 333.200 289.700 ;
        RECT 337.200 290.300 338.000 290.400 ;
        RECT 346.800 290.300 347.600 290.400 ;
        RECT 337.200 289.700 347.600 290.300 ;
        RECT 337.200 289.600 338.000 289.700 ;
        RECT 346.800 289.600 347.600 289.700 ;
        RECT 470.000 290.300 470.800 290.400 ;
        RECT 471.600 290.300 472.400 290.400 ;
        RECT 470.000 289.700 472.400 290.300 ;
        RECT 470.000 289.600 470.800 289.700 ;
        RECT 471.600 289.600 472.400 289.700 ;
        RECT 474.800 290.300 475.600 290.400 ;
        RECT 583.600 290.300 584.400 290.400 ;
        RECT 615.600 290.300 616.400 290.400 ;
        RECT 474.800 289.700 616.400 290.300 ;
        RECT 474.800 289.600 475.600 289.700 ;
        RECT 583.600 289.600 584.400 289.700 ;
        RECT 615.600 289.600 616.400 289.700 ;
        RECT 620.400 290.300 621.200 290.400 ;
        RECT 625.200 290.300 626.000 290.400 ;
        RECT 620.400 289.700 626.000 290.300 ;
        RECT 620.400 289.600 621.200 289.700 ;
        RECT 625.200 289.600 626.000 289.700 ;
        RECT 670.000 290.300 670.800 290.400 ;
        RECT 676.400 290.300 677.200 290.400 ;
        RECT 670.000 289.700 677.200 290.300 ;
        RECT 670.000 289.600 670.800 289.700 ;
        RECT 676.400 289.600 677.200 289.700 ;
        RECT 10.800 288.300 11.600 288.400 ;
        RECT 17.200 288.300 18.000 288.400 ;
        RECT 10.800 287.700 18.000 288.300 ;
        RECT 10.800 287.600 11.600 287.700 ;
        RECT 17.200 287.600 18.000 287.700 ;
        RECT 33.200 288.300 34.000 288.400 ;
        RECT 42.800 288.300 43.600 288.400 ;
        RECT 33.200 287.700 43.600 288.300 ;
        RECT 33.200 287.600 34.000 287.700 ;
        RECT 42.800 287.600 43.600 287.700 ;
        RECT 52.400 288.300 53.200 288.400 ;
        RECT 105.200 288.300 106.000 288.400 ;
        RECT 52.400 287.700 106.000 288.300 ;
        RECT 52.400 287.600 53.200 287.700 ;
        RECT 105.200 287.600 106.000 287.700 ;
        RECT 150.000 288.300 150.800 288.400 ;
        RECT 156.400 288.300 157.200 288.400 ;
        RECT 150.000 287.700 157.200 288.300 ;
        RECT 150.000 287.600 150.800 287.700 ;
        RECT 156.400 287.600 157.200 287.700 ;
        RECT 322.800 288.300 323.600 288.400 ;
        RECT 343.600 288.300 344.400 288.400 ;
        RECT 322.800 287.700 344.400 288.300 ;
        RECT 322.800 287.600 323.600 287.700 ;
        RECT 343.600 287.600 344.400 287.700 ;
        RECT 351.600 288.300 352.400 288.400 ;
        RECT 406.000 288.300 406.800 288.400 ;
        RECT 351.600 287.700 406.800 288.300 ;
        RECT 351.600 287.600 352.400 287.700 ;
        RECT 406.000 287.600 406.800 287.700 ;
        RECT 471.600 288.300 472.400 288.400 ;
        RECT 511.600 288.300 512.400 288.400 ;
        RECT 562.800 288.300 563.600 288.400 ;
        RECT 471.600 287.700 563.600 288.300 ;
        RECT 471.600 287.600 472.400 287.700 ;
        RECT 511.600 287.600 512.400 287.700 ;
        RECT 562.800 287.600 563.600 287.700 ;
        RECT 586.800 288.300 587.600 288.400 ;
        RECT 598.000 288.300 598.800 288.400 ;
        RECT 586.800 287.700 598.800 288.300 ;
        RECT 615.700 288.300 616.300 289.600 ;
        RECT 641.200 288.300 642.000 288.400 ;
        RECT 652.400 288.300 653.200 288.400 ;
        RECT 615.700 287.700 653.200 288.300 ;
        RECT 586.800 287.600 587.600 287.700 ;
        RECT 598.000 287.600 598.800 287.700 ;
        RECT 641.200 287.600 642.000 287.700 ;
        RECT 652.400 287.600 653.200 287.700 ;
        RECT 78.000 286.300 78.800 286.400 ;
        RECT 119.600 286.300 120.400 286.400 ;
        RECT 134.000 286.300 134.800 286.400 ;
        RECT 153.200 286.300 154.000 286.400 ;
        RECT 78.000 285.700 154.000 286.300 ;
        RECT 78.000 285.600 78.800 285.700 ;
        RECT 119.600 285.600 120.400 285.700 ;
        RECT 134.000 285.600 134.800 285.700 ;
        RECT 153.200 285.600 154.000 285.700 ;
        RECT 242.800 286.300 243.600 286.400 ;
        RECT 361.200 286.300 362.000 286.400 ;
        RECT 372.400 286.300 373.200 286.400 ;
        RECT 242.800 285.700 373.200 286.300 ;
        RECT 242.800 285.600 243.600 285.700 ;
        RECT 361.200 285.600 362.000 285.700 ;
        RECT 372.400 285.600 373.200 285.700 ;
        RECT 564.400 286.300 565.200 286.400 ;
        RECT 602.800 286.300 603.600 286.400 ;
        RECT 564.400 285.700 603.600 286.300 ;
        RECT 564.400 285.600 565.200 285.700 ;
        RECT 602.800 285.600 603.600 285.700 ;
        RECT 614.000 286.300 614.800 286.400 ;
        RECT 625.200 286.300 626.000 286.400 ;
        RECT 614.000 285.700 626.000 286.300 ;
        RECT 614.000 285.600 614.800 285.700 ;
        RECT 625.200 285.600 626.000 285.700 ;
        RECT 87.600 284.300 88.400 284.400 ;
        RECT 132.400 284.300 133.200 284.400 ;
        RECT 87.600 283.700 133.200 284.300 ;
        RECT 87.600 283.600 88.400 283.700 ;
        RECT 132.400 283.600 133.200 283.700 ;
        RECT 161.200 284.300 162.000 284.400 ;
        RECT 178.800 284.300 179.600 284.400 ;
        RECT 201.200 284.300 202.000 284.400 ;
        RECT 215.600 284.300 216.400 284.400 ;
        RECT 223.600 284.300 224.400 284.400 ;
        RECT 161.200 283.700 224.400 284.300 ;
        RECT 161.200 283.600 162.000 283.700 ;
        RECT 178.800 283.600 179.600 283.700 ;
        RECT 201.200 283.600 202.000 283.700 ;
        RECT 215.600 283.600 216.400 283.700 ;
        RECT 223.600 283.600 224.400 283.700 ;
        RECT 326.000 284.300 326.800 284.400 ;
        RECT 346.800 284.300 347.600 284.400 ;
        RECT 326.000 283.700 347.600 284.300 ;
        RECT 326.000 283.600 326.800 283.700 ;
        RECT 346.800 283.600 347.600 283.700 ;
        RECT 348.400 284.300 349.200 284.400 ;
        RECT 375.600 284.300 376.400 284.400 ;
        RECT 348.400 283.700 376.400 284.300 ;
        RECT 348.400 283.600 349.200 283.700 ;
        RECT 375.600 283.600 376.400 283.700 ;
        RECT 502.000 284.300 502.800 284.400 ;
        RECT 556.400 284.300 557.200 284.400 ;
        RECT 502.000 283.700 557.200 284.300 ;
        RECT 502.000 283.600 502.800 283.700 ;
        RECT 556.400 283.600 557.200 283.700 ;
        RECT 596.400 284.300 597.200 284.400 ;
        RECT 599.600 284.300 600.400 284.400 ;
        RECT 609.200 284.300 610.000 284.400 ;
        RECT 596.400 283.700 610.000 284.300 ;
        RECT 596.400 283.600 597.200 283.700 ;
        RECT 599.600 283.600 600.400 283.700 ;
        RECT 609.200 283.600 610.000 283.700 ;
        RECT 628.400 284.300 629.200 284.400 ;
        RECT 634.800 284.300 635.600 284.400 ;
        RECT 628.400 283.700 635.600 284.300 ;
        RECT 628.400 283.600 629.200 283.700 ;
        RECT 634.800 283.600 635.600 283.700 ;
        RECT 204.400 282.300 205.200 282.400 ;
        RECT 278.000 282.300 278.800 282.400 ;
        RECT 204.400 281.700 278.800 282.300 ;
        RECT 204.400 281.600 205.200 281.700 ;
        RECT 278.000 281.600 278.800 281.700 ;
        RECT 308.400 282.300 309.200 282.400 ;
        RECT 340.400 282.300 341.200 282.400 ;
        RECT 308.400 281.700 341.200 282.300 ;
        RECT 308.400 281.600 309.200 281.700 ;
        RECT 340.400 281.600 341.200 281.700 ;
        RECT 342.000 282.300 342.800 282.400 ;
        RECT 398.000 282.300 398.800 282.400 ;
        RECT 342.000 281.700 398.800 282.300 ;
        RECT 342.000 281.600 342.800 281.700 ;
        RECT 398.000 281.600 398.800 281.700 ;
        RECT 510.000 282.300 510.800 282.400 ;
        RECT 532.400 282.300 533.200 282.400 ;
        RECT 599.600 282.300 600.400 282.400 ;
        RECT 510.000 281.700 600.400 282.300 ;
        RECT 510.000 281.600 510.800 281.700 ;
        RECT 532.400 281.600 533.200 281.700 ;
        RECT 599.600 281.600 600.400 281.700 ;
        RECT 650.800 282.300 651.600 282.400 ;
        RECT 658.800 282.300 659.600 282.400 ;
        RECT 650.800 281.700 659.600 282.300 ;
        RECT 650.800 281.600 651.600 281.700 ;
        RECT 658.800 281.600 659.600 281.700 ;
        RECT 154.800 280.300 155.600 280.400 ;
        RECT 170.800 280.300 171.600 280.400 ;
        RECT 154.800 279.700 171.600 280.300 ;
        RECT 154.800 279.600 155.600 279.700 ;
        RECT 170.800 279.600 171.600 279.700 ;
        RECT 185.200 280.300 186.000 280.400 ;
        RECT 242.800 280.300 243.600 280.400 ;
        RECT 185.200 279.700 243.600 280.300 ;
        RECT 185.200 279.600 186.000 279.700 ;
        RECT 242.800 279.600 243.600 279.700 ;
        RECT 282.800 280.300 283.600 280.400 ;
        RECT 300.400 280.300 301.200 280.400 ;
        RECT 282.800 279.700 301.200 280.300 ;
        RECT 282.800 279.600 283.600 279.700 ;
        RECT 300.400 279.600 301.200 279.700 ;
        RECT 314.800 280.300 315.600 280.400 ;
        RECT 346.800 280.300 347.600 280.400 ;
        RECT 314.800 279.700 347.600 280.300 ;
        RECT 314.800 279.600 315.600 279.700 ;
        RECT 346.800 279.600 347.600 279.700 ;
        RECT 350.000 279.600 350.800 280.400 ;
        RECT 481.200 280.300 482.000 280.400 ;
        RECT 506.800 280.300 507.600 280.400 ;
        RECT 529.200 280.300 530.000 280.400 ;
        RECT 481.200 279.700 530.000 280.300 ;
        RECT 481.200 279.600 482.000 279.700 ;
        RECT 506.800 279.600 507.600 279.700 ;
        RECT 529.200 279.600 530.000 279.700 ;
        RECT 542.000 280.300 542.800 280.400 ;
        RECT 561.200 280.300 562.000 280.400 ;
        RECT 542.000 279.700 562.000 280.300 ;
        RECT 542.000 279.600 542.800 279.700 ;
        RECT 561.200 279.600 562.000 279.700 ;
        RECT 586.800 280.300 587.600 280.400 ;
        RECT 591.600 280.300 592.400 280.400 ;
        RECT 658.800 280.300 659.600 280.400 ;
        RECT 586.800 279.700 659.600 280.300 ;
        RECT 586.800 279.600 587.600 279.700 ;
        RECT 591.600 279.600 592.400 279.700 ;
        RECT 658.800 279.600 659.600 279.700 ;
        RECT 17.200 278.300 18.000 278.400 ;
        RECT 33.200 278.300 34.000 278.400 ;
        RECT 17.200 277.700 34.000 278.300 ;
        RECT 17.200 277.600 18.000 277.700 ;
        RECT 33.200 277.600 34.000 277.700 ;
        RECT 47.600 278.300 48.400 278.400 ;
        RECT 68.400 278.300 69.200 278.400 ;
        RECT 47.600 277.700 69.200 278.300 ;
        RECT 47.600 277.600 48.400 277.700 ;
        RECT 68.400 277.600 69.200 277.700 ;
        RECT 158.000 277.600 158.800 278.400 ;
        RECT 238.000 278.300 238.800 278.400 ;
        RECT 247.600 278.300 248.400 278.400 ;
        RECT 238.000 277.700 248.400 278.300 ;
        RECT 238.000 277.600 238.800 277.700 ;
        RECT 247.600 277.600 248.400 277.700 ;
        RECT 274.800 278.300 275.600 278.400 ;
        RECT 310.000 278.300 310.800 278.400 ;
        RECT 274.800 277.700 310.800 278.300 ;
        RECT 274.800 277.600 275.600 277.700 ;
        RECT 310.000 277.600 310.800 277.700 ;
        RECT 343.600 278.300 344.400 278.400 ;
        RECT 358.000 278.300 358.800 278.400 ;
        RECT 343.600 277.700 358.800 278.300 ;
        RECT 343.600 277.600 344.400 277.700 ;
        RECT 358.000 277.600 358.800 277.700 ;
        RECT 362.800 278.300 363.600 278.400 ;
        RECT 378.800 278.300 379.600 278.400 ;
        RECT 402.800 278.300 403.600 278.400 ;
        RECT 409.200 278.300 410.000 278.400 ;
        RECT 455.600 278.300 456.400 278.400 ;
        RECT 362.800 277.700 456.400 278.300 ;
        RECT 362.800 277.600 363.600 277.700 ;
        RECT 378.800 277.600 379.600 277.700 ;
        RECT 402.800 277.600 403.600 277.700 ;
        RECT 409.200 277.600 410.000 277.700 ;
        RECT 455.600 277.600 456.400 277.700 ;
        RECT 534.000 278.300 534.800 278.400 ;
        RECT 548.400 278.300 549.200 278.400 ;
        RECT 558.000 278.300 558.800 278.400 ;
        RECT 534.000 277.700 558.800 278.300 ;
        RECT 534.000 277.600 534.800 277.700 ;
        RECT 548.400 277.600 549.200 277.700 ;
        RECT 558.000 277.600 558.800 277.700 ;
        RECT 572.400 278.300 573.200 278.400 ;
        RECT 628.400 278.300 629.200 278.400 ;
        RECT 572.400 277.700 629.200 278.300 ;
        RECT 572.400 277.600 573.200 277.700 ;
        RECT 628.400 277.600 629.200 277.700 ;
        RECT 156.400 276.300 157.200 276.400 ;
        RECT 314.800 276.300 315.600 276.400 ;
        RECT 156.400 275.700 315.600 276.300 ;
        RECT 156.400 275.600 157.200 275.700 ;
        RECT 314.800 275.600 315.600 275.700 ;
        RECT 319.600 276.300 320.400 276.400 ;
        RECT 334.000 276.300 334.800 276.400 ;
        RECT 342.000 276.300 342.800 276.400 ;
        RECT 319.600 275.700 342.800 276.300 ;
        RECT 319.600 275.600 320.400 275.700 ;
        RECT 334.000 275.600 334.800 275.700 ;
        RECT 342.000 275.600 342.800 275.700 ;
        RECT 345.200 276.300 346.000 276.400 ;
        RECT 366.000 276.300 366.800 276.400 ;
        RECT 382.000 276.300 382.800 276.400 ;
        RECT 345.200 275.700 382.800 276.300 ;
        RECT 345.200 275.600 346.000 275.700 ;
        RECT 366.000 275.600 366.800 275.700 ;
        RECT 382.000 275.600 382.800 275.700 ;
        RECT 583.600 276.300 584.400 276.400 ;
        RECT 617.200 276.300 618.000 276.400 ;
        RECT 583.600 275.700 618.000 276.300 ;
        RECT 583.600 275.600 584.400 275.700 ;
        RECT 617.200 275.600 618.000 275.700 ;
        RECT 630.000 276.300 630.800 276.400 ;
        RECT 657.200 276.300 658.000 276.400 ;
        RECT 666.800 276.300 667.600 276.400 ;
        RECT 630.000 275.700 667.600 276.300 ;
        RECT 630.000 275.600 630.800 275.700 ;
        RECT 657.200 275.600 658.000 275.700 ;
        RECT 666.800 275.600 667.600 275.700 ;
        RECT 100.400 274.300 101.200 274.400 ;
        RECT 233.200 274.300 234.000 274.400 ;
        RECT 100.400 273.700 234.000 274.300 ;
        RECT 100.400 273.600 101.200 273.700 ;
        RECT 233.200 273.600 234.000 273.700 ;
        RECT 276.400 274.300 277.200 274.400 ;
        RECT 297.200 274.300 298.000 274.400 ;
        RECT 276.400 273.700 298.000 274.300 ;
        RECT 276.400 273.600 277.200 273.700 ;
        RECT 297.200 273.600 298.000 273.700 ;
        RECT 340.400 274.300 341.200 274.400 ;
        RECT 362.800 274.300 363.600 274.400 ;
        RECT 340.400 273.700 363.600 274.300 ;
        RECT 340.400 273.600 341.200 273.700 ;
        RECT 362.800 273.600 363.600 273.700 ;
        RECT 406.000 274.300 406.800 274.400 ;
        RECT 410.800 274.300 411.600 274.400 ;
        RECT 406.000 273.700 411.600 274.300 ;
        RECT 406.000 273.600 406.800 273.700 ;
        RECT 410.800 273.600 411.600 273.700 ;
        RECT 519.600 274.300 520.400 274.400 ;
        RECT 546.800 274.300 547.600 274.400 ;
        RECT 519.600 273.700 547.600 274.300 ;
        RECT 519.600 273.600 520.400 273.700 ;
        RECT 546.800 273.600 547.600 273.700 ;
        RECT 604.400 274.300 605.200 274.400 ;
        RECT 634.800 274.300 635.600 274.400 ;
        RECT 638.000 274.300 638.800 274.400 ;
        RECT 604.400 273.700 638.800 274.300 ;
        RECT 604.400 273.600 605.200 273.700 ;
        RECT 634.800 273.600 635.600 273.700 ;
        RECT 638.000 273.600 638.800 273.700 ;
        RECT 646.000 274.300 646.800 274.400 ;
        RECT 660.400 274.300 661.200 274.400 ;
        RECT 646.000 273.700 661.200 274.300 ;
        RECT 646.000 273.600 646.800 273.700 ;
        RECT 660.400 273.600 661.200 273.700 ;
        RECT 663.600 274.300 664.400 274.400 ;
        RECT 676.400 274.300 677.200 274.400 ;
        RECT 663.600 273.700 677.200 274.300 ;
        RECT 663.600 273.600 664.400 273.700 ;
        RECT 676.400 273.600 677.200 273.700 ;
        RECT 58.800 272.300 59.600 272.400 ;
        RECT 65.200 272.300 66.000 272.400 ;
        RECT 58.800 271.700 66.000 272.300 ;
        RECT 58.800 271.600 59.600 271.700 ;
        RECT 65.200 271.600 66.000 271.700 ;
        RECT 108.400 272.300 109.200 272.400 ;
        RECT 137.200 272.300 138.000 272.400 ;
        RECT 174.000 272.300 174.800 272.400 ;
        RECT 108.400 271.700 174.800 272.300 ;
        RECT 108.400 271.600 109.200 271.700 ;
        RECT 137.200 271.600 138.000 271.700 ;
        RECT 174.000 271.600 174.800 271.700 ;
        RECT 274.800 272.300 275.600 272.400 ;
        RECT 281.200 272.300 282.000 272.400 ;
        RECT 274.800 271.700 282.000 272.300 ;
        RECT 274.800 271.600 275.600 271.700 ;
        RECT 281.200 271.600 282.000 271.700 ;
        RECT 292.400 271.600 293.200 272.400 ;
        RECT 340.400 272.300 341.200 272.400 ;
        RECT 359.600 272.300 360.400 272.400 ;
        RECT 340.400 271.700 360.400 272.300 ;
        RECT 340.400 271.600 341.200 271.700 ;
        RECT 359.600 271.600 360.400 271.700 ;
        RECT 361.200 272.300 362.000 272.400 ;
        RECT 377.200 272.300 378.000 272.400 ;
        RECT 361.200 271.700 378.000 272.300 ;
        RECT 361.200 271.600 362.000 271.700 ;
        RECT 377.200 271.600 378.000 271.700 ;
        RECT 527.600 272.300 528.400 272.400 ;
        RECT 538.800 272.300 539.600 272.400 ;
        RECT 527.600 271.700 539.600 272.300 ;
        RECT 527.600 271.600 528.400 271.700 ;
        RECT 538.800 271.600 539.600 271.700 ;
        RECT 559.600 272.300 560.400 272.400 ;
        RECT 623.600 272.300 624.400 272.400 ;
        RECT 626.800 272.300 627.600 272.400 ;
        RECT 559.600 271.700 627.600 272.300 ;
        RECT 559.600 271.600 560.400 271.700 ;
        RECT 623.600 271.600 624.400 271.700 ;
        RECT 626.800 271.600 627.600 271.700 ;
        RECT 639.600 272.300 640.400 272.400 ;
        RECT 641.200 272.300 642.000 272.400 ;
        RECT 646.000 272.300 646.800 272.400 ;
        RECT 639.600 271.700 646.800 272.300 ;
        RECT 639.600 271.600 640.400 271.700 ;
        RECT 641.200 271.600 642.000 271.700 ;
        RECT 646.000 271.600 646.800 271.700 ;
        RECT 654.000 272.300 654.800 272.400 ;
        RECT 663.600 272.300 664.400 272.400 ;
        RECT 654.000 271.700 664.400 272.300 ;
        RECT 654.000 271.600 654.800 271.700 ;
        RECT 663.600 271.600 664.400 271.700 ;
        RECT 38.000 270.300 38.800 270.400 ;
        RECT 87.600 270.300 88.400 270.400 ;
        RECT 38.000 269.700 88.400 270.300 ;
        RECT 38.000 269.600 38.800 269.700 ;
        RECT 87.600 269.600 88.400 269.700 ;
        RECT 111.600 270.300 112.400 270.400 ;
        RECT 190.000 270.300 190.800 270.400 ;
        RECT 111.600 269.700 190.800 270.300 ;
        RECT 111.600 269.600 112.400 269.700 ;
        RECT 190.000 269.600 190.800 269.700 ;
        RECT 218.800 270.300 219.600 270.400 ;
        RECT 231.600 270.300 232.400 270.400 ;
        RECT 218.800 269.700 232.400 270.300 ;
        RECT 218.800 269.600 219.600 269.700 ;
        RECT 231.600 269.600 232.400 269.700 ;
        RECT 258.800 270.300 259.600 270.400 ;
        RECT 260.400 270.300 261.200 270.400 ;
        RECT 271.600 270.300 272.400 270.400 ;
        RECT 297.200 270.300 298.000 270.400 ;
        RECT 258.800 269.700 298.000 270.300 ;
        RECT 258.800 269.600 259.600 269.700 ;
        RECT 260.400 269.600 261.200 269.700 ;
        RECT 271.600 269.600 272.400 269.700 ;
        RECT 297.200 269.600 298.000 269.700 ;
        RECT 310.000 270.300 310.800 270.400 ;
        RECT 340.400 270.300 341.200 270.400 ;
        RECT 310.000 269.700 341.200 270.300 ;
        RECT 310.000 269.600 310.800 269.700 ;
        RECT 340.400 269.600 341.200 269.700 ;
        RECT 342.000 270.300 342.800 270.400 ;
        RECT 375.600 270.300 376.400 270.400 ;
        RECT 342.000 269.700 376.400 270.300 ;
        RECT 342.000 269.600 342.800 269.700 ;
        RECT 375.600 269.600 376.400 269.700 ;
        RECT 378.800 270.300 379.600 270.400 ;
        RECT 385.200 270.300 386.000 270.400 ;
        RECT 386.800 270.300 387.600 270.400 ;
        RECT 378.800 269.700 387.600 270.300 ;
        RECT 378.800 269.600 379.600 269.700 ;
        RECT 385.200 269.600 386.000 269.700 ;
        RECT 386.800 269.600 387.600 269.700 ;
        RECT 450.800 270.300 451.600 270.400 ;
        RECT 468.400 270.300 469.200 270.400 ;
        RECT 450.800 269.700 469.200 270.300 ;
        RECT 450.800 269.600 451.600 269.700 ;
        RECT 468.400 269.600 469.200 269.700 ;
        RECT 514.800 270.300 515.600 270.400 ;
        RECT 524.400 270.300 525.200 270.400 ;
        RECT 514.800 269.700 525.200 270.300 ;
        RECT 514.800 269.600 515.600 269.700 ;
        RECT 524.400 269.600 525.200 269.700 ;
        RECT 538.800 270.300 539.600 270.400 ;
        RECT 545.200 270.300 546.000 270.400 ;
        RECT 538.800 269.700 546.000 270.300 ;
        RECT 538.800 269.600 539.600 269.700 ;
        RECT 545.200 269.600 546.000 269.700 ;
        RECT 562.800 270.300 563.600 270.400 ;
        RECT 580.400 270.300 581.200 270.400 ;
        RECT 562.800 269.700 581.200 270.300 ;
        RECT 562.800 269.600 563.600 269.700 ;
        RECT 580.400 269.600 581.200 269.700 ;
        RECT 593.200 270.300 594.000 270.400 ;
        RECT 607.600 270.300 608.400 270.400 ;
        RECT 636.400 270.300 637.200 270.400 ;
        RECT 644.400 270.300 645.200 270.400 ;
        RECT 593.200 269.700 645.200 270.300 ;
        RECT 593.200 269.600 594.000 269.700 ;
        RECT 607.600 269.600 608.400 269.700 ;
        RECT 636.400 269.600 637.200 269.700 ;
        RECT 644.400 269.600 645.200 269.700 ;
        RECT 649.200 270.300 650.000 270.400 ;
        RECT 657.200 270.300 658.000 270.400 ;
        RECT 649.200 269.700 658.000 270.300 ;
        RECT 649.200 269.600 650.000 269.700 ;
        RECT 657.200 269.600 658.000 269.700 ;
        RECT 660.400 270.300 661.200 270.400 ;
        RECT 666.800 270.300 667.600 270.400 ;
        RECT 660.400 269.700 667.600 270.300 ;
        RECT 660.400 269.600 661.200 269.700 ;
        RECT 666.800 269.600 667.600 269.700 ;
        RECT 6.000 268.300 6.800 268.400 ;
        RECT 14.000 268.300 14.800 268.400 ;
        RECT 6.000 267.700 14.800 268.300 ;
        RECT 6.000 267.600 6.800 267.700 ;
        RECT 14.000 267.600 14.800 267.700 ;
        RECT 55.600 268.300 56.400 268.400 ;
        RECT 57.200 268.300 58.000 268.400 ;
        RECT 60.400 268.300 61.200 268.400 ;
        RECT 111.600 268.300 112.400 268.400 ;
        RECT 55.600 267.700 112.400 268.300 ;
        RECT 55.600 267.600 56.400 267.700 ;
        RECT 57.200 267.600 58.000 267.700 ;
        RECT 60.400 267.600 61.200 267.700 ;
        RECT 111.600 267.600 112.400 267.700 ;
        RECT 156.400 268.300 157.200 268.400 ;
        RECT 170.800 268.300 171.600 268.400 ;
        RECT 156.400 267.700 171.600 268.300 ;
        RECT 156.400 267.600 157.200 267.700 ;
        RECT 170.800 267.600 171.600 267.700 ;
        RECT 268.400 268.300 269.200 268.400 ;
        RECT 273.200 268.300 274.000 268.400 ;
        RECT 268.400 267.700 274.000 268.300 ;
        RECT 268.400 267.600 269.200 267.700 ;
        RECT 273.200 267.600 274.000 267.700 ;
        RECT 286.000 267.600 286.800 268.400 ;
        RECT 326.000 268.300 326.800 268.400 ;
        RECT 335.600 268.300 336.400 268.400 ;
        RECT 326.000 267.700 336.400 268.300 ;
        RECT 326.000 267.600 326.800 267.700 ;
        RECT 335.600 267.600 336.400 267.700 ;
        RECT 439.600 268.300 440.400 268.400 ;
        RECT 463.600 268.300 464.400 268.400 ;
        RECT 439.600 267.700 464.400 268.300 ;
        RECT 439.600 267.600 440.400 267.700 ;
        RECT 463.600 267.600 464.400 267.700 ;
        RECT 489.200 268.300 490.000 268.400 ;
        RECT 506.800 268.300 507.600 268.400 ;
        RECT 489.200 267.700 507.600 268.300 ;
        RECT 489.200 267.600 490.000 267.700 ;
        RECT 506.800 267.600 507.600 267.700 ;
        RECT 529.200 268.300 530.000 268.400 ;
        RECT 534.000 268.300 534.800 268.400 ;
        RECT 529.200 267.700 534.800 268.300 ;
        RECT 529.200 267.600 530.000 267.700 ;
        RECT 534.000 267.600 534.800 267.700 ;
        RECT 562.800 268.300 563.600 268.400 ;
        RECT 585.200 268.300 586.000 268.400 ;
        RECT 562.800 267.700 586.000 268.300 ;
        RECT 562.800 267.600 563.600 267.700 ;
        RECT 585.200 267.600 586.000 267.700 ;
        RECT 599.600 268.300 600.400 268.400 ;
        RECT 604.400 268.300 605.200 268.400 ;
        RECT 618.800 268.300 619.600 268.400 ;
        RECT 634.800 268.300 635.600 268.400 ;
        RECT 652.400 268.300 653.200 268.400 ;
        RECT 663.600 268.300 664.400 268.400 ;
        RECT 665.200 268.300 666.000 268.400 ;
        RECT 599.600 267.700 666.000 268.300 ;
        RECT 599.600 267.600 600.400 267.700 ;
        RECT 604.400 267.600 605.200 267.700 ;
        RECT 618.800 267.600 619.600 267.700 ;
        RECT 634.800 267.600 635.600 267.700 ;
        RECT 652.400 267.600 653.200 267.700 ;
        RECT 663.600 267.600 664.400 267.700 ;
        RECT 665.200 267.600 666.000 267.700 ;
        RECT 17.200 266.300 18.000 266.400 ;
        RECT 36.400 266.300 37.200 266.400 ;
        RECT 17.200 265.700 37.200 266.300 ;
        RECT 17.200 265.600 18.000 265.700 ;
        RECT 36.400 265.600 37.200 265.700 ;
        RECT 50.800 266.300 51.600 266.400 ;
        RECT 108.400 266.300 109.200 266.400 ;
        RECT 50.800 265.700 109.200 266.300 ;
        RECT 50.800 265.600 51.600 265.700 ;
        RECT 108.400 265.600 109.200 265.700 ;
        RECT 153.200 266.300 154.000 266.400 ;
        RECT 186.800 266.300 187.600 266.400 ;
        RECT 206.000 266.300 206.800 266.400 ;
        RECT 153.200 265.700 206.800 266.300 ;
        RECT 153.200 265.600 154.000 265.700 ;
        RECT 186.800 265.600 187.600 265.700 ;
        RECT 206.000 265.600 206.800 265.700 ;
        RECT 249.200 266.300 250.000 266.400 ;
        RECT 270.000 266.300 270.800 266.400 ;
        RECT 249.200 265.700 270.800 266.300 ;
        RECT 249.200 265.600 250.000 265.700 ;
        RECT 270.000 265.600 270.800 265.700 ;
        RECT 306.800 266.300 307.600 266.400 ;
        RECT 343.600 266.300 344.400 266.400 ;
        RECT 306.800 265.700 344.400 266.300 ;
        RECT 306.800 265.600 307.600 265.700 ;
        RECT 343.600 265.600 344.400 265.700 ;
        RECT 348.400 266.300 349.200 266.400 ;
        RECT 353.200 266.300 354.000 266.400 ;
        RECT 354.800 266.300 355.600 266.400 ;
        RECT 348.400 265.700 355.600 266.300 ;
        RECT 348.400 265.600 349.200 265.700 ;
        RECT 353.200 265.600 354.000 265.700 ;
        RECT 354.800 265.600 355.600 265.700 ;
        RECT 356.400 266.300 357.200 266.400 ;
        RECT 370.800 266.300 371.600 266.400 ;
        RECT 356.400 265.700 371.600 266.300 ;
        RECT 356.400 265.600 357.200 265.700 ;
        RECT 370.800 265.600 371.600 265.700 ;
        RECT 375.600 266.300 376.400 266.400 ;
        RECT 410.800 266.300 411.600 266.400 ;
        RECT 375.600 265.700 411.600 266.300 ;
        RECT 375.600 265.600 376.400 265.700 ;
        RECT 410.800 265.600 411.600 265.700 ;
        RECT 425.200 266.300 426.000 266.400 ;
        RECT 455.600 266.300 456.400 266.400 ;
        RECT 425.200 265.700 456.400 266.300 ;
        RECT 425.200 265.600 426.000 265.700 ;
        RECT 455.600 265.600 456.400 265.700 ;
        RECT 478.000 266.300 478.800 266.400 ;
        RECT 489.200 266.300 490.000 266.400 ;
        RECT 478.000 265.700 490.000 266.300 ;
        RECT 478.000 265.600 478.800 265.700 ;
        RECT 489.200 265.600 490.000 265.700 ;
        RECT 500.400 266.300 501.200 266.400 ;
        RECT 519.600 266.300 520.400 266.400 ;
        RECT 542.000 266.300 542.800 266.400 ;
        RECT 559.600 266.300 560.400 266.400 ;
        RECT 569.200 266.300 570.000 266.400 ;
        RECT 500.400 265.700 570.000 266.300 ;
        RECT 585.300 266.300 585.900 267.600 ;
        RECT 612.400 266.300 613.200 266.400 ;
        RECT 585.300 265.700 613.200 266.300 ;
        RECT 500.400 265.600 501.200 265.700 ;
        RECT 519.600 265.600 520.400 265.700 ;
        RECT 542.000 265.600 542.800 265.700 ;
        RECT 559.600 265.600 560.400 265.700 ;
        RECT 569.200 265.600 570.000 265.700 ;
        RECT 612.400 265.600 613.200 265.700 ;
        RECT 622.000 266.300 622.800 266.400 ;
        RECT 630.000 266.300 630.800 266.400 ;
        RECT 622.000 265.700 630.800 266.300 ;
        RECT 622.000 265.600 622.800 265.700 ;
        RECT 630.000 265.600 630.800 265.700 ;
        RECT 31.600 264.300 32.400 264.400 ;
        RECT 66.800 264.300 67.600 264.400 ;
        RECT 84.400 264.300 85.200 264.400 ;
        RECT 118.000 264.300 118.800 264.400 ;
        RECT 129.200 264.300 130.000 264.400 ;
        RECT 31.600 263.700 130.000 264.300 ;
        RECT 31.600 263.600 32.400 263.700 ;
        RECT 66.800 263.600 67.600 263.700 ;
        RECT 84.400 263.600 85.200 263.700 ;
        RECT 118.000 263.600 118.800 263.700 ;
        RECT 129.200 263.600 130.000 263.700 ;
        RECT 287.600 264.300 288.400 264.400 ;
        RECT 394.800 264.300 395.600 264.400 ;
        RECT 287.600 263.700 395.600 264.300 ;
        RECT 287.600 263.600 288.400 263.700 ;
        RECT 394.800 263.600 395.600 263.700 ;
        RECT 550.000 264.300 550.800 264.400 ;
        RECT 570.800 264.300 571.600 264.400 ;
        RECT 578.800 264.300 579.600 264.400 ;
        RECT 601.200 264.300 602.000 264.400 ;
        RECT 550.000 263.700 602.000 264.300 ;
        RECT 550.000 263.600 550.800 263.700 ;
        RECT 570.800 263.600 571.600 263.700 ;
        RECT 578.800 263.600 579.600 263.700 ;
        RECT 601.200 263.600 602.000 263.700 ;
        RECT 626.800 264.300 627.600 264.400 ;
        RECT 642.800 264.300 643.600 264.400 ;
        RECT 626.800 263.700 643.600 264.300 ;
        RECT 626.800 263.600 627.600 263.700 ;
        RECT 642.800 263.600 643.600 263.700 ;
        RECT 20.400 262.300 21.200 262.400 ;
        RECT 26.800 262.300 27.600 262.400 ;
        RECT 20.400 261.700 27.600 262.300 ;
        RECT 20.400 261.600 21.200 261.700 ;
        RECT 26.800 261.600 27.600 261.700 ;
        RECT 106.800 262.300 107.600 262.400 ;
        RECT 220.400 262.300 221.200 262.400 ;
        RECT 225.200 262.300 226.000 262.400 ;
        RECT 106.800 261.700 226.000 262.300 ;
        RECT 106.800 261.600 107.600 261.700 ;
        RECT 220.400 261.600 221.200 261.700 ;
        RECT 225.200 261.600 226.000 261.700 ;
        RECT 230.000 262.300 230.800 262.400 ;
        RECT 258.800 262.300 259.600 262.400 ;
        RECT 230.000 261.700 259.600 262.300 ;
        RECT 230.000 261.600 230.800 261.700 ;
        RECT 258.800 261.600 259.600 261.700 ;
        RECT 284.400 262.300 285.200 262.400 ;
        RECT 313.200 262.300 314.000 262.400 ;
        RECT 350.000 262.300 350.800 262.400 ;
        RECT 367.600 262.300 368.400 262.400 ;
        RECT 406.000 262.300 406.800 262.400 ;
        RECT 284.400 261.700 406.800 262.300 ;
        RECT 284.400 261.600 285.200 261.700 ;
        RECT 313.200 261.600 314.000 261.700 ;
        RECT 350.000 261.600 350.800 261.700 ;
        RECT 367.600 261.600 368.400 261.700 ;
        RECT 406.000 261.600 406.800 261.700 ;
        RECT 521.200 262.300 522.000 262.400 ;
        RECT 548.400 262.300 549.200 262.400 ;
        RECT 521.200 261.700 549.200 262.300 ;
        RECT 521.200 261.600 522.000 261.700 ;
        RECT 548.400 261.600 549.200 261.700 ;
        RECT 12.400 260.300 13.200 260.400 ;
        RECT 54.000 260.300 54.800 260.400 ;
        RECT 12.400 259.700 54.800 260.300 ;
        RECT 12.400 259.600 13.200 259.700 ;
        RECT 54.000 259.600 54.800 259.700 ;
        RECT 65.200 260.300 66.000 260.400 ;
        RECT 70.000 260.300 70.800 260.400 ;
        RECT 65.200 259.700 70.800 260.300 ;
        RECT 65.200 259.600 66.000 259.700 ;
        RECT 70.000 259.600 70.800 259.700 ;
        RECT 89.200 260.300 90.000 260.400 ;
        RECT 98.800 260.300 99.600 260.400 ;
        RECT 89.200 259.700 99.600 260.300 ;
        RECT 89.200 259.600 90.000 259.700 ;
        RECT 98.800 259.600 99.600 259.700 ;
        RECT 103.600 260.300 104.400 260.400 ;
        RECT 122.800 260.300 123.600 260.400 ;
        RECT 103.600 259.700 123.600 260.300 ;
        RECT 103.600 259.600 104.400 259.700 ;
        RECT 122.800 259.600 123.600 259.700 ;
        RECT 124.400 260.300 125.200 260.400 ;
        RECT 130.800 260.300 131.600 260.400 ;
        RECT 142.000 260.300 142.800 260.400 ;
        RECT 183.600 260.300 184.400 260.400 ;
        RECT 124.400 259.700 184.400 260.300 ;
        RECT 124.400 259.600 125.200 259.700 ;
        RECT 130.800 259.600 131.600 259.700 ;
        RECT 142.000 259.600 142.800 259.700 ;
        RECT 183.600 259.600 184.400 259.700 ;
        RECT 241.200 260.300 242.000 260.400 ;
        RECT 246.000 260.300 246.800 260.400 ;
        RECT 241.200 259.700 246.800 260.300 ;
        RECT 241.200 259.600 242.000 259.700 ;
        RECT 246.000 259.600 246.800 259.700 ;
        RECT 295.600 259.600 296.400 260.400 ;
        RECT 297.200 260.300 298.000 260.400 ;
        RECT 302.000 260.300 302.800 260.400 ;
        RECT 297.200 259.700 302.800 260.300 ;
        RECT 297.200 259.600 298.000 259.700 ;
        RECT 302.000 259.600 302.800 259.700 ;
        RECT 364.400 260.300 365.200 260.400 ;
        RECT 369.200 260.300 370.000 260.400 ;
        RECT 402.800 260.300 403.600 260.400 ;
        RECT 364.400 259.700 403.600 260.300 ;
        RECT 364.400 259.600 365.200 259.700 ;
        RECT 369.200 259.600 370.000 259.700 ;
        RECT 402.800 259.600 403.600 259.700 ;
        RECT 442.800 260.300 443.600 260.400 ;
        RECT 450.800 260.300 451.600 260.400 ;
        RECT 481.200 260.300 482.000 260.400 ;
        RECT 527.600 260.300 528.400 260.400 ;
        RECT 442.800 259.700 528.400 260.300 ;
        RECT 442.800 259.600 443.600 259.700 ;
        RECT 450.800 259.600 451.600 259.700 ;
        RECT 481.200 259.600 482.000 259.700 ;
        RECT 527.600 259.600 528.400 259.700 ;
        RECT 534.000 260.300 534.800 260.400 ;
        RECT 566.000 260.300 566.800 260.400 ;
        RECT 534.000 259.700 566.800 260.300 ;
        RECT 534.000 259.600 534.800 259.700 ;
        RECT 566.000 259.600 566.800 259.700 ;
        RECT 580.400 260.300 581.200 260.400 ;
        RECT 596.400 260.300 597.200 260.400 ;
        RECT 580.400 259.700 597.200 260.300 ;
        RECT 580.400 259.600 581.200 259.700 ;
        RECT 596.400 259.600 597.200 259.700 ;
        RECT 641.200 260.300 642.000 260.400 ;
        RECT 666.800 260.300 667.600 260.400 ;
        RECT 641.200 259.700 667.600 260.300 ;
        RECT 641.200 259.600 642.000 259.700 ;
        RECT 666.800 259.600 667.600 259.700 ;
        RECT 97.200 258.300 98.000 258.400 ;
        RECT 186.800 258.300 187.600 258.400 ;
        RECT 97.200 257.700 187.600 258.300 ;
        RECT 97.200 257.600 98.000 257.700 ;
        RECT 186.800 257.600 187.600 257.700 ;
        RECT 209.200 258.300 210.000 258.400 ;
        RECT 217.200 258.300 218.000 258.400 ;
        RECT 223.600 258.300 224.400 258.400 ;
        RECT 209.200 257.700 224.400 258.300 ;
        RECT 209.200 257.600 210.000 257.700 ;
        RECT 217.200 257.600 218.000 257.700 ;
        RECT 223.600 257.600 224.400 257.700 ;
        RECT 228.400 258.300 229.200 258.400 ;
        RECT 274.800 258.300 275.600 258.400 ;
        RECT 321.200 258.300 322.000 258.400 ;
        RECT 228.400 257.700 322.000 258.300 ;
        RECT 228.400 257.600 229.200 257.700 ;
        RECT 274.800 257.600 275.600 257.700 ;
        RECT 321.200 257.600 322.000 257.700 ;
        RECT 327.600 258.300 328.400 258.400 ;
        RECT 340.400 258.300 341.200 258.400 ;
        RECT 327.600 257.700 341.200 258.300 ;
        RECT 327.600 257.600 328.400 257.700 ;
        RECT 340.400 257.600 341.200 257.700 ;
        RECT 350.000 258.300 350.800 258.400 ;
        RECT 369.200 258.300 370.000 258.400 ;
        RECT 350.000 257.700 370.000 258.300 ;
        RECT 350.000 257.600 350.800 257.700 ;
        RECT 369.200 257.600 370.000 257.700 ;
        RECT 410.800 258.300 411.600 258.400 ;
        RECT 446.000 258.300 446.800 258.400 ;
        RECT 410.800 257.700 446.800 258.300 ;
        RECT 410.800 257.600 411.600 257.700 ;
        RECT 446.000 257.600 446.800 257.700 ;
        RECT 455.600 257.600 456.400 258.400 ;
        RECT 462.000 258.300 462.800 258.400 ;
        RECT 470.000 258.300 470.800 258.400 ;
        RECT 462.000 257.700 470.800 258.300 ;
        RECT 462.000 257.600 462.800 257.700 ;
        RECT 470.000 257.600 470.800 257.700 ;
        RECT 551.600 258.300 552.400 258.400 ;
        RECT 553.200 258.300 554.000 258.400 ;
        RECT 551.600 257.700 554.000 258.300 ;
        RECT 551.600 257.600 552.400 257.700 ;
        RECT 553.200 257.600 554.000 257.700 ;
        RECT 588.400 258.300 589.200 258.400 ;
        RECT 602.800 258.300 603.600 258.400 ;
        RECT 588.400 257.700 603.600 258.300 ;
        RECT 588.400 257.600 589.200 257.700 ;
        RECT 602.800 257.600 603.600 257.700 ;
        RECT 612.400 258.300 613.200 258.400 ;
        RECT 622.000 258.300 622.800 258.400 ;
        RECT 612.400 257.700 622.800 258.300 ;
        RECT 612.400 257.600 613.200 257.700 ;
        RECT 622.000 257.600 622.800 257.700 ;
        RECT 642.800 258.300 643.600 258.400 ;
        RECT 660.400 258.300 661.200 258.400 ;
        RECT 687.600 258.300 688.400 258.400 ;
        RECT 642.800 257.700 688.400 258.300 ;
        RECT 642.800 257.600 643.600 257.700 ;
        RECT 660.400 257.600 661.200 257.700 ;
        RECT 687.600 257.600 688.400 257.700 ;
        RECT 10.800 256.300 11.600 256.400 ;
        RECT 14.000 256.300 14.800 256.400 ;
        RECT 10.800 255.700 14.800 256.300 ;
        RECT 10.800 255.600 11.600 255.700 ;
        RECT 14.000 255.600 14.800 255.700 ;
        RECT 105.200 256.300 106.000 256.400 ;
        RECT 106.800 256.300 107.600 256.400 ;
        RECT 105.200 255.700 107.600 256.300 ;
        RECT 105.200 255.600 106.000 255.700 ;
        RECT 106.800 255.600 107.600 255.700 ;
        RECT 119.600 256.300 120.400 256.400 ;
        RECT 156.400 256.300 157.200 256.400 ;
        RECT 158.000 256.300 158.800 256.400 ;
        RECT 119.600 255.700 158.800 256.300 ;
        RECT 119.600 255.600 120.400 255.700 ;
        RECT 156.400 255.600 157.200 255.700 ;
        RECT 158.000 255.600 158.800 255.700 ;
        RECT 241.200 256.300 242.000 256.400 ;
        RECT 290.800 256.300 291.600 256.400 ;
        RECT 241.200 255.700 291.600 256.300 ;
        RECT 241.200 255.600 242.000 255.700 ;
        RECT 290.800 255.600 291.600 255.700 ;
        RECT 294.000 256.300 294.800 256.400 ;
        RECT 329.200 256.300 330.000 256.400 ;
        RECT 294.000 255.700 330.000 256.300 ;
        RECT 294.000 255.600 294.800 255.700 ;
        RECT 329.200 255.600 330.000 255.700 ;
        RECT 346.800 256.300 347.600 256.400 ;
        RECT 372.400 256.300 373.200 256.400 ;
        RECT 346.800 255.700 373.200 256.300 ;
        RECT 346.800 255.600 347.600 255.700 ;
        RECT 372.400 255.600 373.200 255.700 ;
        RECT 380.400 256.300 381.200 256.400 ;
        RECT 386.800 256.300 387.600 256.400 ;
        RECT 380.400 255.700 387.600 256.300 ;
        RECT 380.400 255.600 381.200 255.700 ;
        RECT 386.800 255.600 387.600 255.700 ;
        RECT 401.200 256.300 402.000 256.400 ;
        RECT 410.800 256.300 411.600 256.400 ;
        RECT 401.200 255.700 411.600 256.300 ;
        RECT 401.200 255.600 402.000 255.700 ;
        RECT 410.800 255.600 411.600 255.700 ;
        RECT 436.400 256.300 437.200 256.400 ;
        RECT 439.600 256.300 440.400 256.400 ;
        RECT 471.600 256.300 472.400 256.400 ;
        RECT 436.400 255.700 472.400 256.300 ;
        RECT 436.400 255.600 437.200 255.700 ;
        RECT 439.600 255.600 440.400 255.700 ;
        RECT 471.600 255.600 472.400 255.700 ;
        RECT 505.200 256.300 506.000 256.400 ;
        RECT 510.000 256.300 510.800 256.400 ;
        RECT 543.600 256.300 544.400 256.400 ;
        RECT 505.200 255.700 544.400 256.300 ;
        RECT 505.200 255.600 506.000 255.700 ;
        RECT 510.000 255.600 510.800 255.700 ;
        RECT 543.600 255.600 544.400 255.700 ;
        RECT 569.200 256.300 570.000 256.400 ;
        RECT 588.400 256.300 589.200 256.400 ;
        RECT 569.200 255.700 589.200 256.300 ;
        RECT 569.200 255.600 570.000 255.700 ;
        RECT 588.400 255.600 589.200 255.700 ;
        RECT 634.800 256.300 635.600 256.400 ;
        RECT 655.600 256.300 656.400 256.400 ;
        RECT 634.800 255.700 656.400 256.300 ;
        RECT 634.800 255.600 635.600 255.700 ;
        RECT 655.600 255.600 656.400 255.700 ;
        RECT 658.800 256.300 659.600 256.400 ;
        RECT 662.000 256.300 662.800 256.400 ;
        RECT 658.800 255.700 662.800 256.300 ;
        RECT 658.800 255.600 659.600 255.700 ;
        RECT 662.000 255.600 662.800 255.700 ;
        RECT 34.800 254.300 35.600 254.400 ;
        RECT 50.800 254.300 51.600 254.400 ;
        RECT 34.800 253.700 51.600 254.300 ;
        RECT 34.800 253.600 35.600 253.700 ;
        RECT 50.800 253.600 51.600 253.700 ;
        RECT 82.800 254.300 83.600 254.400 ;
        RECT 108.400 254.300 109.200 254.400 ;
        RECT 82.800 253.700 109.200 254.300 ;
        RECT 82.800 253.600 83.600 253.700 ;
        RECT 108.400 253.600 109.200 253.700 ;
        RECT 140.400 254.300 141.200 254.400 ;
        RECT 169.200 254.300 170.000 254.400 ;
        RECT 140.400 253.700 170.000 254.300 ;
        RECT 140.400 253.600 141.200 253.700 ;
        RECT 169.200 253.600 170.000 253.700 ;
        RECT 183.600 254.300 184.400 254.400 ;
        RECT 198.000 254.300 198.800 254.400 ;
        RECT 183.600 253.700 198.800 254.300 ;
        RECT 183.600 253.600 184.400 253.700 ;
        RECT 198.000 253.600 198.800 253.700 ;
        RECT 226.800 254.300 227.600 254.400 ;
        RECT 244.400 254.300 245.200 254.400 ;
        RECT 226.800 253.700 245.200 254.300 ;
        RECT 226.800 253.600 227.600 253.700 ;
        RECT 244.400 253.600 245.200 253.700 ;
        RECT 326.000 254.300 326.800 254.400 ;
        RECT 330.800 254.300 331.600 254.400 ;
        RECT 326.000 253.700 331.600 254.300 ;
        RECT 326.000 253.600 326.800 253.700 ;
        RECT 330.800 253.600 331.600 253.700 ;
        RECT 334.000 254.300 334.800 254.400 ;
        RECT 337.200 254.300 338.000 254.400 ;
        RECT 334.000 253.700 338.000 254.300 ;
        RECT 334.000 253.600 334.800 253.700 ;
        RECT 337.200 253.600 338.000 253.700 ;
        RECT 338.800 254.300 339.600 254.400 ;
        RECT 380.400 254.300 381.200 254.400 ;
        RECT 338.800 253.700 381.200 254.300 ;
        RECT 338.800 253.600 339.600 253.700 ;
        RECT 380.400 253.600 381.200 253.700 ;
        RECT 398.000 254.300 398.800 254.400 ;
        RECT 404.400 254.300 405.200 254.400 ;
        RECT 398.000 253.700 405.200 254.300 ;
        RECT 398.000 253.600 398.800 253.700 ;
        RECT 404.400 253.600 405.200 253.700 ;
        RECT 414.000 254.300 414.800 254.400 ;
        RECT 436.400 254.300 437.200 254.400 ;
        RECT 414.000 253.700 437.200 254.300 ;
        RECT 414.000 253.600 414.800 253.700 ;
        RECT 436.400 253.600 437.200 253.700 ;
        RECT 481.200 254.300 482.000 254.400 ;
        RECT 484.400 254.300 485.200 254.400 ;
        RECT 481.200 253.700 485.200 254.300 ;
        RECT 481.200 253.600 482.000 253.700 ;
        RECT 484.400 253.600 485.200 253.700 ;
        RECT 506.800 254.300 507.600 254.400 ;
        RECT 524.400 254.300 525.200 254.400 ;
        RECT 506.800 253.700 525.200 254.300 ;
        RECT 506.800 253.600 507.600 253.700 ;
        RECT 524.400 253.600 525.200 253.700 ;
        RECT 554.800 254.300 555.600 254.400 ;
        RECT 582.000 254.300 582.800 254.400 ;
        RECT 593.200 254.300 594.000 254.400 ;
        RECT 554.800 253.700 594.000 254.300 ;
        RECT 554.800 253.600 555.600 253.700 ;
        RECT 582.000 253.600 582.800 253.700 ;
        RECT 593.200 253.600 594.000 253.700 ;
        RECT 618.800 254.300 619.600 254.400 ;
        RECT 628.400 254.300 629.200 254.400 ;
        RECT 618.800 253.700 629.200 254.300 ;
        RECT 618.800 253.600 619.600 253.700 ;
        RECT 628.400 253.600 629.200 253.700 ;
        RECT 630.000 254.300 630.800 254.400 ;
        RECT 641.200 254.300 642.000 254.400 ;
        RECT 630.000 253.700 642.000 254.300 ;
        RECT 630.000 253.600 630.800 253.700 ;
        RECT 641.200 253.600 642.000 253.700 ;
        RECT 654.000 254.300 654.800 254.400 ;
        RECT 658.800 254.300 659.600 254.400 ;
        RECT 654.000 253.700 659.600 254.300 ;
        RECT 654.000 253.600 654.800 253.700 ;
        RECT 658.800 253.600 659.600 253.700 ;
        RECT 44.400 252.300 45.200 252.400 ;
        RECT 58.800 252.300 59.600 252.400 ;
        RECT 44.400 251.700 59.600 252.300 ;
        RECT 44.400 251.600 45.200 251.700 ;
        RECT 58.800 251.600 59.600 251.700 ;
        RECT 78.000 252.300 78.800 252.400 ;
        RECT 167.600 252.300 168.400 252.400 ;
        RECT 180.400 252.300 181.200 252.400 ;
        RECT 78.000 251.700 181.200 252.300 ;
        RECT 78.000 251.600 78.800 251.700 ;
        RECT 167.600 251.600 168.400 251.700 ;
        RECT 180.400 251.600 181.200 251.700 ;
        RECT 209.200 252.300 210.000 252.400 ;
        RECT 218.800 252.300 219.600 252.400 ;
        RECT 209.200 251.700 219.600 252.300 ;
        RECT 209.200 251.600 210.000 251.700 ;
        RECT 218.800 251.600 219.600 251.700 ;
        RECT 233.200 252.300 234.000 252.400 ;
        RECT 310.000 252.300 310.800 252.400 ;
        RECT 233.200 251.700 310.800 252.300 ;
        RECT 233.200 251.600 234.000 251.700 ;
        RECT 310.000 251.600 310.800 251.700 ;
        RECT 314.800 252.300 315.600 252.400 ;
        RECT 316.400 252.300 317.200 252.400 ;
        RECT 314.800 251.700 317.200 252.300 ;
        RECT 314.800 251.600 315.600 251.700 ;
        RECT 316.400 251.600 317.200 251.700 ;
        RECT 326.000 252.300 326.800 252.400 ;
        RECT 329.200 252.300 330.000 252.400 ;
        RECT 326.000 251.700 330.000 252.300 ;
        RECT 326.000 251.600 326.800 251.700 ;
        RECT 329.200 251.600 330.000 251.700 ;
        RECT 367.600 252.300 368.400 252.400 ;
        RECT 385.200 252.300 386.000 252.400 ;
        RECT 367.600 251.700 386.000 252.300 ;
        RECT 367.600 251.600 368.400 251.700 ;
        RECT 385.200 251.600 386.000 251.700 ;
        RECT 391.600 252.300 392.400 252.400 ;
        RECT 414.000 252.300 414.800 252.400 ;
        RECT 391.600 251.700 414.800 252.300 ;
        RECT 391.600 251.600 392.400 251.700 ;
        RECT 414.000 251.600 414.800 251.700 ;
        RECT 457.200 252.300 458.000 252.400 ;
        RECT 486.000 252.300 486.800 252.400 ;
        RECT 498.800 252.300 499.600 252.400 ;
        RECT 457.200 251.700 499.600 252.300 ;
        RECT 457.200 251.600 458.000 251.700 ;
        RECT 486.000 251.600 486.800 251.700 ;
        RECT 498.800 251.600 499.600 251.700 ;
        RECT 548.400 252.300 549.200 252.400 ;
        RECT 558.000 252.300 558.800 252.400 ;
        RECT 548.400 251.700 558.800 252.300 ;
        RECT 548.400 251.600 549.200 251.700 ;
        RECT 558.000 251.600 558.800 251.700 ;
        RECT 575.600 252.300 576.400 252.400 ;
        RECT 588.400 252.300 589.200 252.400 ;
        RECT 575.600 251.700 589.200 252.300 ;
        RECT 575.600 251.600 576.400 251.700 ;
        RECT 588.400 251.600 589.200 251.700 ;
        RECT 594.800 252.300 595.600 252.400 ;
        RECT 612.400 252.300 613.200 252.400 ;
        RECT 594.800 251.700 613.200 252.300 ;
        RECT 594.800 251.600 595.600 251.700 ;
        RECT 612.400 251.600 613.200 251.700 ;
        RECT 614.000 252.300 614.800 252.400 ;
        RECT 633.200 252.300 634.000 252.400 ;
        RECT 614.000 251.700 634.000 252.300 ;
        RECT 614.000 251.600 614.800 251.700 ;
        RECT 633.200 251.600 634.000 251.700 ;
        RECT 641.200 252.300 642.000 252.400 ;
        RECT 644.400 252.300 645.200 252.400 ;
        RECT 641.200 251.700 645.200 252.300 ;
        RECT 641.200 251.600 642.000 251.700 ;
        RECT 644.400 251.600 645.200 251.700 ;
        RECT 657.200 252.300 658.000 252.400 ;
        RECT 665.200 252.300 666.000 252.400 ;
        RECT 657.200 251.700 666.000 252.300 ;
        RECT 657.200 251.600 658.000 251.700 ;
        RECT 665.200 251.600 666.000 251.700 ;
        RECT 668.400 252.300 669.200 252.400 ;
        RECT 674.800 252.300 675.600 252.400 ;
        RECT 668.400 251.700 675.600 252.300 ;
        RECT 668.400 251.600 669.200 251.700 ;
        RECT 674.800 251.600 675.600 251.700 ;
        RECT 4.400 250.300 5.200 250.400 ;
        RECT 50.800 250.300 51.600 250.400 ;
        RECT 57.200 250.300 58.000 250.400 ;
        RECT 4.400 249.700 58.000 250.300 ;
        RECT 4.400 249.600 5.200 249.700 ;
        RECT 50.800 249.600 51.600 249.700 ;
        RECT 57.200 249.600 58.000 249.700 ;
        RECT 156.400 250.300 157.200 250.400 ;
        RECT 201.200 250.300 202.000 250.400 ;
        RECT 156.400 249.700 202.000 250.300 ;
        RECT 156.400 249.600 157.200 249.700 ;
        RECT 201.200 249.600 202.000 249.700 ;
        RECT 289.200 250.300 290.000 250.400 ;
        RECT 290.800 250.300 291.600 250.400 ;
        RECT 383.600 250.300 384.400 250.400 ;
        RECT 388.400 250.300 389.200 250.400 ;
        RECT 391.600 250.300 392.400 250.400 ;
        RECT 289.200 249.700 291.600 250.300 ;
        RECT 289.200 249.600 290.000 249.700 ;
        RECT 290.800 249.600 291.600 249.700 ;
        RECT 310.100 249.700 382.700 250.300 ;
        RECT 310.100 248.300 310.700 249.700 ;
        RECT 290.900 247.700 310.700 248.300 ;
        RECT 311.600 248.300 312.400 248.400 ;
        RECT 318.000 248.300 318.800 248.400 ;
        RECT 321.200 248.300 322.000 248.400 ;
        RECT 311.600 247.700 322.000 248.300 ;
        RECT 290.900 246.400 291.500 247.700 ;
        RECT 311.600 247.600 312.400 247.700 ;
        RECT 318.000 247.600 318.800 247.700 ;
        RECT 321.200 247.600 322.000 247.700 ;
        RECT 324.400 248.300 325.200 248.400 ;
        RECT 327.600 248.300 328.400 248.400 ;
        RECT 324.400 247.700 328.400 248.300 ;
        RECT 324.400 247.600 325.200 247.700 ;
        RECT 327.600 247.600 328.400 247.700 ;
        RECT 337.200 248.300 338.000 248.400 ;
        RECT 342.000 248.300 342.800 248.400 ;
        RECT 337.200 247.700 342.800 248.300 ;
        RECT 337.200 247.600 338.000 247.700 ;
        RECT 342.000 247.600 342.800 247.700 ;
        RECT 351.600 248.300 352.400 248.400 ;
        RECT 354.800 248.300 355.600 248.400 ;
        RECT 351.600 247.700 355.600 248.300 ;
        RECT 382.100 248.300 382.700 249.700 ;
        RECT 383.600 249.700 392.400 250.300 ;
        RECT 383.600 249.600 384.400 249.700 ;
        RECT 388.400 249.600 389.200 249.700 ;
        RECT 391.600 249.600 392.400 249.700 ;
        RECT 415.600 250.300 416.400 250.400 ;
        RECT 426.800 250.300 427.600 250.400 ;
        RECT 415.600 249.700 427.600 250.300 ;
        RECT 415.600 249.600 416.400 249.700 ;
        RECT 426.800 249.600 427.600 249.700 ;
        RECT 428.400 250.300 429.200 250.400 ;
        RECT 460.400 250.300 461.200 250.400 ;
        RECT 428.400 249.700 461.200 250.300 ;
        RECT 428.400 249.600 429.200 249.700 ;
        RECT 460.400 249.600 461.200 249.700 ;
        RECT 478.000 250.300 478.800 250.400 ;
        RECT 514.800 250.300 515.600 250.400 ;
        RECT 478.000 249.700 515.600 250.300 ;
        RECT 478.000 249.600 478.800 249.700 ;
        RECT 514.800 249.600 515.600 249.700 ;
        RECT 631.600 250.300 632.400 250.400 ;
        RECT 652.400 250.300 653.200 250.400 ;
        RECT 631.600 249.700 653.200 250.300 ;
        RECT 631.600 249.600 632.400 249.700 ;
        RECT 652.400 249.600 653.200 249.700 ;
        RECT 657.200 250.300 658.000 250.400 ;
        RECT 663.600 250.300 664.400 250.400 ;
        RECT 657.200 249.700 664.400 250.300 ;
        RECT 657.200 249.600 658.000 249.700 ;
        RECT 663.600 249.600 664.400 249.700 ;
        RECT 666.800 250.300 667.600 250.400 ;
        RECT 668.400 250.300 669.200 250.400 ;
        RECT 666.800 249.700 669.200 250.300 ;
        RECT 666.800 249.600 667.600 249.700 ;
        RECT 668.400 249.600 669.200 249.700 ;
        RECT 490.800 248.300 491.600 248.400 ;
        RECT 500.400 248.300 501.200 248.400 ;
        RECT 382.100 247.700 501.200 248.300 ;
        RECT 351.600 247.600 352.400 247.700 ;
        RECT 354.800 247.600 355.600 247.700 ;
        RECT 490.800 247.600 491.600 247.700 ;
        RECT 500.400 247.600 501.200 247.700 ;
        RECT 644.400 248.300 645.200 248.400 ;
        RECT 647.600 248.300 648.400 248.400 ;
        RECT 644.400 247.700 648.400 248.300 ;
        RECT 644.400 247.600 645.200 247.700 ;
        RECT 647.600 247.600 648.400 247.700 ;
        RECT 76.400 246.300 77.200 246.400 ;
        RECT 290.800 246.300 291.600 246.400 ;
        RECT 76.400 245.700 291.600 246.300 ;
        RECT 76.400 245.600 77.200 245.700 ;
        RECT 290.800 245.600 291.600 245.700 ;
        RECT 292.400 246.300 293.200 246.400 ;
        RECT 327.600 246.300 328.400 246.400 ;
        RECT 335.600 246.300 336.400 246.400 ;
        RECT 377.200 246.300 378.000 246.400 ;
        RECT 378.800 246.300 379.600 246.400 ;
        RECT 385.200 246.300 386.000 246.400 ;
        RECT 292.400 245.700 386.000 246.300 ;
        RECT 292.400 245.600 293.200 245.700 ;
        RECT 327.600 245.600 328.400 245.700 ;
        RECT 335.600 245.600 336.400 245.700 ;
        RECT 377.200 245.600 378.000 245.700 ;
        RECT 378.800 245.600 379.600 245.700 ;
        RECT 385.200 245.600 386.000 245.700 ;
        RECT 390.000 246.300 390.800 246.400 ;
        RECT 423.600 246.300 424.400 246.400 ;
        RECT 390.000 245.700 424.400 246.300 ;
        RECT 390.000 245.600 390.800 245.700 ;
        RECT 423.600 245.600 424.400 245.700 ;
        RECT 260.400 244.300 261.200 244.400 ;
        RECT 268.400 244.300 269.200 244.400 ;
        RECT 337.200 244.300 338.000 244.400 ;
        RECT 366.000 244.300 366.800 244.400 ;
        RECT 388.400 244.300 389.200 244.400 ;
        RECT 458.800 244.300 459.600 244.400 ;
        RECT 260.400 243.700 459.600 244.300 ;
        RECT 260.400 243.600 261.200 243.700 ;
        RECT 268.400 243.600 269.200 243.700 ;
        RECT 337.200 243.600 338.000 243.700 ;
        RECT 366.000 243.600 366.800 243.700 ;
        RECT 388.400 243.600 389.200 243.700 ;
        RECT 458.800 243.600 459.600 243.700 ;
        RECT 673.200 244.300 674.000 244.400 ;
        RECT 679.600 244.300 680.400 244.400 ;
        RECT 673.200 243.700 680.400 244.300 ;
        RECT 673.200 243.600 674.000 243.700 ;
        RECT 679.600 243.600 680.400 243.700 ;
        RECT 137.200 242.300 138.000 242.400 ;
        RECT 167.600 242.300 168.400 242.400 ;
        RECT 137.200 241.700 168.400 242.300 ;
        RECT 137.200 241.600 138.000 241.700 ;
        RECT 167.600 241.600 168.400 241.700 ;
        RECT 284.400 242.300 285.200 242.400 ;
        RECT 286.000 242.300 286.800 242.400 ;
        RECT 284.400 241.700 286.800 242.300 ;
        RECT 284.400 241.600 285.200 241.700 ;
        RECT 286.000 241.600 286.800 241.700 ;
        RECT 295.600 241.600 296.400 242.400 ;
        RECT 318.000 242.300 318.800 242.400 ;
        RECT 322.800 242.300 323.600 242.400 ;
        RECT 318.000 241.700 323.600 242.300 ;
        RECT 318.000 241.600 318.800 241.700 ;
        RECT 322.800 241.600 323.600 241.700 ;
        RECT 340.400 242.300 341.200 242.400 ;
        RECT 361.200 242.300 362.000 242.400 ;
        RECT 340.400 241.700 362.000 242.300 ;
        RECT 340.400 241.600 341.200 241.700 ;
        RECT 361.200 241.600 362.000 241.700 ;
        RECT 383.600 242.300 384.400 242.400 ;
        RECT 393.200 242.300 394.000 242.400 ;
        RECT 383.600 241.700 394.000 242.300 ;
        RECT 383.600 241.600 384.400 241.700 ;
        RECT 393.200 241.600 394.000 241.700 ;
        RECT 153.200 240.300 154.000 240.400 ;
        RECT 156.400 240.300 157.200 240.400 ;
        RECT 153.200 239.700 157.200 240.300 ;
        RECT 153.200 239.600 154.000 239.700 ;
        RECT 156.400 239.600 157.200 239.700 ;
        RECT 180.400 240.300 181.200 240.400 ;
        RECT 185.200 240.300 186.000 240.400 ;
        RECT 230.000 240.300 230.800 240.400 ;
        RECT 271.600 240.300 272.400 240.400 ;
        RECT 337.200 240.300 338.000 240.400 ;
        RECT 180.400 239.700 338.000 240.300 ;
        RECT 180.400 239.600 181.200 239.700 ;
        RECT 185.200 239.600 186.000 239.700 ;
        RECT 230.000 239.600 230.800 239.700 ;
        RECT 271.600 239.600 272.400 239.700 ;
        RECT 337.200 239.600 338.000 239.700 ;
        RECT 354.800 240.300 355.600 240.400 ;
        RECT 650.800 240.300 651.600 240.400 ;
        RECT 654.000 240.300 654.800 240.400 ;
        RECT 354.800 239.700 413.100 240.300 ;
        RECT 354.800 239.600 355.600 239.700 ;
        RECT 122.800 238.300 123.600 238.400 ;
        RECT 140.400 238.300 141.200 238.400 ;
        RECT 122.800 237.700 141.200 238.300 ;
        RECT 122.800 237.600 123.600 237.700 ;
        RECT 140.400 237.600 141.200 237.700 ;
        RECT 167.600 238.300 168.400 238.400 ;
        RECT 354.800 238.300 355.600 238.400 ;
        RECT 167.600 237.700 355.600 238.300 ;
        RECT 167.600 237.600 168.400 237.700 ;
        RECT 354.800 237.600 355.600 237.700 ;
        RECT 378.800 238.300 379.600 238.400 ;
        RECT 385.200 238.300 386.000 238.400 ;
        RECT 401.200 238.300 402.000 238.400 ;
        RECT 378.800 237.700 402.000 238.300 ;
        RECT 412.500 238.300 413.100 239.700 ;
        RECT 650.800 239.700 654.800 240.300 ;
        RECT 650.800 239.600 651.600 239.700 ;
        RECT 654.000 239.600 654.800 239.700 ;
        RECT 428.400 238.300 429.200 238.400 ;
        RECT 412.500 237.700 429.200 238.300 ;
        RECT 378.800 237.600 379.600 237.700 ;
        RECT 385.200 237.600 386.000 237.700 ;
        RECT 401.200 237.600 402.000 237.700 ;
        RECT 428.400 237.600 429.200 237.700 ;
        RECT 610.800 238.300 611.600 238.400 ;
        RECT 630.000 238.300 630.800 238.400 ;
        RECT 610.800 237.700 630.800 238.300 ;
        RECT 610.800 237.600 611.600 237.700 ;
        RECT 630.000 237.600 630.800 237.700 ;
        RECT 217.200 236.300 218.000 236.400 ;
        RECT 239.600 236.300 240.400 236.400 ;
        RECT 217.200 235.700 240.400 236.300 ;
        RECT 217.200 235.600 218.000 235.700 ;
        RECT 239.600 235.600 240.400 235.700 ;
        RECT 330.800 236.300 331.600 236.400 ;
        RECT 369.200 236.300 370.000 236.400 ;
        RECT 330.800 235.700 370.000 236.300 ;
        RECT 330.800 235.600 331.600 235.700 ;
        RECT 369.200 235.600 370.000 235.700 ;
        RECT 375.600 236.300 376.400 236.400 ;
        RECT 380.400 236.300 381.200 236.400 ;
        RECT 375.600 235.700 381.200 236.300 ;
        RECT 375.600 235.600 376.400 235.700 ;
        RECT 380.400 235.600 381.200 235.700 ;
        RECT 660.400 236.300 661.200 236.400 ;
        RECT 682.800 236.300 683.600 236.400 ;
        RECT 660.400 235.700 683.600 236.300 ;
        RECT 660.400 235.600 661.200 235.700 ;
        RECT 682.800 235.600 683.600 235.700 ;
        RECT 167.600 234.300 168.400 234.400 ;
        RECT 242.800 234.300 243.600 234.400 ;
        RECT 167.600 233.700 243.600 234.300 ;
        RECT 167.600 233.600 168.400 233.700 ;
        RECT 242.800 233.600 243.600 233.700 ;
        RECT 327.600 234.300 328.400 234.400 ;
        RECT 361.200 234.300 362.000 234.400 ;
        RECT 327.600 233.700 362.000 234.300 ;
        RECT 327.600 233.600 328.400 233.700 ;
        RECT 361.200 233.600 362.000 233.700 ;
        RECT 375.600 234.300 376.400 234.400 ;
        RECT 382.000 234.300 382.800 234.400 ;
        RECT 375.600 233.700 382.800 234.300 ;
        RECT 375.600 233.600 376.400 233.700 ;
        RECT 382.000 233.600 382.800 233.700 ;
        RECT 423.600 234.300 424.400 234.400 ;
        RECT 482.800 234.300 483.600 234.400 ;
        RECT 489.200 234.300 490.000 234.400 ;
        RECT 423.600 233.700 490.000 234.300 ;
        RECT 423.600 233.600 424.400 233.700 ;
        RECT 482.800 233.600 483.600 233.700 ;
        RECT 489.200 233.600 490.000 233.700 ;
        RECT 65.200 232.300 66.000 232.400 ;
        RECT 78.000 232.300 78.800 232.400 ;
        RECT 65.200 231.700 78.800 232.300 ;
        RECT 65.200 231.600 66.000 231.700 ;
        RECT 78.000 231.600 78.800 231.700 ;
        RECT 100.400 232.300 101.200 232.400 ;
        RECT 159.600 232.300 160.400 232.400 ;
        RECT 100.400 231.700 160.400 232.300 ;
        RECT 100.400 231.600 101.200 231.700 ;
        RECT 159.600 231.600 160.400 231.700 ;
        RECT 236.400 232.300 237.200 232.400 ;
        RECT 238.000 232.300 238.800 232.400 ;
        RECT 294.000 232.300 294.800 232.400 ;
        RECT 236.400 231.700 294.800 232.300 ;
        RECT 236.400 231.600 237.200 231.700 ;
        RECT 238.000 231.600 238.800 231.700 ;
        RECT 294.000 231.600 294.800 231.700 ;
        RECT 330.800 232.300 331.600 232.400 ;
        RECT 362.800 232.300 363.600 232.400 ;
        RECT 330.800 231.700 363.600 232.300 ;
        RECT 330.800 231.600 331.600 231.700 ;
        RECT 362.800 231.600 363.600 231.700 ;
        RECT 393.200 232.300 394.000 232.400 ;
        RECT 402.800 232.300 403.600 232.400 ;
        RECT 393.200 231.700 403.600 232.300 ;
        RECT 393.200 231.600 394.000 231.700 ;
        RECT 402.800 231.600 403.600 231.700 ;
        RECT 410.800 232.300 411.600 232.400 ;
        RECT 426.800 232.300 427.600 232.400 ;
        RECT 457.200 232.300 458.000 232.400 ;
        RECT 410.800 231.700 458.000 232.300 ;
        RECT 410.800 231.600 411.600 231.700 ;
        RECT 426.800 231.600 427.600 231.700 ;
        RECT 457.200 231.600 458.000 231.700 ;
        RECT 538.800 232.300 539.600 232.400 ;
        RECT 556.400 232.300 557.200 232.400 ;
        RECT 538.800 231.700 557.200 232.300 ;
        RECT 538.800 231.600 539.600 231.700 ;
        RECT 556.400 231.600 557.200 231.700 ;
        RECT 558.000 232.300 558.800 232.400 ;
        RECT 566.000 232.300 566.800 232.400 ;
        RECT 572.400 232.300 573.200 232.400 ;
        RECT 558.000 231.700 573.200 232.300 ;
        RECT 558.000 231.600 558.800 231.700 ;
        RECT 566.000 231.600 566.800 231.700 ;
        RECT 572.400 231.600 573.200 231.700 ;
        RECT 623.600 232.300 624.400 232.400 ;
        RECT 646.000 232.300 646.800 232.400 ;
        RECT 623.600 231.700 646.800 232.300 ;
        RECT 623.600 231.600 624.400 231.700 ;
        RECT 646.000 231.600 646.800 231.700 ;
        RECT 18.800 230.300 19.600 230.400 ;
        RECT 58.800 230.300 59.600 230.400 ;
        RECT 18.800 229.700 59.600 230.300 ;
        RECT 18.800 229.600 19.600 229.700 ;
        RECT 58.800 229.600 59.600 229.700 ;
        RECT 76.400 230.300 77.200 230.400 ;
        RECT 79.600 230.300 80.400 230.400 ;
        RECT 76.400 229.700 80.400 230.300 ;
        RECT 76.400 229.600 77.200 229.700 ;
        RECT 79.600 229.600 80.400 229.700 ;
        RECT 111.600 230.300 112.400 230.400 ;
        RECT 118.000 230.300 118.800 230.400 ;
        RECT 148.400 230.300 149.200 230.400 ;
        RECT 111.600 229.700 149.200 230.300 ;
        RECT 111.600 229.600 112.400 229.700 ;
        RECT 118.000 229.600 118.800 229.700 ;
        RECT 148.400 229.600 149.200 229.700 ;
        RECT 207.600 230.300 208.400 230.400 ;
        RECT 233.200 230.300 234.000 230.400 ;
        RECT 207.600 229.700 234.000 230.300 ;
        RECT 207.600 229.600 208.400 229.700 ;
        RECT 233.200 229.600 234.000 229.700 ;
        RECT 270.000 230.300 270.800 230.400 ;
        RECT 287.600 230.300 288.400 230.400 ;
        RECT 290.800 230.300 291.600 230.400 ;
        RECT 270.000 229.700 291.600 230.300 ;
        RECT 270.000 229.600 270.800 229.700 ;
        RECT 287.600 229.600 288.400 229.700 ;
        RECT 290.800 229.600 291.600 229.700 ;
        RECT 300.400 230.300 301.200 230.400 ;
        RECT 306.800 230.300 307.600 230.400 ;
        RECT 313.200 230.300 314.000 230.400 ;
        RECT 300.400 229.700 314.000 230.300 ;
        RECT 300.400 229.600 301.200 229.700 ;
        RECT 306.800 229.600 307.600 229.700 ;
        RECT 313.200 229.600 314.000 229.700 ;
        RECT 316.400 230.300 317.200 230.400 ;
        RECT 364.400 230.300 365.200 230.400 ;
        RECT 316.400 229.700 365.200 230.300 ;
        RECT 316.400 229.600 317.200 229.700 ;
        RECT 364.400 229.600 365.200 229.700 ;
        RECT 372.400 230.300 373.200 230.400 ;
        RECT 385.200 230.300 386.000 230.400 ;
        RECT 390.000 230.300 390.800 230.400 ;
        RECT 372.400 229.700 390.800 230.300 ;
        RECT 372.400 229.600 373.200 229.700 ;
        RECT 385.200 229.600 386.000 229.700 ;
        RECT 390.000 229.600 390.800 229.700 ;
        RECT 550.000 230.300 550.800 230.400 ;
        RECT 585.200 230.300 586.000 230.400 ;
        RECT 550.000 229.700 586.000 230.300 ;
        RECT 550.000 229.600 550.800 229.700 ;
        RECT 585.200 229.600 586.000 229.700 ;
        RECT 607.600 230.300 608.400 230.400 ;
        RECT 620.400 230.300 621.200 230.400 ;
        RECT 633.200 230.300 634.000 230.400 ;
        RECT 607.600 229.700 634.000 230.300 ;
        RECT 607.600 229.600 608.400 229.700 ;
        RECT 620.400 229.600 621.200 229.700 ;
        RECT 633.200 229.600 634.000 229.700 ;
        RECT 674.800 230.300 675.600 230.400 ;
        RECT 686.000 230.300 686.800 230.400 ;
        RECT 674.800 229.700 686.800 230.300 ;
        RECT 674.800 229.600 675.600 229.700 ;
        RECT 686.000 229.600 686.800 229.700 ;
        RECT 42.800 228.300 43.600 228.400 ;
        RECT 57.200 228.300 58.000 228.400 ;
        RECT 42.800 227.700 58.000 228.300 ;
        RECT 42.800 227.600 43.600 227.700 ;
        RECT 57.200 227.600 58.000 227.700 ;
        RECT 70.000 228.300 70.800 228.400 ;
        RECT 74.800 228.300 75.600 228.400 ;
        RECT 127.600 228.300 128.400 228.400 ;
        RECT 135.600 228.300 136.400 228.400 ;
        RECT 70.000 227.700 136.400 228.300 ;
        RECT 70.000 227.600 70.800 227.700 ;
        RECT 74.800 227.600 75.600 227.700 ;
        RECT 127.600 227.600 128.400 227.700 ;
        RECT 135.600 227.600 136.400 227.700 ;
        RECT 159.600 228.300 160.400 228.400 ;
        RECT 175.600 228.300 176.400 228.400 ;
        RECT 159.600 227.700 176.400 228.300 ;
        RECT 159.600 227.600 160.400 227.700 ;
        RECT 175.600 227.600 176.400 227.700 ;
        RECT 228.400 228.300 229.200 228.400 ;
        RECT 233.200 228.300 234.000 228.400 ;
        RECT 319.600 228.300 320.400 228.400 ;
        RECT 228.400 227.700 320.400 228.300 ;
        RECT 228.400 227.600 229.200 227.700 ;
        RECT 233.200 227.600 234.000 227.700 ;
        RECT 319.600 227.600 320.400 227.700 ;
        RECT 350.000 228.300 350.800 228.400 ;
        RECT 356.400 228.300 357.200 228.400 ;
        RECT 350.000 227.700 357.200 228.300 ;
        RECT 350.000 227.600 350.800 227.700 ;
        RECT 356.400 227.600 357.200 227.700 ;
        RECT 366.000 228.300 366.800 228.400 ;
        RECT 370.800 228.300 371.600 228.400 ;
        RECT 366.000 227.700 371.600 228.300 ;
        RECT 366.000 227.600 366.800 227.700 ;
        RECT 370.800 227.600 371.600 227.700 ;
        RECT 383.600 228.300 384.400 228.400 ;
        RECT 385.200 228.300 386.000 228.400 ;
        RECT 383.600 227.700 386.000 228.300 ;
        RECT 383.600 227.600 384.400 227.700 ;
        RECT 385.200 227.600 386.000 227.700 ;
        RECT 399.600 228.300 400.400 228.400 ;
        RECT 431.600 228.300 432.400 228.400 ;
        RECT 399.600 227.700 432.400 228.300 ;
        RECT 399.600 227.600 400.400 227.700 ;
        RECT 431.600 227.600 432.400 227.700 ;
        RECT 466.800 228.300 467.600 228.400 ;
        RECT 492.400 228.300 493.200 228.400 ;
        RECT 466.800 227.700 493.200 228.300 ;
        RECT 466.800 227.600 467.600 227.700 ;
        RECT 492.400 227.600 493.200 227.700 ;
        RECT 514.800 228.300 515.600 228.400 ;
        RECT 529.200 228.300 530.000 228.400 ;
        RECT 514.800 227.700 530.000 228.300 ;
        RECT 514.800 227.600 515.600 227.700 ;
        RECT 529.200 227.600 530.000 227.700 ;
        RECT 540.400 228.300 541.200 228.400 ;
        RECT 556.400 228.300 557.200 228.400 ;
        RECT 540.400 227.700 557.200 228.300 ;
        RECT 540.400 227.600 541.200 227.700 ;
        RECT 556.400 227.600 557.200 227.700 ;
        RECT 559.600 228.300 560.400 228.400 ;
        RECT 567.600 228.300 568.400 228.400 ;
        RECT 559.600 227.700 568.400 228.300 ;
        RECT 559.600 227.600 560.400 227.700 ;
        RECT 567.600 227.600 568.400 227.700 ;
        RECT 18.800 226.300 19.600 226.400 ;
        RECT 23.600 226.300 24.400 226.400 ;
        RECT 18.800 225.700 24.400 226.300 ;
        RECT 18.800 225.600 19.600 225.700 ;
        RECT 23.600 225.600 24.400 225.700 ;
        RECT 62.000 226.300 62.800 226.400 ;
        RECT 66.800 226.300 67.600 226.400 ;
        RECT 62.000 225.700 67.600 226.300 ;
        RECT 62.000 225.600 62.800 225.700 ;
        RECT 66.800 225.600 67.600 225.700 ;
        RECT 119.600 226.300 120.400 226.400 ;
        RECT 130.800 226.300 131.600 226.400 ;
        RECT 119.600 225.700 131.600 226.300 ;
        RECT 119.600 225.600 120.400 225.700 ;
        RECT 130.800 225.600 131.600 225.700 ;
        RECT 134.000 226.300 134.800 226.400 ;
        RECT 158.000 226.300 158.800 226.400 ;
        RECT 174.000 226.300 174.800 226.400 ;
        RECT 134.000 225.700 174.800 226.300 ;
        RECT 134.000 225.600 134.800 225.700 ;
        RECT 158.000 225.600 158.800 225.700 ;
        RECT 174.000 225.600 174.800 225.700 ;
        RECT 204.400 226.300 205.200 226.400 ;
        RECT 241.200 226.300 242.000 226.400 ;
        RECT 204.400 225.700 242.000 226.300 ;
        RECT 204.400 225.600 205.200 225.700 ;
        RECT 241.200 225.600 242.000 225.700 ;
        RECT 286.000 225.600 286.800 226.400 ;
        RECT 294.000 226.300 294.800 226.400 ;
        RECT 313.200 226.300 314.000 226.400 ;
        RECT 324.400 226.300 325.200 226.400 ;
        RECT 294.000 225.700 325.200 226.300 ;
        RECT 294.000 225.600 294.800 225.700 ;
        RECT 313.200 225.600 314.000 225.700 ;
        RECT 324.400 225.600 325.200 225.700 ;
        RECT 402.800 226.300 403.600 226.400 ;
        RECT 423.600 226.300 424.400 226.400 ;
        RECT 402.800 225.700 424.400 226.300 ;
        RECT 402.800 225.600 403.600 225.700 ;
        RECT 423.600 225.600 424.400 225.700 ;
        RECT 425.200 226.300 426.000 226.400 ;
        RECT 436.400 226.300 437.200 226.400 ;
        RECT 425.200 225.700 437.200 226.300 ;
        RECT 425.200 225.600 426.000 225.700 ;
        RECT 436.400 225.600 437.200 225.700 ;
        RECT 486.000 226.300 486.800 226.400 ;
        RECT 500.400 226.300 501.200 226.400 ;
        RECT 486.000 225.700 501.200 226.300 ;
        RECT 486.000 225.600 486.800 225.700 ;
        RECT 500.400 225.600 501.200 225.700 ;
        RECT 534.000 226.300 534.800 226.400 ;
        RECT 542.000 226.300 542.800 226.400 ;
        RECT 546.800 226.300 547.600 226.400 ;
        RECT 554.800 226.300 555.600 226.400 ;
        RECT 561.200 226.300 562.000 226.400 ;
        RECT 534.000 225.700 562.000 226.300 ;
        RECT 534.000 225.600 534.800 225.700 ;
        RECT 542.000 225.600 542.800 225.700 ;
        RECT 546.800 225.600 547.600 225.700 ;
        RECT 554.800 225.600 555.600 225.700 ;
        RECT 561.200 225.600 562.000 225.700 ;
        RECT 52.400 224.300 53.200 224.400 ;
        RECT 70.000 224.300 70.800 224.400 ;
        RECT 52.400 223.700 70.800 224.300 ;
        RECT 52.400 223.600 53.200 223.700 ;
        RECT 70.000 223.600 70.800 223.700 ;
        RECT 103.600 224.300 104.400 224.400 ;
        RECT 156.400 224.300 157.200 224.400 ;
        RECT 103.600 223.700 157.200 224.300 ;
        RECT 103.600 223.600 104.400 223.700 ;
        RECT 156.400 223.600 157.200 223.700 ;
        RECT 174.000 224.300 174.800 224.400 ;
        RECT 180.400 224.300 181.200 224.400 ;
        RECT 174.000 223.700 181.200 224.300 ;
        RECT 174.000 223.600 174.800 223.700 ;
        RECT 180.400 223.600 181.200 223.700 ;
        RECT 234.800 224.300 235.600 224.400 ;
        RECT 242.800 224.300 243.600 224.400 ;
        RECT 273.200 224.300 274.000 224.400 ;
        RECT 234.800 223.700 274.000 224.300 ;
        RECT 234.800 223.600 235.600 223.700 ;
        RECT 242.800 223.600 243.600 223.700 ;
        RECT 273.200 223.600 274.000 223.700 ;
        RECT 302.000 224.300 302.800 224.400 ;
        RECT 308.400 224.300 309.200 224.400 ;
        RECT 302.000 223.700 309.200 224.300 ;
        RECT 302.000 223.600 302.800 223.700 ;
        RECT 308.400 223.600 309.200 223.700 ;
        RECT 343.600 224.300 344.400 224.400 ;
        RECT 348.400 224.300 349.200 224.400 ;
        RECT 343.600 223.700 349.200 224.300 ;
        RECT 343.600 223.600 344.400 223.700 ;
        RECT 348.400 223.600 349.200 223.700 ;
        RECT 375.600 224.300 376.400 224.400 ;
        RECT 380.400 224.300 381.200 224.400 ;
        RECT 375.600 223.700 381.200 224.300 ;
        RECT 375.600 223.600 376.400 223.700 ;
        RECT 380.400 223.600 381.200 223.700 ;
        RECT 593.200 224.300 594.000 224.400 ;
        RECT 626.800 224.300 627.600 224.400 ;
        RECT 628.400 224.300 629.200 224.400 ;
        RECT 646.000 224.300 646.800 224.400 ;
        RECT 668.400 224.300 669.200 224.400 ;
        RECT 593.200 223.700 669.200 224.300 ;
        RECT 593.200 223.600 594.000 223.700 ;
        RECT 626.800 223.600 627.600 223.700 ;
        RECT 628.400 223.600 629.200 223.700 ;
        RECT 646.000 223.600 646.800 223.700 ;
        RECT 668.400 223.600 669.200 223.700 ;
        RECT 135.600 222.300 136.400 222.400 ;
        RECT 138.800 222.300 139.600 222.400 ;
        RECT 135.600 221.700 139.600 222.300 ;
        RECT 135.600 221.600 136.400 221.700 ;
        RECT 138.800 221.600 139.600 221.700 ;
        RECT 158.000 222.300 158.800 222.400 ;
        RECT 188.400 222.300 189.200 222.400 ;
        RECT 234.800 222.300 235.600 222.400 ;
        RECT 158.000 221.700 235.600 222.300 ;
        RECT 158.000 221.600 158.800 221.700 ;
        RECT 188.400 221.600 189.200 221.700 ;
        RECT 234.800 221.600 235.600 221.700 ;
        RECT 273.200 222.300 274.000 222.400 ;
        RECT 321.200 222.300 322.000 222.400 ;
        RECT 367.600 222.300 368.400 222.400 ;
        RECT 273.200 221.700 368.400 222.300 ;
        RECT 273.200 221.600 274.000 221.700 ;
        RECT 321.200 221.600 322.000 221.700 ;
        RECT 367.600 221.600 368.400 221.700 ;
        RECT 372.400 222.300 373.200 222.400 ;
        RECT 394.800 222.300 395.600 222.400 ;
        RECT 372.400 221.700 395.600 222.300 ;
        RECT 372.400 221.600 373.200 221.700 ;
        RECT 394.800 221.600 395.600 221.700 ;
        RECT 506.800 222.300 507.600 222.400 ;
        RECT 511.600 222.300 512.400 222.400 ;
        RECT 506.800 221.700 512.400 222.300 ;
        RECT 506.800 221.600 507.600 221.700 ;
        RECT 511.600 221.600 512.400 221.700 ;
        RECT 586.800 222.300 587.600 222.400 ;
        RECT 596.400 222.300 597.200 222.400 ;
        RECT 586.800 221.700 597.200 222.300 ;
        RECT 586.800 221.600 587.600 221.700 ;
        RECT 596.400 221.600 597.200 221.700 ;
        RECT 642.800 222.300 643.600 222.400 ;
        RECT 649.200 222.300 650.000 222.400 ;
        RECT 642.800 221.700 650.000 222.300 ;
        RECT 642.800 221.600 643.600 221.700 ;
        RECT 649.200 221.600 650.000 221.700 ;
        RECT 73.200 220.300 74.000 220.400 ;
        RECT 81.200 220.300 82.000 220.400 ;
        RECT 73.200 219.700 82.000 220.300 ;
        RECT 73.200 219.600 74.000 219.700 ;
        RECT 81.200 219.600 82.000 219.700 ;
        RECT 134.000 220.300 134.800 220.400 ;
        RECT 138.800 220.300 139.600 220.400 ;
        RECT 134.000 219.700 139.600 220.300 ;
        RECT 134.000 219.600 134.800 219.700 ;
        RECT 138.800 219.600 139.600 219.700 ;
        RECT 236.400 220.300 237.200 220.400 ;
        RECT 239.600 220.300 240.400 220.400 ;
        RECT 236.400 219.700 240.400 220.300 ;
        RECT 236.400 219.600 237.200 219.700 ;
        RECT 239.600 219.600 240.400 219.700 ;
        RECT 318.000 220.300 318.800 220.400 ;
        RECT 375.600 220.300 376.400 220.400 ;
        RECT 318.000 219.700 376.400 220.300 ;
        RECT 318.000 219.600 318.800 219.700 ;
        RECT 375.600 219.600 376.400 219.700 ;
        RECT 377.200 220.300 378.000 220.400 ;
        RECT 401.200 220.300 402.000 220.400 ;
        RECT 377.200 219.700 402.000 220.300 ;
        RECT 377.200 219.600 378.000 219.700 ;
        RECT 401.200 219.600 402.000 219.700 ;
        RECT 404.400 220.300 405.200 220.400 ;
        RECT 410.800 220.300 411.600 220.400 ;
        RECT 404.400 219.700 411.600 220.300 ;
        RECT 404.400 219.600 405.200 219.700 ;
        RECT 410.800 219.600 411.600 219.700 ;
        RECT 2.800 218.300 3.600 218.400 ;
        RECT 26.800 218.300 27.600 218.400 ;
        RECT 39.600 218.300 40.400 218.400 ;
        RECT 78.000 218.300 78.800 218.400 ;
        RECT 87.600 218.300 88.400 218.400 ;
        RECT 2.800 217.700 88.400 218.300 ;
        RECT 2.800 217.600 3.600 217.700 ;
        RECT 26.800 217.600 27.600 217.700 ;
        RECT 39.600 217.600 40.400 217.700 ;
        RECT 78.000 217.600 78.800 217.700 ;
        RECT 87.600 217.600 88.400 217.700 ;
        RECT 154.800 218.300 155.600 218.400 ;
        RECT 158.000 218.300 158.800 218.400 ;
        RECT 154.800 217.700 158.800 218.300 ;
        RECT 154.800 217.600 155.600 217.700 ;
        RECT 158.000 217.600 158.800 217.700 ;
        RECT 231.600 218.300 232.400 218.400 ;
        RECT 236.400 218.300 237.200 218.400 ;
        RECT 231.600 217.700 237.200 218.300 ;
        RECT 231.600 217.600 232.400 217.700 ;
        RECT 236.400 217.600 237.200 217.700 ;
        RECT 250.800 218.300 251.600 218.400 ;
        RECT 302.000 218.300 302.800 218.400 ;
        RECT 250.800 217.700 302.800 218.300 ;
        RECT 250.800 217.600 251.600 217.700 ;
        RECT 302.000 217.600 302.800 217.700 ;
        RECT 310.000 218.300 310.800 218.400 ;
        RECT 330.800 218.300 331.600 218.400 ;
        RECT 310.000 217.700 331.600 218.300 ;
        RECT 375.700 218.300 376.300 219.600 ;
        RECT 390.000 218.300 390.800 218.400 ;
        RECT 375.700 217.700 390.800 218.300 ;
        RECT 310.000 217.600 310.800 217.700 ;
        RECT 330.800 217.600 331.600 217.700 ;
        RECT 390.000 217.600 390.800 217.700 ;
        RECT 470.000 218.300 470.800 218.400 ;
        RECT 503.600 218.300 504.400 218.400 ;
        RECT 518.000 218.300 518.800 218.400 ;
        RECT 470.000 217.700 518.800 218.300 ;
        RECT 470.000 217.600 470.800 217.700 ;
        RECT 503.600 217.600 504.400 217.700 ;
        RECT 518.000 217.600 518.800 217.700 ;
        RECT 527.600 218.300 528.400 218.400 ;
        RECT 580.400 218.300 581.200 218.400 ;
        RECT 527.600 217.700 581.200 218.300 ;
        RECT 527.600 217.600 528.400 217.700 ;
        RECT 580.400 217.600 581.200 217.700 ;
        RECT 14.000 216.300 14.800 216.400 ;
        RECT 49.200 216.300 50.000 216.400 ;
        RECT 58.800 216.300 59.600 216.400 ;
        RECT 106.800 216.300 107.600 216.400 ;
        RECT 108.400 216.300 109.200 216.400 ;
        RECT 135.600 216.300 136.400 216.400 ;
        RECT 150.000 216.300 150.800 216.400 ;
        RECT 14.000 215.700 96.300 216.300 ;
        RECT 14.000 215.600 14.800 215.700 ;
        RECT 49.200 215.600 50.000 215.700 ;
        RECT 58.800 215.600 59.600 215.700 ;
        RECT 95.700 214.400 96.300 215.700 ;
        RECT 106.800 215.700 150.800 216.300 ;
        RECT 106.800 215.600 107.600 215.700 ;
        RECT 108.400 215.600 109.200 215.700 ;
        RECT 135.600 215.600 136.400 215.700 ;
        RECT 150.000 215.600 150.800 215.700 ;
        RECT 156.400 216.300 157.200 216.400 ;
        RECT 170.800 216.300 171.600 216.400 ;
        RECT 156.400 215.700 171.600 216.300 ;
        RECT 156.400 215.600 157.200 215.700 ;
        RECT 170.800 215.600 171.600 215.700 ;
        RECT 183.600 216.300 184.400 216.400 ;
        RECT 215.600 216.300 216.400 216.400 ;
        RECT 183.600 215.700 216.400 216.300 ;
        RECT 183.600 215.600 184.400 215.700 ;
        RECT 215.600 215.600 216.400 215.700 ;
        RECT 258.800 216.300 259.600 216.400 ;
        RECT 260.400 216.300 261.200 216.400 ;
        RECT 258.800 215.700 261.200 216.300 ;
        RECT 258.800 215.600 259.600 215.700 ;
        RECT 260.400 215.600 261.200 215.700 ;
        RECT 281.200 216.300 282.000 216.400 ;
        RECT 289.200 216.300 290.000 216.400 ;
        RECT 281.200 215.700 290.000 216.300 ;
        RECT 281.200 215.600 282.000 215.700 ;
        RECT 289.200 215.600 290.000 215.700 ;
        RECT 294.000 216.300 294.800 216.400 ;
        RECT 298.800 216.300 299.600 216.400 ;
        RECT 294.000 215.700 299.600 216.300 ;
        RECT 294.000 215.600 294.800 215.700 ;
        RECT 298.800 215.600 299.600 215.700 ;
        RECT 305.200 216.300 306.000 216.400 ;
        RECT 334.000 216.300 334.800 216.400 ;
        RECT 305.200 215.700 334.800 216.300 ;
        RECT 305.200 215.600 306.000 215.700 ;
        RECT 334.000 215.600 334.800 215.700 ;
        RECT 337.200 216.300 338.000 216.400 ;
        RECT 342.000 216.300 342.800 216.400 ;
        RECT 337.200 215.700 342.800 216.300 ;
        RECT 337.200 215.600 338.000 215.700 ;
        RECT 342.000 215.600 342.800 215.700 ;
        RECT 423.600 216.300 424.400 216.400 ;
        RECT 450.800 216.300 451.600 216.400 ;
        RECT 466.800 216.300 467.600 216.400 ;
        RECT 423.600 215.700 467.600 216.300 ;
        RECT 423.600 215.600 424.400 215.700 ;
        RECT 450.800 215.600 451.600 215.700 ;
        RECT 466.800 215.600 467.600 215.700 ;
        RECT 470.000 216.300 470.800 216.400 ;
        RECT 537.200 216.300 538.000 216.400 ;
        RECT 470.000 215.700 538.000 216.300 ;
        RECT 470.000 215.600 470.800 215.700 ;
        RECT 537.200 215.600 538.000 215.700 ;
        RECT 548.400 216.300 549.200 216.400 ;
        RECT 564.400 216.300 565.200 216.400 ;
        RECT 548.400 215.700 565.200 216.300 ;
        RECT 548.400 215.600 549.200 215.700 ;
        RECT 564.400 215.600 565.200 215.700 ;
        RECT 655.600 216.300 656.400 216.400 ;
        RECT 662.000 216.300 662.800 216.400 ;
        RECT 655.600 215.700 662.800 216.300 ;
        RECT 655.600 215.600 656.400 215.700 ;
        RECT 662.000 215.600 662.800 215.700 ;
        RECT 9.200 214.300 10.000 214.400 ;
        RECT 23.600 214.300 24.400 214.400 ;
        RECT 9.200 213.700 24.400 214.300 ;
        RECT 9.200 213.600 10.000 213.700 ;
        RECT 23.600 213.600 24.400 213.700 ;
        RECT 95.600 214.300 96.400 214.400 ;
        RECT 124.400 214.300 125.200 214.400 ;
        RECT 95.600 213.700 125.200 214.300 ;
        RECT 95.600 213.600 96.400 213.700 ;
        RECT 124.400 213.600 125.200 213.700 ;
        RECT 183.600 214.300 184.400 214.400 ;
        RECT 190.000 214.300 190.800 214.400 ;
        RECT 183.600 213.700 190.800 214.300 ;
        RECT 183.600 213.600 184.400 213.700 ;
        RECT 190.000 213.600 190.800 213.700 ;
        RECT 201.200 214.300 202.000 214.400 ;
        RECT 226.800 214.300 227.600 214.400 ;
        RECT 201.200 213.700 227.600 214.300 ;
        RECT 201.200 213.600 202.000 213.700 ;
        RECT 226.800 213.600 227.600 213.700 ;
        RECT 231.600 214.300 232.400 214.400 ;
        RECT 238.000 214.300 238.800 214.400 ;
        RECT 231.600 213.700 238.800 214.300 ;
        RECT 231.600 213.600 232.400 213.700 ;
        RECT 238.000 213.600 238.800 213.700 ;
        RECT 295.600 214.300 296.400 214.400 ;
        RECT 303.600 214.300 304.400 214.400 ;
        RECT 295.600 213.700 304.400 214.300 ;
        RECT 295.600 213.600 296.400 213.700 ;
        RECT 303.600 213.600 304.400 213.700 ;
        RECT 321.200 214.300 322.000 214.400 ;
        RECT 345.200 214.300 346.000 214.400 ;
        RECT 321.200 213.700 346.000 214.300 ;
        RECT 321.200 213.600 322.000 213.700 ;
        RECT 345.200 213.600 346.000 213.700 ;
        RECT 359.600 214.300 360.400 214.400 ;
        RECT 375.600 214.300 376.400 214.400 ;
        RECT 359.600 213.700 376.400 214.300 ;
        RECT 359.600 213.600 360.400 213.700 ;
        RECT 375.600 213.600 376.400 213.700 ;
        RECT 388.400 214.300 389.200 214.400 ;
        RECT 391.600 214.300 392.400 214.400 ;
        RECT 396.400 214.300 397.200 214.400 ;
        RECT 388.400 213.700 397.200 214.300 ;
        RECT 388.400 213.600 389.200 213.700 ;
        RECT 391.600 213.600 392.400 213.700 ;
        RECT 396.400 213.600 397.200 213.700 ;
        RECT 420.400 214.300 421.200 214.400 ;
        RECT 476.400 214.300 477.200 214.400 ;
        RECT 420.400 213.700 477.200 214.300 ;
        RECT 420.400 213.600 421.200 213.700 ;
        RECT 476.400 213.600 477.200 213.700 ;
        RECT 500.400 214.300 501.200 214.400 ;
        RECT 543.600 214.300 544.400 214.400 ;
        RECT 500.400 213.700 544.400 214.300 ;
        RECT 500.400 213.600 501.200 213.700 ;
        RECT 543.600 213.600 544.400 213.700 ;
        RECT 545.200 214.300 546.000 214.400 ;
        RECT 548.400 214.300 549.200 214.400 ;
        RECT 545.200 213.700 549.200 214.300 ;
        RECT 545.200 213.600 546.000 213.700 ;
        RECT 548.400 213.600 549.200 213.700 ;
        RECT 551.600 214.300 552.400 214.400 ;
        RECT 554.800 214.300 555.600 214.400 ;
        RECT 551.600 213.700 555.600 214.300 ;
        RECT 551.600 213.600 552.400 213.700 ;
        RECT 554.800 213.600 555.600 213.700 ;
        RECT 566.000 214.300 566.800 214.400 ;
        RECT 577.200 214.300 578.000 214.400 ;
        RECT 590.000 214.300 590.800 214.400 ;
        RECT 566.000 213.700 590.800 214.300 ;
        RECT 566.000 213.600 566.800 213.700 ;
        RECT 577.200 213.600 578.000 213.700 ;
        RECT 590.000 213.600 590.800 213.700 ;
        RECT 599.600 214.300 600.400 214.400 ;
        RECT 607.600 214.300 608.400 214.400 ;
        RECT 599.600 213.700 608.400 214.300 ;
        RECT 599.600 213.600 600.400 213.700 ;
        RECT 607.600 213.600 608.400 213.700 ;
        RECT 610.800 214.300 611.600 214.400 ;
        RECT 631.600 214.300 632.400 214.400 ;
        RECT 610.800 213.700 632.400 214.300 ;
        RECT 610.800 213.600 611.600 213.700 ;
        RECT 631.600 213.600 632.400 213.700 ;
        RECT 646.000 214.300 646.800 214.400 ;
        RECT 665.200 214.300 666.000 214.400 ;
        RECT 646.000 213.700 666.000 214.300 ;
        RECT 646.000 213.600 646.800 213.700 ;
        RECT 665.200 213.600 666.000 213.700 ;
        RECT 138.800 212.300 139.600 212.400 ;
        RECT 226.800 212.300 227.600 212.400 ;
        RECT 231.700 212.300 232.300 213.600 ;
        RECT 138.800 211.700 232.300 212.300 ;
        RECT 249.200 212.300 250.000 212.400 ;
        RECT 255.600 212.300 256.400 212.400 ;
        RECT 273.200 212.300 274.000 212.400 ;
        RECT 249.200 211.700 274.000 212.300 ;
        RECT 138.800 211.600 139.600 211.700 ;
        RECT 226.800 211.600 227.600 211.700 ;
        RECT 249.200 211.600 250.000 211.700 ;
        RECT 255.600 211.600 256.400 211.700 ;
        RECT 273.200 211.600 274.000 211.700 ;
        RECT 298.800 212.300 299.600 212.400 ;
        RECT 310.000 212.300 310.800 212.400 ;
        RECT 327.600 212.300 328.400 212.400 ;
        RECT 298.800 211.700 328.400 212.300 ;
        RECT 298.800 211.600 299.600 211.700 ;
        RECT 310.000 211.600 310.800 211.700 ;
        RECT 327.600 211.600 328.400 211.700 ;
        RECT 332.400 212.300 333.200 212.400 ;
        RECT 337.200 212.300 338.000 212.400 ;
        RECT 332.400 211.700 338.000 212.300 ;
        RECT 332.400 211.600 333.200 211.700 ;
        RECT 337.200 211.600 338.000 211.700 ;
        RECT 342.000 212.300 342.800 212.400 ;
        RECT 391.600 212.300 392.400 212.400 ;
        RECT 342.000 211.700 392.400 212.300 ;
        RECT 342.000 211.600 342.800 211.700 ;
        RECT 391.600 211.600 392.400 211.700 ;
        RECT 396.400 212.300 397.200 212.400 ;
        RECT 433.200 212.300 434.000 212.400 ;
        RECT 442.800 212.300 443.600 212.400 ;
        RECT 450.800 212.300 451.600 212.400 ;
        RECT 396.400 211.700 451.600 212.300 ;
        RECT 396.400 211.600 397.200 211.700 ;
        RECT 433.200 211.600 434.000 211.700 ;
        RECT 442.800 211.600 443.600 211.700 ;
        RECT 450.800 211.600 451.600 211.700 ;
        RECT 545.200 212.300 546.000 212.400 ;
        RECT 569.200 212.300 570.000 212.400 ;
        RECT 545.200 211.700 570.000 212.300 ;
        RECT 545.200 211.600 546.000 211.700 ;
        RECT 569.200 211.600 570.000 211.700 ;
        RECT 578.800 212.300 579.600 212.400 ;
        RECT 598.000 212.300 598.800 212.400 ;
        RECT 599.600 212.300 600.400 212.400 ;
        RECT 612.400 212.300 613.200 212.400 ;
        RECT 578.800 211.700 613.200 212.300 ;
        RECT 578.800 211.600 579.600 211.700 ;
        RECT 598.000 211.600 598.800 211.700 ;
        RECT 599.600 211.600 600.400 211.700 ;
        RECT 612.400 211.600 613.200 211.700 ;
        RECT 655.600 212.300 656.400 212.400 ;
        RECT 658.800 212.300 659.600 212.400 ;
        RECT 671.600 212.300 672.400 212.400 ;
        RECT 655.600 211.700 672.400 212.300 ;
        RECT 655.600 211.600 656.400 211.700 ;
        RECT 658.800 211.600 659.600 211.700 ;
        RECT 671.600 211.600 672.400 211.700 ;
        RECT 238.000 210.300 238.800 210.400 ;
        RECT 257.200 210.300 258.000 210.400 ;
        RECT 278.000 210.300 278.800 210.400 ;
        RECT 238.000 209.700 278.800 210.300 ;
        RECT 238.000 209.600 238.800 209.700 ;
        RECT 257.200 209.600 258.000 209.700 ;
        RECT 278.000 209.600 278.800 209.700 ;
        RECT 303.600 210.300 304.400 210.400 ;
        RECT 306.800 210.300 307.600 210.400 ;
        RECT 303.600 209.700 307.600 210.300 ;
        RECT 303.600 209.600 304.400 209.700 ;
        RECT 306.800 209.600 307.600 209.700 ;
        RECT 313.200 210.300 314.000 210.400 ;
        RECT 346.800 210.300 347.600 210.400 ;
        RECT 350.000 210.300 350.800 210.400 ;
        RECT 313.200 209.700 350.800 210.300 ;
        RECT 313.200 209.600 314.000 209.700 ;
        RECT 346.800 209.600 347.600 209.700 ;
        RECT 350.000 209.600 350.800 209.700 ;
        RECT 479.600 210.300 480.400 210.400 ;
        RECT 489.200 210.300 490.000 210.400 ;
        RECT 479.600 209.700 490.000 210.300 ;
        RECT 479.600 209.600 480.400 209.700 ;
        RECT 489.200 209.600 490.000 209.700 ;
        RECT 527.600 210.300 528.400 210.400 ;
        RECT 556.400 210.300 557.200 210.400 ;
        RECT 527.600 209.700 557.200 210.300 ;
        RECT 527.600 209.600 528.400 209.700 ;
        RECT 556.400 209.600 557.200 209.700 ;
        RECT 567.600 210.300 568.400 210.400 ;
        RECT 578.800 210.300 579.600 210.400 ;
        RECT 567.600 209.700 579.600 210.300 ;
        RECT 567.600 209.600 568.400 209.700 ;
        RECT 578.800 209.600 579.600 209.700 ;
        RECT 593.200 210.300 594.000 210.400 ;
        RECT 602.800 210.300 603.600 210.400 ;
        RECT 593.200 209.700 603.600 210.300 ;
        RECT 593.200 209.600 594.000 209.700 ;
        RECT 602.800 209.600 603.600 209.700 ;
        RECT 254.000 208.300 254.800 208.400 ;
        RECT 335.600 208.300 336.400 208.400 ;
        RECT 254.000 207.700 336.400 208.300 ;
        RECT 254.000 207.600 254.800 207.700 ;
        RECT 335.600 207.600 336.400 207.700 ;
        RECT 401.200 208.300 402.000 208.400 ;
        RECT 426.800 208.300 427.600 208.400 ;
        RECT 401.200 207.700 427.600 208.300 ;
        RECT 401.200 207.600 402.000 207.700 ;
        RECT 426.800 207.600 427.600 207.700 ;
        RECT 436.400 208.300 437.200 208.400 ;
        RECT 439.600 208.300 440.400 208.400 ;
        RECT 436.400 207.700 440.400 208.300 ;
        RECT 436.400 207.600 437.200 207.700 ;
        RECT 439.600 207.600 440.400 207.700 ;
        RECT 529.200 208.300 530.000 208.400 ;
        RECT 551.600 208.300 552.400 208.400 ;
        RECT 529.200 207.700 552.400 208.300 ;
        RECT 529.200 207.600 530.000 207.700 ;
        RECT 551.600 207.600 552.400 207.700 ;
        RECT 554.800 208.300 555.600 208.400 ;
        RECT 601.200 208.300 602.000 208.400 ;
        RECT 554.800 207.700 602.000 208.300 ;
        RECT 554.800 207.600 555.600 207.700 ;
        RECT 601.200 207.600 602.000 207.700 ;
        RECT 300.400 206.300 301.200 206.400 ;
        RECT 303.600 206.300 304.400 206.400 ;
        RECT 300.400 205.700 304.400 206.300 ;
        RECT 300.400 205.600 301.200 205.700 ;
        RECT 303.600 205.600 304.400 205.700 ;
        RECT 334.000 206.300 334.800 206.400 ;
        RECT 396.400 206.300 397.200 206.400 ;
        RECT 334.000 205.700 397.200 206.300 ;
        RECT 334.000 205.600 334.800 205.700 ;
        RECT 396.400 205.600 397.200 205.700 ;
        RECT 526.000 206.300 526.800 206.400 ;
        RECT 534.000 206.300 534.800 206.400 ;
        RECT 526.000 205.700 534.800 206.300 ;
        RECT 526.000 205.600 526.800 205.700 ;
        RECT 534.000 205.600 534.800 205.700 ;
        RECT 679.600 206.300 680.400 206.400 ;
        RECT 686.000 206.300 686.800 206.400 ;
        RECT 679.600 205.700 686.800 206.300 ;
        RECT 679.600 205.600 680.400 205.700 ;
        RECT 686.000 205.600 686.800 205.700 ;
        RECT 10.800 204.300 11.600 204.400 ;
        RECT 42.800 204.300 43.600 204.400 ;
        RECT 68.400 204.300 69.200 204.400 ;
        RECT 10.800 203.700 69.200 204.300 ;
        RECT 10.800 203.600 11.600 203.700 ;
        RECT 42.800 203.600 43.600 203.700 ;
        RECT 68.400 203.600 69.200 203.700 ;
        RECT 338.800 204.300 339.600 204.400 ;
        RECT 402.800 204.300 403.600 204.400 ;
        RECT 338.800 203.700 403.600 204.300 ;
        RECT 338.800 203.600 339.600 203.700 ;
        RECT 402.800 203.600 403.600 203.700 ;
        RECT 9.200 202.300 10.000 202.400 ;
        RECT 14.000 202.300 14.800 202.400 ;
        RECT 9.200 201.700 14.800 202.300 ;
        RECT 9.200 201.600 10.000 201.700 ;
        RECT 14.000 201.600 14.800 201.700 ;
        RECT 439.600 202.300 440.400 202.400 ;
        RECT 494.000 202.300 494.800 202.400 ;
        RECT 439.600 201.700 494.800 202.300 ;
        RECT 439.600 201.600 440.400 201.700 ;
        RECT 494.000 201.600 494.800 201.700 ;
        RECT 503.600 202.300 504.400 202.400 ;
        RECT 506.800 202.300 507.600 202.400 ;
        RECT 503.600 201.700 507.600 202.300 ;
        RECT 503.600 201.600 504.400 201.700 ;
        RECT 506.800 201.600 507.600 201.700 ;
        RECT 252.400 200.300 253.200 200.400 ;
        RECT 255.600 200.300 256.400 200.400 ;
        RECT 270.000 200.300 270.800 200.400 ;
        RECT 278.000 200.300 278.800 200.400 ;
        RECT 252.400 199.700 278.800 200.300 ;
        RECT 252.400 199.600 253.200 199.700 ;
        RECT 255.600 199.600 256.400 199.700 ;
        RECT 270.000 199.600 270.800 199.700 ;
        RECT 278.000 199.600 278.800 199.700 ;
        RECT 281.200 200.300 282.000 200.400 ;
        RECT 322.800 200.300 323.600 200.400 ;
        RECT 281.200 199.700 323.600 200.300 ;
        RECT 281.200 199.600 282.000 199.700 ;
        RECT 322.800 199.600 323.600 199.700 ;
        RECT 679.600 200.300 680.400 200.400 ;
        RECT 682.800 200.300 683.600 200.400 ;
        RECT 679.600 199.700 683.600 200.300 ;
        RECT 679.600 199.600 680.400 199.700 ;
        RECT 682.800 199.600 683.600 199.700 ;
        RECT 63.600 198.300 64.400 198.400 ;
        RECT 209.200 198.300 210.000 198.400 ;
        RECT 63.600 197.700 210.000 198.300 ;
        RECT 63.600 197.600 64.400 197.700 ;
        RECT 209.200 197.600 210.000 197.700 ;
        RECT 324.400 198.300 325.200 198.400 ;
        RECT 358.000 198.300 358.800 198.400 ;
        RECT 324.400 197.700 358.800 198.300 ;
        RECT 324.400 197.600 325.200 197.700 ;
        RECT 358.000 197.600 358.800 197.700 ;
        RECT 375.600 198.300 376.400 198.400 ;
        RECT 380.400 198.300 381.200 198.400 ;
        RECT 375.600 197.700 381.200 198.300 ;
        RECT 375.600 197.600 376.400 197.700 ;
        RECT 380.400 197.600 381.200 197.700 ;
        RECT 382.000 198.300 382.800 198.400 ;
        RECT 417.200 198.300 418.000 198.400 ;
        RECT 382.000 197.700 418.000 198.300 ;
        RECT 382.000 197.600 382.800 197.700 ;
        RECT 417.200 197.600 418.000 197.700 ;
        RECT 426.800 198.300 427.600 198.400 ;
        RECT 428.400 198.300 429.200 198.400 ;
        RECT 426.800 197.700 429.200 198.300 ;
        RECT 426.800 197.600 427.600 197.700 ;
        RECT 428.400 197.600 429.200 197.700 ;
        RECT 446.000 198.300 446.800 198.400 ;
        RECT 466.800 198.300 467.600 198.400 ;
        RECT 446.000 197.700 467.600 198.300 ;
        RECT 446.000 197.600 446.800 197.700 ;
        RECT 466.800 197.600 467.600 197.700 ;
        RECT 618.800 198.300 619.600 198.400 ;
        RECT 634.800 198.300 635.600 198.400 ;
        RECT 618.800 197.700 635.600 198.300 ;
        RECT 618.800 197.600 619.600 197.700 ;
        RECT 634.800 197.600 635.600 197.700 ;
        RECT 652.400 198.300 653.200 198.400 ;
        RECT 682.800 198.300 683.600 198.400 ;
        RECT 652.400 197.700 683.600 198.300 ;
        RECT 652.400 197.600 653.200 197.700 ;
        RECT 682.800 197.600 683.600 197.700 ;
        RECT 49.200 196.300 50.000 196.400 ;
        RECT 105.200 196.300 106.000 196.400 ;
        RECT 49.200 195.700 106.000 196.300 ;
        RECT 49.200 195.600 50.000 195.700 ;
        RECT 105.200 195.600 106.000 195.700 ;
        RECT 180.400 196.300 181.200 196.400 ;
        RECT 226.800 196.300 227.600 196.400 ;
        RECT 370.800 196.300 371.600 196.400 ;
        RECT 465.200 196.300 466.000 196.400 ;
        RECT 180.400 195.700 466.000 196.300 ;
        RECT 180.400 195.600 181.200 195.700 ;
        RECT 226.800 195.600 227.600 195.700 ;
        RECT 370.800 195.600 371.600 195.700 ;
        RECT 465.200 195.600 466.000 195.700 ;
        RECT 466.800 196.300 467.600 196.400 ;
        RECT 518.000 196.300 518.800 196.400 ;
        RECT 522.800 196.300 523.600 196.400 ;
        RECT 466.800 195.700 523.600 196.300 ;
        RECT 466.800 195.600 467.600 195.700 ;
        RECT 518.000 195.600 518.800 195.700 ;
        RECT 522.800 195.600 523.600 195.700 ;
        RECT 582.000 196.300 582.800 196.400 ;
        RECT 636.400 196.300 637.200 196.400 ;
        RECT 582.000 195.700 637.200 196.300 ;
        RECT 582.000 195.600 582.800 195.700 ;
        RECT 636.400 195.600 637.200 195.700 ;
        RECT 647.600 196.300 648.400 196.400 ;
        RECT 654.000 196.300 654.800 196.400 ;
        RECT 647.600 195.700 654.800 196.300 ;
        RECT 647.600 195.600 648.400 195.700 ;
        RECT 654.000 195.600 654.800 195.700 ;
        RECT 663.600 195.600 664.400 196.400 ;
        RECT 57.200 194.300 58.000 194.400 ;
        RECT 79.600 194.300 80.400 194.400 ;
        RECT 57.200 193.700 80.400 194.300 ;
        RECT 57.200 193.600 58.000 193.700 ;
        RECT 79.600 193.600 80.400 193.700 ;
        RECT 372.400 194.300 373.200 194.400 ;
        RECT 375.600 194.300 376.400 194.400 ;
        RECT 372.400 193.700 376.400 194.300 ;
        RECT 372.400 193.600 373.200 193.700 ;
        RECT 375.600 193.600 376.400 193.700 ;
        RECT 390.000 194.300 390.800 194.400 ;
        RECT 398.000 194.300 398.800 194.400 ;
        RECT 404.400 194.300 405.200 194.400 ;
        RECT 390.000 193.700 405.200 194.300 ;
        RECT 390.000 193.600 390.800 193.700 ;
        RECT 398.000 193.600 398.800 193.700 ;
        RECT 404.400 193.600 405.200 193.700 ;
        RECT 436.400 194.300 437.200 194.400 ;
        RECT 481.200 194.300 482.000 194.400 ;
        RECT 495.600 194.300 496.400 194.400 ;
        RECT 436.400 193.700 496.400 194.300 ;
        RECT 436.400 193.600 437.200 193.700 ;
        RECT 481.200 193.600 482.000 193.700 ;
        RECT 495.600 193.600 496.400 193.700 ;
        RECT 559.600 194.300 560.400 194.400 ;
        RECT 578.800 194.300 579.600 194.400 ;
        RECT 559.600 193.700 579.600 194.300 ;
        RECT 559.600 193.600 560.400 193.700 ;
        RECT 578.800 193.600 579.600 193.700 ;
        RECT 622.000 194.300 622.800 194.400 ;
        RECT 631.600 194.300 632.400 194.400 ;
        RECT 639.600 194.300 640.400 194.400 ;
        RECT 650.800 194.300 651.600 194.400 ;
        RECT 622.000 193.700 640.400 194.300 ;
        RECT 622.000 193.600 622.800 193.700 ;
        RECT 631.600 193.600 632.400 193.700 ;
        RECT 639.600 193.600 640.400 193.700 ;
        RECT 642.900 193.700 651.600 194.300 ;
        RECT 9.200 192.300 10.000 192.400 ;
        RECT 50.800 192.300 51.600 192.400 ;
        RECT 9.200 191.700 51.600 192.300 ;
        RECT 9.200 191.600 10.000 191.700 ;
        RECT 50.800 191.600 51.600 191.700 ;
        RECT 71.600 192.300 72.400 192.400 ;
        RECT 76.400 192.300 77.200 192.400 ;
        RECT 71.600 191.700 77.200 192.300 ;
        RECT 71.600 191.600 72.400 191.700 ;
        RECT 76.400 191.600 77.200 191.700 ;
        RECT 82.800 192.300 83.600 192.400 ;
        RECT 140.400 192.300 141.200 192.400 ;
        RECT 82.800 191.700 141.200 192.300 ;
        RECT 82.800 191.600 83.600 191.700 ;
        RECT 140.400 191.600 141.200 191.700 ;
        RECT 210.800 192.300 211.600 192.400 ;
        RECT 238.000 192.300 238.800 192.400 ;
        RECT 210.800 191.700 238.800 192.300 ;
        RECT 210.800 191.600 211.600 191.700 ;
        RECT 238.000 191.600 238.800 191.700 ;
        RECT 330.800 192.300 331.600 192.400 ;
        RECT 340.400 192.300 341.200 192.400 ;
        RECT 330.800 191.700 341.200 192.300 ;
        RECT 330.800 191.600 331.600 191.700 ;
        RECT 340.400 191.600 341.200 191.700 ;
        RECT 346.800 192.300 347.600 192.400 ;
        RECT 375.600 192.300 376.400 192.400 ;
        RECT 382.000 192.300 382.800 192.400 ;
        RECT 346.800 191.700 382.800 192.300 ;
        RECT 346.800 191.600 347.600 191.700 ;
        RECT 375.600 191.600 376.400 191.700 ;
        RECT 382.000 191.600 382.800 191.700 ;
        RECT 393.200 192.300 394.000 192.400 ;
        RECT 401.200 192.300 402.000 192.400 ;
        RECT 393.200 191.700 402.000 192.300 ;
        RECT 393.200 191.600 394.000 191.700 ;
        RECT 401.200 191.600 402.000 191.700 ;
        RECT 436.400 192.300 437.200 192.400 ;
        RECT 455.600 192.300 456.400 192.400 ;
        RECT 436.400 191.700 456.400 192.300 ;
        RECT 436.400 191.600 437.200 191.700 ;
        RECT 455.600 191.600 456.400 191.700 ;
        RECT 465.200 192.300 466.000 192.400 ;
        RECT 484.400 192.300 485.200 192.400 ;
        RECT 487.600 192.300 488.400 192.400 ;
        RECT 465.200 191.700 488.400 192.300 ;
        RECT 465.200 191.600 466.000 191.700 ;
        RECT 484.400 191.600 485.200 191.700 ;
        RECT 487.600 191.600 488.400 191.700 ;
        RECT 575.600 192.300 576.400 192.400 ;
        RECT 598.000 192.300 598.800 192.400 ;
        RECT 575.600 191.700 598.800 192.300 ;
        RECT 575.600 191.600 576.400 191.700 ;
        RECT 598.000 191.600 598.800 191.700 ;
        RECT 620.400 192.300 621.200 192.400 ;
        RECT 628.400 192.300 629.200 192.400 ;
        RECT 620.400 191.700 629.200 192.300 ;
        RECT 620.400 191.600 621.200 191.700 ;
        RECT 628.400 191.600 629.200 191.700 ;
        RECT 630.000 192.300 630.800 192.400 ;
        RECT 642.900 192.300 643.500 193.700 ;
        RECT 650.800 193.600 651.600 193.700 ;
        RECT 657.200 194.300 658.000 194.400 ;
        RECT 671.600 194.300 672.400 194.400 ;
        RECT 657.200 193.700 672.400 194.300 ;
        RECT 657.200 193.600 658.000 193.700 ;
        RECT 671.600 193.600 672.400 193.700 ;
        RECT 676.400 194.300 677.200 194.400 ;
        RECT 678.000 194.300 678.800 194.400 ;
        RECT 676.400 193.700 678.800 194.300 ;
        RECT 676.400 193.600 677.200 193.700 ;
        RECT 678.000 193.600 678.800 193.700 ;
        RECT 630.000 191.700 643.500 192.300 ;
        RECT 644.400 192.300 645.200 192.400 ;
        RECT 649.200 192.300 650.000 192.400 ;
        RECT 676.400 192.300 677.200 192.400 ;
        RECT 644.400 191.700 677.200 192.300 ;
        RECT 630.000 191.600 630.800 191.700 ;
        RECT 644.400 191.600 645.200 191.700 ;
        RECT 649.200 191.600 650.000 191.700 ;
        RECT 676.400 191.600 677.200 191.700 ;
        RECT 6.000 190.300 6.800 190.400 ;
        RECT 7.600 190.300 8.400 190.400 ;
        RECT 63.600 190.300 64.400 190.400 ;
        RECT 6.000 189.700 64.400 190.300 ;
        RECT 6.000 189.600 6.800 189.700 ;
        RECT 7.600 189.600 8.400 189.700 ;
        RECT 63.600 189.600 64.400 189.700 ;
        RECT 70.000 190.300 70.800 190.400 ;
        RECT 73.200 190.300 74.000 190.400 ;
        RECT 70.000 189.700 74.000 190.300 ;
        RECT 70.000 189.600 70.800 189.700 ;
        RECT 73.200 189.600 74.000 189.700 ;
        RECT 90.800 189.600 91.600 190.400 ;
        RECT 150.000 190.300 150.800 190.400 ;
        RECT 164.400 190.300 165.200 190.400 ;
        RECT 150.000 189.700 165.200 190.300 ;
        RECT 150.000 189.600 150.800 189.700 ;
        RECT 164.400 189.600 165.200 189.700 ;
        RECT 214.000 190.300 214.800 190.400 ;
        RECT 217.200 190.300 218.000 190.400 ;
        RECT 225.200 190.300 226.000 190.400 ;
        RECT 214.000 189.700 226.000 190.300 ;
        RECT 214.000 189.600 214.800 189.700 ;
        RECT 217.200 189.600 218.000 189.700 ;
        RECT 225.200 189.600 226.000 189.700 ;
        RECT 300.400 190.300 301.200 190.400 ;
        RECT 310.000 190.300 310.800 190.400 ;
        RECT 300.400 189.700 310.800 190.300 ;
        RECT 300.400 189.600 301.200 189.700 ;
        RECT 310.000 189.600 310.800 189.700 ;
        RECT 319.600 190.300 320.400 190.400 ;
        RECT 340.400 190.300 341.200 190.400 ;
        RECT 319.600 189.700 341.200 190.300 ;
        RECT 319.600 189.600 320.400 189.700 ;
        RECT 340.400 189.600 341.200 189.700 ;
        RECT 345.200 190.300 346.000 190.400 ;
        RECT 383.600 190.300 384.400 190.400 ;
        RECT 345.200 189.700 384.400 190.300 ;
        RECT 345.200 189.600 346.000 189.700 ;
        RECT 383.600 189.600 384.400 189.700 ;
        RECT 402.800 190.300 403.600 190.400 ;
        RECT 404.400 190.300 405.200 190.400 ;
        RECT 402.800 189.700 405.200 190.300 ;
        RECT 402.800 189.600 403.600 189.700 ;
        RECT 404.400 189.600 405.200 189.700 ;
        RECT 417.200 190.300 418.000 190.400 ;
        RECT 462.000 190.300 462.800 190.400 ;
        RECT 417.200 189.700 462.800 190.300 ;
        RECT 417.200 189.600 418.000 189.700 ;
        RECT 462.000 189.600 462.800 189.700 ;
        RECT 465.200 190.300 466.000 190.400 ;
        RECT 468.400 190.300 469.200 190.400 ;
        RECT 465.200 189.700 469.200 190.300 ;
        RECT 465.200 189.600 466.000 189.700 ;
        RECT 468.400 189.600 469.200 189.700 ;
        RECT 476.400 190.300 477.200 190.400 ;
        RECT 487.600 190.300 488.400 190.400 ;
        RECT 476.400 189.700 488.400 190.300 ;
        RECT 476.400 189.600 477.200 189.700 ;
        RECT 487.600 189.600 488.400 189.700 ;
        RECT 545.200 190.300 546.000 190.400 ;
        RECT 561.200 190.300 562.000 190.400 ;
        RECT 545.200 189.700 562.000 190.300 ;
        RECT 545.200 189.600 546.000 189.700 ;
        RECT 561.200 189.600 562.000 189.700 ;
        RECT 564.400 190.300 565.200 190.400 ;
        RECT 577.200 190.300 578.000 190.400 ;
        RECT 564.400 189.700 578.000 190.300 ;
        RECT 564.400 189.600 565.200 189.700 ;
        RECT 577.200 189.600 578.000 189.700 ;
        RECT 588.400 190.300 589.200 190.400 ;
        RECT 609.200 190.300 610.000 190.400 ;
        RECT 588.400 189.700 610.000 190.300 ;
        RECT 588.400 189.600 589.200 189.700 ;
        RECT 609.200 189.600 610.000 189.700 ;
        RECT 623.600 190.300 624.400 190.400 ;
        RECT 665.200 190.300 666.000 190.400 ;
        RECT 623.600 189.700 666.000 190.300 ;
        RECT 623.600 189.600 624.400 189.700 ;
        RECT 665.200 189.600 666.000 189.700 ;
        RECT 671.600 190.300 672.400 190.400 ;
        RECT 687.600 190.300 688.400 190.400 ;
        RECT 671.600 189.700 688.400 190.300 ;
        RECT 671.600 189.600 672.400 189.700 ;
        RECT 687.600 189.600 688.400 189.700 ;
        RECT 15.600 188.300 16.400 188.400 ;
        RECT 17.200 188.300 18.000 188.400 ;
        RECT 15.600 187.700 18.000 188.300 ;
        RECT 15.600 187.600 16.400 187.700 ;
        RECT 17.200 187.600 18.000 187.700 ;
        RECT 55.600 188.300 56.400 188.400 ;
        RECT 60.400 188.300 61.200 188.400 ;
        RECT 55.600 187.700 61.200 188.300 ;
        RECT 55.600 187.600 56.400 187.700 ;
        RECT 60.400 187.600 61.200 187.700 ;
        RECT 65.200 188.300 66.000 188.400 ;
        RECT 78.000 188.300 78.800 188.400 ;
        RECT 84.400 188.300 85.200 188.400 ;
        RECT 108.400 188.300 109.200 188.400 ;
        RECT 119.600 188.300 120.400 188.400 ;
        RECT 65.200 187.700 120.400 188.300 ;
        RECT 65.200 187.600 66.000 187.700 ;
        RECT 78.000 187.600 78.800 187.700 ;
        RECT 84.400 187.600 85.200 187.700 ;
        RECT 108.400 187.600 109.200 187.700 ;
        RECT 119.600 187.600 120.400 187.700 ;
        RECT 142.000 188.300 142.800 188.400 ;
        RECT 220.400 188.300 221.200 188.400 ;
        RECT 230.000 188.300 230.800 188.400 ;
        RECT 142.000 187.700 230.800 188.300 ;
        RECT 142.000 187.600 142.800 187.700 ;
        RECT 220.400 187.600 221.200 187.700 ;
        RECT 230.000 187.600 230.800 187.700 ;
        RECT 260.400 188.300 261.200 188.400 ;
        RECT 289.200 188.300 290.000 188.400 ;
        RECT 260.400 187.700 290.000 188.300 ;
        RECT 260.400 187.600 261.200 187.700 ;
        RECT 289.200 187.600 290.000 187.700 ;
        RECT 338.800 188.300 339.600 188.400 ;
        RECT 350.000 188.300 350.800 188.400 ;
        RECT 338.800 187.700 350.800 188.300 ;
        RECT 338.800 187.600 339.600 187.700 ;
        RECT 350.000 187.600 350.800 187.700 ;
        RECT 361.200 188.300 362.000 188.400 ;
        RECT 369.200 188.300 370.000 188.400 ;
        RECT 372.400 188.300 373.200 188.400 ;
        RECT 361.200 187.700 373.200 188.300 ;
        RECT 361.200 187.600 362.000 187.700 ;
        RECT 369.200 187.600 370.000 187.700 ;
        RECT 372.400 187.600 373.200 187.700 ;
        RECT 407.600 188.300 408.400 188.400 ;
        RECT 420.400 188.300 421.200 188.400 ;
        RECT 436.400 188.300 437.200 188.400 ;
        RECT 407.600 187.700 437.200 188.300 ;
        RECT 407.600 187.600 408.400 187.700 ;
        RECT 420.400 187.600 421.200 187.700 ;
        RECT 436.400 187.600 437.200 187.700 ;
        RECT 446.000 188.300 446.800 188.400 ;
        RECT 465.200 188.300 466.000 188.400 ;
        RECT 446.000 187.700 466.000 188.300 ;
        RECT 446.000 187.600 446.800 187.700 ;
        RECT 465.200 187.600 466.000 187.700 ;
        RECT 468.400 188.300 469.200 188.400 ;
        RECT 516.400 188.300 517.200 188.400 ;
        RECT 468.400 187.700 517.200 188.300 ;
        RECT 468.400 187.600 469.200 187.700 ;
        RECT 516.400 187.600 517.200 187.700 ;
        RECT 519.600 188.300 520.400 188.400 ;
        RECT 545.200 188.300 546.000 188.400 ;
        RECT 519.600 187.700 546.000 188.300 ;
        RECT 519.600 187.600 520.400 187.700 ;
        RECT 545.200 187.600 546.000 187.700 ;
        RECT 569.200 188.300 570.000 188.400 ;
        RECT 596.400 188.300 597.200 188.400 ;
        RECT 617.200 188.300 618.000 188.400 ;
        RECT 569.200 187.700 618.000 188.300 ;
        RECT 569.200 187.600 570.000 187.700 ;
        RECT 596.400 187.600 597.200 187.700 ;
        RECT 617.200 187.600 618.000 187.700 ;
        RECT 625.200 188.300 626.000 188.400 ;
        RECT 630.000 188.300 630.800 188.400 ;
        RECT 625.200 187.700 630.800 188.300 ;
        RECT 625.200 187.600 626.000 187.700 ;
        RECT 630.000 187.600 630.800 187.700 ;
        RECT 631.600 188.300 632.400 188.400 ;
        RECT 647.600 188.300 648.400 188.400 ;
        RECT 676.400 188.300 677.200 188.400 ;
        RECT 631.600 187.700 677.200 188.300 ;
        RECT 631.600 187.600 632.400 187.700 ;
        RECT 647.600 187.600 648.400 187.700 ;
        RECT 676.400 187.600 677.200 187.700 ;
        RECT 9.200 186.300 10.000 186.400 ;
        RECT 30.000 186.300 30.800 186.400 ;
        RECT 9.200 185.700 30.800 186.300 ;
        RECT 9.200 185.600 10.000 185.700 ;
        RECT 30.000 185.600 30.800 185.700 ;
        RECT 33.200 186.300 34.000 186.400 ;
        RECT 47.600 186.300 48.400 186.400 ;
        RECT 33.200 185.700 48.400 186.300 ;
        RECT 33.200 185.600 34.000 185.700 ;
        RECT 47.600 185.600 48.400 185.700 ;
        RECT 62.000 186.300 62.800 186.400 ;
        RECT 70.000 186.300 70.800 186.400 ;
        RECT 62.000 185.700 70.800 186.300 ;
        RECT 62.000 185.600 62.800 185.700 ;
        RECT 70.000 185.600 70.800 185.700 ;
        RECT 92.400 186.300 93.200 186.400 ;
        RECT 122.800 186.300 123.600 186.400 ;
        RECT 92.400 185.700 123.600 186.300 ;
        RECT 92.400 185.600 93.200 185.700 ;
        RECT 122.800 185.600 123.600 185.700 ;
        RECT 170.800 186.300 171.600 186.400 ;
        RECT 199.600 186.300 200.400 186.400 ;
        RECT 170.800 185.700 200.400 186.300 ;
        RECT 170.800 185.600 171.600 185.700 ;
        RECT 199.600 185.600 200.400 185.700 ;
        RECT 202.800 186.300 203.600 186.400 ;
        RECT 212.400 186.300 213.200 186.400 ;
        RECT 202.800 185.700 213.200 186.300 ;
        RECT 202.800 185.600 203.600 185.700 ;
        RECT 212.400 185.600 213.200 185.700 ;
        RECT 223.600 186.300 224.400 186.400 ;
        RECT 249.200 186.300 250.000 186.400 ;
        RECT 223.600 185.700 250.000 186.300 ;
        RECT 223.600 185.600 224.400 185.700 ;
        RECT 249.200 185.600 250.000 185.700 ;
        RECT 305.200 186.300 306.000 186.400 ;
        RECT 308.400 186.300 309.200 186.400 ;
        RECT 305.200 185.700 309.200 186.300 ;
        RECT 305.200 185.600 306.000 185.700 ;
        RECT 308.400 185.600 309.200 185.700 ;
        RECT 322.800 186.300 323.600 186.400 ;
        RECT 356.400 186.300 357.200 186.400 ;
        RECT 322.800 185.700 357.200 186.300 ;
        RECT 322.800 185.600 323.600 185.700 ;
        RECT 356.400 185.600 357.200 185.700 ;
        RECT 396.400 186.300 397.200 186.400 ;
        RECT 401.200 186.300 402.000 186.400 ;
        RECT 396.400 185.700 402.000 186.300 ;
        RECT 396.400 185.600 397.200 185.700 ;
        RECT 401.200 185.600 402.000 185.700 ;
        RECT 433.200 186.300 434.000 186.400 ;
        RECT 444.400 186.300 445.200 186.400 ;
        RECT 470.000 186.300 470.800 186.400 ;
        RECT 433.200 185.700 470.800 186.300 ;
        RECT 433.200 185.600 434.000 185.700 ;
        RECT 444.400 185.600 445.200 185.700 ;
        RECT 470.000 185.600 470.800 185.700 ;
        RECT 516.400 186.300 517.200 186.400 ;
        RECT 524.400 186.300 525.200 186.400 ;
        RECT 526.000 186.300 526.800 186.400 ;
        RECT 516.400 185.700 526.800 186.300 ;
        RECT 516.400 185.600 517.200 185.700 ;
        RECT 524.400 185.600 525.200 185.700 ;
        RECT 526.000 185.600 526.800 185.700 ;
        RECT 558.000 186.300 558.800 186.400 ;
        RECT 585.200 186.300 586.000 186.400 ;
        RECT 590.000 186.300 590.800 186.400 ;
        RECT 558.000 185.700 590.800 186.300 ;
        RECT 558.000 185.600 558.800 185.700 ;
        RECT 585.200 185.600 586.000 185.700 ;
        RECT 590.000 185.600 590.800 185.700 ;
        RECT 598.000 186.300 598.800 186.400 ;
        RECT 612.400 186.300 613.200 186.400 ;
        RECT 660.400 186.300 661.200 186.400 ;
        RECT 598.000 185.700 661.200 186.300 ;
        RECT 598.000 185.600 598.800 185.700 ;
        RECT 612.400 185.600 613.200 185.700 ;
        RECT 660.400 185.600 661.200 185.700 ;
        RECT 663.600 186.300 664.400 186.400 ;
        RECT 666.800 186.300 667.600 186.400 ;
        RECT 670.000 186.300 670.800 186.400 ;
        RECT 663.600 185.700 670.800 186.300 ;
        RECT 663.600 185.600 664.400 185.700 ;
        RECT 666.800 185.600 667.600 185.700 ;
        RECT 670.000 185.600 670.800 185.700 ;
        RECT 14.000 183.600 14.800 184.400 ;
        RECT 174.000 184.300 174.800 184.400 ;
        RECT 183.600 184.300 184.400 184.400 ;
        RECT 199.700 184.300 200.300 185.600 ;
        RECT 246.000 184.300 246.800 184.400 ;
        RECT 174.000 183.700 198.700 184.300 ;
        RECT 199.700 183.700 246.800 184.300 ;
        RECT 174.000 183.600 174.800 183.700 ;
        RECT 183.600 183.600 184.400 183.700 ;
        RECT 17.200 182.300 18.000 182.400 ;
        RECT 58.800 182.300 59.600 182.400 ;
        RECT 17.200 181.700 59.600 182.300 ;
        RECT 17.200 181.600 18.000 181.700 ;
        RECT 58.800 181.600 59.600 181.700 ;
        RECT 169.200 182.300 170.000 182.400 ;
        RECT 188.400 182.300 189.200 182.400 ;
        RECT 169.200 181.700 189.200 182.300 ;
        RECT 198.100 182.300 198.700 183.700 ;
        RECT 246.000 183.600 246.800 183.700 ;
        RECT 369.200 184.300 370.000 184.400 ;
        RECT 383.600 184.300 384.400 184.400 ;
        RECT 369.200 183.700 384.400 184.300 ;
        RECT 369.200 183.600 370.000 183.700 ;
        RECT 383.600 183.600 384.400 183.700 ;
        RECT 410.800 184.300 411.600 184.400 ;
        RECT 412.400 184.300 413.200 184.400 ;
        RECT 474.800 184.300 475.600 184.400 ;
        RECT 410.800 183.700 475.600 184.300 ;
        RECT 410.800 183.600 411.600 183.700 ;
        RECT 412.400 183.600 413.200 183.700 ;
        RECT 474.800 183.600 475.600 183.700 ;
        RECT 518.000 184.300 518.800 184.400 ;
        RECT 530.800 184.300 531.600 184.400 ;
        RECT 518.000 183.700 531.600 184.300 ;
        RECT 518.000 183.600 518.800 183.700 ;
        RECT 530.800 183.600 531.600 183.700 ;
        RECT 532.400 184.300 533.200 184.400 ;
        RECT 537.200 184.300 538.000 184.400 ;
        RECT 532.400 183.700 538.000 184.300 ;
        RECT 532.400 183.600 533.200 183.700 ;
        RECT 537.200 183.600 538.000 183.700 ;
        RECT 556.400 184.300 557.200 184.400 ;
        RECT 562.800 184.300 563.600 184.400 ;
        RECT 556.400 183.700 563.600 184.300 ;
        RECT 556.400 183.600 557.200 183.700 ;
        RECT 562.800 183.600 563.600 183.700 ;
        RECT 567.600 184.300 568.400 184.400 ;
        RECT 582.000 184.300 582.800 184.400 ;
        RECT 567.600 183.700 582.800 184.300 ;
        RECT 567.600 183.600 568.400 183.700 ;
        RECT 582.000 183.600 582.800 183.700 ;
        RECT 591.600 184.300 592.400 184.400 ;
        RECT 598.000 184.300 598.800 184.400 ;
        RECT 591.600 183.700 598.800 184.300 ;
        RECT 591.600 183.600 592.400 183.700 ;
        RECT 598.000 183.600 598.800 183.700 ;
        RECT 615.600 184.300 616.400 184.400 ;
        RECT 618.800 184.300 619.600 184.400 ;
        RECT 615.600 183.700 619.600 184.300 ;
        RECT 615.600 183.600 616.400 183.700 ;
        RECT 618.800 183.600 619.600 183.700 ;
        RECT 650.800 184.300 651.600 184.400 ;
        RECT 678.000 184.300 678.800 184.400 ;
        RECT 650.800 183.700 678.800 184.300 ;
        RECT 650.800 183.600 651.600 183.700 ;
        RECT 678.000 183.600 678.800 183.700 ;
        RECT 206.000 182.300 206.800 182.400 ;
        RECT 198.100 181.700 206.800 182.300 ;
        RECT 169.200 181.600 170.000 181.700 ;
        RECT 188.400 181.600 189.200 181.700 ;
        RECT 206.000 181.600 206.800 181.700 ;
        RECT 354.800 182.300 355.600 182.400 ;
        RECT 367.600 182.300 368.400 182.400 ;
        RECT 407.600 182.300 408.400 182.400 ;
        RECT 354.800 181.700 408.400 182.300 ;
        RECT 354.800 181.600 355.600 181.700 ;
        RECT 367.600 181.600 368.400 181.700 ;
        RECT 407.600 181.600 408.400 181.700 ;
        RECT 447.600 182.300 448.400 182.400 ;
        RECT 452.400 182.300 453.200 182.400 ;
        RECT 447.600 181.700 453.200 182.300 ;
        RECT 447.600 181.600 448.400 181.700 ;
        RECT 452.400 181.600 453.200 181.700 ;
        RECT 458.800 182.300 459.600 182.400 ;
        RECT 489.200 182.300 490.000 182.400 ;
        RECT 458.800 181.700 490.000 182.300 ;
        RECT 458.800 181.600 459.600 181.700 ;
        RECT 489.200 181.600 490.000 181.700 ;
        RECT 521.200 182.300 522.000 182.400 ;
        RECT 530.800 182.300 531.600 182.400 ;
        RECT 554.800 182.300 555.600 182.400 ;
        RECT 521.200 181.700 555.600 182.300 ;
        RECT 521.200 181.600 522.000 181.700 ;
        RECT 530.800 181.600 531.600 181.700 ;
        RECT 554.800 181.600 555.600 181.700 ;
        RECT 612.400 182.300 613.200 182.400 ;
        RECT 622.000 182.300 622.800 182.400 ;
        RECT 612.400 181.700 622.800 182.300 ;
        RECT 612.400 181.600 613.200 181.700 ;
        RECT 622.000 181.600 622.800 181.700 ;
        RECT 636.400 182.300 637.200 182.400 ;
        RECT 660.400 182.300 661.200 182.400 ;
        RECT 636.400 181.700 661.200 182.300 ;
        RECT 636.400 181.600 637.200 181.700 ;
        RECT 660.400 181.600 661.200 181.700 ;
        RECT 662.000 182.300 662.800 182.400 ;
        RECT 665.200 182.300 666.000 182.400 ;
        RECT 662.000 181.700 666.000 182.300 ;
        RECT 662.000 181.600 662.800 181.700 ;
        RECT 665.200 181.600 666.000 181.700 ;
        RECT 673.200 182.300 674.000 182.400 ;
        RECT 682.800 182.300 683.600 182.400 ;
        RECT 673.200 181.700 683.600 182.300 ;
        RECT 673.200 181.600 674.000 181.700 ;
        RECT 682.800 181.600 683.600 181.700 ;
        RECT 154.800 180.300 155.600 180.400 ;
        RECT 217.200 180.300 218.000 180.400 ;
        RECT 154.800 179.700 218.000 180.300 ;
        RECT 154.800 179.600 155.600 179.700 ;
        RECT 217.200 179.600 218.000 179.700 ;
        RECT 335.600 180.300 336.400 180.400 ;
        RECT 340.400 180.300 341.200 180.400 ;
        RECT 366.000 180.300 366.800 180.400 ;
        RECT 377.200 180.300 378.000 180.400 ;
        RECT 409.200 180.300 410.000 180.400 ;
        RECT 335.600 179.700 410.000 180.300 ;
        RECT 335.600 179.600 336.400 179.700 ;
        RECT 340.400 179.600 341.200 179.700 ;
        RECT 366.000 179.600 366.800 179.700 ;
        RECT 377.200 179.600 378.000 179.700 ;
        RECT 409.200 179.600 410.000 179.700 ;
        RECT 513.200 180.300 514.000 180.400 ;
        RECT 532.400 180.300 533.200 180.400 ;
        RECT 513.200 179.700 533.200 180.300 ;
        RECT 513.200 179.600 514.000 179.700 ;
        RECT 532.400 179.600 533.200 179.700 ;
        RECT 641.200 180.300 642.000 180.400 ;
        RECT 655.600 180.300 656.400 180.400 ;
        RECT 658.800 180.300 659.600 180.400 ;
        RECT 641.200 179.700 659.600 180.300 ;
        RECT 641.200 179.600 642.000 179.700 ;
        RECT 655.600 179.600 656.400 179.700 ;
        RECT 658.800 179.600 659.600 179.700 ;
        RECT 674.800 180.300 675.600 180.400 ;
        RECT 684.400 180.300 685.200 180.400 ;
        RECT 674.800 179.700 685.200 180.300 ;
        RECT 674.800 179.600 675.600 179.700 ;
        RECT 684.400 179.600 685.200 179.700 ;
        RECT 52.400 178.300 53.200 178.400 ;
        RECT 79.600 178.300 80.400 178.400 ;
        RECT 52.400 177.700 80.400 178.300 ;
        RECT 52.400 177.600 53.200 177.700 ;
        RECT 79.600 177.600 80.400 177.700 ;
        RECT 118.000 178.300 118.800 178.400 ;
        RECT 258.800 178.300 259.600 178.400 ;
        RECT 270.000 178.300 270.800 178.400 ;
        RECT 353.200 178.300 354.000 178.400 ;
        RECT 412.400 178.300 413.200 178.400 ;
        RECT 118.000 177.700 270.800 178.300 ;
        RECT 118.000 177.600 118.800 177.700 ;
        RECT 258.800 177.600 259.600 177.700 ;
        RECT 270.000 177.600 270.800 177.700 ;
        RECT 271.700 177.700 413.200 178.300 ;
        RECT 17.200 176.300 18.000 176.400 ;
        RECT 33.200 176.300 34.000 176.400 ;
        RECT 38.000 176.300 38.800 176.400 ;
        RECT 17.200 175.700 38.800 176.300 ;
        RECT 17.200 175.600 18.000 175.700 ;
        RECT 33.200 175.600 34.000 175.700 ;
        RECT 38.000 175.600 38.800 175.700 ;
        RECT 63.600 176.300 64.400 176.400 ;
        RECT 70.000 176.300 70.800 176.400 ;
        RECT 63.600 175.700 70.800 176.300 ;
        RECT 63.600 175.600 64.400 175.700 ;
        RECT 70.000 175.600 70.800 175.700 ;
        RECT 134.000 176.300 134.800 176.400 ;
        RECT 140.400 176.300 141.200 176.400 ;
        RECT 134.000 175.700 141.200 176.300 ;
        RECT 134.000 175.600 134.800 175.700 ;
        RECT 140.400 175.600 141.200 175.700 ;
        RECT 150.000 176.300 150.800 176.400 ;
        RECT 158.000 176.300 158.800 176.400 ;
        RECT 150.000 175.700 158.800 176.300 ;
        RECT 150.000 175.600 150.800 175.700 ;
        RECT 158.000 175.600 158.800 175.700 ;
        RECT 161.200 176.300 162.000 176.400 ;
        RECT 169.200 176.300 170.000 176.400 ;
        RECT 198.000 176.300 198.800 176.400 ;
        RECT 161.200 175.700 198.800 176.300 ;
        RECT 161.200 175.600 162.000 175.700 ;
        RECT 169.200 175.600 170.000 175.700 ;
        RECT 198.000 175.600 198.800 175.700 ;
        RECT 209.200 176.300 210.000 176.400 ;
        RECT 265.200 176.300 266.000 176.400 ;
        RECT 271.700 176.300 272.300 177.700 ;
        RECT 353.200 177.600 354.000 177.700 ;
        RECT 412.400 177.600 413.200 177.700 ;
        RECT 436.400 178.300 437.200 178.400 ;
        RECT 458.800 178.300 459.600 178.400 ;
        RECT 436.400 177.700 459.600 178.300 ;
        RECT 436.400 177.600 437.200 177.700 ;
        RECT 458.800 177.600 459.600 177.700 ;
        RECT 506.800 178.300 507.600 178.400 ;
        RECT 521.200 178.300 522.000 178.400 ;
        RECT 540.400 178.300 541.200 178.400 ;
        RECT 506.800 177.700 541.200 178.300 ;
        RECT 506.800 177.600 507.600 177.700 ;
        RECT 521.200 177.600 522.000 177.700 ;
        RECT 540.400 177.600 541.200 177.700 ;
        RECT 577.200 178.300 578.000 178.400 ;
        RECT 586.800 178.300 587.600 178.400 ;
        RECT 577.200 177.700 587.600 178.300 ;
        RECT 577.200 177.600 578.000 177.700 ;
        RECT 586.800 177.600 587.600 177.700 ;
        RECT 646.000 178.300 646.800 178.400 ;
        RECT 663.600 178.300 664.400 178.400 ;
        RECT 646.000 177.700 664.400 178.300 ;
        RECT 646.000 177.600 646.800 177.700 ;
        RECT 663.600 177.600 664.400 177.700 ;
        RECT 666.800 178.300 667.600 178.400 ;
        RECT 671.600 178.300 672.400 178.400 ;
        RECT 666.800 177.700 672.400 178.300 ;
        RECT 666.800 177.600 667.600 177.700 ;
        RECT 671.600 177.600 672.400 177.700 ;
        RECT 209.200 175.700 272.300 176.300 ;
        RECT 314.800 176.300 315.600 176.400 ;
        RECT 337.200 176.300 338.000 176.400 ;
        RECT 314.800 175.700 338.000 176.300 ;
        RECT 209.200 175.600 210.000 175.700 ;
        RECT 265.200 175.600 266.000 175.700 ;
        RECT 314.800 175.600 315.600 175.700 ;
        RECT 337.200 175.600 338.000 175.700 ;
        RECT 406.000 176.300 406.800 176.400 ;
        RECT 450.800 176.300 451.600 176.400 ;
        RECT 406.000 175.700 451.600 176.300 ;
        RECT 406.000 175.600 406.800 175.700 ;
        RECT 450.800 175.600 451.600 175.700 ;
        RECT 484.400 175.600 485.200 176.400 ;
        RECT 490.800 176.300 491.600 176.400 ;
        RECT 542.000 176.300 542.800 176.400 ;
        RECT 490.800 175.700 542.800 176.300 ;
        RECT 490.800 175.600 491.600 175.700 ;
        RECT 542.000 175.600 542.800 175.700 ;
        RECT 554.800 176.300 555.600 176.400 ;
        RECT 578.800 176.300 579.600 176.400 ;
        RECT 598.000 176.300 598.800 176.400 ;
        RECT 554.800 175.700 598.800 176.300 ;
        RECT 554.800 175.600 555.600 175.700 ;
        RECT 578.800 175.600 579.600 175.700 ;
        RECT 598.000 175.600 598.800 175.700 ;
        RECT 614.000 176.300 614.800 176.400 ;
        RECT 617.200 176.300 618.000 176.400 ;
        RECT 614.000 175.700 618.000 176.300 ;
        RECT 614.000 175.600 614.800 175.700 ;
        RECT 617.200 175.600 618.000 175.700 ;
        RECT 623.600 176.300 624.400 176.400 ;
        RECT 630.000 176.300 630.800 176.400 ;
        RECT 623.600 175.700 630.800 176.300 ;
        RECT 623.600 175.600 624.400 175.700 ;
        RECT 630.000 175.600 630.800 175.700 ;
        RECT 658.800 176.300 659.600 176.400 ;
        RECT 679.600 176.300 680.400 176.400 ;
        RECT 658.800 175.700 680.400 176.300 ;
        RECT 658.800 175.600 659.600 175.700 ;
        RECT 679.600 175.600 680.400 175.700 ;
        RECT 6.000 174.300 6.800 174.400 ;
        RECT 14.000 174.300 14.800 174.400 ;
        RECT 6.000 173.700 14.800 174.300 ;
        RECT 6.000 173.600 6.800 173.700 ;
        RECT 14.000 173.600 14.800 173.700 ;
        RECT 30.000 174.300 30.800 174.400 ;
        RECT 58.800 174.300 59.600 174.400 ;
        RECT 65.200 174.300 66.000 174.400 ;
        RECT 30.000 173.700 66.000 174.300 ;
        RECT 30.000 173.600 30.800 173.700 ;
        RECT 58.800 173.600 59.600 173.700 ;
        RECT 65.200 173.600 66.000 173.700 ;
        RECT 68.400 174.300 69.200 174.400 ;
        RECT 89.200 174.300 90.000 174.400 ;
        RECT 68.400 173.700 90.000 174.300 ;
        RECT 68.400 173.600 69.200 173.700 ;
        RECT 89.200 173.600 90.000 173.700 ;
        RECT 137.200 174.300 138.000 174.400 ;
        RECT 166.000 174.300 166.800 174.400 ;
        RECT 194.800 174.300 195.600 174.400 ;
        RECT 202.800 174.300 203.600 174.400 ;
        RECT 204.400 174.300 205.200 174.400 ;
        RECT 137.200 173.700 158.700 174.300 ;
        RECT 137.200 173.600 138.000 173.700 ;
        RECT 158.100 172.400 158.700 173.700 ;
        RECT 166.000 173.700 205.200 174.300 ;
        RECT 166.000 173.600 166.800 173.700 ;
        RECT 194.800 173.600 195.600 173.700 ;
        RECT 202.800 173.600 203.600 173.700 ;
        RECT 204.400 173.600 205.200 173.700 ;
        RECT 209.200 174.300 210.000 174.400 ;
        RECT 214.000 174.300 214.800 174.400 ;
        RECT 255.600 174.300 256.400 174.400 ;
        RECT 263.600 174.300 264.400 174.400 ;
        RECT 209.200 173.700 264.400 174.300 ;
        RECT 209.200 173.600 210.000 173.700 ;
        RECT 214.000 173.600 214.800 173.700 ;
        RECT 255.600 173.600 256.400 173.700 ;
        RECT 263.600 173.600 264.400 173.700 ;
        RECT 279.600 174.300 280.400 174.400 ;
        RECT 284.400 174.300 285.200 174.400 ;
        RECT 279.600 173.700 285.200 174.300 ;
        RECT 279.600 173.600 280.400 173.700 ;
        RECT 284.400 173.600 285.200 173.700 ;
        RECT 313.200 174.300 314.000 174.400 ;
        RECT 318.000 174.300 318.800 174.400 ;
        RECT 346.800 174.300 347.600 174.400 ;
        RECT 313.200 173.700 347.600 174.300 ;
        RECT 313.200 173.600 314.000 173.700 ;
        RECT 318.000 173.600 318.800 173.700 ;
        RECT 346.800 173.600 347.600 173.700 ;
        RECT 386.800 174.300 387.600 174.400 ;
        RECT 394.800 174.300 395.600 174.400 ;
        RECT 386.800 173.700 395.600 174.300 ;
        RECT 386.800 173.600 387.600 173.700 ;
        RECT 394.800 173.600 395.600 173.700 ;
        RECT 458.800 174.300 459.600 174.400 ;
        RECT 554.800 174.300 555.600 174.400 ;
        RECT 458.800 173.700 555.600 174.300 ;
        RECT 458.800 173.600 459.600 173.700 ;
        RECT 554.800 173.600 555.600 173.700 ;
        RECT 607.600 174.300 608.400 174.400 ;
        RECT 652.400 174.300 653.200 174.400 ;
        RECT 671.600 174.300 672.400 174.400 ;
        RECT 607.600 173.700 672.400 174.300 ;
        RECT 607.600 173.600 608.400 173.700 ;
        RECT 652.400 173.600 653.200 173.700 ;
        RECT 671.600 173.600 672.400 173.700 ;
        RECT 674.800 174.300 675.600 174.400 ;
        RECT 681.200 174.300 682.000 174.400 ;
        RECT 674.800 173.700 682.000 174.300 ;
        RECT 674.800 173.600 675.600 173.700 ;
        RECT 681.200 173.600 682.000 173.700 ;
        RECT 25.200 172.300 26.000 172.400 ;
        RECT 79.600 172.300 80.400 172.400 ;
        RECT 25.200 171.700 80.400 172.300 ;
        RECT 25.200 171.600 26.000 171.700 ;
        RECT 79.600 171.600 80.400 171.700 ;
        RECT 119.600 172.300 120.400 172.400 ;
        RECT 122.800 172.300 123.600 172.400 ;
        RECT 146.800 172.300 147.600 172.400 ;
        RECT 156.400 172.300 157.200 172.400 ;
        RECT 119.600 171.700 157.200 172.300 ;
        RECT 119.600 171.600 120.400 171.700 ;
        RECT 122.800 171.600 123.600 171.700 ;
        RECT 146.800 171.600 147.600 171.700 ;
        RECT 156.400 171.600 157.200 171.700 ;
        RECT 158.000 172.300 158.800 172.400 ;
        RECT 167.600 172.300 168.400 172.400 ;
        RECT 158.000 171.700 168.400 172.300 ;
        RECT 158.000 171.600 158.800 171.700 ;
        RECT 167.600 171.600 168.400 171.700 ;
        RECT 185.200 172.300 186.000 172.400 ;
        RECT 188.400 172.300 189.200 172.400 ;
        RECT 185.200 171.700 189.200 172.300 ;
        RECT 185.200 171.600 186.000 171.700 ;
        RECT 188.400 171.600 189.200 171.700 ;
        RECT 250.800 172.300 251.600 172.400 ;
        RECT 274.800 172.300 275.600 172.400 ;
        RECT 250.800 171.700 275.600 172.300 ;
        RECT 250.800 171.600 251.600 171.700 ;
        RECT 274.800 171.600 275.600 171.700 ;
        RECT 316.400 172.300 317.200 172.400 ;
        RECT 321.200 172.300 322.000 172.400 ;
        RECT 316.400 171.700 322.000 172.300 ;
        RECT 316.400 171.600 317.200 171.700 ;
        RECT 321.200 171.600 322.000 171.700 ;
        RECT 447.600 172.300 448.400 172.400 ;
        RECT 457.200 172.300 458.000 172.400 ;
        RECT 447.600 171.700 458.000 172.300 ;
        RECT 447.600 171.600 448.400 171.700 ;
        RECT 457.200 171.600 458.000 171.700 ;
        RECT 463.600 172.300 464.400 172.400 ;
        RECT 473.200 172.300 474.000 172.400 ;
        RECT 482.800 172.300 483.600 172.400 ;
        RECT 463.600 171.700 483.600 172.300 ;
        RECT 463.600 171.600 464.400 171.700 ;
        RECT 473.200 171.600 474.000 171.700 ;
        RECT 482.800 171.600 483.600 171.700 ;
        RECT 500.400 172.300 501.200 172.400 ;
        RECT 508.400 172.300 509.200 172.400 ;
        RECT 500.400 171.700 509.200 172.300 ;
        RECT 500.400 171.600 501.200 171.700 ;
        RECT 508.400 171.600 509.200 171.700 ;
        RECT 559.600 172.300 560.400 172.400 ;
        RECT 582.000 172.300 582.800 172.400 ;
        RECT 559.600 171.700 582.800 172.300 ;
        RECT 559.600 171.600 560.400 171.700 ;
        RECT 582.000 171.600 582.800 171.700 ;
        RECT 594.800 172.300 595.600 172.400 ;
        RECT 615.600 172.300 616.400 172.400 ;
        RECT 594.800 171.700 616.400 172.300 ;
        RECT 594.800 171.600 595.600 171.700 ;
        RECT 615.600 171.600 616.400 171.700 ;
        RECT 626.800 172.300 627.600 172.400 ;
        RECT 639.600 172.300 640.400 172.400 ;
        RECT 626.800 171.700 640.400 172.300 ;
        RECT 626.800 171.600 627.600 171.700 ;
        RECT 639.600 171.600 640.400 171.700 ;
        RECT 642.800 172.300 643.600 172.400 ;
        RECT 674.800 172.300 675.600 172.400 ;
        RECT 642.800 171.700 675.600 172.300 ;
        RECT 642.800 171.600 643.600 171.700 ;
        RECT 674.800 171.600 675.600 171.700 ;
        RECT 52.400 170.300 53.200 170.400 ;
        RECT 55.600 170.300 56.400 170.400 ;
        RECT 62.000 170.300 62.800 170.400 ;
        RECT 52.400 169.700 62.800 170.300 ;
        RECT 52.400 169.600 53.200 169.700 ;
        RECT 55.600 169.600 56.400 169.700 ;
        RECT 62.000 169.600 62.800 169.700 ;
        RECT 65.200 170.300 66.000 170.400 ;
        RECT 74.800 170.300 75.600 170.400 ;
        RECT 108.400 170.300 109.200 170.400 ;
        RECT 118.000 170.300 118.800 170.400 ;
        RECT 65.200 169.700 118.800 170.300 ;
        RECT 65.200 169.600 66.000 169.700 ;
        RECT 74.800 169.600 75.600 169.700 ;
        RECT 108.400 169.600 109.200 169.700 ;
        RECT 118.000 169.600 118.800 169.700 ;
        RECT 124.400 170.300 125.200 170.400 ;
        RECT 148.400 170.300 149.200 170.400 ;
        RECT 124.400 169.700 149.200 170.300 ;
        RECT 124.400 169.600 125.200 169.700 ;
        RECT 148.400 169.600 149.200 169.700 ;
        RECT 153.200 170.300 154.000 170.400 ;
        RECT 178.800 170.300 179.600 170.400 ;
        RECT 153.200 169.700 179.600 170.300 ;
        RECT 153.200 169.600 154.000 169.700 ;
        RECT 178.800 169.600 179.600 169.700 ;
        RECT 180.400 170.300 181.200 170.400 ;
        RECT 186.800 170.300 187.600 170.400 ;
        RECT 190.000 170.300 190.800 170.400 ;
        RECT 180.400 169.700 190.800 170.300 ;
        RECT 180.400 169.600 181.200 169.700 ;
        RECT 186.800 169.600 187.600 169.700 ;
        RECT 190.000 169.600 190.800 169.700 ;
        RECT 255.600 170.300 256.400 170.400 ;
        RECT 313.200 170.300 314.000 170.400 ;
        RECT 255.600 169.700 314.000 170.300 ;
        RECT 255.600 169.600 256.400 169.700 ;
        RECT 313.200 169.600 314.000 169.700 ;
        RECT 322.800 170.300 323.600 170.400 ;
        RECT 343.600 170.300 344.400 170.400 ;
        RECT 356.400 170.300 357.200 170.400 ;
        RECT 322.800 169.700 357.200 170.300 ;
        RECT 322.800 169.600 323.600 169.700 ;
        RECT 343.600 169.600 344.400 169.700 ;
        RECT 356.400 169.600 357.200 169.700 ;
        RECT 526.000 170.300 526.800 170.400 ;
        RECT 534.000 170.300 534.800 170.400 ;
        RECT 556.400 170.300 557.200 170.400 ;
        RECT 562.800 170.300 563.600 170.400 ;
        RECT 526.000 169.700 563.600 170.300 ;
        RECT 526.000 169.600 526.800 169.700 ;
        RECT 534.000 169.600 534.800 169.700 ;
        RECT 556.400 169.600 557.200 169.700 ;
        RECT 562.800 169.600 563.600 169.700 ;
        RECT 582.000 170.300 582.800 170.400 ;
        RECT 583.600 170.300 584.400 170.400 ;
        RECT 582.000 169.700 584.400 170.300 ;
        RECT 582.000 169.600 582.800 169.700 ;
        RECT 583.600 169.600 584.400 169.700 ;
        RECT 591.600 170.300 592.400 170.400 ;
        RECT 618.800 170.300 619.600 170.400 ;
        RECT 628.400 170.300 629.200 170.400 ;
        RECT 591.600 169.700 629.200 170.300 ;
        RECT 591.600 169.600 592.400 169.700 ;
        RECT 618.800 169.600 619.600 169.700 ;
        RECT 628.400 169.600 629.200 169.700 ;
        RECT 636.400 170.300 637.200 170.400 ;
        RECT 646.000 170.300 646.800 170.400 ;
        RECT 636.400 169.700 646.800 170.300 ;
        RECT 636.400 169.600 637.200 169.700 ;
        RECT 646.000 169.600 646.800 169.700 ;
        RECT 33.200 168.300 34.000 168.400 ;
        RECT 55.600 168.300 56.400 168.400 ;
        RECT 33.200 167.700 56.400 168.300 ;
        RECT 33.200 167.600 34.000 167.700 ;
        RECT 55.600 167.600 56.400 167.700 ;
        RECT 121.200 168.300 122.000 168.400 ;
        RECT 151.600 168.300 152.400 168.400 ;
        RECT 121.200 167.700 152.400 168.300 ;
        RECT 121.200 167.600 122.000 167.700 ;
        RECT 151.600 167.600 152.400 167.700 ;
        RECT 154.800 168.300 155.600 168.400 ;
        RECT 174.000 168.300 174.800 168.400 ;
        RECT 154.800 167.700 174.800 168.300 ;
        RECT 154.800 167.600 155.600 167.700 ;
        RECT 174.000 167.600 174.800 167.700 ;
        RECT 182.000 168.300 182.800 168.400 ;
        RECT 202.800 168.300 203.600 168.400 ;
        RECT 182.000 167.700 203.600 168.300 ;
        RECT 182.000 167.600 182.800 167.700 ;
        RECT 202.800 167.600 203.600 167.700 ;
        RECT 401.200 168.300 402.000 168.400 ;
        RECT 422.000 168.300 422.800 168.400 ;
        RECT 401.200 167.700 422.800 168.300 ;
        RECT 401.200 167.600 402.000 167.700 ;
        RECT 422.000 167.600 422.800 167.700 ;
        RECT 503.600 168.300 504.400 168.400 ;
        RECT 519.600 168.300 520.400 168.400 ;
        RECT 546.800 168.300 547.600 168.400 ;
        RECT 503.600 167.700 547.600 168.300 ;
        RECT 503.600 167.600 504.400 167.700 ;
        RECT 519.600 167.600 520.400 167.700 ;
        RECT 546.800 167.600 547.600 167.700 ;
        RECT 604.400 168.300 605.200 168.400 ;
        RECT 623.600 168.300 624.400 168.400 ;
        RECT 604.400 167.700 624.400 168.300 ;
        RECT 604.400 167.600 605.200 167.700 ;
        RECT 623.600 167.600 624.400 167.700 ;
        RECT 638.000 168.300 638.800 168.400 ;
        RECT 649.200 168.300 650.000 168.400 ;
        RECT 638.000 167.700 650.000 168.300 ;
        RECT 638.000 167.600 638.800 167.700 ;
        RECT 649.200 167.600 650.000 167.700 ;
        RECT 679.600 168.300 680.400 168.400 ;
        RECT 682.800 168.300 683.600 168.400 ;
        RECT 679.600 167.700 683.600 168.300 ;
        RECT 679.600 167.600 680.400 167.700 ;
        RECT 682.800 167.600 683.600 167.700 ;
        RECT 42.800 166.300 43.600 166.400 ;
        RECT 111.600 166.300 112.400 166.400 ;
        RECT 42.800 165.700 112.400 166.300 ;
        RECT 42.800 165.600 43.600 165.700 ;
        RECT 111.600 165.600 112.400 165.700 ;
        RECT 518.000 166.300 518.800 166.400 ;
        RECT 567.600 166.300 568.400 166.400 ;
        RECT 518.000 165.700 568.400 166.300 ;
        RECT 518.000 165.600 518.800 165.700 ;
        RECT 567.600 165.600 568.400 165.700 ;
        RECT 580.400 166.300 581.200 166.400 ;
        RECT 602.800 166.300 603.600 166.400 ;
        RECT 626.800 166.300 627.600 166.400 ;
        RECT 580.400 165.700 627.600 166.300 ;
        RECT 580.400 165.600 581.200 165.700 ;
        RECT 602.800 165.600 603.600 165.700 ;
        RECT 626.800 165.600 627.600 165.700 ;
        RECT 90.800 163.600 91.600 164.400 ;
        RECT 114.800 164.300 115.600 164.400 ;
        RECT 124.400 164.300 125.200 164.400 ;
        RECT 143.600 164.300 144.400 164.400 ;
        RECT 148.400 164.300 149.200 164.400 ;
        RECT 114.800 163.700 149.200 164.300 ;
        RECT 114.800 163.600 115.600 163.700 ;
        RECT 124.400 163.600 125.200 163.700 ;
        RECT 143.600 163.600 144.400 163.700 ;
        RECT 148.400 163.600 149.200 163.700 ;
        RECT 150.000 164.300 150.800 164.400 ;
        RECT 177.200 164.300 178.000 164.400 ;
        RECT 183.600 164.300 184.400 164.400 ;
        RECT 215.600 164.300 216.400 164.400 ;
        RECT 150.000 163.700 216.400 164.300 ;
        RECT 150.000 163.600 150.800 163.700 ;
        RECT 177.200 163.600 178.000 163.700 ;
        RECT 183.600 163.600 184.400 163.700 ;
        RECT 215.600 163.600 216.400 163.700 ;
        RECT 295.600 164.300 296.400 164.400 ;
        RECT 329.200 164.300 330.000 164.400 ;
        RECT 295.600 163.700 330.000 164.300 ;
        RECT 295.600 163.600 296.400 163.700 ;
        RECT 329.200 163.600 330.000 163.700 ;
        RECT 454.000 164.300 454.800 164.400 ;
        RECT 465.200 164.300 466.000 164.400 ;
        RECT 454.000 163.700 466.000 164.300 ;
        RECT 454.000 163.600 454.800 163.700 ;
        RECT 465.200 163.600 466.000 163.700 ;
        RECT 486.000 164.300 486.800 164.400 ;
        RECT 503.600 164.300 504.400 164.400 ;
        RECT 486.000 163.700 504.400 164.300 ;
        RECT 486.000 163.600 486.800 163.700 ;
        RECT 503.600 163.600 504.400 163.700 ;
        RECT 529.200 164.300 530.000 164.400 ;
        RECT 545.200 164.300 546.000 164.400 ;
        RECT 580.400 164.300 581.200 164.400 ;
        RECT 529.200 163.700 581.200 164.300 ;
        RECT 529.200 163.600 530.000 163.700 ;
        RECT 545.200 163.600 546.000 163.700 ;
        RECT 580.400 163.600 581.200 163.700 ;
        RECT 582.000 164.300 582.800 164.400 ;
        RECT 594.800 164.300 595.600 164.400 ;
        RECT 582.000 163.700 595.600 164.300 ;
        RECT 582.000 163.600 582.800 163.700 ;
        RECT 594.800 163.600 595.600 163.700 ;
        RECT 606.000 164.300 606.800 164.400 ;
        RECT 609.200 164.300 610.000 164.400 ;
        RECT 606.000 163.700 610.000 164.300 ;
        RECT 606.000 163.600 606.800 163.700 ;
        RECT 609.200 163.600 610.000 163.700 ;
        RECT 670.000 164.300 670.800 164.400 ;
        RECT 676.400 164.300 677.200 164.400 ;
        RECT 670.000 163.700 677.200 164.300 ;
        RECT 670.000 163.600 670.800 163.700 ;
        RECT 676.400 163.600 677.200 163.700 ;
        RECT 9.200 162.300 10.000 162.400 ;
        RECT 14.000 162.300 14.800 162.400 ;
        RECT 9.200 161.700 14.800 162.300 ;
        RECT 9.200 161.600 10.000 161.700 ;
        RECT 14.000 161.600 14.800 161.700 ;
        RECT 41.200 162.300 42.000 162.400 ;
        RECT 54.000 162.300 54.800 162.400 ;
        RECT 87.600 162.300 88.400 162.400 ;
        RECT 41.200 161.700 88.400 162.300 ;
        RECT 41.200 161.600 42.000 161.700 ;
        RECT 54.000 161.600 54.800 161.700 ;
        RECT 87.600 161.600 88.400 161.700 ;
        RECT 233.200 162.300 234.000 162.400 ;
        RECT 238.000 162.300 238.800 162.400 ;
        RECT 233.200 161.700 238.800 162.300 ;
        RECT 233.200 161.600 234.000 161.700 ;
        RECT 238.000 161.600 238.800 161.700 ;
        RECT 497.200 162.300 498.000 162.400 ;
        RECT 506.800 162.300 507.600 162.400 ;
        RECT 497.200 161.700 507.600 162.300 ;
        RECT 497.200 161.600 498.000 161.700 ;
        RECT 506.800 161.600 507.600 161.700 ;
        RECT 540.400 162.300 541.200 162.400 ;
        RECT 546.800 162.300 547.600 162.400 ;
        RECT 540.400 161.700 547.600 162.300 ;
        RECT 540.400 161.600 541.200 161.700 ;
        RECT 546.800 161.600 547.600 161.700 ;
        RECT 577.200 162.300 578.000 162.400 ;
        RECT 585.200 162.300 586.000 162.400 ;
        RECT 577.200 161.700 586.000 162.300 ;
        RECT 577.200 161.600 578.000 161.700 ;
        RECT 585.200 161.600 586.000 161.700 ;
        RECT 681.200 162.300 682.000 162.400 ;
        RECT 684.400 162.300 685.200 162.400 ;
        RECT 681.200 161.700 685.200 162.300 ;
        RECT 681.200 161.600 682.000 161.700 ;
        RECT 684.400 161.600 685.200 161.700 ;
        RECT 142.000 160.300 142.800 160.400 ;
        RECT 154.800 160.300 155.600 160.400 ;
        RECT 142.000 159.700 155.600 160.300 ;
        RECT 142.000 159.600 142.800 159.700 ;
        RECT 154.800 159.600 155.600 159.700 ;
        RECT 161.200 160.300 162.000 160.400 ;
        RECT 166.000 160.300 166.800 160.400 ;
        RECT 161.200 159.700 166.800 160.300 ;
        RECT 161.200 159.600 162.000 159.700 ;
        RECT 166.000 159.600 166.800 159.700 ;
        RECT 457.200 160.300 458.000 160.400 ;
        RECT 458.800 160.300 459.600 160.400 ;
        RECT 457.200 159.700 459.600 160.300 ;
        RECT 457.200 159.600 458.000 159.700 ;
        RECT 458.800 159.600 459.600 159.700 ;
        RECT 494.000 160.300 494.800 160.400 ;
        RECT 508.400 160.300 509.200 160.400 ;
        RECT 534.000 160.300 534.800 160.400 ;
        RECT 543.600 160.300 544.400 160.400 ;
        RECT 494.000 159.700 544.400 160.300 ;
        RECT 494.000 159.600 494.800 159.700 ;
        RECT 508.400 159.600 509.200 159.700 ;
        RECT 534.000 159.600 534.800 159.700 ;
        RECT 543.600 159.600 544.400 159.700 ;
        RECT 561.200 160.300 562.000 160.400 ;
        RECT 588.400 160.300 589.200 160.400 ;
        RECT 561.200 159.700 589.200 160.300 ;
        RECT 561.200 159.600 562.000 159.700 ;
        RECT 588.400 159.600 589.200 159.700 ;
        RECT 593.200 159.600 594.000 160.400 ;
        RECT 626.800 160.300 627.600 160.400 ;
        RECT 655.600 160.300 656.400 160.400 ;
        RECT 626.800 159.700 656.400 160.300 ;
        RECT 626.800 159.600 627.600 159.700 ;
        RECT 655.600 159.600 656.400 159.700 ;
        RECT 28.400 158.300 29.200 158.400 ;
        RECT 36.400 158.300 37.200 158.400 ;
        RECT 122.800 158.300 123.600 158.400 ;
        RECT 28.400 157.700 123.600 158.300 ;
        RECT 28.400 157.600 29.200 157.700 ;
        RECT 36.400 157.600 37.200 157.700 ;
        RECT 122.800 157.600 123.600 157.700 ;
        RECT 132.400 158.300 133.200 158.400 ;
        RECT 138.800 158.300 139.600 158.400 ;
        RECT 132.400 157.700 139.600 158.300 ;
        RECT 132.400 157.600 133.200 157.700 ;
        RECT 138.800 157.600 139.600 157.700 ;
        RECT 399.600 158.300 400.400 158.400 ;
        RECT 428.400 158.300 429.200 158.400 ;
        RECT 399.600 157.700 429.200 158.300 ;
        RECT 399.600 157.600 400.400 157.700 ;
        RECT 428.400 157.600 429.200 157.700 ;
        RECT 511.600 158.300 512.400 158.400 ;
        RECT 599.600 158.300 600.400 158.400 ;
        RECT 633.200 158.300 634.000 158.400 ;
        RECT 649.200 158.300 650.000 158.400 ;
        RECT 511.600 157.700 650.000 158.300 ;
        RECT 511.600 157.600 512.400 157.700 ;
        RECT 599.600 157.600 600.400 157.700 ;
        RECT 633.200 157.600 634.000 157.700 ;
        RECT 649.200 157.600 650.000 157.700 ;
        RECT 44.400 156.300 45.200 156.400 ;
        RECT 73.200 156.300 74.000 156.400 ;
        RECT 44.400 155.700 74.000 156.300 ;
        RECT 44.400 155.600 45.200 155.700 ;
        RECT 73.200 155.600 74.000 155.700 ;
        RECT 79.600 156.300 80.400 156.400 ;
        RECT 134.000 156.300 134.800 156.400 ;
        RECT 162.800 156.300 163.600 156.400 ;
        RECT 170.800 156.300 171.600 156.400 ;
        RECT 79.600 155.700 171.600 156.300 ;
        RECT 79.600 155.600 80.400 155.700 ;
        RECT 134.000 155.600 134.800 155.700 ;
        RECT 162.800 155.600 163.600 155.700 ;
        RECT 170.800 155.600 171.600 155.700 ;
        RECT 193.200 156.300 194.000 156.400 ;
        RECT 196.400 156.300 197.200 156.400 ;
        RECT 193.200 155.700 197.200 156.300 ;
        RECT 193.200 155.600 194.000 155.700 ;
        RECT 196.400 155.600 197.200 155.700 ;
        RECT 473.200 156.300 474.000 156.400 ;
        RECT 484.400 156.300 485.200 156.400 ;
        RECT 473.200 155.700 485.200 156.300 ;
        RECT 473.200 155.600 474.000 155.700 ;
        RECT 484.400 155.600 485.200 155.700 ;
        RECT 537.200 156.300 538.000 156.400 ;
        RECT 550.000 156.300 550.800 156.400 ;
        RECT 537.200 155.700 550.800 156.300 ;
        RECT 537.200 155.600 538.000 155.700 ;
        RECT 550.000 155.600 550.800 155.700 ;
        RECT 558.000 156.300 558.800 156.400 ;
        RECT 574.000 156.300 574.800 156.400 ;
        RECT 558.000 155.700 574.800 156.300 ;
        RECT 558.000 155.600 558.800 155.700 ;
        RECT 574.000 155.600 574.800 155.700 ;
        RECT 578.800 156.300 579.600 156.400 ;
        RECT 641.200 156.300 642.000 156.400 ;
        RECT 578.800 155.700 642.000 156.300 ;
        RECT 578.800 155.600 579.600 155.700 ;
        RECT 641.200 155.600 642.000 155.700 ;
        RECT 647.600 156.300 648.400 156.400 ;
        RECT 668.400 156.300 669.200 156.400 ;
        RECT 647.600 155.700 669.200 156.300 ;
        RECT 647.600 155.600 648.400 155.700 ;
        RECT 668.400 155.600 669.200 155.700 ;
        RECT 94.000 154.300 94.800 154.400 ;
        RECT 68.500 153.700 94.800 154.300 ;
        RECT 68.500 152.400 69.100 153.700 ;
        RECT 94.000 153.600 94.800 153.700 ;
        RECT 127.600 154.300 128.400 154.400 ;
        RECT 159.600 154.300 160.400 154.400 ;
        RECT 194.800 154.300 195.600 154.400 ;
        RECT 206.000 154.300 206.800 154.400 ;
        RECT 127.600 153.700 206.800 154.300 ;
        RECT 127.600 153.600 128.400 153.700 ;
        RECT 159.600 153.600 160.400 153.700 ;
        RECT 194.800 153.600 195.600 153.700 ;
        RECT 206.000 153.600 206.800 153.700 ;
        RECT 209.200 154.300 210.000 154.400 ;
        RECT 217.200 154.300 218.000 154.400 ;
        RECT 209.200 153.700 218.000 154.300 ;
        RECT 209.200 153.600 210.000 153.700 ;
        RECT 217.200 153.600 218.000 153.700 ;
        RECT 311.600 154.300 312.400 154.400 ;
        RECT 345.200 154.300 346.000 154.400 ;
        RECT 356.400 154.300 357.200 154.400 ;
        RECT 311.600 153.700 357.200 154.300 ;
        RECT 311.600 153.600 312.400 153.700 ;
        RECT 345.200 153.600 346.000 153.700 ;
        RECT 356.400 153.600 357.200 153.700 ;
        RECT 436.400 154.300 437.200 154.400 ;
        RECT 545.200 154.300 546.000 154.400 ;
        RECT 436.400 153.700 546.000 154.300 ;
        RECT 436.400 153.600 437.200 153.700 ;
        RECT 545.200 153.600 546.000 153.700 ;
        RECT 585.200 154.300 586.000 154.400 ;
        RECT 594.800 154.300 595.600 154.400 ;
        RECT 585.200 153.700 595.600 154.300 ;
        RECT 585.200 153.600 586.000 153.700 ;
        RECT 594.800 153.600 595.600 153.700 ;
        RECT 614.000 154.300 614.800 154.400 ;
        RECT 622.000 154.300 622.800 154.400 ;
        RECT 614.000 153.700 622.800 154.300 ;
        RECT 614.000 153.600 614.800 153.700 ;
        RECT 622.000 153.600 622.800 153.700 ;
        RECT 646.000 154.300 646.800 154.400 ;
        RECT 654.000 154.300 654.800 154.400 ;
        RECT 646.000 153.700 654.800 154.300 ;
        RECT 646.000 153.600 646.800 153.700 ;
        RECT 654.000 153.600 654.800 153.700 ;
        RECT 655.600 154.300 656.400 154.400 ;
        RECT 670.000 154.300 670.800 154.400 ;
        RECT 682.800 154.300 683.600 154.400 ;
        RECT 655.600 153.700 683.600 154.300 ;
        RECT 655.600 153.600 656.400 153.700 ;
        RECT 670.000 153.600 670.800 153.700 ;
        RECT 682.800 153.600 683.600 153.700 ;
        RECT 2.800 152.300 3.600 152.400 ;
        RECT 10.800 152.300 11.600 152.400 ;
        RECT 33.200 152.300 34.000 152.400 ;
        RECT 2.800 151.700 34.000 152.300 ;
        RECT 2.800 151.600 3.600 151.700 ;
        RECT 10.800 151.600 11.600 151.700 ;
        RECT 33.200 151.600 34.000 151.700 ;
        RECT 34.800 152.300 35.600 152.400 ;
        RECT 41.200 152.300 42.000 152.400 ;
        RECT 34.800 151.700 42.000 152.300 ;
        RECT 34.800 151.600 35.600 151.700 ;
        RECT 41.200 151.600 42.000 151.700 ;
        RECT 49.200 152.300 50.000 152.400 ;
        RECT 52.400 152.300 53.200 152.400 ;
        RECT 49.200 151.700 53.200 152.300 ;
        RECT 49.200 151.600 50.000 151.700 ;
        RECT 52.400 151.600 53.200 151.700 ;
        RECT 58.800 152.300 59.600 152.400 ;
        RECT 68.400 152.300 69.200 152.400 ;
        RECT 58.800 151.700 69.200 152.300 ;
        RECT 58.800 151.600 59.600 151.700 ;
        RECT 68.400 151.600 69.200 151.700 ;
        RECT 86.000 152.300 86.800 152.400 ;
        RECT 103.600 152.300 104.400 152.400 ;
        RECT 119.600 152.300 120.400 152.400 ;
        RECT 201.200 152.300 202.000 152.400 ;
        RECT 86.000 151.700 120.400 152.300 ;
        RECT 86.000 151.600 86.800 151.700 ;
        RECT 103.600 151.600 104.400 151.700 ;
        RECT 119.600 151.600 120.400 151.700 ;
        RECT 191.700 151.700 202.000 152.300 ;
        RECT 191.700 150.400 192.300 151.700 ;
        RECT 201.200 151.600 202.000 151.700 ;
        RECT 215.600 152.300 216.400 152.400 ;
        RECT 246.000 152.300 246.800 152.400 ;
        RECT 215.600 151.700 246.800 152.300 ;
        RECT 215.600 151.600 216.400 151.700 ;
        RECT 246.000 151.600 246.800 151.700 ;
        RECT 306.800 152.300 307.600 152.400 ;
        RECT 319.600 152.300 320.400 152.400 ;
        RECT 306.800 151.700 320.400 152.300 ;
        RECT 306.800 151.600 307.600 151.700 ;
        RECT 319.600 151.600 320.400 151.700 ;
        RECT 345.200 152.300 346.000 152.400 ;
        RECT 351.600 152.300 352.400 152.400 ;
        RECT 345.200 151.700 352.400 152.300 ;
        RECT 345.200 151.600 346.000 151.700 ;
        RECT 351.600 151.600 352.400 151.700 ;
        RECT 521.200 152.300 522.000 152.400 ;
        RECT 530.800 152.300 531.600 152.400 ;
        RECT 521.200 151.700 531.600 152.300 ;
        RECT 521.200 151.600 522.000 151.700 ;
        RECT 530.800 151.600 531.600 151.700 ;
        RECT 537.200 152.300 538.000 152.400 ;
        RECT 542.000 152.300 542.800 152.400 ;
        RECT 537.200 151.700 542.800 152.300 ;
        RECT 537.200 151.600 538.000 151.700 ;
        RECT 542.000 151.600 542.800 151.700 ;
        RECT 564.400 152.300 565.200 152.400 ;
        RECT 574.000 152.300 574.800 152.400 ;
        RECT 564.400 151.700 574.800 152.300 ;
        RECT 564.400 151.600 565.200 151.700 ;
        RECT 574.000 151.600 574.800 151.700 ;
        RECT 580.400 152.300 581.200 152.400 ;
        RECT 593.200 152.300 594.000 152.400 ;
        RECT 630.000 152.300 630.800 152.400 ;
        RECT 646.100 152.300 646.700 153.600 ;
        RECT 580.400 151.700 589.100 152.300 ;
        RECT 580.400 151.600 581.200 151.700 ;
        RECT 14.000 150.300 14.800 150.400 ;
        RECT 52.400 150.300 53.200 150.400 ;
        RECT 14.000 149.700 53.200 150.300 ;
        RECT 14.000 149.600 14.800 149.700 ;
        RECT 52.400 149.600 53.200 149.700 ;
        RECT 55.600 150.300 56.400 150.400 ;
        RECT 63.600 150.300 64.400 150.400 ;
        RECT 55.600 149.700 64.400 150.300 ;
        RECT 55.600 149.600 56.400 149.700 ;
        RECT 63.600 149.600 64.400 149.700 ;
        RECT 66.800 150.300 67.600 150.400 ;
        RECT 105.200 150.300 106.000 150.400 ;
        RECT 66.800 149.700 106.000 150.300 ;
        RECT 66.800 149.600 67.600 149.700 ;
        RECT 105.200 149.600 106.000 149.700 ;
        RECT 146.800 150.300 147.600 150.400 ;
        RECT 151.600 150.300 152.400 150.400 ;
        RECT 146.800 149.700 152.400 150.300 ;
        RECT 146.800 149.600 147.600 149.700 ;
        RECT 151.600 149.600 152.400 149.700 ;
        RECT 154.800 150.300 155.600 150.400 ;
        RECT 167.600 150.300 168.400 150.400 ;
        RECT 154.800 149.700 168.400 150.300 ;
        RECT 154.800 149.600 155.600 149.700 ;
        RECT 167.600 149.600 168.400 149.700 ;
        RECT 174.000 150.300 174.800 150.400 ;
        RECT 191.600 150.300 192.400 150.400 ;
        RECT 174.000 149.700 192.400 150.300 ;
        RECT 174.000 149.600 174.800 149.700 ;
        RECT 191.600 149.600 192.400 149.700 ;
        RECT 196.400 150.300 197.200 150.400 ;
        RECT 209.200 150.300 210.000 150.400 ;
        RECT 196.400 149.700 210.000 150.300 ;
        RECT 196.400 149.600 197.200 149.700 ;
        RECT 209.200 149.600 210.000 149.700 ;
        RECT 212.400 150.300 213.200 150.400 ;
        RECT 228.400 150.300 229.200 150.400 ;
        RECT 212.400 149.700 229.200 150.300 ;
        RECT 212.400 149.600 213.200 149.700 ;
        RECT 228.400 149.600 229.200 149.700 ;
        RECT 238.000 150.300 238.800 150.400 ;
        RECT 247.600 150.300 248.400 150.400 ;
        RECT 260.400 150.300 261.200 150.400 ;
        RECT 238.000 149.700 261.200 150.300 ;
        RECT 238.000 149.600 238.800 149.700 ;
        RECT 247.600 149.600 248.400 149.700 ;
        RECT 260.400 149.600 261.200 149.700 ;
        RECT 380.400 150.300 381.200 150.400 ;
        RECT 386.800 150.300 387.600 150.400 ;
        RECT 380.400 149.700 387.600 150.300 ;
        RECT 380.400 149.600 381.200 149.700 ;
        RECT 386.800 149.600 387.600 149.700 ;
        RECT 407.600 150.300 408.400 150.400 ;
        RECT 441.200 150.300 442.000 150.400 ;
        RECT 407.600 149.700 442.000 150.300 ;
        RECT 407.600 149.600 408.400 149.700 ;
        RECT 441.200 149.600 442.000 149.700 ;
        RECT 462.000 150.300 462.800 150.400 ;
        RECT 479.600 150.300 480.400 150.400 ;
        RECT 462.000 149.700 480.400 150.300 ;
        RECT 462.000 149.600 462.800 149.700 ;
        RECT 479.600 149.600 480.400 149.700 ;
        RECT 514.800 150.300 515.600 150.400 ;
        RECT 518.000 150.300 518.800 150.400 ;
        RECT 514.800 149.700 518.800 150.300 ;
        RECT 514.800 149.600 515.600 149.700 ;
        RECT 518.000 149.600 518.800 149.700 ;
        RECT 519.600 150.300 520.400 150.400 ;
        RECT 538.800 150.300 539.600 150.400 ;
        RECT 542.000 150.300 542.800 150.400 ;
        RECT 519.600 149.700 542.800 150.300 ;
        RECT 519.600 149.600 520.400 149.700 ;
        RECT 538.800 149.600 539.600 149.700 ;
        RECT 542.000 149.600 542.800 149.700 ;
        RECT 545.200 150.300 546.000 150.400 ;
        RECT 562.800 150.300 563.600 150.400 ;
        RECT 545.200 149.700 563.600 150.300 ;
        RECT 545.200 149.600 546.000 149.700 ;
        RECT 562.800 149.600 563.600 149.700 ;
        RECT 567.600 150.300 568.400 150.400 ;
        RECT 582.000 150.300 582.800 150.400 ;
        RECT 567.600 149.700 582.800 150.300 ;
        RECT 567.600 149.600 568.400 149.700 ;
        RECT 582.000 149.600 582.800 149.700 ;
        RECT 583.600 150.300 584.400 150.400 ;
        RECT 585.200 150.300 586.000 150.400 ;
        RECT 583.600 149.700 586.000 150.300 ;
        RECT 588.500 150.300 589.100 151.700 ;
        RECT 593.200 151.700 646.700 152.300 ;
        RECT 593.200 151.600 594.000 151.700 ;
        RECT 630.000 151.600 630.800 151.700 ;
        RECT 663.600 151.600 664.400 152.400 ;
        RECT 671.600 152.300 672.400 152.400 ;
        RECT 678.000 152.300 678.800 152.400 ;
        RECT 671.600 151.700 678.800 152.300 ;
        RECT 671.600 151.600 672.400 151.700 ;
        RECT 678.000 151.600 678.800 151.700 ;
        RECT 620.400 150.300 621.200 150.400 ;
        RECT 622.000 150.300 622.800 150.400 ;
        RECT 628.400 150.300 629.200 150.400 ;
        RECT 588.500 149.700 629.200 150.300 ;
        RECT 583.600 149.600 584.400 149.700 ;
        RECT 585.200 149.600 586.000 149.700 ;
        RECT 620.400 149.600 621.200 149.700 ;
        RECT 622.000 149.600 622.800 149.700 ;
        RECT 628.400 149.600 629.200 149.700 ;
        RECT 650.800 150.300 651.600 150.400 ;
        RECT 660.400 150.300 661.200 150.400 ;
        RECT 650.800 149.700 661.200 150.300 ;
        RECT 650.800 149.600 651.600 149.700 ;
        RECT 660.400 149.600 661.200 149.700 ;
        RECT 668.400 150.300 669.200 150.400 ;
        RECT 679.600 150.300 680.400 150.400 ;
        RECT 668.400 149.700 680.400 150.300 ;
        RECT 668.400 149.600 669.200 149.700 ;
        RECT 679.600 149.600 680.400 149.700 ;
        RECT 17.200 148.300 18.000 148.400 ;
        RECT 18.800 148.300 19.600 148.400 ;
        RECT 23.600 148.300 24.400 148.400 ;
        RECT 30.000 148.300 30.800 148.400 ;
        RECT 17.200 147.700 30.800 148.300 ;
        RECT 17.200 147.600 18.000 147.700 ;
        RECT 18.800 147.600 19.600 147.700 ;
        RECT 23.600 147.600 24.400 147.700 ;
        RECT 30.000 147.600 30.800 147.700 ;
        RECT 31.600 148.300 32.400 148.400 ;
        RECT 34.800 148.300 35.600 148.400 ;
        RECT 31.600 147.700 35.600 148.300 ;
        RECT 31.600 147.600 32.400 147.700 ;
        RECT 34.800 147.600 35.600 147.700 ;
        RECT 39.600 148.300 40.400 148.400 ;
        RECT 42.800 148.300 43.600 148.400 ;
        RECT 39.600 147.700 43.600 148.300 ;
        RECT 39.600 147.600 40.400 147.700 ;
        RECT 42.800 147.600 43.600 147.700 ;
        RECT 90.800 148.300 91.600 148.400 ;
        RECT 121.200 148.300 122.000 148.400 ;
        RECT 90.800 147.700 122.000 148.300 ;
        RECT 90.800 147.600 91.600 147.700 ;
        RECT 121.200 147.600 122.000 147.700 ;
        RECT 138.800 148.300 139.600 148.400 ;
        RECT 150.000 148.300 150.800 148.400 ;
        RECT 138.800 147.700 150.800 148.300 ;
        RECT 138.800 147.600 139.600 147.700 ;
        RECT 150.000 147.600 150.800 147.700 ;
        RECT 158.000 148.300 158.800 148.400 ;
        RECT 185.200 148.300 186.000 148.400 ;
        RECT 158.000 147.700 186.000 148.300 ;
        RECT 158.000 147.600 158.800 147.700 ;
        RECT 185.200 147.600 186.000 147.700 ;
        RECT 202.800 148.300 203.600 148.400 ;
        RECT 214.000 148.300 214.800 148.400 ;
        RECT 202.800 147.700 214.800 148.300 ;
        RECT 202.800 147.600 203.600 147.700 ;
        RECT 214.000 147.600 214.800 147.700 ;
        RECT 242.800 148.300 243.600 148.400 ;
        RECT 249.200 148.300 250.000 148.400 ;
        RECT 242.800 147.700 250.000 148.300 ;
        RECT 242.800 147.600 243.600 147.700 ;
        RECT 249.200 147.600 250.000 147.700 ;
        RECT 303.600 148.300 304.400 148.400 ;
        RECT 305.200 148.300 306.000 148.400 ;
        RECT 303.600 147.700 306.000 148.300 ;
        RECT 303.600 147.600 304.400 147.700 ;
        RECT 305.200 147.600 306.000 147.700 ;
        RECT 450.800 148.300 451.600 148.400 ;
        RECT 466.800 148.300 467.600 148.400 ;
        RECT 450.800 147.700 467.600 148.300 ;
        RECT 450.800 147.600 451.600 147.700 ;
        RECT 466.800 147.600 467.600 147.700 ;
        RECT 508.400 148.300 509.200 148.400 ;
        RECT 527.600 148.300 528.400 148.400 ;
        RECT 556.400 148.300 557.200 148.400 ;
        RECT 508.400 147.700 557.200 148.300 ;
        RECT 508.400 147.600 509.200 147.700 ;
        RECT 527.600 147.600 528.400 147.700 ;
        RECT 556.400 147.600 557.200 147.700 ;
        RECT 569.200 148.300 570.000 148.400 ;
        RECT 580.400 148.300 581.200 148.400 ;
        RECT 569.200 147.700 581.200 148.300 ;
        RECT 569.200 147.600 570.000 147.700 ;
        RECT 580.400 147.600 581.200 147.700 ;
        RECT 591.600 148.300 592.400 148.400 ;
        RECT 606.000 148.300 606.800 148.400 ;
        RECT 591.600 147.700 606.800 148.300 ;
        RECT 591.600 147.600 592.400 147.700 ;
        RECT 606.000 147.600 606.800 147.700 ;
        RECT 31.600 146.300 32.400 146.400 ;
        RECT 41.200 146.300 42.000 146.400 ;
        RECT 62.000 146.300 62.800 146.400 ;
        RECT 31.600 145.700 62.800 146.300 ;
        RECT 31.600 145.600 32.400 145.700 ;
        RECT 41.200 145.600 42.000 145.700 ;
        RECT 62.000 145.600 62.800 145.700 ;
        RECT 74.800 146.300 75.600 146.400 ;
        RECT 92.400 146.300 93.200 146.400 ;
        RECT 74.800 145.700 93.200 146.300 ;
        RECT 74.800 145.600 75.600 145.700 ;
        RECT 92.400 145.600 93.200 145.700 ;
        RECT 100.400 146.300 101.200 146.400 ;
        RECT 118.000 146.300 118.800 146.400 ;
        RECT 129.200 146.300 130.000 146.400 ;
        RECT 100.400 145.700 130.000 146.300 ;
        RECT 100.400 145.600 101.200 145.700 ;
        RECT 118.000 145.600 118.800 145.700 ;
        RECT 129.200 145.600 130.000 145.700 ;
        RECT 148.400 146.300 149.200 146.400 ;
        RECT 156.400 146.300 157.200 146.400 ;
        RECT 182.000 146.300 182.800 146.400 ;
        RECT 148.400 145.700 182.800 146.300 ;
        RECT 148.400 145.600 149.200 145.700 ;
        RECT 156.400 145.600 157.200 145.700 ;
        RECT 182.000 145.600 182.800 145.700 ;
        RECT 218.800 146.300 219.600 146.400 ;
        RECT 233.200 146.300 234.000 146.400 ;
        RECT 273.200 146.300 274.000 146.400 ;
        RECT 287.600 146.300 288.400 146.400 ;
        RECT 218.800 145.700 288.400 146.300 ;
        RECT 218.800 145.600 219.600 145.700 ;
        RECT 233.200 145.600 234.000 145.700 ;
        RECT 273.200 145.600 274.000 145.700 ;
        RECT 287.600 145.600 288.400 145.700 ;
        RECT 303.600 146.300 304.400 146.400 ;
        RECT 326.000 146.300 326.800 146.400 ;
        RECT 303.600 145.700 326.800 146.300 ;
        RECT 303.600 145.600 304.400 145.700 ;
        RECT 326.000 145.600 326.800 145.700 ;
        RECT 329.200 146.300 330.000 146.400 ;
        RECT 340.400 146.300 341.200 146.400 ;
        RECT 329.200 145.700 341.200 146.300 ;
        RECT 329.200 145.600 330.000 145.700 ;
        RECT 340.400 145.600 341.200 145.700 ;
        RECT 415.600 146.300 416.400 146.400 ;
        RECT 425.200 146.300 426.000 146.400 ;
        RECT 415.600 145.700 426.000 146.300 ;
        RECT 415.600 145.600 416.400 145.700 ;
        RECT 425.200 145.600 426.000 145.700 ;
        RECT 470.000 146.300 470.800 146.400 ;
        RECT 474.800 146.300 475.600 146.400 ;
        RECT 510.000 146.300 510.800 146.400 ;
        RECT 470.000 145.700 510.800 146.300 ;
        RECT 470.000 145.600 470.800 145.700 ;
        RECT 474.800 145.600 475.600 145.700 ;
        RECT 510.000 145.600 510.800 145.700 ;
        RECT 532.400 146.300 533.200 146.400 ;
        RECT 548.400 146.300 549.200 146.400 ;
        RECT 532.400 145.700 549.200 146.300 ;
        RECT 532.400 145.600 533.200 145.700 ;
        RECT 548.400 145.600 549.200 145.700 ;
        RECT 554.800 146.300 555.600 146.400 ;
        RECT 569.300 146.300 569.900 147.600 ;
        RECT 554.800 145.700 569.900 146.300 ;
        RECT 591.600 146.300 592.400 146.400 ;
        RECT 593.200 146.300 594.000 146.400 ;
        RECT 591.600 145.700 594.000 146.300 ;
        RECT 554.800 145.600 555.600 145.700 ;
        RECT 591.600 145.600 592.400 145.700 ;
        RECT 593.200 145.600 594.000 145.700 ;
        RECT 596.400 146.300 597.200 146.400 ;
        RECT 625.200 146.300 626.000 146.400 ;
        RECT 596.400 145.700 626.000 146.300 ;
        RECT 596.400 145.600 597.200 145.700 ;
        RECT 625.200 145.600 626.000 145.700 ;
        RECT 642.800 146.300 643.600 146.400 ;
        RECT 646.000 146.300 646.800 146.400 ;
        RECT 657.200 146.300 658.000 146.400 ;
        RECT 670.000 146.300 670.800 146.400 ;
        RECT 642.800 145.700 670.800 146.300 ;
        RECT 642.800 145.600 643.600 145.700 ;
        RECT 646.000 145.600 646.800 145.700 ;
        RECT 657.200 145.600 658.000 145.700 ;
        RECT 670.000 145.600 670.800 145.700 ;
        RECT 54.000 144.300 54.800 144.400 ;
        RECT 71.600 144.300 72.400 144.400 ;
        RECT 82.800 144.300 83.600 144.400 ;
        RECT 54.000 143.700 83.600 144.300 ;
        RECT 54.000 143.600 54.800 143.700 ;
        RECT 71.600 143.600 72.400 143.700 ;
        RECT 82.800 143.600 83.600 143.700 ;
        RECT 151.600 144.300 152.400 144.400 ;
        RECT 159.600 144.300 160.400 144.400 ;
        RECT 151.600 143.700 160.400 144.300 ;
        RECT 151.600 143.600 152.400 143.700 ;
        RECT 159.600 143.600 160.400 143.700 ;
        RECT 162.800 144.300 163.600 144.400 ;
        RECT 174.000 144.300 174.800 144.400 ;
        RECT 162.800 143.700 174.800 144.300 ;
        RECT 162.800 143.600 163.600 143.700 ;
        RECT 174.000 143.600 174.800 143.700 ;
        RECT 220.400 144.300 221.200 144.400 ;
        RECT 241.200 144.300 242.000 144.400 ;
        RECT 252.400 144.300 253.200 144.400 ;
        RECT 265.200 144.300 266.000 144.400 ;
        RECT 220.400 143.700 253.200 144.300 ;
        RECT 220.400 143.600 221.200 143.700 ;
        RECT 241.200 143.600 242.000 143.700 ;
        RECT 252.400 143.600 253.200 143.700 ;
        RECT 257.300 143.700 266.000 144.300 ;
        RECT 52.400 142.300 53.200 142.400 ;
        RECT 73.200 142.300 74.000 142.400 ;
        RECT 81.200 142.300 82.000 142.400 ;
        RECT 86.000 142.300 86.800 142.400 ;
        RECT 105.200 142.300 106.000 142.400 ;
        RECT 127.600 142.300 128.400 142.400 ;
        RECT 52.400 141.700 128.400 142.300 ;
        RECT 52.400 141.600 53.200 141.700 ;
        RECT 73.200 141.600 74.000 141.700 ;
        RECT 81.200 141.600 82.000 141.700 ;
        RECT 86.000 141.600 86.800 141.700 ;
        RECT 105.200 141.600 106.000 141.700 ;
        RECT 127.600 141.600 128.400 141.700 ;
        RECT 153.200 142.300 154.000 142.400 ;
        RECT 161.200 142.300 162.000 142.400 ;
        RECT 167.600 142.300 168.400 142.400 ;
        RECT 153.200 141.700 168.400 142.300 ;
        RECT 153.200 141.600 154.000 141.700 ;
        RECT 161.200 141.600 162.000 141.700 ;
        RECT 167.600 141.600 168.400 141.700 ;
        RECT 177.200 142.300 178.000 142.400 ;
        RECT 194.800 142.300 195.600 142.400 ;
        RECT 177.200 141.700 195.600 142.300 ;
        RECT 177.200 141.600 178.000 141.700 ;
        RECT 194.800 141.600 195.600 141.700 ;
        RECT 239.600 142.300 240.400 142.400 ;
        RECT 257.300 142.300 257.900 143.700 ;
        RECT 265.200 143.600 266.000 143.700 ;
        RECT 567.600 144.300 568.400 144.400 ;
        RECT 590.000 144.300 590.800 144.400 ;
        RECT 596.400 144.300 597.200 144.400 ;
        RECT 567.600 143.700 579.500 144.300 ;
        RECT 567.600 143.600 568.400 143.700 ;
        RECT 239.600 141.700 257.900 142.300 ;
        RECT 239.600 141.600 240.400 141.700 ;
        RECT 279.600 141.600 280.400 142.400 ;
        RECT 289.200 142.300 290.000 142.400 ;
        RECT 305.200 142.300 306.000 142.400 ;
        RECT 289.200 141.700 306.000 142.300 ;
        RECT 289.200 141.600 290.000 141.700 ;
        RECT 305.200 141.600 306.000 141.700 ;
        RECT 367.600 142.300 368.400 142.400 ;
        RECT 375.600 142.300 376.400 142.400 ;
        RECT 399.600 142.300 400.400 142.400 ;
        RECT 410.800 142.300 411.600 142.400 ;
        RECT 433.200 142.300 434.000 142.400 ;
        RECT 367.600 141.700 434.000 142.300 ;
        RECT 367.600 141.600 368.400 141.700 ;
        RECT 375.600 141.600 376.400 141.700 ;
        RECT 399.600 141.600 400.400 141.700 ;
        RECT 410.800 141.600 411.600 141.700 ;
        RECT 433.200 141.600 434.000 141.700 ;
        RECT 454.000 142.300 454.800 142.400 ;
        RECT 457.200 142.300 458.000 142.400 ;
        RECT 492.400 142.300 493.200 142.400 ;
        RECT 454.000 141.700 493.200 142.300 ;
        RECT 578.900 142.300 579.500 143.700 ;
        RECT 590.000 143.700 597.200 144.300 ;
        RECT 590.000 143.600 590.800 143.700 ;
        RECT 596.400 143.600 597.200 143.700 ;
        RECT 614.000 142.300 614.800 142.400 ;
        RECT 578.900 141.700 614.800 142.300 ;
        RECT 454.000 141.600 454.800 141.700 ;
        RECT 457.200 141.600 458.000 141.700 ;
        RECT 492.400 141.600 493.200 141.700 ;
        RECT 614.000 141.600 614.800 141.700 ;
        RECT 639.600 142.300 640.400 142.400 ;
        RECT 647.600 142.300 648.400 142.400 ;
        RECT 639.600 141.700 648.400 142.300 ;
        RECT 639.600 141.600 640.400 141.700 ;
        RECT 647.600 141.600 648.400 141.700 ;
        RECT 50.800 140.300 51.600 140.400 ;
        RECT 68.400 140.300 69.200 140.400 ;
        RECT 50.800 139.700 69.200 140.300 ;
        RECT 50.800 139.600 51.600 139.700 ;
        RECT 68.400 139.600 69.200 139.700 ;
        RECT 175.600 140.300 176.400 140.400 ;
        RECT 186.800 140.300 187.600 140.400 ;
        RECT 175.600 139.700 187.600 140.300 ;
        RECT 175.600 139.600 176.400 139.700 ;
        RECT 186.800 139.600 187.600 139.700 ;
        RECT 236.400 140.300 237.200 140.400 ;
        RECT 242.800 140.300 243.600 140.400 ;
        RECT 236.400 139.700 243.600 140.300 ;
        RECT 236.400 139.600 237.200 139.700 ;
        RECT 242.800 139.600 243.600 139.700 ;
        RECT 284.400 140.300 285.200 140.400 ;
        RECT 286.000 140.300 286.800 140.400 ;
        RECT 302.000 140.300 302.800 140.400 ;
        RECT 284.400 139.700 302.800 140.300 ;
        RECT 284.400 139.600 285.200 139.700 ;
        RECT 286.000 139.600 286.800 139.700 ;
        RECT 302.000 139.600 302.800 139.700 ;
        RECT 414.000 140.300 414.800 140.400 ;
        RECT 434.800 140.300 435.600 140.400 ;
        RECT 414.000 139.700 435.600 140.300 ;
        RECT 414.000 139.600 414.800 139.700 ;
        RECT 434.800 139.600 435.600 139.700 ;
        RECT 548.400 140.300 549.200 140.400 ;
        RECT 553.200 140.300 554.000 140.400 ;
        RECT 548.400 139.700 554.000 140.300 ;
        RECT 548.400 139.600 549.200 139.700 ;
        RECT 553.200 139.600 554.000 139.700 ;
        RECT 588.400 140.300 589.200 140.400 ;
        RECT 596.400 140.300 597.200 140.400 ;
        RECT 588.400 139.700 597.200 140.300 ;
        RECT 588.400 139.600 589.200 139.700 ;
        RECT 596.400 139.600 597.200 139.700 ;
        RECT 599.600 140.300 600.400 140.400 ;
        RECT 609.200 140.300 610.000 140.400 ;
        RECT 599.600 139.700 610.000 140.300 ;
        RECT 599.600 139.600 600.400 139.700 ;
        RECT 609.200 139.600 610.000 139.700 ;
        RECT 636.400 140.300 637.200 140.400 ;
        RECT 644.400 140.300 645.200 140.400 ;
        RECT 636.400 139.700 645.200 140.300 ;
        RECT 636.400 139.600 637.200 139.700 ;
        RECT 644.400 139.600 645.200 139.700 ;
        RECT 7.600 138.300 8.400 138.400 ;
        RECT 26.800 138.300 27.600 138.400 ;
        RECT 7.600 137.700 27.600 138.300 ;
        RECT 7.600 137.600 8.400 137.700 ;
        RECT 26.800 137.600 27.600 137.700 ;
        RECT 49.200 138.300 50.000 138.400 ;
        RECT 66.800 138.300 67.600 138.400 ;
        RECT 49.200 137.700 67.600 138.300 ;
        RECT 49.200 137.600 50.000 137.700 ;
        RECT 66.800 137.600 67.600 137.700 ;
        RECT 71.600 138.300 72.400 138.400 ;
        RECT 138.800 138.300 139.600 138.400 ;
        RECT 71.600 137.700 139.600 138.300 ;
        RECT 71.600 137.600 72.400 137.700 ;
        RECT 138.800 137.600 139.600 137.700 ;
        RECT 159.600 138.300 160.400 138.400 ;
        RECT 255.600 138.300 256.400 138.400 ;
        RECT 159.600 137.700 256.400 138.300 ;
        RECT 159.600 137.600 160.400 137.700 ;
        RECT 255.600 137.600 256.400 137.700 ;
        RECT 268.400 138.300 269.200 138.400 ;
        RECT 274.800 138.300 275.600 138.400 ;
        RECT 268.400 137.700 275.600 138.300 ;
        RECT 268.400 137.600 269.200 137.700 ;
        RECT 274.800 137.600 275.600 137.700 ;
        RECT 378.800 138.300 379.600 138.400 ;
        RECT 394.800 138.300 395.600 138.400 ;
        RECT 431.600 138.300 432.400 138.400 ;
        RECT 378.800 137.700 432.400 138.300 ;
        RECT 378.800 137.600 379.600 137.700 ;
        RECT 394.800 137.600 395.600 137.700 ;
        RECT 431.600 137.600 432.400 137.700 ;
        RECT 546.800 138.300 547.600 138.400 ;
        RECT 561.200 138.300 562.000 138.400 ;
        RECT 588.400 138.300 589.200 138.400 ;
        RECT 604.400 138.300 605.200 138.400 ;
        RECT 625.200 138.300 626.000 138.400 ;
        RECT 546.800 137.700 569.900 138.300 ;
        RECT 546.800 137.600 547.600 137.700 ;
        RECT 561.200 137.600 562.000 137.700 ;
        RECT 60.400 136.300 61.200 136.400 ;
        RECT 76.400 136.300 77.200 136.400 ;
        RECT 60.400 135.700 77.200 136.300 ;
        RECT 60.400 135.600 61.200 135.700 ;
        RECT 76.400 135.600 77.200 135.700 ;
        RECT 108.400 136.300 109.200 136.400 ;
        RECT 154.800 136.300 155.600 136.400 ;
        RECT 108.400 135.700 155.600 136.300 ;
        RECT 108.400 135.600 109.200 135.700 ;
        RECT 154.800 135.600 155.600 135.700 ;
        RECT 186.800 136.300 187.600 136.400 ;
        RECT 196.400 136.300 197.200 136.400 ;
        RECT 186.800 135.700 197.200 136.300 ;
        RECT 186.800 135.600 187.600 135.700 ;
        RECT 196.400 135.600 197.200 135.700 ;
        RECT 246.000 136.300 246.800 136.400 ;
        RECT 252.400 136.300 253.200 136.400 ;
        RECT 274.800 136.300 275.600 136.400 ;
        RECT 289.200 136.300 290.000 136.400 ;
        RECT 246.000 135.700 290.000 136.300 ;
        RECT 246.000 135.600 246.800 135.700 ;
        RECT 252.400 135.600 253.200 135.700 ;
        RECT 274.800 135.600 275.600 135.700 ;
        RECT 289.200 135.600 290.000 135.700 ;
        RECT 295.600 135.600 296.400 136.400 ;
        RECT 305.200 136.300 306.000 136.400 ;
        RECT 311.600 136.300 312.400 136.400 ;
        RECT 305.200 135.700 312.400 136.300 ;
        RECT 305.200 135.600 306.000 135.700 ;
        RECT 311.600 135.600 312.400 135.700 ;
        RECT 425.200 136.300 426.000 136.400 ;
        RECT 438.000 136.300 438.800 136.400 ;
        RECT 425.200 135.700 438.800 136.300 ;
        RECT 425.200 135.600 426.000 135.700 ;
        RECT 438.000 135.600 438.800 135.700 ;
        RECT 492.400 136.300 493.200 136.400 ;
        RECT 506.800 136.300 507.600 136.400 ;
        RECT 492.400 135.700 507.600 136.300 ;
        RECT 492.400 135.600 493.200 135.700 ;
        RECT 506.800 135.600 507.600 135.700 ;
        RECT 516.400 136.300 517.200 136.400 ;
        RECT 519.600 136.300 520.400 136.400 ;
        RECT 516.400 135.700 520.400 136.300 ;
        RECT 516.400 135.600 517.200 135.700 ;
        RECT 519.600 135.600 520.400 135.700 ;
        RECT 540.400 136.300 541.200 136.400 ;
        RECT 553.200 136.300 554.000 136.400 ;
        RECT 567.600 136.300 568.400 136.400 ;
        RECT 540.400 135.700 568.400 136.300 ;
        RECT 569.300 136.300 569.900 137.700 ;
        RECT 588.400 137.700 626.000 138.300 ;
        RECT 588.400 137.600 589.200 137.700 ;
        RECT 604.400 137.600 605.200 137.700 ;
        RECT 625.200 137.600 626.000 137.700 ;
        RECT 657.200 138.300 658.000 138.400 ;
        RECT 671.600 138.300 672.400 138.400 ;
        RECT 657.200 137.700 672.400 138.300 ;
        RECT 657.200 137.600 658.000 137.700 ;
        RECT 671.600 137.600 672.400 137.700 ;
        RECT 601.200 136.300 602.000 136.400 ;
        RECT 657.200 136.300 658.000 136.400 ;
        RECT 569.300 135.700 658.000 136.300 ;
        RECT 540.400 135.600 541.200 135.700 ;
        RECT 553.200 135.600 554.000 135.700 ;
        RECT 567.600 135.600 568.400 135.700 ;
        RECT 601.200 135.600 602.000 135.700 ;
        RECT 657.200 135.600 658.000 135.700 ;
        RECT 26.800 134.300 27.600 134.400 ;
        RECT 34.800 134.300 35.600 134.400 ;
        RECT 54.000 134.300 54.800 134.400 ;
        RECT 26.800 133.700 54.800 134.300 ;
        RECT 26.800 133.600 27.600 133.700 ;
        RECT 34.800 133.600 35.600 133.700 ;
        RECT 54.000 133.600 54.800 133.700 ;
        RECT 63.600 134.300 64.400 134.400 ;
        RECT 74.800 134.300 75.600 134.400 ;
        RECT 63.600 133.700 75.600 134.300 ;
        RECT 63.600 133.600 64.400 133.700 ;
        RECT 74.800 133.600 75.600 133.700 ;
        RECT 90.800 134.300 91.600 134.400 ;
        RECT 111.600 134.300 112.400 134.400 ;
        RECT 90.800 133.700 112.400 134.300 ;
        RECT 90.800 133.600 91.600 133.700 ;
        RECT 111.600 133.600 112.400 133.700 ;
        RECT 122.800 134.300 123.600 134.400 ;
        RECT 161.200 134.300 162.000 134.400 ;
        RECT 122.800 133.700 162.000 134.300 ;
        RECT 122.800 133.600 123.600 133.700 ;
        RECT 161.200 133.600 162.000 133.700 ;
        RECT 178.800 134.300 179.600 134.400 ;
        RECT 194.800 134.300 195.600 134.400 ;
        RECT 178.800 133.700 195.600 134.300 ;
        RECT 178.800 133.600 179.600 133.700 ;
        RECT 194.800 133.600 195.600 133.700 ;
        RECT 279.600 134.300 280.400 134.400 ;
        RECT 305.200 134.300 306.000 134.400 ;
        RECT 279.600 133.700 306.000 134.300 ;
        RECT 279.600 133.600 280.400 133.700 ;
        RECT 305.200 133.600 306.000 133.700 ;
        RECT 391.600 134.300 392.400 134.400 ;
        RECT 454.000 134.300 454.800 134.400 ;
        RECT 476.400 134.300 477.200 134.400 ;
        RECT 391.600 133.700 433.900 134.300 ;
        RECT 391.600 133.600 392.400 133.700 ;
        RECT 433.300 132.400 433.900 133.700 ;
        RECT 454.000 133.700 477.200 134.300 ;
        RECT 454.000 133.600 454.800 133.700 ;
        RECT 476.400 133.600 477.200 133.700 ;
        RECT 489.200 134.300 490.000 134.400 ;
        RECT 526.000 134.300 526.800 134.400 ;
        RECT 489.200 133.700 526.800 134.300 ;
        RECT 489.200 133.600 490.000 133.700 ;
        RECT 526.000 133.600 526.800 133.700 ;
        RECT 542.000 134.300 542.800 134.400 ;
        RECT 543.600 134.300 544.400 134.400 ;
        RECT 606.000 134.300 606.800 134.400 ;
        RECT 612.400 134.300 613.200 134.400 ;
        RECT 542.000 133.700 613.200 134.300 ;
        RECT 542.000 133.600 542.800 133.700 ;
        RECT 543.600 133.600 544.400 133.700 ;
        RECT 606.000 133.600 606.800 133.700 ;
        RECT 612.400 133.600 613.200 133.700 ;
        RECT 617.200 134.300 618.000 134.400 ;
        RECT 633.200 134.300 634.000 134.400 ;
        RECT 617.200 133.700 634.000 134.300 ;
        RECT 617.200 133.600 618.000 133.700 ;
        RECT 633.200 133.600 634.000 133.700 ;
        RECT 646.000 134.300 646.800 134.400 ;
        RECT 650.800 134.300 651.600 134.400 ;
        RECT 654.000 134.300 654.800 134.400 ;
        RECT 646.000 133.700 654.800 134.300 ;
        RECT 646.000 133.600 646.800 133.700 ;
        RECT 650.800 133.600 651.600 133.700 ;
        RECT 654.000 133.600 654.800 133.700 ;
        RECT 12.400 132.300 13.200 132.400 ;
        RECT 38.000 132.300 38.800 132.400 ;
        RECT 12.400 131.700 38.800 132.300 ;
        RECT 12.400 131.600 13.200 131.700 ;
        RECT 38.000 131.600 38.800 131.700 ;
        RECT 39.600 132.300 40.400 132.400 ;
        RECT 58.800 132.300 59.600 132.400 ;
        RECT 39.600 131.700 59.600 132.300 ;
        RECT 39.600 131.600 40.400 131.700 ;
        RECT 58.800 131.600 59.600 131.700 ;
        RECT 66.800 132.300 67.600 132.400 ;
        RECT 92.400 132.300 93.200 132.400 ;
        RECT 66.800 131.700 93.200 132.300 ;
        RECT 66.800 131.600 67.600 131.700 ;
        RECT 92.400 131.600 93.200 131.700 ;
        RECT 98.800 132.300 99.600 132.400 ;
        RECT 100.400 132.300 101.200 132.400 ;
        RECT 98.800 131.700 101.200 132.300 ;
        RECT 98.800 131.600 99.600 131.700 ;
        RECT 100.400 131.600 101.200 131.700 ;
        RECT 126.000 132.300 126.800 132.400 ;
        RECT 143.600 132.300 144.400 132.400 ;
        RECT 126.000 131.700 144.400 132.300 ;
        RECT 126.000 131.600 126.800 131.700 ;
        RECT 143.600 131.600 144.400 131.700 ;
        RECT 148.400 132.300 149.200 132.400 ;
        RECT 156.400 132.300 157.200 132.400 ;
        RECT 148.400 131.700 157.200 132.300 ;
        RECT 148.400 131.600 149.200 131.700 ;
        RECT 156.400 131.600 157.200 131.700 ;
        RECT 191.600 132.300 192.400 132.400 ;
        RECT 193.200 132.300 194.000 132.400 ;
        RECT 191.600 131.700 194.000 132.300 ;
        RECT 191.600 131.600 192.400 131.700 ;
        RECT 193.200 131.600 194.000 131.700 ;
        RECT 255.600 132.300 256.400 132.400 ;
        RECT 271.600 132.300 272.400 132.400 ;
        RECT 273.200 132.300 274.000 132.400 ;
        RECT 255.600 131.700 274.000 132.300 ;
        RECT 255.600 131.600 256.400 131.700 ;
        RECT 271.600 131.600 272.400 131.700 ;
        RECT 273.200 131.600 274.000 131.700 ;
        RECT 287.600 132.300 288.400 132.400 ;
        RECT 295.600 132.300 296.400 132.400 ;
        RECT 287.600 131.700 296.400 132.300 ;
        RECT 287.600 131.600 288.400 131.700 ;
        RECT 295.600 131.600 296.400 131.700 ;
        RECT 375.600 132.300 376.400 132.400 ;
        RECT 402.800 132.300 403.600 132.400 ;
        RECT 375.600 131.700 403.600 132.300 ;
        RECT 375.600 131.600 376.400 131.700 ;
        RECT 402.800 131.600 403.600 131.700 ;
        RECT 433.200 132.300 434.000 132.400 ;
        RECT 436.400 132.300 437.200 132.400 ;
        RECT 433.200 131.700 437.200 132.300 ;
        RECT 433.200 131.600 434.000 131.700 ;
        RECT 436.400 131.600 437.200 131.700 ;
        RECT 441.200 132.300 442.000 132.400 ;
        RECT 444.400 132.300 445.200 132.400 ;
        RECT 441.200 131.700 445.200 132.300 ;
        RECT 441.200 131.600 442.000 131.700 ;
        RECT 444.400 131.600 445.200 131.700 ;
        RECT 506.800 132.300 507.600 132.400 ;
        RECT 514.800 132.300 515.600 132.400 ;
        RECT 506.800 131.700 515.600 132.300 ;
        RECT 506.800 131.600 507.600 131.700 ;
        RECT 514.800 131.600 515.600 131.700 ;
        RECT 530.800 132.300 531.600 132.400 ;
        RECT 546.800 132.300 547.600 132.400 ;
        RECT 530.800 131.700 547.600 132.300 ;
        RECT 530.800 131.600 531.600 131.700 ;
        RECT 546.800 131.600 547.600 131.700 ;
        RECT 550.000 132.300 550.800 132.400 ;
        RECT 559.600 132.300 560.400 132.400 ;
        RECT 550.000 131.700 560.400 132.300 ;
        RECT 550.000 131.600 550.800 131.700 ;
        RECT 559.600 131.600 560.400 131.700 ;
        RECT 567.600 132.300 568.400 132.400 ;
        RECT 586.800 132.300 587.600 132.400 ;
        RECT 567.600 131.700 587.600 132.300 ;
        RECT 567.600 131.600 568.400 131.700 ;
        RECT 586.800 131.600 587.600 131.700 ;
        RECT 593.200 132.300 594.000 132.400 ;
        RECT 596.400 132.300 597.200 132.400 ;
        RECT 593.200 131.700 597.200 132.300 ;
        RECT 593.200 131.600 594.000 131.700 ;
        RECT 596.400 131.600 597.200 131.700 ;
        RECT 601.200 132.300 602.000 132.400 ;
        RECT 612.400 132.300 613.200 132.400 ;
        RECT 601.200 131.700 613.200 132.300 ;
        RECT 601.200 131.600 602.000 131.700 ;
        RECT 612.400 131.600 613.200 131.700 ;
        RECT 620.400 132.300 621.200 132.400 ;
        RECT 638.000 132.300 638.800 132.400 ;
        RECT 620.400 131.700 638.800 132.300 ;
        RECT 620.400 131.600 621.200 131.700 ;
        RECT 638.000 131.600 638.800 131.700 ;
        RECT 652.400 132.300 653.200 132.400 ;
        RECT 665.200 132.300 666.000 132.400 ;
        RECT 652.400 131.700 666.000 132.300 ;
        RECT 652.400 131.600 653.200 131.700 ;
        RECT 665.200 131.600 666.000 131.700 ;
        RECT 668.400 132.300 669.200 132.400 ;
        RECT 679.600 132.300 680.400 132.400 ;
        RECT 668.400 131.700 680.400 132.300 ;
        RECT 668.400 131.600 669.200 131.700 ;
        RECT 679.600 131.600 680.400 131.700 ;
        RECT 23.600 130.300 24.400 130.400 ;
        RECT 26.800 130.300 27.600 130.400 ;
        RECT 23.600 129.700 27.600 130.300 ;
        RECT 23.600 129.600 24.400 129.700 ;
        RECT 26.800 129.600 27.600 129.700 ;
        RECT 50.800 130.300 51.600 130.400 ;
        RECT 57.200 130.300 58.000 130.400 ;
        RECT 71.600 130.300 72.400 130.400 ;
        RECT 50.800 129.700 72.400 130.300 ;
        RECT 50.800 129.600 51.600 129.700 ;
        RECT 57.200 129.600 58.000 129.700 ;
        RECT 71.600 129.600 72.400 129.700 ;
        RECT 76.400 130.300 77.200 130.400 ;
        RECT 158.000 130.300 158.800 130.400 ;
        RECT 76.400 129.700 158.800 130.300 ;
        RECT 76.400 129.600 77.200 129.700 ;
        RECT 158.000 129.600 158.800 129.700 ;
        RECT 172.400 130.300 173.200 130.400 ;
        RECT 177.200 130.300 178.000 130.400 ;
        RECT 172.400 129.700 178.000 130.300 ;
        RECT 172.400 129.600 173.200 129.700 ;
        RECT 177.200 129.600 178.000 129.700 ;
        RECT 260.400 130.300 261.200 130.400 ;
        RECT 290.800 130.300 291.600 130.400 ;
        RECT 260.400 129.700 291.600 130.300 ;
        RECT 260.400 129.600 261.200 129.700 ;
        RECT 290.800 129.600 291.600 129.700 ;
        RECT 294.000 130.300 294.800 130.400 ;
        RECT 297.200 130.300 298.000 130.400 ;
        RECT 294.000 129.700 298.000 130.300 ;
        RECT 294.000 129.600 294.800 129.700 ;
        RECT 297.200 129.600 298.000 129.700 ;
        RECT 300.400 130.300 301.200 130.400 ;
        RECT 308.400 130.300 309.200 130.400 ;
        RECT 300.400 129.700 309.200 130.300 ;
        RECT 300.400 129.600 301.200 129.700 ;
        RECT 308.400 129.600 309.200 129.700 ;
        RECT 534.000 130.300 534.800 130.400 ;
        RECT 540.400 130.300 541.200 130.400 ;
        RECT 572.400 130.300 573.200 130.400 ;
        RECT 534.000 129.700 573.200 130.300 ;
        RECT 534.000 129.600 534.800 129.700 ;
        RECT 540.400 129.600 541.200 129.700 ;
        RECT 572.400 129.600 573.200 129.700 ;
        RECT 590.000 130.300 590.800 130.400 ;
        RECT 596.400 130.300 597.200 130.400 ;
        RECT 590.000 129.700 597.200 130.300 ;
        RECT 590.000 129.600 590.800 129.700 ;
        RECT 596.400 129.600 597.200 129.700 ;
        RECT 599.600 130.300 600.400 130.400 ;
        RECT 610.800 130.300 611.600 130.400 ;
        RECT 599.600 129.700 611.600 130.300 ;
        RECT 599.600 129.600 600.400 129.700 ;
        RECT 610.800 129.600 611.600 129.700 ;
        RECT 617.200 130.300 618.000 130.400 ;
        RECT 620.400 130.300 621.200 130.400 ;
        RECT 617.200 129.700 621.200 130.300 ;
        RECT 617.200 129.600 618.000 129.700 ;
        RECT 620.400 129.600 621.200 129.700 ;
        RECT 641.200 130.300 642.000 130.400 ;
        RECT 660.400 130.300 661.200 130.400 ;
        RECT 641.200 129.700 661.200 130.300 ;
        RECT 641.200 129.600 642.000 129.700 ;
        RECT 660.400 129.600 661.200 129.700 ;
        RECT 666.800 130.300 667.600 130.400 ;
        RECT 668.400 130.300 669.200 130.400 ;
        RECT 666.800 129.700 669.200 130.300 ;
        RECT 666.800 129.600 667.600 129.700 ;
        RECT 668.400 129.600 669.200 129.700 ;
        RECT 38.000 128.300 38.800 128.400 ;
        RECT 122.800 128.300 123.600 128.400 ;
        RECT 38.000 127.700 123.600 128.300 ;
        RECT 38.000 127.600 38.800 127.700 ;
        RECT 122.800 127.600 123.600 127.700 ;
        RECT 124.400 128.300 125.200 128.400 ;
        RECT 146.800 128.300 147.600 128.400 ;
        RECT 124.400 127.700 147.600 128.300 ;
        RECT 124.400 127.600 125.200 127.700 ;
        RECT 146.800 127.600 147.600 127.700 ;
        RECT 159.600 128.300 160.400 128.400 ;
        RECT 185.200 128.300 186.000 128.400 ;
        RECT 199.600 128.300 200.400 128.400 ;
        RECT 244.400 128.300 245.200 128.400 ;
        RECT 159.600 127.700 245.200 128.300 ;
        RECT 159.600 127.600 160.400 127.700 ;
        RECT 185.200 127.600 186.000 127.700 ;
        RECT 199.600 127.600 200.400 127.700 ;
        RECT 244.400 127.600 245.200 127.700 ;
        RECT 276.400 128.300 277.200 128.400 ;
        RECT 279.600 128.300 280.400 128.400 ;
        RECT 276.400 127.700 280.400 128.300 ;
        RECT 276.400 127.600 277.200 127.700 ;
        RECT 279.600 127.600 280.400 127.700 ;
        RECT 294.000 128.300 294.800 128.400 ;
        RECT 327.600 128.300 328.400 128.400 ;
        RECT 294.000 127.700 328.400 128.300 ;
        RECT 294.000 127.600 294.800 127.700 ;
        RECT 327.600 127.600 328.400 127.700 ;
        RECT 518.000 128.300 518.800 128.400 ;
        RECT 550.000 128.300 550.800 128.400 ;
        RECT 518.000 127.700 550.800 128.300 ;
        RECT 518.000 127.600 518.800 127.700 ;
        RECT 550.000 127.600 550.800 127.700 ;
        RECT 556.400 128.300 557.200 128.400 ;
        RECT 582.000 128.300 582.800 128.400 ;
        RECT 593.200 128.300 594.000 128.400 ;
        RECT 556.400 127.700 594.000 128.300 ;
        RECT 556.400 127.600 557.200 127.700 ;
        RECT 582.000 127.600 582.800 127.700 ;
        RECT 593.200 127.600 594.000 127.700 ;
        RECT 598.000 128.300 598.800 128.400 ;
        RECT 644.400 128.300 645.200 128.400 ;
        RECT 598.000 127.700 645.200 128.300 ;
        RECT 598.000 127.600 598.800 127.700 ;
        RECT 644.400 127.600 645.200 127.700 ;
        RECT 132.400 126.300 133.200 126.400 ;
        RECT 28.500 125.700 133.200 126.300 ;
        RECT 28.500 124.400 29.100 125.700 ;
        RECT 132.400 125.600 133.200 125.700 ;
        RECT 134.000 126.300 134.800 126.400 ;
        RECT 174.000 126.300 174.800 126.400 ;
        RECT 134.000 125.700 174.800 126.300 ;
        RECT 134.000 125.600 134.800 125.700 ;
        RECT 174.000 125.600 174.800 125.700 ;
        RECT 196.400 126.300 197.200 126.400 ;
        RECT 302.000 126.300 302.800 126.400 ;
        RECT 196.400 125.700 302.800 126.300 ;
        RECT 196.400 125.600 197.200 125.700 ;
        RECT 302.000 125.600 302.800 125.700 ;
        RECT 335.600 126.300 336.400 126.400 ;
        RECT 342.000 126.300 342.800 126.400 ;
        RECT 335.600 125.700 342.800 126.300 ;
        RECT 335.600 125.600 336.400 125.700 ;
        RECT 342.000 125.600 342.800 125.700 ;
        RECT 423.600 126.300 424.400 126.400 ;
        RECT 433.200 126.300 434.000 126.400 ;
        RECT 423.600 125.700 434.000 126.300 ;
        RECT 423.600 125.600 424.400 125.700 ;
        RECT 433.200 125.600 434.000 125.700 ;
        RECT 594.800 126.300 595.600 126.400 ;
        RECT 623.600 126.300 624.400 126.400 ;
        RECT 594.800 125.700 624.400 126.300 ;
        RECT 594.800 125.600 595.600 125.700 ;
        RECT 623.600 125.600 624.400 125.700 ;
        RECT 18.800 124.300 19.600 124.400 ;
        RECT 28.400 124.300 29.200 124.400 ;
        RECT 18.800 123.700 29.200 124.300 ;
        RECT 18.800 123.600 19.600 123.700 ;
        RECT 28.400 123.600 29.200 123.700 ;
        RECT 102.000 124.300 102.800 124.400 ;
        RECT 103.600 124.300 104.400 124.400 ;
        RECT 134.100 124.300 134.700 125.600 ;
        RECT 102.000 123.700 134.700 124.300 ;
        RECT 142.000 124.300 142.800 124.400 ;
        RECT 148.400 124.300 149.200 124.400 ;
        RECT 169.200 124.300 170.000 124.400 ;
        RECT 142.000 123.700 170.000 124.300 ;
        RECT 102.000 123.600 102.800 123.700 ;
        RECT 103.600 123.600 104.400 123.700 ;
        RECT 142.000 123.600 142.800 123.700 ;
        RECT 148.400 123.600 149.200 123.700 ;
        RECT 169.200 123.600 170.000 123.700 ;
        RECT 174.000 124.300 174.800 124.400 ;
        RECT 190.000 124.300 190.800 124.400 ;
        RECT 202.800 124.300 203.600 124.400 ;
        RECT 174.000 123.700 203.600 124.300 ;
        RECT 174.000 123.600 174.800 123.700 ;
        RECT 190.000 123.600 190.800 123.700 ;
        RECT 202.800 123.600 203.600 123.700 ;
        RECT 230.000 124.300 230.800 124.400 ;
        RECT 236.400 124.300 237.200 124.400 ;
        RECT 241.200 124.300 242.000 124.400 ;
        RECT 230.000 123.700 237.200 124.300 ;
        RECT 230.000 123.600 230.800 123.700 ;
        RECT 236.400 123.600 237.200 123.700 ;
        RECT 239.700 123.700 242.000 124.300 ;
        RECT 212.400 122.300 213.200 122.400 ;
        RECT 239.700 122.300 240.300 123.700 ;
        RECT 241.200 123.600 242.000 123.700 ;
        RECT 244.400 124.300 245.200 124.400 ;
        RECT 250.800 124.300 251.600 124.400 ;
        RECT 244.400 123.700 251.600 124.300 ;
        RECT 244.400 123.600 245.200 123.700 ;
        RECT 250.800 123.600 251.600 123.700 ;
        RECT 383.600 124.300 384.400 124.400 ;
        RECT 401.200 124.300 402.000 124.400 ;
        RECT 383.600 123.700 402.000 124.300 ;
        RECT 383.600 123.600 384.400 123.700 ;
        RECT 401.200 123.600 402.000 123.700 ;
        RECT 537.200 124.300 538.000 124.400 ;
        RECT 564.400 124.300 565.200 124.400 ;
        RECT 631.600 124.300 632.400 124.400 ;
        RECT 634.800 124.300 635.600 124.400 ;
        RECT 537.200 123.700 635.600 124.300 ;
        RECT 537.200 123.600 538.000 123.700 ;
        RECT 564.400 123.600 565.200 123.700 ;
        RECT 631.600 123.600 632.400 123.700 ;
        RECT 634.800 123.600 635.600 123.700 ;
        RECT 681.200 124.300 682.000 124.400 ;
        RECT 684.400 124.300 685.200 124.400 ;
        RECT 681.200 123.700 685.200 124.300 ;
        RECT 681.200 123.600 682.000 123.700 ;
        RECT 684.400 123.600 685.200 123.700 ;
        RECT 282.800 122.300 283.600 122.400 ;
        RECT 212.400 121.700 240.300 122.300 ;
        RECT 241.300 121.700 283.600 122.300 ;
        RECT 212.400 121.600 213.200 121.700 ;
        RECT 241.300 120.400 241.900 121.700 ;
        RECT 282.800 121.600 283.600 121.700 ;
        RECT 364.400 122.300 365.200 122.400 ;
        RECT 409.200 122.300 410.000 122.400 ;
        RECT 364.400 121.700 410.000 122.300 ;
        RECT 364.400 121.600 365.200 121.700 ;
        RECT 409.200 121.600 410.000 121.700 ;
        RECT 572.400 122.300 573.200 122.400 ;
        RECT 620.400 122.300 621.200 122.400 ;
        RECT 641.200 122.300 642.000 122.400 ;
        RECT 572.400 121.700 642.000 122.300 ;
        RECT 572.400 121.600 573.200 121.700 ;
        RECT 620.400 121.600 621.200 121.700 ;
        RECT 641.200 121.600 642.000 121.700 ;
        RECT 46.000 120.300 46.800 120.400 ;
        RECT 52.400 120.300 53.200 120.400 ;
        RECT 46.000 119.700 53.200 120.300 ;
        RECT 46.000 119.600 46.800 119.700 ;
        RECT 52.400 119.600 53.200 119.700 ;
        RECT 143.600 120.300 144.400 120.400 ;
        RECT 175.600 120.300 176.400 120.400 ;
        RECT 143.600 119.700 176.400 120.300 ;
        RECT 143.600 119.600 144.400 119.700 ;
        RECT 175.600 119.600 176.400 119.700 ;
        RECT 199.600 120.300 200.400 120.400 ;
        RECT 222.000 120.300 222.800 120.400 ;
        RECT 199.600 119.700 222.800 120.300 ;
        RECT 199.600 119.600 200.400 119.700 ;
        RECT 222.000 119.600 222.800 119.700 ;
        RECT 223.600 120.300 224.400 120.400 ;
        RECT 241.200 120.300 242.000 120.400 ;
        RECT 223.600 119.700 242.000 120.300 ;
        RECT 223.600 119.600 224.400 119.700 ;
        RECT 241.200 119.600 242.000 119.700 ;
        RECT 249.200 120.300 250.000 120.400 ;
        RECT 252.400 120.300 253.200 120.400 ;
        RECT 295.600 120.300 296.400 120.400 ;
        RECT 297.200 120.300 298.000 120.400 ;
        RECT 306.800 120.300 307.600 120.400 ;
        RECT 318.000 120.300 318.800 120.400 ;
        RECT 342.000 120.300 342.800 120.400 ;
        RECT 249.200 119.700 342.800 120.300 ;
        RECT 249.200 119.600 250.000 119.700 ;
        RECT 252.400 119.600 253.200 119.700 ;
        RECT 295.600 119.600 296.400 119.700 ;
        RECT 297.200 119.600 298.000 119.700 ;
        RECT 306.800 119.600 307.600 119.700 ;
        RECT 318.000 119.600 318.800 119.700 ;
        RECT 342.000 119.600 342.800 119.700 ;
        RECT 351.600 120.300 352.400 120.400 ;
        RECT 364.400 120.300 365.200 120.400 ;
        RECT 351.600 119.700 365.200 120.300 ;
        RECT 351.600 119.600 352.400 119.700 ;
        RECT 364.400 119.600 365.200 119.700 ;
        RECT 388.400 120.300 389.200 120.400 ;
        RECT 391.600 120.300 392.400 120.400 ;
        RECT 399.600 120.300 400.400 120.400 ;
        RECT 388.400 119.700 400.400 120.300 ;
        RECT 388.400 119.600 389.200 119.700 ;
        RECT 391.600 119.600 392.400 119.700 ;
        RECT 399.600 119.600 400.400 119.700 ;
        RECT 530.800 120.300 531.600 120.400 ;
        RECT 551.600 120.300 552.400 120.400 ;
        RECT 578.800 120.300 579.600 120.400 ;
        RECT 599.600 120.300 600.400 120.400 ;
        RECT 530.800 119.700 600.400 120.300 ;
        RECT 530.800 119.600 531.600 119.700 ;
        RECT 551.600 119.600 552.400 119.700 ;
        RECT 578.800 119.600 579.600 119.700 ;
        RECT 599.600 119.600 600.400 119.700 ;
        RECT 634.800 120.300 635.600 120.400 ;
        RECT 638.000 120.300 638.800 120.400 ;
        RECT 674.800 120.300 675.600 120.400 ;
        RECT 634.800 119.700 675.600 120.300 ;
        RECT 634.800 119.600 635.600 119.700 ;
        RECT 638.000 119.600 638.800 119.700 ;
        RECT 674.800 119.600 675.600 119.700 ;
        RECT 98.800 118.300 99.600 118.400 ;
        RECT 106.800 118.300 107.600 118.400 ;
        RECT 98.800 117.700 107.600 118.300 ;
        RECT 98.800 117.600 99.600 117.700 ;
        RECT 106.800 117.600 107.600 117.700 ;
        RECT 118.000 118.300 118.800 118.400 ;
        RECT 122.800 118.300 123.600 118.400 ;
        RECT 118.000 117.700 123.600 118.300 ;
        RECT 118.000 117.600 118.800 117.700 ;
        RECT 122.800 117.600 123.600 117.700 ;
        RECT 126.000 118.300 126.800 118.400 ;
        RECT 167.600 118.300 168.400 118.400 ;
        RECT 126.000 117.700 168.400 118.300 ;
        RECT 126.000 117.600 126.800 117.700 ;
        RECT 167.600 117.600 168.400 117.700 ;
        RECT 218.800 118.300 219.600 118.400 ;
        RECT 236.400 118.300 237.200 118.400 ;
        RECT 218.800 117.700 237.200 118.300 ;
        RECT 218.800 117.600 219.600 117.700 ;
        RECT 236.400 117.600 237.200 117.700 ;
        RECT 238.000 118.300 238.800 118.400 ;
        RECT 242.800 118.300 243.600 118.400 ;
        RECT 238.000 117.700 243.600 118.300 ;
        RECT 238.000 117.600 238.800 117.700 ;
        RECT 242.800 117.600 243.600 117.700 ;
        RECT 350.000 118.300 350.800 118.400 ;
        RECT 393.200 118.300 394.000 118.400 ;
        RECT 404.400 118.300 405.200 118.400 ;
        RECT 415.600 118.300 416.400 118.400 ;
        RECT 428.400 118.300 429.200 118.400 ;
        RECT 350.000 117.700 429.200 118.300 ;
        RECT 350.000 117.600 350.800 117.700 ;
        RECT 393.200 117.600 394.000 117.700 ;
        RECT 404.400 117.600 405.200 117.700 ;
        RECT 415.600 117.600 416.400 117.700 ;
        RECT 428.400 117.600 429.200 117.700 ;
        RECT 439.600 118.300 440.400 118.400 ;
        RECT 449.200 118.300 450.000 118.400 ;
        RECT 439.600 117.700 450.000 118.300 ;
        RECT 439.600 117.600 440.400 117.700 ;
        RECT 449.200 117.600 450.000 117.700 ;
        RECT 465.200 118.300 466.000 118.400 ;
        RECT 474.800 118.300 475.600 118.400 ;
        RECT 586.800 118.300 587.600 118.400 ;
        RECT 465.200 117.700 587.600 118.300 ;
        RECT 465.200 117.600 466.000 117.700 ;
        RECT 474.800 117.600 475.600 117.700 ;
        RECT 586.800 117.600 587.600 117.700 ;
        RECT 626.800 118.300 627.600 118.400 ;
        RECT 639.600 118.300 640.400 118.400 ;
        RECT 626.800 117.700 640.400 118.300 ;
        RECT 626.800 117.600 627.600 117.700 ;
        RECT 639.600 117.600 640.400 117.700 ;
        RECT 98.800 116.300 99.600 116.400 ;
        RECT 162.800 116.300 163.600 116.400 ;
        RECT 177.200 116.300 178.000 116.400 ;
        RECT 98.800 115.700 178.000 116.300 ;
        RECT 98.800 115.600 99.600 115.700 ;
        RECT 162.800 115.600 163.600 115.700 ;
        RECT 177.200 115.600 178.000 115.700 ;
        RECT 182.000 116.300 182.800 116.400 ;
        RECT 260.400 116.300 261.200 116.400 ;
        RECT 182.000 115.700 261.200 116.300 ;
        RECT 182.000 115.600 182.800 115.700 ;
        RECT 260.400 115.600 261.200 115.700 ;
        RECT 385.200 116.300 386.000 116.400 ;
        RECT 412.400 116.300 413.200 116.400 ;
        RECT 425.200 116.300 426.000 116.400 ;
        RECT 385.200 115.700 426.000 116.300 ;
        RECT 385.200 115.600 386.000 115.700 ;
        RECT 412.400 115.600 413.200 115.700 ;
        RECT 425.200 115.600 426.000 115.700 ;
        RECT 442.800 116.300 443.600 116.400 ;
        RECT 471.600 116.300 472.400 116.400 ;
        RECT 482.800 116.300 483.600 116.400 ;
        RECT 442.800 115.700 483.600 116.300 ;
        RECT 442.800 115.600 443.600 115.700 ;
        RECT 471.600 115.600 472.400 115.700 ;
        RECT 482.800 115.600 483.600 115.700 ;
        RECT 522.800 116.300 523.600 116.400 ;
        RECT 526.000 116.300 526.800 116.400 ;
        RECT 537.200 116.300 538.000 116.400 ;
        RECT 522.800 115.700 538.000 116.300 ;
        RECT 522.800 115.600 523.600 115.700 ;
        RECT 526.000 115.600 526.800 115.700 ;
        RECT 537.200 115.600 538.000 115.700 ;
        RECT 558.000 116.300 558.800 116.400 ;
        RECT 566.000 116.300 566.800 116.400 ;
        RECT 580.400 116.300 581.200 116.400 ;
        RECT 585.200 116.300 586.000 116.400 ;
        RECT 596.400 116.300 597.200 116.400 ;
        RECT 558.000 115.700 597.200 116.300 ;
        RECT 558.000 115.600 558.800 115.700 ;
        RECT 566.000 115.600 566.800 115.700 ;
        RECT 580.400 115.600 581.200 115.700 ;
        RECT 585.200 115.600 586.000 115.700 ;
        RECT 596.400 115.600 597.200 115.700 ;
        RECT 604.400 116.300 605.200 116.400 ;
        RECT 630.000 116.300 630.800 116.400 ;
        RECT 638.000 116.300 638.800 116.400 ;
        RECT 604.400 115.700 638.800 116.300 ;
        RECT 604.400 115.600 605.200 115.700 ;
        RECT 630.000 115.600 630.800 115.700 ;
        RECT 638.000 115.600 638.800 115.700 ;
        RECT 652.400 116.300 653.200 116.400 ;
        RECT 654.000 116.300 654.800 116.400 ;
        RECT 652.400 115.700 654.800 116.300 ;
        RECT 652.400 115.600 653.200 115.700 ;
        RECT 654.000 115.600 654.800 115.700 ;
        RECT 66.800 114.300 67.600 114.400 ;
        RECT 78.000 114.300 78.800 114.400 ;
        RECT 81.200 114.300 82.000 114.400 ;
        RECT 66.800 113.700 82.000 114.300 ;
        RECT 66.800 113.600 67.600 113.700 ;
        RECT 78.000 113.600 78.800 113.700 ;
        RECT 81.200 113.600 82.000 113.700 ;
        RECT 121.200 114.300 122.000 114.400 ;
        RECT 238.000 114.300 238.800 114.400 ;
        RECT 239.600 114.300 240.400 114.400 ;
        RECT 121.200 113.700 128.300 114.300 ;
        RECT 121.200 113.600 122.000 113.700 ;
        RECT 127.700 112.400 128.300 113.700 ;
        RECT 238.000 113.700 240.400 114.300 ;
        RECT 238.000 113.600 238.800 113.700 ;
        RECT 239.600 113.600 240.400 113.700 ;
        RECT 257.200 114.300 258.000 114.400 ;
        RECT 258.800 114.300 259.600 114.400 ;
        RECT 268.400 114.300 269.200 114.400 ;
        RECT 257.200 113.700 269.200 114.300 ;
        RECT 257.200 113.600 258.000 113.700 ;
        RECT 258.800 113.600 259.600 113.700 ;
        RECT 268.400 113.600 269.200 113.700 ;
        RECT 308.400 114.300 309.200 114.400 ;
        RECT 322.800 114.300 323.600 114.400 ;
        RECT 329.200 114.300 330.000 114.400 ;
        RECT 308.400 113.700 330.000 114.300 ;
        RECT 308.400 113.600 309.200 113.700 ;
        RECT 322.800 113.600 323.600 113.700 ;
        RECT 329.200 113.600 330.000 113.700 ;
        RECT 410.800 114.300 411.600 114.400 ;
        RECT 479.600 114.300 480.400 114.400 ;
        RECT 526.000 114.300 526.800 114.400 ;
        RECT 410.800 113.700 526.800 114.300 ;
        RECT 410.800 113.600 411.600 113.700 ;
        RECT 479.600 113.600 480.400 113.700 ;
        RECT 526.000 113.600 526.800 113.700 ;
        RECT 550.000 114.300 550.800 114.400 ;
        RECT 561.200 114.300 562.000 114.400 ;
        RECT 550.000 113.700 562.000 114.300 ;
        RECT 550.000 113.600 550.800 113.700 ;
        RECT 561.200 113.600 562.000 113.700 ;
        RECT 583.600 114.300 584.400 114.400 ;
        RECT 590.000 114.300 590.800 114.400 ;
        RECT 583.600 113.700 590.800 114.300 ;
        RECT 583.600 113.600 584.400 113.700 ;
        RECT 590.000 113.600 590.800 113.700 ;
        RECT 617.200 114.300 618.000 114.400 ;
        RECT 625.200 114.300 626.000 114.400 ;
        RECT 617.200 113.700 626.000 114.300 ;
        RECT 617.200 113.600 618.000 113.700 ;
        RECT 625.200 113.600 626.000 113.700 ;
        RECT 628.400 114.300 629.200 114.400 ;
        RECT 634.800 114.300 635.600 114.400 ;
        RECT 628.400 113.700 635.600 114.300 ;
        RECT 628.400 113.600 629.200 113.700 ;
        RECT 634.800 113.600 635.600 113.700 ;
        RECT 652.400 114.300 653.200 114.400 ;
        RECT 657.200 114.300 658.000 114.400 ;
        RECT 652.400 113.700 658.000 114.300 ;
        RECT 652.400 113.600 653.200 113.700 ;
        RECT 657.200 113.600 658.000 113.700 ;
        RECT 2.800 112.300 3.600 112.400 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 2.800 111.700 6.800 112.300 ;
        RECT 2.800 111.600 3.600 111.700 ;
        RECT 6.000 111.600 6.800 111.700 ;
        RECT 22.000 112.300 22.800 112.400 ;
        RECT 25.200 112.300 26.000 112.400 ;
        RECT 22.000 111.700 26.000 112.300 ;
        RECT 22.000 111.600 22.800 111.700 ;
        RECT 25.200 111.600 26.000 111.700 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 55.600 112.300 56.400 112.400 ;
        RECT 76.400 112.300 77.200 112.400 ;
        RECT 55.600 111.700 77.200 112.300 ;
        RECT 55.600 111.600 56.400 111.700 ;
        RECT 76.400 111.600 77.200 111.700 ;
        RECT 87.600 112.300 88.400 112.400 ;
        RECT 102.000 112.300 102.800 112.400 ;
        RECT 87.600 111.700 102.800 112.300 ;
        RECT 87.600 111.600 88.400 111.700 ;
        RECT 102.000 111.600 102.800 111.700 ;
        RECT 105.200 112.300 106.000 112.400 ;
        RECT 111.600 112.300 112.400 112.400 ;
        RECT 105.200 111.700 112.400 112.300 ;
        RECT 105.200 111.600 106.000 111.700 ;
        RECT 111.600 111.600 112.400 111.700 ;
        RECT 114.800 112.300 115.600 112.400 ;
        RECT 121.200 112.300 122.000 112.400 ;
        RECT 114.800 111.700 122.000 112.300 ;
        RECT 114.800 111.600 115.600 111.700 ;
        RECT 121.200 111.600 122.000 111.700 ;
        RECT 126.000 112.300 126.800 112.400 ;
        RECT 127.600 112.300 128.400 112.400 ;
        RECT 148.400 112.300 149.200 112.400 ;
        RECT 126.000 111.700 149.200 112.300 ;
        RECT 126.000 111.600 126.800 111.700 ;
        RECT 127.600 111.600 128.400 111.700 ;
        RECT 148.400 111.600 149.200 111.700 ;
        RECT 174.000 112.300 174.800 112.400 ;
        RECT 178.800 112.300 179.600 112.400 ;
        RECT 174.000 111.700 179.600 112.300 ;
        RECT 174.000 111.600 174.800 111.700 ;
        RECT 178.800 111.600 179.600 111.700 ;
        RECT 190.000 111.600 190.800 112.400 ;
        RECT 193.200 112.300 194.000 112.400 ;
        RECT 196.400 112.300 197.200 112.400 ;
        RECT 193.200 111.700 197.200 112.300 ;
        RECT 193.200 111.600 194.000 111.700 ;
        RECT 196.400 111.600 197.200 111.700 ;
        RECT 207.600 112.300 208.400 112.400 ;
        RECT 222.000 112.300 222.800 112.400 ;
        RECT 207.600 111.700 222.800 112.300 ;
        RECT 207.600 111.600 208.400 111.700 ;
        RECT 222.000 111.600 222.800 111.700 ;
        RECT 239.600 112.300 240.400 112.400 ;
        RECT 249.200 112.300 250.000 112.400 ;
        RECT 239.600 111.700 250.000 112.300 ;
        RECT 239.600 111.600 240.400 111.700 ;
        RECT 249.200 111.600 250.000 111.700 ;
        RECT 321.200 112.300 322.000 112.400 ;
        RECT 326.000 112.300 326.800 112.400 ;
        RECT 321.200 111.700 326.800 112.300 ;
        RECT 321.200 111.600 322.000 111.700 ;
        RECT 326.000 111.600 326.800 111.700 ;
        RECT 463.600 112.300 464.400 112.400 ;
        RECT 519.600 112.300 520.400 112.400 ;
        RECT 521.200 112.300 522.000 112.400 ;
        RECT 463.600 111.700 522.000 112.300 ;
        RECT 463.600 111.600 464.400 111.700 ;
        RECT 519.600 111.600 520.400 111.700 ;
        RECT 521.200 111.600 522.000 111.700 ;
        RECT 526.000 112.300 526.800 112.400 ;
        RECT 542.000 112.300 542.800 112.400 ;
        RECT 526.000 111.700 542.800 112.300 ;
        RECT 526.000 111.600 526.800 111.700 ;
        RECT 542.000 111.600 542.800 111.700 ;
        RECT 543.600 112.300 544.400 112.400 ;
        RECT 551.600 112.300 552.400 112.400 ;
        RECT 543.600 111.700 552.400 112.300 ;
        RECT 543.600 111.600 544.400 111.700 ;
        RECT 551.600 111.600 552.400 111.700 ;
        RECT 553.200 112.300 554.000 112.400 ;
        RECT 558.000 112.300 558.800 112.400 ;
        RECT 553.200 111.700 558.800 112.300 ;
        RECT 553.200 111.600 554.000 111.700 ;
        RECT 558.000 111.600 558.800 111.700 ;
        RECT 562.800 112.300 563.600 112.400 ;
        RECT 580.400 112.300 581.200 112.400 ;
        RECT 601.200 112.300 602.000 112.400 ;
        RECT 666.800 112.300 667.600 112.400 ;
        RECT 679.600 112.300 680.400 112.400 ;
        RECT 562.800 111.700 680.400 112.300 ;
        RECT 562.800 111.600 563.600 111.700 ;
        RECT 580.400 111.600 581.200 111.700 ;
        RECT 601.200 111.600 602.000 111.700 ;
        RECT 666.800 111.600 667.600 111.700 ;
        RECT 679.600 111.600 680.400 111.700 ;
        RECT 15.600 110.300 16.400 110.400 ;
        RECT 26.800 110.300 27.600 110.400 ;
        RECT 33.200 110.300 34.000 110.400 ;
        RECT 60.400 110.300 61.200 110.400 ;
        RECT 15.600 109.700 61.200 110.300 ;
        RECT 15.600 109.600 16.400 109.700 ;
        RECT 26.800 109.600 27.600 109.700 ;
        RECT 33.200 109.600 34.000 109.700 ;
        RECT 60.400 109.600 61.200 109.700 ;
        RECT 66.800 110.300 67.600 110.400 ;
        RECT 71.600 110.300 72.400 110.400 ;
        RECT 66.800 109.700 72.400 110.300 ;
        RECT 66.800 109.600 67.600 109.700 ;
        RECT 71.600 109.600 72.400 109.700 ;
        RECT 95.600 110.300 96.400 110.400 ;
        RECT 102.000 110.300 102.800 110.400 ;
        RECT 95.600 109.700 102.800 110.300 ;
        RECT 95.600 109.600 96.400 109.700 ;
        RECT 102.000 109.600 102.800 109.700 ;
        RECT 106.800 110.300 107.600 110.400 ;
        RECT 124.400 110.300 125.200 110.400 ;
        RECT 106.800 109.700 125.200 110.300 ;
        RECT 106.800 109.600 107.600 109.700 ;
        RECT 124.400 109.600 125.200 109.700 ;
        RECT 138.800 110.300 139.600 110.400 ;
        RECT 146.800 110.300 147.600 110.400 ;
        RECT 138.800 109.700 147.600 110.300 ;
        RECT 138.800 109.600 139.600 109.700 ;
        RECT 146.800 109.600 147.600 109.700 ;
        RECT 150.000 110.300 150.800 110.400 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 150.000 109.700 157.200 110.300 ;
        RECT 150.000 109.600 150.800 109.700 ;
        RECT 156.400 109.600 157.200 109.700 ;
        RECT 175.600 110.300 176.400 110.400 ;
        RECT 193.200 110.300 194.000 110.400 ;
        RECT 199.600 110.300 200.400 110.400 ;
        RECT 175.600 109.700 200.400 110.300 ;
        RECT 175.600 109.600 176.400 109.700 ;
        RECT 193.200 109.600 194.000 109.700 ;
        RECT 199.600 109.600 200.400 109.700 ;
        RECT 202.800 110.300 203.600 110.400 ;
        RECT 217.200 110.300 218.000 110.400 ;
        RECT 202.800 109.700 218.000 110.300 ;
        RECT 202.800 109.600 203.600 109.700 ;
        RECT 217.200 109.600 218.000 109.700 ;
        RECT 218.800 110.300 219.600 110.400 ;
        RECT 226.800 110.300 227.600 110.400 ;
        RECT 218.800 109.700 227.600 110.300 ;
        RECT 218.800 109.600 219.600 109.700 ;
        RECT 226.800 109.600 227.600 109.700 ;
        RECT 302.000 110.300 302.800 110.400 ;
        RECT 305.200 110.300 306.000 110.400 ;
        RECT 308.400 110.300 309.200 110.400 ;
        RECT 302.000 109.700 309.200 110.300 ;
        RECT 302.000 109.600 302.800 109.700 ;
        RECT 305.200 109.600 306.000 109.700 ;
        RECT 308.400 109.600 309.200 109.700 ;
        RECT 369.200 110.300 370.000 110.400 ;
        RECT 372.400 110.300 373.200 110.400 ;
        RECT 369.200 109.700 373.200 110.300 ;
        RECT 369.200 109.600 370.000 109.700 ;
        RECT 372.400 109.600 373.200 109.700 ;
        RECT 399.600 110.300 400.400 110.400 ;
        RECT 406.000 110.300 406.800 110.400 ;
        RECT 426.800 110.300 427.600 110.400 ;
        RECT 399.600 109.700 427.600 110.300 ;
        RECT 399.600 109.600 400.400 109.700 ;
        RECT 406.000 109.600 406.800 109.700 ;
        RECT 426.800 109.600 427.600 109.700 ;
        RECT 454.000 110.300 454.800 110.400 ;
        RECT 458.800 110.300 459.600 110.400 ;
        RECT 454.000 109.700 459.600 110.300 ;
        RECT 454.000 109.600 454.800 109.700 ;
        RECT 458.800 109.600 459.600 109.700 ;
        RECT 511.600 110.300 512.400 110.400 ;
        RECT 516.400 110.300 517.200 110.400 ;
        RECT 511.600 109.700 517.200 110.300 ;
        RECT 511.600 109.600 512.400 109.700 ;
        RECT 516.400 109.600 517.200 109.700 ;
        RECT 537.200 110.300 538.000 110.400 ;
        RECT 583.600 110.300 584.400 110.400 ;
        RECT 537.200 109.700 584.400 110.300 ;
        RECT 537.200 109.600 538.000 109.700 ;
        RECT 583.600 109.600 584.400 109.700 ;
        RECT 586.800 110.300 587.600 110.400 ;
        RECT 591.600 110.300 592.400 110.400 ;
        RECT 586.800 109.700 592.400 110.300 ;
        RECT 586.800 109.600 587.600 109.700 ;
        RECT 591.600 109.600 592.400 109.700 ;
        RECT 634.800 109.600 635.600 110.400 ;
        RECT 647.600 110.300 648.400 110.400 ;
        RECT 660.400 110.300 661.200 110.400 ;
        RECT 647.600 109.700 661.200 110.300 ;
        RECT 647.600 109.600 648.400 109.700 ;
        RECT 660.400 109.600 661.200 109.700 ;
        RECT 678.000 110.300 678.800 110.400 ;
        RECT 681.200 110.300 682.000 110.400 ;
        RECT 687.600 110.300 688.400 110.400 ;
        RECT 678.000 109.700 688.400 110.300 ;
        RECT 678.000 109.600 678.800 109.700 ;
        RECT 681.200 109.600 682.000 109.700 ;
        RECT 687.600 109.600 688.400 109.700 ;
        RECT 25.200 108.300 26.000 108.400 ;
        RECT 42.800 108.300 43.600 108.400 ;
        RECT 25.200 107.700 43.600 108.300 ;
        RECT 25.200 107.600 26.000 107.700 ;
        RECT 42.800 107.600 43.600 107.700 ;
        RECT 47.600 108.300 48.400 108.400 ;
        RECT 50.800 108.300 51.600 108.400 ;
        RECT 70.000 108.300 70.800 108.400 ;
        RECT 47.600 107.700 51.600 108.300 ;
        RECT 47.600 107.600 48.400 107.700 ;
        RECT 50.800 107.600 51.600 107.700 ;
        RECT 68.500 107.700 70.800 108.300 ;
        RECT 34.800 106.300 35.600 106.400 ;
        RECT 68.500 106.300 69.100 107.700 ;
        RECT 70.000 107.600 70.800 107.700 ;
        RECT 87.600 108.300 88.400 108.400 ;
        RECT 153.200 108.300 154.000 108.400 ;
        RECT 87.600 107.700 154.000 108.300 ;
        RECT 87.600 107.600 88.400 107.700 ;
        RECT 153.200 107.600 154.000 107.700 ;
        RECT 172.400 108.300 173.200 108.400 ;
        RECT 188.400 108.300 189.200 108.400 ;
        RECT 172.400 107.700 189.200 108.300 ;
        RECT 172.400 107.600 173.200 107.700 ;
        RECT 188.400 107.600 189.200 107.700 ;
        RECT 193.200 108.300 194.000 108.400 ;
        RECT 201.200 108.300 202.000 108.400 ;
        RECT 238.000 108.300 238.800 108.400 ;
        RECT 193.200 107.700 238.800 108.300 ;
        RECT 193.200 107.600 194.000 107.700 ;
        RECT 201.200 107.600 202.000 107.700 ;
        RECT 238.000 107.600 238.800 107.700 ;
        RECT 266.800 108.300 267.600 108.400 ;
        RECT 287.600 108.300 288.400 108.400 ;
        RECT 266.800 107.700 288.400 108.300 ;
        RECT 266.800 107.600 267.600 107.700 ;
        RECT 287.600 107.600 288.400 107.700 ;
        RECT 311.600 108.300 312.400 108.400 ;
        RECT 316.400 108.300 317.200 108.400 ;
        RECT 311.600 107.700 317.200 108.300 ;
        RECT 311.600 107.600 312.400 107.700 ;
        RECT 316.400 107.600 317.200 107.700 ;
        RECT 327.600 108.300 328.400 108.400 ;
        RECT 348.400 108.300 349.200 108.400 ;
        RECT 327.600 107.700 349.200 108.300 ;
        RECT 327.600 107.600 328.400 107.700 ;
        RECT 348.400 107.600 349.200 107.700 ;
        RECT 383.600 108.300 384.400 108.400 ;
        RECT 398.000 108.300 398.800 108.400 ;
        RECT 383.600 107.700 398.800 108.300 ;
        RECT 383.600 107.600 384.400 107.700 ;
        RECT 398.000 107.600 398.800 107.700 ;
        RECT 402.800 108.300 403.600 108.400 ;
        RECT 407.600 108.300 408.400 108.400 ;
        RECT 402.800 107.700 408.400 108.300 ;
        RECT 402.800 107.600 403.600 107.700 ;
        RECT 407.600 107.600 408.400 107.700 ;
        RECT 417.200 108.300 418.000 108.400 ;
        RECT 430.000 108.300 430.800 108.400 ;
        RECT 417.200 107.700 430.800 108.300 ;
        RECT 417.200 107.600 418.000 107.700 ;
        RECT 430.000 107.600 430.800 107.700 ;
        RECT 450.800 108.300 451.600 108.400 ;
        RECT 466.800 108.300 467.600 108.400 ;
        RECT 450.800 107.700 467.600 108.300 ;
        RECT 450.800 107.600 451.600 107.700 ;
        RECT 466.800 107.600 467.600 107.700 ;
        RECT 470.000 108.300 470.800 108.400 ;
        RECT 476.400 108.300 477.200 108.400 ;
        RECT 470.000 107.700 477.200 108.300 ;
        RECT 470.000 107.600 470.800 107.700 ;
        RECT 476.400 107.600 477.200 107.700 ;
        RECT 481.200 108.300 482.000 108.400 ;
        RECT 502.000 108.300 502.800 108.400 ;
        RECT 481.200 107.700 502.800 108.300 ;
        RECT 481.200 107.600 482.000 107.700 ;
        RECT 502.000 107.600 502.800 107.700 ;
        RECT 532.400 108.300 533.200 108.400 ;
        RECT 542.000 108.300 542.800 108.400 ;
        RECT 532.400 107.700 542.800 108.300 ;
        RECT 532.400 107.600 533.200 107.700 ;
        RECT 542.000 107.600 542.800 107.700 ;
        RECT 545.200 108.300 546.000 108.400 ;
        RECT 553.200 108.300 554.000 108.400 ;
        RECT 545.200 107.700 554.000 108.300 ;
        RECT 545.200 107.600 546.000 107.700 ;
        RECT 553.200 107.600 554.000 107.700 ;
        RECT 554.800 108.300 555.600 108.400 ;
        RECT 559.600 108.300 560.400 108.400 ;
        RECT 574.000 108.300 574.800 108.400 ;
        RECT 585.200 108.300 586.000 108.400 ;
        RECT 594.800 108.300 595.600 108.400 ;
        RECT 554.800 107.700 595.600 108.300 ;
        RECT 554.800 107.600 555.600 107.700 ;
        RECT 559.600 107.600 560.400 107.700 ;
        RECT 574.000 107.600 574.800 107.700 ;
        RECT 585.200 107.600 586.000 107.700 ;
        RECT 594.800 107.600 595.600 107.700 ;
        RECT 599.600 108.300 600.400 108.400 ;
        RECT 630.000 108.300 630.800 108.400 ;
        RECT 599.600 107.700 630.800 108.300 ;
        RECT 599.600 107.600 600.400 107.700 ;
        RECT 630.000 107.600 630.800 107.700 ;
        RECT 634.800 108.300 635.600 108.400 ;
        RECT 673.200 108.300 674.000 108.400 ;
        RECT 634.800 107.700 674.000 108.300 ;
        RECT 634.800 107.600 635.600 107.700 ;
        RECT 673.200 107.600 674.000 107.700 ;
        RECT 34.800 105.700 69.100 106.300 ;
        RECT 34.800 105.600 35.600 105.700 ;
        RECT 1.200 104.300 2.000 104.400 ;
        RECT 6.000 104.300 6.800 104.400 ;
        RECT 1.200 103.700 6.800 104.300 ;
        RECT 68.500 104.300 69.100 105.700 ;
        RECT 70.000 106.300 70.800 106.400 ;
        RECT 79.600 106.300 80.400 106.400 ;
        RECT 100.400 106.300 101.200 106.400 ;
        RECT 70.000 105.700 101.200 106.300 ;
        RECT 70.000 105.600 70.800 105.700 ;
        RECT 79.600 105.600 80.400 105.700 ;
        RECT 100.400 105.600 101.200 105.700 ;
        RECT 102.000 106.300 102.800 106.400 ;
        RECT 103.600 106.300 104.400 106.400 ;
        RECT 102.000 105.700 104.400 106.300 ;
        RECT 102.000 105.600 102.800 105.700 ;
        RECT 103.600 105.600 104.400 105.700 ;
        RECT 134.000 106.300 134.800 106.400 ;
        RECT 180.400 106.300 181.200 106.400 ;
        RECT 134.000 105.700 181.200 106.300 ;
        RECT 134.000 105.600 134.800 105.700 ;
        RECT 180.400 105.600 181.200 105.700 ;
        RECT 186.800 106.300 187.600 106.400 ;
        RECT 194.800 106.300 195.600 106.400 ;
        RECT 186.800 105.700 195.600 106.300 ;
        RECT 186.800 105.600 187.600 105.700 ;
        RECT 194.800 105.600 195.600 105.700 ;
        RECT 217.200 106.300 218.000 106.400 ;
        RECT 220.400 106.300 221.200 106.400 ;
        RECT 225.200 106.300 226.000 106.400 ;
        RECT 255.600 106.300 256.400 106.400 ;
        RECT 217.200 105.700 256.400 106.300 ;
        RECT 217.200 105.600 218.000 105.700 ;
        RECT 220.400 105.600 221.200 105.700 ;
        RECT 225.200 105.600 226.000 105.700 ;
        RECT 255.600 105.600 256.400 105.700 ;
        RECT 284.400 106.300 285.200 106.400 ;
        RECT 324.400 106.300 325.200 106.400 ;
        RECT 345.200 106.300 346.000 106.400 ;
        RECT 361.200 106.300 362.000 106.400 ;
        RECT 380.400 106.300 381.200 106.400 ;
        RECT 383.600 106.300 384.400 106.400 ;
        RECT 284.400 105.700 384.400 106.300 ;
        RECT 284.400 105.600 285.200 105.700 ;
        RECT 324.400 105.600 325.200 105.700 ;
        RECT 345.200 105.600 346.000 105.700 ;
        RECT 361.200 105.600 362.000 105.700 ;
        RECT 380.400 105.600 381.200 105.700 ;
        RECT 383.600 105.600 384.400 105.700 ;
        RECT 425.200 106.300 426.000 106.400 ;
        RECT 441.200 106.300 442.000 106.400 ;
        RECT 457.200 106.300 458.000 106.400 ;
        RECT 484.400 106.300 485.200 106.400 ;
        RECT 498.800 106.300 499.600 106.400 ;
        RECT 529.200 106.300 530.000 106.400 ;
        RECT 425.200 105.700 530.000 106.300 ;
        RECT 425.200 105.600 426.000 105.700 ;
        RECT 441.200 105.600 442.000 105.700 ;
        RECT 457.200 105.600 458.000 105.700 ;
        RECT 484.400 105.600 485.200 105.700 ;
        RECT 498.800 105.600 499.600 105.700 ;
        RECT 529.200 105.600 530.000 105.700 ;
        RECT 588.400 106.300 589.200 106.400 ;
        RECT 612.400 106.300 613.200 106.400 ;
        RECT 588.400 105.700 613.200 106.300 ;
        RECT 588.400 105.600 589.200 105.700 ;
        RECT 612.400 105.600 613.200 105.700 ;
        RECT 623.600 106.300 624.400 106.400 ;
        RECT 638.000 106.300 638.800 106.400 ;
        RECT 647.600 106.300 648.400 106.400 ;
        RECT 623.600 105.700 648.400 106.300 ;
        RECT 623.600 105.600 624.400 105.700 ;
        RECT 638.000 105.600 638.800 105.700 ;
        RECT 647.600 105.600 648.400 105.700 ;
        RECT 126.000 104.300 126.800 104.400 ;
        RECT 137.200 104.300 138.000 104.400 ;
        RECT 68.500 103.700 138.000 104.300 ;
        RECT 1.200 103.600 2.000 103.700 ;
        RECT 6.000 103.600 6.800 103.700 ;
        RECT 126.000 103.600 126.800 103.700 ;
        RECT 137.200 103.600 138.000 103.700 ;
        RECT 143.600 104.300 144.400 104.400 ;
        RECT 158.000 104.300 158.800 104.400 ;
        RECT 231.600 104.300 232.400 104.400 ;
        RECT 242.800 104.300 243.600 104.400 ;
        RECT 143.600 103.700 158.800 104.300 ;
        RECT 143.600 103.600 144.400 103.700 ;
        RECT 158.000 103.600 158.800 103.700 ;
        RECT 225.300 103.700 243.600 104.300 ;
        RECT 225.300 102.400 225.900 103.700 ;
        RECT 231.600 103.600 232.400 103.700 ;
        RECT 242.800 103.600 243.600 103.700 ;
        RECT 524.400 104.300 525.200 104.400 ;
        RECT 546.800 104.300 547.600 104.400 ;
        RECT 562.800 104.300 563.600 104.400 ;
        RECT 577.200 104.300 578.000 104.400 ;
        RECT 583.600 104.300 584.400 104.400 ;
        RECT 524.400 103.700 584.400 104.300 ;
        RECT 524.400 103.600 525.200 103.700 ;
        RECT 546.800 103.600 547.600 103.700 ;
        RECT 562.800 103.600 563.600 103.700 ;
        RECT 577.200 103.600 578.000 103.700 ;
        RECT 583.600 103.600 584.400 103.700 ;
        RECT 590.000 104.300 590.800 104.400 ;
        RECT 601.200 104.300 602.000 104.400 ;
        RECT 590.000 103.700 602.000 104.300 ;
        RECT 590.000 103.600 590.800 103.700 ;
        RECT 601.200 103.600 602.000 103.700 ;
        RECT 630.000 104.300 630.800 104.400 ;
        RECT 681.200 104.300 682.000 104.400 ;
        RECT 630.000 103.700 682.000 104.300 ;
        RECT 630.000 103.600 630.800 103.700 ;
        RECT 681.200 103.600 682.000 103.700 ;
        RECT 42.800 102.300 43.600 102.400 ;
        RECT 94.000 102.300 94.800 102.400 ;
        RECT 98.800 102.300 99.600 102.400 ;
        RECT 42.800 101.700 99.600 102.300 ;
        RECT 42.800 101.600 43.600 101.700 ;
        RECT 94.000 101.600 94.800 101.700 ;
        RECT 98.800 101.600 99.600 101.700 ;
        RECT 100.400 102.300 101.200 102.400 ;
        RECT 121.200 102.300 122.000 102.400 ;
        RECT 145.200 102.300 146.000 102.400 ;
        RECT 225.200 102.300 226.000 102.400 ;
        RECT 100.400 101.700 226.000 102.300 ;
        RECT 100.400 101.600 101.200 101.700 ;
        RECT 121.200 101.600 122.000 101.700 ;
        RECT 145.200 101.600 146.000 101.700 ;
        RECT 225.200 101.600 226.000 101.700 ;
        RECT 230.000 102.300 230.800 102.400 ;
        RECT 233.200 102.300 234.000 102.400 ;
        RECT 230.000 101.700 234.000 102.300 ;
        RECT 230.000 101.600 230.800 101.700 ;
        RECT 233.200 101.600 234.000 101.700 ;
        RECT 292.400 102.300 293.200 102.400 ;
        RECT 295.600 102.300 296.400 102.400 ;
        RECT 316.400 102.300 317.200 102.400 ;
        RECT 292.400 101.700 317.200 102.300 ;
        RECT 292.400 101.600 293.200 101.700 ;
        RECT 295.600 101.600 296.400 101.700 ;
        RECT 316.400 101.600 317.200 101.700 ;
        RECT 506.800 102.300 507.600 102.400 ;
        RECT 548.400 102.300 549.200 102.400 ;
        RECT 556.400 102.300 557.200 102.400 ;
        RECT 506.800 101.700 557.200 102.300 ;
        RECT 506.800 101.600 507.600 101.700 ;
        RECT 548.400 101.600 549.200 101.700 ;
        RECT 556.400 101.600 557.200 101.700 ;
        RECT 610.800 102.300 611.600 102.400 ;
        RECT 615.600 102.300 616.400 102.400 ;
        RECT 610.800 101.700 616.400 102.300 ;
        RECT 610.800 101.600 611.600 101.700 ;
        RECT 615.600 101.600 616.400 101.700 ;
        RECT 31.600 100.300 32.400 100.400 ;
        RECT 42.800 100.300 43.600 100.400 ;
        RECT 31.600 99.700 43.600 100.300 ;
        RECT 31.600 99.600 32.400 99.700 ;
        RECT 42.800 99.600 43.600 99.700 ;
        RECT 79.600 100.300 80.400 100.400 ;
        RECT 127.600 100.300 128.400 100.400 ;
        RECT 79.600 99.700 128.400 100.300 ;
        RECT 79.600 99.600 80.400 99.700 ;
        RECT 127.600 99.600 128.400 99.700 ;
        RECT 223.600 100.300 224.400 100.400 ;
        RECT 239.600 100.300 240.400 100.400 ;
        RECT 223.600 99.700 240.400 100.300 ;
        RECT 223.600 99.600 224.400 99.700 ;
        RECT 239.600 99.600 240.400 99.700 ;
        RECT 358.000 100.300 358.800 100.400 ;
        RECT 364.400 100.300 365.200 100.400 ;
        RECT 358.000 99.700 365.200 100.300 ;
        RECT 358.000 99.600 358.800 99.700 ;
        RECT 364.400 99.600 365.200 99.700 ;
        RECT 430.000 100.300 430.800 100.400 ;
        RECT 452.400 100.300 453.200 100.400 ;
        RECT 460.400 100.300 461.200 100.400 ;
        RECT 465.200 100.300 466.000 100.400 ;
        RECT 430.000 99.700 466.000 100.300 ;
        RECT 430.000 99.600 430.800 99.700 ;
        RECT 452.400 99.600 453.200 99.700 ;
        RECT 460.400 99.600 461.200 99.700 ;
        RECT 465.200 99.600 466.000 99.700 ;
        RECT 490.800 100.300 491.600 100.400 ;
        RECT 495.600 100.300 496.400 100.400 ;
        RECT 490.800 99.700 496.400 100.300 ;
        RECT 490.800 99.600 491.600 99.700 ;
        RECT 495.600 99.600 496.400 99.700 ;
        RECT 609.200 100.300 610.000 100.400 ;
        RECT 622.000 100.300 622.800 100.400 ;
        RECT 609.200 99.700 622.800 100.300 ;
        RECT 609.200 99.600 610.000 99.700 ;
        RECT 622.000 99.600 622.800 99.700 ;
        RECT 641.200 100.300 642.000 100.400 ;
        RECT 642.800 100.300 643.600 100.400 ;
        RECT 641.200 99.700 643.600 100.300 ;
        RECT 641.200 99.600 642.000 99.700 ;
        RECT 642.800 99.600 643.600 99.700 ;
        RECT 682.800 99.600 683.600 100.400 ;
        RECT 26.800 98.300 27.600 98.400 ;
        RECT 38.000 98.300 38.800 98.400 ;
        RECT 26.800 97.700 38.800 98.300 ;
        RECT 26.800 97.600 27.600 97.700 ;
        RECT 38.000 97.600 38.800 97.700 ;
        RECT 42.800 98.300 43.600 98.400 ;
        RECT 46.000 98.300 46.800 98.400 ;
        RECT 42.800 97.700 46.800 98.300 ;
        RECT 42.800 97.600 43.600 97.700 ;
        RECT 46.000 97.600 46.800 97.700 ;
        RECT 52.400 98.300 53.200 98.400 ;
        RECT 58.800 98.300 59.600 98.400 ;
        RECT 52.400 97.700 59.600 98.300 ;
        RECT 52.400 97.600 53.200 97.700 ;
        RECT 58.800 97.600 59.600 97.700 ;
        RECT 110.000 98.300 110.800 98.400 ;
        RECT 130.800 98.300 131.600 98.400 ;
        RECT 178.800 98.300 179.600 98.400 ;
        RECT 110.000 97.700 179.600 98.300 ;
        RECT 110.000 97.600 110.800 97.700 ;
        RECT 130.800 97.600 131.600 97.700 ;
        RECT 178.800 97.600 179.600 97.700 ;
        RECT 428.400 98.300 429.200 98.400 ;
        RECT 450.800 98.300 451.600 98.400 ;
        RECT 428.400 97.700 451.600 98.300 ;
        RECT 428.400 97.600 429.200 97.700 ;
        RECT 450.800 97.600 451.600 97.700 ;
        RECT 465.200 98.300 466.000 98.400 ;
        RECT 471.600 98.300 472.400 98.400 ;
        RECT 465.200 97.700 472.400 98.300 ;
        RECT 465.200 97.600 466.000 97.700 ;
        RECT 471.600 97.600 472.400 97.700 ;
        RECT 473.200 98.300 474.000 98.400 ;
        RECT 518.000 98.300 518.800 98.400 ;
        RECT 473.200 97.700 518.800 98.300 ;
        RECT 473.200 97.600 474.000 97.700 ;
        RECT 518.000 97.600 518.800 97.700 ;
        RECT 583.600 98.300 584.400 98.400 ;
        RECT 604.400 98.300 605.200 98.400 ;
        RECT 625.200 98.300 626.000 98.400 ;
        RECT 583.600 97.700 626.000 98.300 ;
        RECT 642.900 98.300 643.500 99.600 ;
        RECT 686.000 98.300 686.800 98.400 ;
        RECT 642.900 97.700 686.800 98.300 ;
        RECT 583.600 97.600 584.400 97.700 ;
        RECT 604.400 97.600 605.200 97.700 ;
        RECT 625.200 97.600 626.000 97.700 ;
        RECT 686.000 97.600 686.800 97.700 ;
        RECT 22.000 96.300 22.800 96.400 ;
        RECT 36.400 96.300 37.200 96.400 ;
        RECT 22.000 95.700 37.200 96.300 ;
        RECT 22.000 95.600 22.800 95.700 ;
        RECT 36.400 95.600 37.200 95.700 ;
        RECT 47.600 96.300 48.400 96.400 ;
        RECT 65.200 96.300 66.000 96.400 ;
        RECT 71.600 96.300 72.400 96.400 ;
        RECT 90.800 96.300 91.600 96.400 ;
        RECT 47.600 95.700 91.600 96.300 ;
        RECT 47.600 95.600 48.400 95.700 ;
        RECT 65.200 95.600 66.000 95.700 ;
        RECT 71.600 95.600 72.400 95.700 ;
        RECT 90.800 95.600 91.600 95.700 ;
        RECT 100.400 96.300 101.200 96.400 ;
        RECT 118.000 96.300 118.800 96.400 ;
        RECT 100.400 95.700 118.800 96.300 ;
        RECT 100.400 95.600 101.200 95.700 ;
        RECT 118.000 95.600 118.800 95.700 ;
        RECT 137.200 96.300 138.000 96.400 ;
        RECT 175.600 96.300 176.400 96.400 ;
        RECT 137.200 95.700 176.400 96.300 ;
        RECT 137.200 95.600 138.000 95.700 ;
        RECT 175.600 95.600 176.400 95.700 ;
        RECT 210.800 96.300 211.600 96.400 ;
        RECT 217.200 96.300 218.000 96.400 ;
        RECT 231.600 96.300 232.400 96.400 ;
        RECT 238.000 96.300 238.800 96.400 ;
        RECT 210.800 95.700 238.800 96.300 ;
        RECT 210.800 95.600 211.600 95.700 ;
        RECT 217.200 95.600 218.000 95.700 ;
        RECT 231.600 95.600 232.400 95.700 ;
        RECT 238.000 95.600 238.800 95.700 ;
        RECT 295.600 96.300 296.400 96.400 ;
        RECT 311.600 96.300 312.400 96.400 ;
        RECT 342.000 96.300 342.800 96.400 ;
        RECT 295.600 95.700 342.800 96.300 ;
        RECT 295.600 95.600 296.400 95.700 ;
        RECT 311.600 95.600 312.400 95.700 ;
        RECT 342.000 95.600 342.800 95.700 ;
        RECT 390.000 96.300 390.800 96.400 ;
        RECT 428.400 96.300 429.200 96.400 ;
        RECT 390.000 95.700 429.200 96.300 ;
        RECT 390.000 95.600 390.800 95.700 ;
        RECT 428.400 95.600 429.200 95.700 ;
        RECT 457.200 96.300 458.000 96.400 ;
        RECT 458.800 96.300 459.600 96.400 ;
        RECT 457.200 95.700 459.600 96.300 ;
        RECT 457.200 95.600 458.000 95.700 ;
        RECT 458.800 95.600 459.600 95.700 ;
        RECT 474.800 96.300 475.600 96.400 ;
        RECT 487.600 96.300 488.400 96.400 ;
        RECT 474.800 95.700 488.400 96.300 ;
        RECT 474.800 95.600 475.600 95.700 ;
        RECT 487.600 95.600 488.400 95.700 ;
        RECT 503.600 95.600 504.400 96.400 ;
        RECT 535.600 95.600 536.400 96.400 ;
        RECT 564.400 96.300 565.200 96.400 ;
        RECT 575.600 96.300 576.400 96.400 ;
        RECT 564.400 95.700 576.400 96.300 ;
        RECT 564.400 95.600 565.200 95.700 ;
        RECT 575.600 95.600 576.400 95.700 ;
        RECT 580.400 96.300 581.200 96.400 ;
        RECT 583.600 96.300 584.400 96.400 ;
        RECT 580.400 95.700 584.400 96.300 ;
        RECT 580.400 95.600 581.200 95.700 ;
        RECT 583.600 95.600 584.400 95.700 ;
        RECT 599.600 96.300 600.400 96.400 ;
        RECT 612.400 96.300 613.200 96.400 ;
        RECT 657.200 96.300 658.000 96.400 ;
        RECT 658.800 96.300 659.600 96.400 ;
        RECT 599.600 95.700 651.500 96.300 ;
        RECT 599.600 95.600 600.400 95.700 ;
        RECT 612.400 95.600 613.200 95.700 ;
        RECT 650.900 94.400 651.500 95.700 ;
        RECT 657.200 95.700 659.600 96.300 ;
        RECT 657.200 95.600 658.000 95.700 ;
        RECT 658.800 95.600 659.600 95.700 ;
        RECT 9.200 94.300 10.000 94.400 ;
        RECT 23.600 94.300 24.400 94.400 ;
        RECT 9.200 93.700 24.400 94.300 ;
        RECT 9.200 93.600 10.000 93.700 ;
        RECT 23.600 93.600 24.400 93.700 ;
        RECT 30.000 93.600 30.800 94.400 ;
        RECT 54.000 94.300 54.800 94.400 ;
        RECT 63.600 94.300 64.400 94.400 ;
        RECT 54.000 93.700 64.400 94.300 ;
        RECT 54.000 93.600 54.800 93.700 ;
        RECT 63.600 93.600 64.400 93.700 ;
        RECT 97.200 94.300 98.000 94.400 ;
        RECT 134.000 94.300 134.800 94.400 ;
        RECT 97.200 93.700 134.800 94.300 ;
        RECT 97.200 93.600 98.000 93.700 ;
        RECT 134.000 93.600 134.800 93.700 ;
        RECT 135.600 94.300 136.400 94.400 ;
        RECT 143.600 94.300 144.400 94.400 ;
        RECT 135.600 93.700 144.400 94.300 ;
        RECT 135.600 93.600 136.400 93.700 ;
        RECT 143.600 93.600 144.400 93.700 ;
        RECT 146.800 94.300 147.600 94.400 ;
        RECT 172.400 94.300 173.200 94.400 ;
        RECT 146.800 93.700 173.200 94.300 ;
        RECT 146.800 93.600 147.600 93.700 ;
        RECT 172.400 93.600 173.200 93.700 ;
        RECT 196.400 94.300 197.200 94.400 ;
        RECT 204.400 94.300 205.200 94.400 ;
        RECT 196.400 93.700 205.200 94.300 ;
        RECT 196.400 93.600 197.200 93.700 ;
        RECT 204.400 93.600 205.200 93.700 ;
        RECT 247.600 93.600 248.400 94.400 ;
        RECT 249.200 94.300 250.000 94.400 ;
        RECT 274.800 94.300 275.600 94.400 ;
        RECT 249.200 93.700 275.600 94.300 ;
        RECT 249.200 93.600 250.000 93.700 ;
        RECT 274.800 93.600 275.600 93.700 ;
        RECT 305.200 94.300 306.000 94.400 ;
        RECT 327.600 94.300 328.400 94.400 ;
        RECT 305.200 93.700 328.400 94.300 ;
        RECT 305.200 93.600 306.000 93.700 ;
        RECT 327.600 93.600 328.400 93.700 ;
        RECT 380.400 94.300 381.200 94.400 ;
        RECT 391.600 94.300 392.400 94.400 ;
        RECT 380.400 93.700 392.400 94.300 ;
        RECT 380.400 93.600 381.200 93.700 ;
        RECT 391.600 93.600 392.400 93.700 ;
        RECT 412.400 94.300 413.200 94.400 ;
        RECT 442.800 94.300 443.600 94.400 ;
        RECT 412.400 93.700 443.600 94.300 ;
        RECT 412.400 93.600 413.200 93.700 ;
        RECT 442.800 93.600 443.600 93.700 ;
        RECT 458.800 94.300 459.600 94.400 ;
        RECT 502.000 94.300 502.800 94.400 ;
        RECT 508.400 94.300 509.200 94.400 ;
        RECT 510.000 94.300 510.800 94.400 ;
        RECT 518.000 94.300 518.800 94.400 ;
        RECT 458.800 93.700 518.800 94.300 ;
        RECT 458.800 93.600 459.600 93.700 ;
        RECT 502.000 93.600 502.800 93.700 ;
        RECT 508.400 93.600 509.200 93.700 ;
        RECT 510.000 93.600 510.800 93.700 ;
        RECT 518.000 93.600 518.800 93.700 ;
        RECT 561.200 94.300 562.000 94.400 ;
        RECT 567.600 94.300 568.400 94.400 ;
        RECT 561.200 93.700 568.400 94.300 ;
        RECT 561.200 93.600 562.000 93.700 ;
        RECT 567.600 93.600 568.400 93.700 ;
        RECT 618.800 94.300 619.600 94.400 ;
        RECT 623.600 94.300 624.400 94.400 ;
        RECT 618.800 93.700 624.400 94.300 ;
        RECT 618.800 93.600 619.600 93.700 ;
        RECT 623.600 93.600 624.400 93.700 ;
        RECT 630.000 94.300 630.800 94.400 ;
        RECT 636.400 94.300 637.200 94.400 ;
        RECT 644.400 94.300 645.200 94.400 ;
        RECT 630.000 93.700 645.200 94.300 ;
        RECT 630.000 93.600 630.800 93.700 ;
        RECT 636.400 93.600 637.200 93.700 ;
        RECT 644.400 93.600 645.200 93.700 ;
        RECT 650.800 94.300 651.600 94.400 ;
        RECT 657.200 94.300 658.000 94.400 ;
        RECT 650.800 93.700 658.000 94.300 ;
        RECT 650.800 93.600 651.600 93.700 ;
        RECT 657.200 93.600 658.000 93.700 ;
        RECT 1.200 92.300 2.000 92.400 ;
        RECT 17.200 92.300 18.000 92.400 ;
        RECT 1.200 91.700 18.000 92.300 ;
        RECT 1.200 91.600 2.000 91.700 ;
        RECT 17.200 91.600 18.000 91.700 ;
        RECT 20.400 92.300 21.200 92.400 ;
        RECT 38.000 92.300 38.800 92.400 ;
        RECT 41.200 92.300 42.000 92.400 ;
        RECT 20.400 91.700 42.000 92.300 ;
        RECT 20.400 91.600 21.200 91.700 ;
        RECT 38.000 91.600 38.800 91.700 ;
        RECT 41.200 91.600 42.000 91.700 ;
        RECT 54.000 92.300 54.800 92.400 ;
        RECT 68.400 92.300 69.200 92.400 ;
        RECT 54.000 91.700 69.200 92.300 ;
        RECT 54.000 91.600 54.800 91.700 ;
        RECT 68.400 91.600 69.200 91.700 ;
        RECT 92.400 92.300 93.200 92.400 ;
        RECT 103.600 92.300 104.400 92.400 ;
        RECT 135.600 92.300 136.400 92.400 ;
        RECT 145.200 92.300 146.000 92.400 ;
        RECT 92.400 91.700 102.700 92.300 ;
        RECT 92.400 91.600 93.200 91.700 ;
        RECT 14.000 90.300 14.800 90.400 ;
        RECT 17.200 90.300 18.000 90.400 ;
        RECT 100.400 90.300 101.200 90.400 ;
        RECT 14.000 89.700 101.200 90.300 ;
        RECT 102.100 90.300 102.700 91.700 ;
        RECT 103.600 91.700 146.000 92.300 ;
        RECT 103.600 91.600 104.400 91.700 ;
        RECT 135.600 91.600 136.400 91.700 ;
        RECT 145.200 91.600 146.000 91.700 ;
        RECT 162.800 92.300 163.600 92.400 ;
        RECT 193.200 92.300 194.000 92.400 ;
        RECT 162.800 91.700 194.000 92.300 ;
        RECT 162.800 91.600 163.600 91.700 ;
        RECT 193.200 91.600 194.000 91.700 ;
        RECT 382.000 92.300 382.800 92.400 ;
        RECT 393.200 92.300 394.000 92.400 ;
        RECT 382.000 91.700 394.000 92.300 ;
        RECT 382.000 91.600 382.800 91.700 ;
        RECT 393.200 91.600 394.000 91.700 ;
        RECT 394.800 92.300 395.600 92.400 ;
        RECT 401.200 92.300 402.000 92.400 ;
        RECT 450.800 92.300 451.600 92.400 ;
        RECT 460.400 92.300 461.200 92.400 ;
        RECT 394.800 91.700 411.500 92.300 ;
        RECT 394.800 91.600 395.600 91.700 ;
        RECT 401.200 91.600 402.000 91.700 ;
        RECT 111.600 90.300 112.400 90.400 ;
        RECT 102.100 89.700 112.400 90.300 ;
        RECT 14.000 89.600 14.800 89.700 ;
        RECT 17.200 89.600 18.000 89.700 ;
        RECT 100.400 89.600 101.200 89.700 ;
        RECT 111.600 89.600 112.400 89.700 ;
        RECT 122.800 90.300 123.600 90.400 ;
        RECT 134.000 90.300 134.800 90.400 ;
        RECT 122.800 89.700 134.800 90.300 ;
        RECT 122.800 89.600 123.600 89.700 ;
        RECT 134.000 89.600 134.800 89.700 ;
        RECT 143.600 90.300 144.400 90.400 ;
        RECT 156.400 90.300 157.200 90.400 ;
        RECT 143.600 89.700 157.200 90.300 ;
        RECT 143.600 89.600 144.400 89.700 ;
        RECT 156.400 89.600 157.200 89.700 ;
        RECT 302.000 90.300 302.800 90.400 ;
        RECT 308.400 90.300 309.200 90.400 ;
        RECT 302.000 89.700 309.200 90.300 ;
        RECT 302.000 89.600 302.800 89.700 ;
        RECT 308.400 89.600 309.200 89.700 ;
        RECT 386.800 90.300 387.600 90.400 ;
        RECT 404.400 90.300 405.200 90.400 ;
        RECT 409.200 90.300 410.000 90.400 ;
        RECT 386.800 89.700 410.000 90.300 ;
        RECT 410.900 90.300 411.500 91.700 ;
        RECT 450.800 91.700 461.200 92.300 ;
        RECT 450.800 91.600 451.600 91.700 ;
        RECT 460.400 91.600 461.200 91.700 ;
        RECT 551.600 92.300 552.400 92.400 ;
        RECT 564.400 92.300 565.200 92.400 ;
        RECT 572.400 92.300 573.200 92.400 ;
        RECT 551.600 91.700 573.200 92.300 ;
        RECT 551.600 91.600 552.400 91.700 ;
        RECT 564.400 91.600 565.200 91.700 ;
        RECT 572.400 91.600 573.200 91.700 ;
        RECT 574.000 92.300 574.800 92.400 ;
        RECT 602.800 92.300 603.600 92.400 ;
        RECT 574.000 91.700 603.600 92.300 ;
        RECT 574.000 91.600 574.800 91.700 ;
        RECT 602.800 91.600 603.600 91.700 ;
        RECT 610.800 92.300 611.600 92.400 ;
        RECT 620.400 92.300 621.200 92.400 ;
        RECT 610.800 91.700 621.200 92.300 ;
        RECT 610.800 91.600 611.600 91.700 ;
        RECT 620.400 91.600 621.200 91.700 ;
        RECT 630.000 92.300 630.800 92.400 ;
        RECT 634.800 92.300 635.600 92.400 ;
        RECT 630.000 91.700 635.600 92.300 ;
        RECT 630.000 91.600 630.800 91.700 ;
        RECT 634.800 91.600 635.600 91.700 ;
        RECT 636.400 92.300 637.200 92.400 ;
        RECT 646.000 92.300 646.800 92.400 ;
        RECT 636.400 91.700 646.800 92.300 ;
        RECT 636.400 91.600 637.200 91.700 ;
        RECT 646.000 91.600 646.800 91.700 ;
        RECT 535.600 90.300 536.400 90.400 ;
        RECT 410.900 89.700 536.400 90.300 ;
        RECT 386.800 89.600 387.600 89.700 ;
        RECT 404.400 89.600 405.200 89.700 ;
        RECT 409.200 89.600 410.000 89.700 ;
        RECT 535.600 89.600 536.400 89.700 ;
        RECT 537.200 90.300 538.000 90.400 ;
        RECT 553.200 90.300 554.000 90.400 ;
        RECT 537.200 89.700 554.000 90.300 ;
        RECT 537.200 89.600 538.000 89.700 ;
        RECT 553.200 89.600 554.000 89.700 ;
        RECT 559.600 90.300 560.400 90.400 ;
        RECT 562.800 90.300 563.600 90.400 ;
        RECT 559.600 89.700 563.600 90.300 ;
        RECT 559.600 89.600 560.400 89.700 ;
        RECT 562.800 89.600 563.600 89.700 ;
        RECT 596.400 90.300 597.200 90.400 ;
        RECT 620.400 90.300 621.200 90.400 ;
        RECT 596.400 89.700 621.200 90.300 ;
        RECT 596.400 89.600 597.200 89.700 ;
        RECT 620.400 89.600 621.200 89.700 ;
        RECT 23.600 88.300 24.400 88.400 ;
        RECT 39.600 88.300 40.400 88.400 ;
        RECT 23.600 87.700 40.400 88.300 ;
        RECT 23.600 87.600 24.400 87.700 ;
        RECT 39.600 87.600 40.400 87.700 ;
        RECT 52.400 88.300 53.200 88.400 ;
        RECT 82.800 88.300 83.600 88.400 ;
        RECT 52.400 87.700 83.600 88.300 ;
        RECT 52.400 87.600 53.200 87.700 ;
        RECT 82.800 87.600 83.600 87.700 ;
        RECT 92.400 88.300 93.200 88.400 ;
        RECT 97.200 88.300 98.000 88.400 ;
        RECT 92.400 87.700 98.000 88.300 ;
        RECT 92.400 87.600 93.200 87.700 ;
        RECT 97.200 87.600 98.000 87.700 ;
        RECT 130.800 88.300 131.600 88.400 ;
        RECT 138.800 88.300 139.600 88.400 ;
        RECT 130.800 87.700 139.600 88.300 ;
        RECT 130.800 87.600 131.600 87.700 ;
        RECT 138.800 87.600 139.600 87.700 ;
        RECT 148.400 88.300 149.200 88.400 ;
        RECT 174.000 88.300 174.800 88.400 ;
        RECT 183.600 88.300 184.400 88.400 ;
        RECT 148.400 87.700 184.400 88.300 ;
        RECT 148.400 87.600 149.200 87.700 ;
        RECT 174.000 87.600 174.800 87.700 ;
        RECT 183.600 87.600 184.400 87.700 ;
        RECT 438.000 88.300 438.800 88.400 ;
        RECT 439.600 88.300 440.400 88.400 ;
        RECT 476.400 88.300 477.200 88.400 ;
        RECT 438.000 87.700 477.200 88.300 ;
        RECT 438.000 87.600 438.800 87.700 ;
        RECT 439.600 87.600 440.400 87.700 ;
        RECT 476.400 87.600 477.200 87.700 ;
        RECT 527.600 88.300 528.400 88.400 ;
        RECT 553.200 88.300 554.000 88.400 ;
        RECT 527.600 87.700 554.000 88.300 ;
        RECT 527.600 87.600 528.400 87.700 ;
        RECT 553.200 87.600 554.000 87.700 ;
        RECT 617.200 88.300 618.000 88.400 ;
        RECT 670.000 88.300 670.800 88.400 ;
        RECT 617.200 87.700 670.800 88.300 ;
        RECT 617.200 87.600 618.000 87.700 ;
        RECT 670.000 87.600 670.800 87.700 ;
        RECT 26.800 86.300 27.600 86.400 ;
        RECT 50.800 86.300 51.600 86.400 ;
        RECT 57.200 86.300 58.000 86.400 ;
        RECT 26.800 85.700 58.000 86.300 ;
        RECT 26.800 85.600 27.600 85.700 ;
        RECT 50.800 85.600 51.600 85.700 ;
        RECT 57.200 85.600 58.000 85.700 ;
        RECT 58.800 86.300 59.600 86.400 ;
        RECT 129.200 86.300 130.000 86.400 ;
        RECT 132.400 86.300 133.200 86.400 ;
        RECT 177.200 86.300 178.000 86.400 ;
        RECT 182.000 86.300 182.800 86.400 ;
        RECT 58.800 85.700 182.800 86.300 ;
        RECT 58.800 85.600 59.600 85.700 ;
        RECT 129.200 85.600 130.000 85.700 ;
        RECT 132.400 85.600 133.200 85.700 ;
        RECT 177.200 85.600 178.000 85.700 ;
        RECT 182.000 85.600 182.800 85.700 ;
        RECT 522.800 86.300 523.600 86.400 ;
        RECT 567.600 86.300 568.400 86.400 ;
        RECT 522.800 85.700 568.400 86.300 ;
        RECT 522.800 85.600 523.600 85.700 ;
        RECT 567.600 85.600 568.400 85.700 ;
        RECT 41.200 84.300 42.000 84.400 ;
        RECT 55.600 84.300 56.400 84.400 ;
        RECT 86.000 84.300 86.800 84.400 ;
        RECT 90.800 84.300 91.600 84.400 ;
        RECT 41.200 83.700 91.600 84.300 ;
        RECT 41.200 83.600 42.000 83.700 ;
        RECT 55.600 83.600 56.400 83.700 ;
        RECT 86.000 83.600 86.800 83.700 ;
        RECT 90.800 83.600 91.600 83.700 ;
        RECT 110.000 84.300 110.800 84.400 ;
        RECT 127.600 84.300 128.400 84.400 ;
        RECT 110.000 83.700 128.400 84.300 ;
        RECT 110.000 83.600 110.800 83.700 ;
        RECT 127.600 83.600 128.400 83.700 ;
        RECT 129.200 84.300 130.000 84.400 ;
        RECT 135.600 84.300 136.400 84.400 ;
        RECT 129.200 83.700 136.400 84.300 ;
        RECT 129.200 83.600 130.000 83.700 ;
        RECT 135.600 83.600 136.400 83.700 ;
        RECT 138.800 84.300 139.600 84.400 ;
        RECT 169.200 84.300 170.000 84.400 ;
        RECT 138.800 83.700 170.000 84.300 ;
        RECT 138.800 83.600 139.600 83.700 ;
        RECT 169.200 83.600 170.000 83.700 ;
        RECT 238.000 84.300 238.800 84.400 ;
        RECT 249.200 84.300 250.000 84.400 ;
        RECT 238.000 83.700 250.000 84.300 ;
        RECT 238.000 83.600 238.800 83.700 ;
        RECT 249.200 83.600 250.000 83.700 ;
        RECT 457.200 84.300 458.000 84.400 ;
        RECT 641.200 84.300 642.000 84.400 ;
        RECT 457.200 83.700 642.000 84.300 ;
        RECT 457.200 83.600 458.000 83.700 ;
        RECT 641.200 83.600 642.000 83.700 ;
        RECT 676.400 84.300 677.200 84.400 ;
        RECT 682.800 84.300 683.600 84.400 ;
        RECT 676.400 83.700 683.600 84.300 ;
        RECT 676.400 83.600 677.200 83.700 ;
        RECT 682.800 83.600 683.600 83.700 ;
        RECT 87.600 82.300 88.400 82.400 ;
        RECT 97.200 82.300 98.000 82.400 ;
        RECT 87.600 81.700 98.000 82.300 ;
        RECT 87.600 81.600 88.400 81.700 ;
        RECT 97.200 81.600 98.000 81.700 ;
        RECT 143.600 82.300 144.400 82.400 ;
        RECT 150.000 82.300 150.800 82.400 ;
        RECT 143.600 81.700 150.800 82.300 ;
        RECT 143.600 81.600 144.400 81.700 ;
        RECT 150.000 81.600 150.800 81.700 ;
        RECT 175.600 82.300 176.400 82.400 ;
        RECT 186.800 82.300 187.600 82.400 ;
        RECT 305.200 82.300 306.000 82.400 ;
        RECT 321.200 82.300 322.000 82.400 ;
        RECT 175.600 81.700 187.600 82.300 ;
        RECT 175.600 81.600 176.400 81.700 ;
        RECT 186.800 81.600 187.600 81.700 ;
        RECT 257.300 81.700 322.000 82.300 ;
        RECT 127.600 80.300 128.400 80.400 ;
        RECT 154.800 80.300 155.600 80.400 ;
        RECT 127.600 79.700 155.600 80.300 ;
        RECT 127.600 79.600 128.400 79.700 ;
        RECT 154.800 79.600 155.600 79.700 ;
        RECT 162.800 80.300 163.600 80.400 ;
        RECT 257.300 80.300 257.900 81.700 ;
        RECT 305.200 81.600 306.000 81.700 ;
        RECT 321.200 81.600 322.000 81.700 ;
        RECT 446.000 82.300 446.800 82.400 ;
        RECT 556.400 82.300 557.200 82.400 ;
        RECT 446.000 81.700 557.200 82.300 ;
        RECT 446.000 81.600 446.800 81.700 ;
        RECT 556.400 81.600 557.200 81.700 ;
        RECT 567.600 82.300 568.400 82.400 ;
        RECT 569.200 82.300 570.000 82.400 ;
        RECT 567.600 81.700 570.000 82.300 ;
        RECT 567.600 81.600 568.400 81.700 ;
        RECT 569.200 81.600 570.000 81.700 ;
        RECT 572.400 82.300 573.200 82.400 ;
        RECT 590.000 82.300 590.800 82.400 ;
        RECT 572.400 81.700 590.800 82.300 ;
        RECT 572.400 81.600 573.200 81.700 ;
        RECT 590.000 81.600 590.800 81.700 ;
        RECT 162.800 79.700 257.900 80.300 ;
        RECT 258.800 80.300 259.600 80.400 ;
        RECT 260.400 80.300 261.200 80.400 ;
        RECT 258.800 79.700 261.200 80.300 ;
        RECT 162.800 79.600 163.600 79.700 ;
        RECT 258.800 79.600 259.600 79.700 ;
        RECT 260.400 79.600 261.200 79.700 ;
        RECT 271.600 80.300 272.400 80.400 ;
        RECT 278.000 80.300 278.800 80.400 ;
        RECT 271.600 79.700 278.800 80.300 ;
        RECT 271.600 79.600 272.400 79.700 ;
        RECT 278.000 79.600 278.800 79.700 ;
        RECT 558.000 80.300 558.800 80.400 ;
        RECT 617.200 80.300 618.000 80.400 ;
        RECT 558.000 79.700 618.000 80.300 ;
        RECT 558.000 79.600 558.800 79.700 ;
        RECT 617.200 79.600 618.000 79.700 ;
        RECT 142.000 77.600 142.800 78.400 ;
        RECT 238.000 78.300 238.800 78.400 ;
        RECT 268.400 78.300 269.200 78.400 ;
        RECT 238.000 77.700 269.200 78.300 ;
        RECT 238.000 77.600 238.800 77.700 ;
        RECT 268.400 77.600 269.200 77.700 ;
        RECT 556.400 78.300 557.200 78.400 ;
        RECT 582.000 78.300 582.800 78.400 ;
        RECT 556.400 77.700 582.800 78.300 ;
        RECT 556.400 77.600 557.200 77.700 ;
        RECT 582.000 77.600 582.800 77.700 ;
        RECT 622.000 78.300 622.800 78.400 ;
        RECT 633.200 78.300 634.000 78.400 ;
        RECT 622.000 77.700 634.000 78.300 ;
        RECT 622.000 77.600 622.800 77.700 ;
        RECT 633.200 77.600 634.000 77.700 ;
        RECT 663.600 78.300 664.400 78.400 ;
        RECT 666.800 78.300 667.600 78.400 ;
        RECT 663.600 77.700 667.600 78.300 ;
        RECT 663.600 77.600 664.400 77.700 ;
        RECT 666.800 77.600 667.600 77.700 ;
        RECT 86.000 76.300 86.800 76.400 ;
        RECT 140.400 76.300 141.200 76.400 ;
        RECT 86.000 75.700 141.200 76.300 ;
        RECT 86.000 75.600 86.800 75.700 ;
        RECT 140.400 75.600 141.200 75.700 ;
        RECT 172.400 76.300 173.200 76.400 ;
        RECT 175.600 76.300 176.400 76.400 ;
        RECT 172.400 75.700 176.400 76.300 ;
        RECT 172.400 75.600 173.200 75.700 ;
        RECT 175.600 75.600 176.400 75.700 ;
        RECT 260.400 76.300 261.200 76.400 ;
        RECT 263.600 76.300 264.400 76.400 ;
        RECT 260.400 75.700 264.400 76.300 ;
        RECT 260.400 75.600 261.200 75.700 ;
        RECT 263.600 75.600 264.400 75.700 ;
        RECT 542.000 76.300 542.800 76.400 ;
        RECT 580.400 76.300 581.200 76.400 ;
        RECT 542.000 75.700 581.200 76.300 ;
        RECT 542.000 75.600 542.800 75.700 ;
        RECT 580.400 75.600 581.200 75.700 ;
        RECT 582.000 76.300 582.800 76.400 ;
        RECT 586.800 76.300 587.600 76.400 ;
        RECT 612.400 76.300 613.200 76.400 ;
        RECT 625.200 76.300 626.000 76.400 ;
        RECT 582.000 75.700 626.000 76.300 ;
        RECT 582.000 75.600 582.800 75.700 ;
        RECT 586.800 75.600 587.600 75.700 ;
        RECT 612.400 75.600 613.200 75.700 ;
        RECT 625.200 75.600 626.000 75.700 ;
        RECT 670.000 76.300 670.800 76.400 ;
        RECT 684.400 76.300 685.200 76.400 ;
        RECT 670.000 75.700 685.200 76.300 ;
        RECT 670.000 75.600 670.800 75.700 ;
        RECT 684.400 75.600 685.200 75.700 ;
        RECT 142.000 74.300 142.800 74.400 ;
        RECT 156.400 74.300 157.200 74.400 ;
        RECT 34.900 73.700 142.800 74.300 ;
        RECT 34.900 72.400 35.500 73.700 ;
        RECT 142.000 73.600 142.800 73.700 ;
        RECT 145.300 73.700 157.200 74.300 ;
        RECT 18.800 72.300 19.600 72.400 ;
        RECT 25.200 72.300 26.000 72.400 ;
        RECT 34.800 72.300 35.600 72.400 ;
        RECT 18.800 71.700 35.600 72.300 ;
        RECT 18.800 71.600 19.600 71.700 ;
        RECT 25.200 71.600 26.000 71.700 ;
        RECT 34.800 71.600 35.600 71.700 ;
        RECT 38.000 72.300 38.800 72.400 ;
        RECT 42.800 72.300 43.600 72.400 ;
        RECT 38.000 71.700 43.600 72.300 ;
        RECT 38.000 71.600 38.800 71.700 ;
        RECT 42.800 71.600 43.600 71.700 ;
        RECT 46.000 72.300 46.800 72.400 ;
        RECT 73.200 72.300 74.000 72.400 ;
        RECT 46.000 71.700 74.000 72.300 ;
        RECT 46.000 71.600 46.800 71.700 ;
        RECT 73.200 71.600 74.000 71.700 ;
        RECT 90.800 72.300 91.600 72.400 ;
        RECT 94.000 72.300 94.800 72.400 ;
        RECT 126.000 72.300 126.800 72.400 ;
        RECT 90.800 71.700 126.800 72.300 ;
        RECT 90.800 71.600 91.600 71.700 ;
        RECT 94.000 71.600 94.800 71.700 ;
        RECT 126.000 71.600 126.800 71.700 ;
        RECT 132.400 72.300 133.200 72.400 ;
        RECT 145.300 72.300 145.900 73.700 ;
        RECT 156.400 73.600 157.200 73.700 ;
        RECT 169.200 74.300 170.000 74.400 ;
        RECT 231.600 74.300 232.400 74.400 ;
        RECT 290.800 74.300 291.600 74.400 ;
        RECT 169.200 73.700 291.600 74.300 ;
        RECT 169.200 73.600 170.000 73.700 ;
        RECT 231.600 73.600 232.400 73.700 ;
        RECT 290.800 73.600 291.600 73.700 ;
        RECT 300.400 74.300 301.200 74.400 ;
        RECT 314.800 74.300 315.600 74.400 ;
        RECT 334.000 74.300 334.800 74.400 ;
        RECT 300.400 73.700 334.800 74.300 ;
        RECT 300.400 73.600 301.200 73.700 ;
        RECT 314.800 73.600 315.600 73.700 ;
        RECT 334.000 73.600 334.800 73.700 ;
        RECT 353.200 74.300 354.000 74.400 ;
        RECT 361.200 74.300 362.000 74.400 ;
        RECT 353.200 73.700 362.000 74.300 ;
        RECT 353.200 73.600 354.000 73.700 ;
        RECT 361.200 73.600 362.000 73.700 ;
        RECT 377.200 74.300 378.000 74.400 ;
        RECT 390.000 74.300 390.800 74.400 ;
        RECT 377.200 73.700 390.800 74.300 ;
        RECT 377.200 73.600 378.000 73.700 ;
        RECT 390.000 73.600 390.800 73.700 ;
        RECT 396.400 74.300 397.200 74.400 ;
        RECT 465.200 74.300 466.000 74.400 ;
        RECT 396.400 73.700 466.000 74.300 ;
        RECT 396.400 73.600 397.200 73.700 ;
        RECT 465.200 73.600 466.000 73.700 ;
        RECT 502.000 74.300 502.800 74.400 ;
        RECT 513.200 74.300 514.000 74.400 ;
        RECT 502.000 73.700 514.000 74.300 ;
        RECT 502.000 73.600 502.800 73.700 ;
        RECT 513.200 73.600 514.000 73.700 ;
        RECT 577.200 74.300 578.000 74.400 ;
        RECT 583.600 74.300 584.400 74.400 ;
        RECT 577.200 73.700 584.400 74.300 ;
        RECT 577.200 73.600 578.000 73.700 ;
        RECT 583.600 73.600 584.400 73.700 ;
        RECT 585.200 74.300 586.000 74.400 ;
        RECT 610.800 74.300 611.600 74.400 ;
        RECT 623.600 74.300 624.400 74.400 ;
        RECT 642.800 74.300 643.600 74.400 ;
        RECT 644.400 74.300 645.200 74.400 ;
        RECT 585.200 73.700 624.400 74.300 ;
        RECT 585.200 73.600 586.000 73.700 ;
        RECT 610.800 73.600 611.600 73.700 ;
        RECT 623.600 73.600 624.400 73.700 ;
        RECT 630.100 73.700 645.200 74.300 ;
        RECT 630.100 72.400 630.700 73.700 ;
        RECT 642.800 73.600 643.600 73.700 ;
        RECT 644.400 73.600 645.200 73.700 ;
        RECT 679.600 74.300 680.400 74.400 ;
        RECT 684.400 74.300 685.200 74.400 ;
        RECT 679.600 73.700 685.200 74.300 ;
        RECT 679.600 73.600 680.400 73.700 ;
        RECT 684.400 73.600 685.200 73.700 ;
        RECT 132.400 71.700 145.900 72.300 ;
        RECT 146.800 72.300 147.600 72.400 ;
        RECT 153.200 72.300 154.000 72.400 ;
        RECT 146.800 71.700 154.000 72.300 ;
        RECT 132.400 71.600 133.200 71.700 ;
        RECT 146.800 71.600 147.600 71.700 ;
        RECT 153.200 71.600 154.000 71.700 ;
        RECT 159.600 72.300 160.400 72.400 ;
        RECT 166.000 72.300 166.800 72.400 ;
        RECT 172.400 72.300 173.200 72.400 ;
        RECT 159.600 71.700 173.200 72.300 ;
        RECT 159.600 71.600 160.400 71.700 ;
        RECT 166.000 71.600 166.800 71.700 ;
        RECT 172.400 71.600 173.200 71.700 ;
        RECT 175.600 72.300 176.400 72.400 ;
        RECT 185.200 72.300 186.000 72.400 ;
        RECT 175.600 71.700 186.000 72.300 ;
        RECT 175.600 71.600 176.400 71.700 ;
        RECT 185.200 71.600 186.000 71.700 ;
        RECT 193.200 71.600 194.000 72.400 ;
        RECT 343.600 72.300 344.400 72.400 ;
        RECT 350.000 72.300 350.800 72.400 ;
        RECT 343.600 71.700 350.800 72.300 ;
        RECT 343.600 71.600 344.400 71.700 ;
        RECT 350.000 71.600 350.800 71.700 ;
        RECT 398.000 72.300 398.800 72.400 ;
        RECT 404.400 72.300 405.200 72.400 ;
        RECT 398.000 71.700 405.200 72.300 ;
        RECT 398.000 71.600 398.800 71.700 ;
        RECT 404.400 71.600 405.200 71.700 ;
        RECT 478.000 72.300 478.800 72.400 ;
        RECT 508.400 72.300 509.200 72.400 ;
        RECT 478.000 71.700 509.200 72.300 ;
        RECT 478.000 71.600 478.800 71.700 ;
        RECT 508.400 71.600 509.200 71.700 ;
        RECT 518.000 72.300 518.800 72.400 ;
        RECT 538.800 72.300 539.600 72.400 ;
        RECT 518.000 71.700 539.600 72.300 ;
        RECT 518.000 71.600 518.800 71.700 ;
        RECT 538.800 71.600 539.600 71.700 ;
        RECT 543.600 72.300 544.400 72.400 ;
        RECT 569.200 72.300 570.000 72.400 ;
        RECT 601.200 72.300 602.000 72.400 ;
        RECT 543.600 71.700 563.500 72.300 ;
        RECT 543.600 71.600 544.400 71.700 ;
        RECT 20.400 69.600 21.200 70.400 ;
        RECT 30.000 70.300 30.800 70.400 ;
        RECT 38.000 70.300 38.800 70.400 ;
        RECT 30.000 69.700 38.800 70.300 ;
        RECT 30.000 69.600 30.800 69.700 ;
        RECT 38.000 69.600 38.800 69.700 ;
        RECT 50.800 70.300 51.600 70.400 ;
        RECT 60.400 70.300 61.200 70.400 ;
        RECT 50.800 69.700 61.200 70.300 ;
        RECT 50.800 69.600 51.600 69.700 ;
        RECT 60.400 69.600 61.200 69.700 ;
        RECT 102.000 70.300 102.800 70.400 ;
        RECT 114.800 70.300 115.600 70.400 ;
        RECT 102.000 69.700 115.600 70.300 ;
        RECT 102.000 69.600 102.800 69.700 ;
        RECT 114.800 69.600 115.600 69.700 ;
        RECT 127.600 70.300 128.400 70.400 ;
        RECT 137.200 70.300 138.000 70.400 ;
        RECT 127.600 69.700 138.000 70.300 ;
        RECT 127.600 69.600 128.400 69.700 ;
        RECT 137.200 69.600 138.000 69.700 ;
        RECT 140.400 70.300 141.200 70.400 ;
        RECT 162.800 70.300 163.600 70.400 ;
        RECT 140.400 69.700 163.600 70.300 ;
        RECT 140.400 69.600 141.200 69.700 ;
        RECT 162.800 69.600 163.600 69.700 ;
        RECT 170.800 70.300 171.600 70.400 ;
        RECT 174.000 70.300 174.800 70.400 ;
        RECT 170.800 69.700 174.800 70.300 ;
        RECT 170.800 69.600 171.600 69.700 ;
        RECT 174.000 69.600 174.800 69.700 ;
        RECT 183.600 70.300 184.400 70.400 ;
        RECT 193.200 70.300 194.000 70.400 ;
        RECT 183.600 69.700 194.000 70.300 ;
        RECT 183.600 69.600 184.400 69.700 ;
        RECT 193.200 69.600 194.000 69.700 ;
        RECT 223.600 70.300 224.400 70.400 ;
        RECT 230.000 70.300 230.800 70.400 ;
        RECT 273.200 70.300 274.000 70.400 ;
        RECT 289.200 70.300 290.000 70.400 ;
        RECT 223.600 69.700 290.000 70.300 ;
        RECT 223.600 69.600 224.400 69.700 ;
        RECT 230.000 69.600 230.800 69.700 ;
        RECT 273.200 69.600 274.000 69.700 ;
        RECT 289.200 69.600 290.000 69.700 ;
        RECT 294.000 70.300 294.800 70.400 ;
        RECT 298.800 70.300 299.600 70.400 ;
        RECT 294.000 69.700 299.600 70.300 ;
        RECT 294.000 69.600 294.800 69.700 ;
        RECT 298.800 69.600 299.600 69.700 ;
        RECT 399.600 70.300 400.400 70.400 ;
        RECT 431.600 70.300 432.400 70.400 ;
        RECT 399.600 69.700 432.400 70.300 ;
        RECT 399.600 69.600 400.400 69.700 ;
        RECT 431.600 69.600 432.400 69.700 ;
        RECT 449.200 70.300 450.000 70.400 ;
        RECT 454.000 70.300 454.800 70.400 ;
        RECT 449.200 69.700 454.800 70.300 ;
        RECT 449.200 69.600 450.000 69.700 ;
        RECT 454.000 69.600 454.800 69.700 ;
        RECT 535.600 70.300 536.400 70.400 ;
        RECT 538.800 70.300 539.600 70.400 ;
        RECT 535.600 69.700 539.600 70.300 ;
        RECT 535.600 69.600 536.400 69.700 ;
        RECT 538.800 69.600 539.600 69.700 ;
        RECT 540.400 70.300 541.200 70.400 ;
        RECT 542.000 70.300 542.800 70.400 ;
        RECT 540.400 69.700 542.800 70.300 ;
        RECT 540.400 69.600 541.200 69.700 ;
        RECT 542.000 69.600 542.800 69.700 ;
        RECT 553.200 70.300 554.000 70.400 ;
        RECT 561.200 70.300 562.000 70.400 ;
        RECT 553.200 69.700 562.000 70.300 ;
        RECT 562.900 70.300 563.500 71.700 ;
        RECT 569.200 71.700 602.000 72.300 ;
        RECT 569.200 71.600 570.000 71.700 ;
        RECT 601.200 71.600 602.000 71.700 ;
        RECT 626.800 72.300 627.600 72.400 ;
        RECT 630.000 72.300 630.800 72.400 ;
        RECT 626.800 71.700 630.800 72.300 ;
        RECT 626.800 71.600 627.600 71.700 ;
        RECT 630.000 71.600 630.800 71.700 ;
        RECT 646.000 72.300 646.800 72.400 ;
        RECT 663.600 72.300 664.400 72.400 ;
        RECT 646.000 71.700 664.400 72.300 ;
        RECT 646.000 71.600 646.800 71.700 ;
        RECT 663.600 71.600 664.400 71.700 ;
        RECT 585.200 70.300 586.000 70.400 ;
        RECT 562.900 69.700 586.000 70.300 ;
        RECT 553.200 69.600 554.000 69.700 ;
        RECT 561.200 69.600 562.000 69.700 ;
        RECT 585.200 69.600 586.000 69.700 ;
        RECT 634.800 70.300 635.600 70.400 ;
        RECT 639.600 70.300 640.400 70.400 ;
        RECT 634.800 69.700 640.400 70.300 ;
        RECT 634.800 69.600 635.600 69.700 ;
        RECT 639.600 69.600 640.400 69.700 ;
        RECT 642.800 70.300 643.600 70.400 ;
        RECT 652.400 70.300 653.200 70.400 ;
        RECT 642.800 69.700 653.200 70.300 ;
        RECT 642.800 69.600 643.600 69.700 ;
        RECT 652.400 69.600 653.200 69.700 ;
        RECT 654.000 70.300 654.800 70.400 ;
        RECT 666.800 70.300 667.600 70.400 ;
        RECT 654.000 69.700 667.600 70.300 ;
        RECT 654.000 69.600 654.800 69.700 ;
        RECT 666.800 69.600 667.600 69.700 ;
        RECT 6.000 68.300 6.800 68.400 ;
        RECT 31.600 68.300 32.400 68.400 ;
        RECT 47.600 68.300 48.400 68.400 ;
        RECT 63.600 68.300 64.400 68.400 ;
        RECT 6.000 67.700 64.400 68.300 ;
        RECT 6.000 67.600 6.800 67.700 ;
        RECT 31.600 67.600 32.400 67.700 ;
        RECT 47.600 67.600 48.400 67.700 ;
        RECT 63.600 67.600 64.400 67.700 ;
        RECT 106.800 68.300 107.600 68.400 ;
        RECT 122.800 68.300 123.600 68.400 ;
        RECT 106.800 67.700 123.600 68.300 ;
        RECT 106.800 67.600 107.600 67.700 ;
        RECT 122.800 67.600 123.600 67.700 ;
        RECT 143.600 68.300 144.400 68.400 ;
        RECT 172.400 68.300 173.200 68.400 ;
        RECT 202.800 68.300 203.600 68.400 ;
        RECT 143.600 67.700 171.500 68.300 ;
        RECT 143.600 67.600 144.400 67.700 ;
        RECT 170.900 66.400 171.500 67.700 ;
        RECT 172.400 67.700 203.600 68.300 ;
        RECT 172.400 67.600 173.200 67.700 ;
        RECT 202.800 67.600 203.600 67.700 ;
        RECT 204.400 68.300 205.200 68.400 ;
        RECT 212.400 68.300 213.200 68.400 ;
        RECT 289.200 68.300 290.000 68.400 ;
        RECT 204.400 67.700 290.000 68.300 ;
        RECT 204.400 67.600 205.200 67.700 ;
        RECT 212.400 67.600 213.200 67.700 ;
        RECT 289.200 67.600 290.000 67.700 ;
        RECT 295.600 68.300 296.400 68.400 ;
        RECT 306.800 68.300 307.600 68.400 ;
        RECT 295.600 67.700 307.600 68.300 ;
        RECT 295.600 67.600 296.400 67.700 ;
        RECT 306.800 67.600 307.600 67.700 ;
        RECT 532.400 68.300 533.200 68.400 ;
        RECT 671.600 68.300 672.400 68.400 ;
        RECT 673.200 68.300 674.000 68.400 ;
        RECT 532.400 67.700 674.000 68.300 ;
        RECT 532.400 67.600 533.200 67.700 ;
        RECT 671.600 67.600 672.400 67.700 ;
        RECT 673.200 67.600 674.000 67.700 ;
        RECT 9.200 66.300 10.000 66.400 ;
        RECT 26.800 66.300 27.600 66.400 ;
        RECT 9.200 65.700 27.600 66.300 ;
        RECT 9.200 65.600 10.000 65.700 ;
        RECT 26.800 65.600 27.600 65.700 ;
        RECT 113.200 66.300 114.000 66.400 ;
        RECT 132.400 66.300 133.200 66.400 ;
        RECT 113.200 65.700 133.200 66.300 ;
        RECT 113.200 65.600 114.000 65.700 ;
        RECT 132.400 65.600 133.200 65.700 ;
        RECT 153.200 66.300 154.000 66.400 ;
        RECT 161.200 66.300 162.000 66.400 ;
        RECT 153.200 65.700 162.000 66.300 ;
        RECT 153.200 65.600 154.000 65.700 ;
        RECT 161.200 65.600 162.000 65.700 ;
        RECT 170.800 66.300 171.600 66.400 ;
        RECT 180.400 66.300 181.200 66.400 ;
        RECT 190.000 66.300 190.800 66.400 ;
        RECT 191.600 66.300 192.400 66.400 ;
        RECT 170.800 65.700 192.400 66.300 ;
        RECT 170.800 65.600 171.600 65.700 ;
        RECT 180.400 65.600 181.200 65.700 ;
        RECT 190.000 65.600 190.800 65.700 ;
        RECT 191.600 65.600 192.400 65.700 ;
        RECT 206.000 66.300 206.800 66.400 ;
        RECT 226.800 66.300 227.600 66.400 ;
        RECT 239.600 66.300 240.400 66.400 ;
        RECT 206.000 65.700 240.400 66.300 ;
        RECT 206.000 65.600 206.800 65.700 ;
        RECT 226.800 65.600 227.600 65.700 ;
        RECT 239.600 65.600 240.400 65.700 ;
        RECT 249.200 66.300 250.000 66.400 ;
        RECT 252.400 66.300 253.200 66.400 ;
        RECT 249.200 65.700 253.200 66.300 ;
        RECT 249.200 65.600 250.000 65.700 ;
        RECT 252.400 65.600 253.200 65.700 ;
        RECT 292.400 66.300 293.200 66.400 ;
        RECT 314.800 66.300 315.600 66.400 ;
        RECT 292.400 65.700 315.600 66.300 ;
        RECT 292.400 65.600 293.200 65.700 ;
        RECT 314.800 65.600 315.600 65.700 ;
        RECT 462.000 66.300 462.800 66.400 ;
        RECT 468.400 66.300 469.200 66.400 ;
        RECT 462.000 65.700 469.200 66.300 ;
        RECT 462.000 65.600 462.800 65.700 ;
        RECT 468.400 65.600 469.200 65.700 ;
        RECT 497.200 66.300 498.000 66.400 ;
        RECT 503.600 66.300 504.400 66.400 ;
        RECT 511.600 66.300 512.400 66.400 ;
        RECT 497.200 65.700 512.400 66.300 ;
        RECT 497.200 65.600 498.000 65.700 ;
        RECT 503.600 65.600 504.400 65.700 ;
        RECT 511.600 65.600 512.400 65.700 ;
        RECT 558.000 65.600 558.800 66.400 ;
        RECT 567.600 66.300 568.400 66.400 ;
        RECT 602.800 66.300 603.600 66.400 ;
        RECT 567.600 65.700 603.600 66.300 ;
        RECT 567.600 65.600 568.400 65.700 ;
        RECT 602.800 65.600 603.600 65.700 ;
        RECT 654.000 66.300 654.800 66.400 ;
        RECT 668.400 66.300 669.200 66.400 ;
        RECT 654.000 65.700 669.200 66.300 ;
        RECT 654.000 65.600 654.800 65.700 ;
        RECT 668.400 65.600 669.200 65.700 ;
        RECT 671.600 66.300 672.400 66.400 ;
        RECT 673.200 66.300 674.000 66.400 ;
        RECT 671.600 65.700 674.000 66.300 ;
        RECT 671.600 65.600 672.400 65.700 ;
        RECT 673.200 65.600 674.000 65.700 ;
        RECT 20.400 64.300 21.200 64.400 ;
        RECT 52.400 64.300 53.200 64.400 ;
        RECT 20.400 63.700 53.200 64.300 ;
        RECT 20.400 63.600 21.200 63.700 ;
        RECT 52.400 63.600 53.200 63.700 ;
        RECT 66.800 64.300 67.600 64.400 ;
        RECT 111.600 64.300 112.400 64.400 ;
        RECT 66.800 63.700 112.400 64.300 ;
        RECT 66.800 63.600 67.600 63.700 ;
        RECT 111.600 63.600 112.400 63.700 ;
        RECT 119.600 64.300 120.400 64.400 ;
        RECT 122.800 64.300 123.600 64.400 ;
        RECT 119.600 63.700 123.600 64.300 ;
        RECT 119.600 63.600 120.400 63.700 ;
        RECT 122.800 63.600 123.600 63.700 ;
        RECT 159.600 64.300 160.400 64.400 ;
        RECT 276.400 64.300 277.200 64.400 ;
        RECT 287.600 64.300 288.400 64.400 ;
        RECT 305.200 64.300 306.000 64.400 ;
        RECT 159.600 63.700 286.700 64.300 ;
        RECT 159.600 63.600 160.400 63.700 ;
        RECT 276.400 63.600 277.200 63.700 ;
        RECT 57.200 62.300 58.000 62.400 ;
        RECT 65.200 62.300 66.000 62.400 ;
        RECT 82.800 62.300 83.600 62.400 ;
        RECT 87.600 62.300 88.400 62.400 ;
        RECT 57.200 61.700 88.400 62.300 ;
        RECT 57.200 61.600 58.000 61.700 ;
        RECT 65.200 61.600 66.000 61.700 ;
        RECT 82.800 61.600 83.600 61.700 ;
        RECT 87.600 61.600 88.400 61.700 ;
        RECT 89.200 62.300 90.000 62.400 ;
        RECT 126.000 62.300 126.800 62.400 ;
        RECT 89.200 61.700 126.800 62.300 ;
        RECT 89.200 61.600 90.000 61.700 ;
        RECT 126.000 61.600 126.800 61.700 ;
        RECT 234.800 62.300 235.600 62.400 ;
        RECT 252.400 62.300 253.200 62.400 ;
        RECT 234.800 61.700 253.200 62.300 ;
        RECT 286.100 62.300 286.700 63.700 ;
        RECT 287.600 63.700 306.000 64.300 ;
        RECT 287.600 63.600 288.400 63.700 ;
        RECT 305.200 63.600 306.000 63.700 ;
        RECT 335.600 64.300 336.400 64.400 ;
        RECT 369.200 64.300 370.000 64.400 ;
        RECT 335.600 63.700 370.000 64.300 ;
        RECT 335.600 63.600 336.400 63.700 ;
        RECT 369.200 63.600 370.000 63.700 ;
        RECT 535.600 64.300 536.400 64.400 ;
        RECT 542.000 64.300 542.800 64.400 ;
        RECT 551.600 64.300 552.400 64.400 ;
        RECT 535.600 63.700 552.400 64.300 ;
        RECT 535.600 63.600 536.400 63.700 ;
        RECT 542.000 63.600 542.800 63.700 ;
        RECT 551.600 63.600 552.400 63.700 ;
        RECT 609.200 64.300 610.000 64.400 ;
        RECT 636.400 64.300 637.200 64.400 ;
        RECT 639.600 64.300 640.400 64.400 ;
        RECT 609.200 63.700 640.400 64.300 ;
        RECT 609.200 63.600 610.000 63.700 ;
        RECT 636.400 63.600 637.200 63.700 ;
        RECT 639.600 63.600 640.400 63.700 ;
        RECT 298.800 62.300 299.600 62.400 ;
        RECT 286.100 61.700 299.600 62.300 ;
        RECT 234.800 61.600 235.600 61.700 ;
        RECT 252.400 61.600 253.200 61.700 ;
        RECT 298.800 61.600 299.600 61.700 ;
        RECT 348.400 62.300 349.200 62.400 ;
        RECT 372.400 62.300 373.200 62.400 ;
        RECT 348.400 61.700 373.200 62.300 ;
        RECT 348.400 61.600 349.200 61.700 ;
        RECT 372.400 61.600 373.200 61.700 ;
        RECT 450.800 62.300 451.600 62.400 ;
        RECT 559.600 62.300 560.400 62.400 ;
        RECT 450.800 61.700 560.400 62.300 ;
        RECT 450.800 61.600 451.600 61.700 ;
        RECT 559.600 61.600 560.400 61.700 ;
        RECT 583.600 62.300 584.400 62.400 ;
        RECT 599.600 62.300 600.400 62.400 ;
        RECT 583.600 61.700 600.400 62.300 ;
        RECT 583.600 61.600 584.400 61.700 ;
        RECT 599.600 61.600 600.400 61.700 ;
        RECT 614.000 62.300 614.800 62.400 ;
        RECT 636.400 62.300 637.200 62.400 ;
        RECT 614.000 61.700 637.200 62.300 ;
        RECT 614.000 61.600 614.800 61.700 ;
        RECT 636.400 61.600 637.200 61.700 ;
        RECT 50.800 60.300 51.600 60.400 ;
        RECT 58.800 60.300 59.600 60.400 ;
        RECT 50.800 59.700 59.600 60.300 ;
        RECT 50.800 59.600 51.600 59.700 ;
        RECT 58.800 59.600 59.600 59.700 ;
        RECT 110.000 60.300 110.800 60.400 ;
        RECT 113.200 60.300 114.000 60.400 ;
        RECT 110.000 59.700 114.000 60.300 ;
        RECT 110.000 59.600 110.800 59.700 ;
        RECT 113.200 59.600 114.000 59.700 ;
        RECT 378.800 60.300 379.600 60.400 ;
        RECT 394.800 60.300 395.600 60.400 ;
        RECT 378.800 59.700 395.600 60.300 ;
        RECT 378.800 59.600 379.600 59.700 ;
        RECT 394.800 59.600 395.600 59.700 ;
        RECT 418.800 60.300 419.600 60.400 ;
        RECT 446.000 60.300 446.800 60.400 ;
        RECT 418.800 59.700 446.800 60.300 ;
        RECT 418.800 59.600 419.600 59.700 ;
        RECT 446.000 59.600 446.800 59.700 ;
        RECT 474.800 60.300 475.600 60.400 ;
        RECT 481.200 60.300 482.000 60.400 ;
        RECT 474.800 59.700 482.000 60.300 ;
        RECT 474.800 59.600 475.600 59.700 ;
        RECT 481.200 59.600 482.000 59.700 ;
        RECT 567.600 60.300 568.400 60.400 ;
        RECT 569.200 60.300 570.000 60.400 ;
        RECT 567.600 59.700 570.000 60.300 ;
        RECT 567.600 59.600 568.400 59.700 ;
        RECT 569.200 59.600 570.000 59.700 ;
        RECT 580.400 60.300 581.200 60.400 ;
        RECT 593.200 60.300 594.000 60.400 ;
        RECT 580.400 59.700 594.000 60.300 ;
        RECT 580.400 59.600 581.200 59.700 ;
        RECT 593.200 59.600 594.000 59.700 ;
        RECT 612.400 59.600 613.200 60.400 ;
        RECT 49.200 58.300 50.000 58.400 ;
        RECT 84.400 58.300 85.200 58.400 ;
        RECT 49.200 57.700 85.200 58.300 ;
        RECT 49.200 57.600 50.000 57.700 ;
        RECT 84.400 57.600 85.200 57.700 ;
        RECT 94.000 58.300 94.800 58.400 ;
        RECT 130.800 58.300 131.600 58.400 ;
        RECT 94.000 57.700 131.600 58.300 ;
        RECT 94.000 57.600 94.800 57.700 ;
        RECT 130.800 57.600 131.600 57.700 ;
        RECT 150.000 58.300 150.800 58.400 ;
        RECT 164.400 58.300 165.200 58.400 ;
        RECT 150.000 57.700 165.200 58.300 ;
        RECT 150.000 57.600 150.800 57.700 ;
        RECT 164.400 57.600 165.200 57.700 ;
        RECT 255.600 58.300 256.400 58.400 ;
        RECT 297.200 58.300 298.000 58.400 ;
        RECT 306.800 58.300 307.600 58.400 ;
        RECT 255.600 57.700 307.600 58.300 ;
        RECT 255.600 57.600 256.400 57.700 ;
        RECT 297.200 57.600 298.000 57.700 ;
        RECT 306.800 57.600 307.600 57.700 ;
        RECT 359.600 58.300 360.400 58.400 ;
        RECT 386.800 58.300 387.600 58.400 ;
        RECT 359.600 57.700 387.600 58.300 ;
        RECT 359.600 57.600 360.400 57.700 ;
        RECT 386.800 57.600 387.600 57.700 ;
        RECT 399.600 58.300 400.400 58.400 ;
        RECT 447.600 58.300 448.400 58.400 ;
        RECT 399.600 57.700 448.400 58.300 ;
        RECT 399.600 57.600 400.400 57.700 ;
        RECT 447.600 57.600 448.400 57.700 ;
        RECT 490.800 58.300 491.600 58.400 ;
        RECT 502.000 58.300 502.800 58.400 ;
        RECT 551.600 58.300 552.400 58.400 ;
        RECT 558.000 58.300 558.800 58.400 ;
        RECT 490.800 57.700 502.800 58.300 ;
        RECT 490.800 57.600 491.600 57.700 ;
        RECT 502.000 57.600 502.800 57.700 ;
        RECT 529.300 57.700 558.800 58.300 ;
        RECT 529.300 56.400 529.900 57.700 ;
        RECT 551.600 57.600 552.400 57.700 ;
        RECT 558.000 57.600 558.800 57.700 ;
        RECT 582.000 57.600 582.800 58.400 ;
        RECT 588.400 58.300 589.200 58.400 ;
        RECT 599.600 58.300 600.400 58.400 ;
        RECT 588.400 57.700 600.400 58.300 ;
        RECT 588.400 57.600 589.200 57.700 ;
        RECT 599.600 57.600 600.400 57.700 ;
        RECT 678.000 58.300 678.800 58.400 ;
        RECT 679.600 58.300 680.400 58.400 ;
        RECT 678.000 57.700 680.400 58.300 ;
        RECT 678.000 57.600 678.800 57.700 ;
        RECT 679.600 57.600 680.400 57.700 ;
        RECT 20.400 56.300 21.200 56.400 ;
        RECT 22.000 56.300 22.800 56.400 ;
        RECT 20.400 55.700 22.800 56.300 ;
        RECT 20.400 55.600 21.200 55.700 ;
        RECT 22.000 55.600 22.800 55.700 ;
        RECT 30.000 56.300 30.800 56.400 ;
        RECT 41.200 56.300 42.000 56.400 ;
        RECT 30.000 55.700 42.000 56.300 ;
        RECT 30.000 55.600 30.800 55.700 ;
        RECT 41.200 55.600 42.000 55.700 ;
        RECT 54.000 56.300 54.800 56.400 ;
        RECT 94.000 56.300 94.800 56.400 ;
        RECT 54.000 55.700 94.800 56.300 ;
        RECT 54.000 55.600 54.800 55.700 ;
        RECT 94.000 55.600 94.800 55.700 ;
        RECT 113.200 56.300 114.000 56.400 ;
        RECT 122.800 56.300 123.600 56.400 ;
        RECT 113.200 55.700 123.600 56.300 ;
        RECT 113.200 55.600 114.000 55.700 ;
        RECT 122.800 55.600 123.600 55.700 ;
        RECT 126.000 56.300 126.800 56.400 ;
        RECT 140.400 56.300 141.200 56.400 ;
        RECT 126.000 55.700 141.200 56.300 ;
        RECT 126.000 55.600 126.800 55.700 ;
        RECT 140.400 55.600 141.200 55.700 ;
        RECT 193.200 56.300 194.000 56.400 ;
        RECT 214.000 56.300 214.800 56.400 ;
        RECT 215.600 56.300 216.400 56.400 ;
        RECT 193.200 55.700 216.400 56.300 ;
        RECT 193.200 55.600 194.000 55.700 ;
        RECT 214.000 55.600 214.800 55.700 ;
        RECT 215.600 55.600 216.400 55.700 ;
        RECT 247.600 56.300 248.400 56.400 ;
        RECT 257.200 56.300 258.000 56.400 ;
        RECT 295.600 56.300 296.400 56.400 ;
        RECT 247.600 55.700 296.400 56.300 ;
        RECT 247.600 55.600 248.400 55.700 ;
        RECT 257.200 55.600 258.000 55.700 ;
        RECT 295.600 55.600 296.400 55.700 ;
        RECT 302.000 56.300 302.800 56.400 ;
        RECT 310.000 56.300 310.800 56.400 ;
        RECT 302.000 55.700 310.800 56.300 ;
        RECT 302.000 55.600 302.800 55.700 ;
        RECT 310.000 55.600 310.800 55.700 ;
        RECT 332.400 56.300 333.200 56.400 ;
        RECT 375.600 56.300 376.400 56.400 ;
        RECT 415.600 56.300 416.400 56.400 ;
        RECT 428.400 56.300 429.200 56.400 ;
        RECT 332.400 55.700 429.200 56.300 ;
        RECT 332.400 55.600 333.200 55.700 ;
        RECT 375.600 55.600 376.400 55.700 ;
        RECT 415.600 55.600 416.400 55.700 ;
        RECT 428.400 55.600 429.200 55.700 ;
        RECT 505.200 56.300 506.000 56.400 ;
        RECT 518.000 56.300 518.800 56.400 ;
        RECT 505.200 55.700 518.800 56.300 ;
        RECT 505.200 55.600 506.000 55.700 ;
        RECT 518.000 55.600 518.800 55.700 ;
        RECT 519.600 56.300 520.400 56.400 ;
        RECT 529.200 56.300 530.000 56.400 ;
        RECT 519.600 55.700 530.000 56.300 ;
        RECT 519.600 55.600 520.400 55.700 ;
        RECT 529.200 55.600 530.000 55.700 ;
        RECT 540.400 56.300 541.200 56.400 ;
        RECT 567.600 56.300 568.400 56.400 ;
        RECT 540.400 55.700 568.400 56.300 ;
        RECT 582.100 56.300 582.700 57.600 ;
        RECT 594.800 56.300 595.600 56.400 ;
        RECT 582.100 55.700 595.600 56.300 ;
        RECT 540.400 55.600 541.200 55.700 ;
        RECT 567.600 55.600 568.400 55.700 ;
        RECT 594.800 55.600 595.600 55.700 ;
        RECT 626.800 56.300 627.600 56.400 ;
        RECT 654.000 56.300 654.800 56.400 ;
        RECT 626.800 55.700 654.800 56.300 ;
        RECT 626.800 55.600 627.600 55.700 ;
        RECT 654.000 55.600 654.800 55.700 ;
        RECT 673.200 56.300 674.000 56.400 ;
        RECT 686.000 56.300 686.800 56.400 ;
        RECT 673.200 55.700 686.800 56.300 ;
        RECT 673.200 55.600 674.000 55.700 ;
        RECT 686.000 55.600 686.800 55.700 ;
        RECT 9.200 54.300 10.000 54.400 ;
        RECT 26.800 54.300 27.600 54.400 ;
        RECT 9.200 53.700 27.600 54.300 ;
        RECT 9.200 53.600 10.000 53.700 ;
        RECT 26.800 53.600 27.600 53.700 ;
        RECT 30.000 54.300 30.800 54.400 ;
        RECT 36.400 54.300 37.200 54.400 ;
        RECT 30.000 53.700 37.200 54.300 ;
        RECT 30.000 53.600 30.800 53.700 ;
        RECT 36.400 53.600 37.200 53.700 ;
        RECT 44.400 54.300 45.200 54.400 ;
        RECT 92.400 54.300 93.200 54.400 ;
        RECT 118.000 54.300 118.800 54.400 ;
        RECT 130.800 54.300 131.600 54.400 ;
        RECT 44.400 53.700 91.500 54.300 ;
        RECT 44.400 53.600 45.200 53.700 ;
        RECT 22.000 52.300 22.800 52.400 ;
        RECT 54.000 52.300 54.800 52.400 ;
        RECT 22.000 51.700 54.800 52.300 ;
        RECT 22.000 51.600 22.800 51.700 ;
        RECT 54.000 51.600 54.800 51.700 ;
        RECT 60.400 52.300 61.200 52.400 ;
        RECT 70.000 52.300 70.800 52.400 ;
        RECT 60.400 51.700 70.800 52.300 ;
        RECT 90.900 52.300 91.500 53.700 ;
        RECT 92.400 53.700 131.600 54.300 ;
        RECT 92.400 53.600 93.200 53.700 ;
        RECT 118.000 53.600 118.800 53.700 ;
        RECT 130.800 53.600 131.600 53.700 ;
        RECT 276.400 54.300 277.200 54.400 ;
        RECT 297.200 54.300 298.000 54.400 ;
        RECT 276.400 53.700 298.000 54.300 ;
        RECT 276.400 53.600 277.200 53.700 ;
        RECT 297.200 53.600 298.000 53.700 ;
        RECT 390.000 54.300 390.800 54.400 ;
        RECT 393.200 54.300 394.000 54.400 ;
        RECT 401.200 54.300 402.000 54.400 ;
        RECT 390.000 53.700 402.000 54.300 ;
        RECT 390.000 53.600 390.800 53.700 ;
        RECT 393.200 53.600 394.000 53.700 ;
        RECT 401.200 53.600 402.000 53.700 ;
        RECT 441.200 54.300 442.000 54.400 ;
        RECT 442.800 54.300 443.600 54.400 ;
        RECT 441.200 53.700 443.600 54.300 ;
        RECT 441.200 53.600 442.000 53.700 ;
        RECT 442.800 53.600 443.600 53.700 ;
        RECT 449.200 54.300 450.000 54.400 ;
        RECT 454.000 54.300 454.800 54.400 ;
        RECT 457.200 54.300 458.000 54.400 ;
        RECT 449.200 53.700 458.000 54.300 ;
        RECT 449.200 53.600 450.000 53.700 ;
        RECT 454.000 53.600 454.800 53.700 ;
        RECT 457.200 53.600 458.000 53.700 ;
        RECT 471.600 54.300 472.400 54.400 ;
        RECT 492.400 54.300 493.200 54.400 ;
        RECT 471.600 53.700 493.200 54.300 ;
        RECT 471.600 53.600 472.400 53.700 ;
        RECT 492.400 53.600 493.200 53.700 ;
        RECT 510.000 54.300 510.800 54.400 ;
        RECT 524.400 54.300 525.200 54.400 ;
        RECT 510.000 53.700 525.200 54.300 ;
        RECT 510.000 53.600 510.800 53.700 ;
        RECT 524.400 53.600 525.200 53.700 ;
        RECT 538.800 54.300 539.600 54.400 ;
        RECT 543.600 54.300 544.400 54.400 ;
        RECT 538.800 53.700 544.400 54.300 ;
        RECT 538.800 53.600 539.600 53.700 ;
        RECT 543.600 53.600 544.400 53.700 ;
        RECT 561.200 54.300 562.000 54.400 ;
        RECT 580.400 54.300 581.200 54.400 ;
        RECT 585.200 54.300 586.000 54.400 ;
        RECT 561.200 53.700 586.000 54.300 ;
        RECT 561.200 53.600 562.000 53.700 ;
        RECT 580.400 53.600 581.200 53.700 ;
        RECT 585.200 53.600 586.000 53.700 ;
        RECT 598.000 54.300 598.800 54.400 ;
        RECT 618.800 54.300 619.600 54.400 ;
        RECT 628.400 54.300 629.200 54.400 ;
        RECT 634.800 54.300 635.600 54.400 ;
        RECT 598.000 53.700 635.600 54.300 ;
        RECT 598.000 53.600 598.800 53.700 ;
        RECT 618.800 53.600 619.600 53.700 ;
        RECT 628.400 53.600 629.200 53.700 ;
        RECT 634.800 53.600 635.600 53.700 ;
        RECT 636.400 54.300 637.200 54.400 ;
        RECT 642.800 54.300 643.600 54.400 ;
        RECT 636.400 53.700 643.600 54.300 ;
        RECT 636.400 53.600 637.200 53.700 ;
        RECT 642.800 53.600 643.600 53.700 ;
        RECT 646.000 54.300 646.800 54.400 ;
        RECT 650.800 54.300 651.600 54.400 ;
        RECT 646.000 53.700 651.600 54.300 ;
        RECT 646.000 53.600 646.800 53.700 ;
        RECT 650.800 53.600 651.600 53.700 ;
        RECT 660.400 54.300 661.200 54.400 ;
        RECT 666.800 54.300 667.600 54.400 ;
        RECT 660.400 53.700 667.600 54.300 ;
        RECT 660.400 53.600 661.200 53.700 ;
        RECT 666.800 53.600 667.600 53.700 ;
        RECT 668.400 54.300 669.200 54.400 ;
        RECT 687.600 54.300 688.400 54.400 ;
        RECT 668.400 53.700 688.400 54.300 ;
        RECT 668.400 53.600 669.200 53.700 ;
        RECT 687.600 53.600 688.400 53.700 ;
        RECT 95.600 52.300 96.400 52.400 ;
        RECT 105.200 52.300 106.000 52.400 ;
        RECT 90.900 51.700 106.000 52.300 ;
        RECT 60.400 51.600 61.200 51.700 ;
        RECT 70.000 51.600 70.800 51.700 ;
        RECT 95.600 51.600 96.400 51.700 ;
        RECT 105.200 51.600 106.000 51.700 ;
        RECT 119.600 52.300 120.400 52.400 ;
        RECT 132.400 52.300 133.200 52.400 ;
        RECT 119.600 51.700 133.200 52.300 ;
        RECT 119.600 51.600 120.400 51.700 ;
        RECT 132.400 51.600 133.200 51.700 ;
        RECT 138.800 52.300 139.600 52.400 ;
        RECT 148.400 52.300 149.200 52.400 ;
        RECT 151.600 52.300 152.400 52.400 ;
        RECT 138.800 51.700 152.400 52.300 ;
        RECT 138.800 51.600 139.600 51.700 ;
        RECT 148.400 51.600 149.200 51.700 ;
        RECT 151.600 51.600 152.400 51.700 ;
        RECT 158.000 52.300 158.800 52.400 ;
        RECT 162.800 52.300 163.600 52.400 ;
        RECT 158.000 51.700 163.600 52.300 ;
        RECT 158.000 51.600 158.800 51.700 ;
        RECT 162.800 51.600 163.600 51.700 ;
        RECT 164.400 52.300 165.200 52.400 ;
        RECT 182.000 52.300 182.800 52.400 ;
        RECT 164.400 51.700 182.800 52.300 ;
        RECT 164.400 51.600 165.200 51.700 ;
        RECT 182.000 51.600 182.800 51.700 ;
        RECT 260.400 52.300 261.200 52.400 ;
        RECT 266.800 52.300 267.600 52.400 ;
        RECT 260.400 51.700 267.600 52.300 ;
        RECT 260.400 51.600 261.200 51.700 ;
        RECT 266.800 51.600 267.600 51.700 ;
        RECT 358.000 52.300 358.800 52.400 ;
        RECT 367.600 52.300 368.400 52.400 ;
        RECT 358.000 51.700 368.400 52.300 ;
        RECT 358.000 51.600 358.800 51.700 ;
        RECT 367.600 51.600 368.400 51.700 ;
        RECT 428.400 52.300 429.200 52.400 ;
        RECT 439.600 52.300 440.400 52.400 ;
        RECT 428.400 51.700 440.400 52.300 ;
        RECT 428.400 51.600 429.200 51.700 ;
        RECT 439.600 51.600 440.400 51.700 ;
        RECT 455.600 52.300 456.400 52.400 ;
        RECT 462.000 52.300 462.800 52.400 ;
        RECT 455.600 51.700 462.800 52.300 ;
        RECT 455.600 51.600 456.400 51.700 ;
        RECT 462.000 51.600 462.800 51.700 ;
        RECT 494.000 52.300 494.800 52.400 ;
        RECT 500.400 52.300 501.200 52.400 ;
        RECT 494.000 51.700 501.200 52.300 ;
        RECT 494.000 51.600 494.800 51.700 ;
        RECT 500.400 51.600 501.200 51.700 ;
        RECT 503.600 52.300 504.400 52.400 ;
        RECT 514.800 52.300 515.600 52.400 ;
        RECT 503.600 51.700 515.600 52.300 ;
        RECT 503.600 51.600 504.400 51.700 ;
        RECT 514.800 51.600 515.600 51.700 ;
        RECT 522.800 52.300 523.600 52.400 ;
        RECT 529.200 52.300 530.000 52.400 ;
        RECT 522.800 51.700 530.000 52.300 ;
        RECT 522.800 51.600 523.600 51.700 ;
        RECT 529.200 51.600 530.000 51.700 ;
        RECT 530.800 52.300 531.600 52.400 ;
        RECT 553.200 52.300 554.000 52.400 ;
        RECT 530.800 51.700 554.000 52.300 ;
        RECT 530.800 51.600 531.600 51.700 ;
        RECT 553.200 51.600 554.000 51.700 ;
        RECT 558.000 52.300 558.800 52.400 ;
        RECT 596.400 52.300 597.200 52.400 ;
        RECT 558.000 51.700 597.200 52.300 ;
        RECT 558.000 51.600 558.800 51.700 ;
        RECT 596.400 51.600 597.200 51.700 ;
        RECT 602.800 52.300 603.600 52.400 ;
        RECT 625.200 52.300 626.000 52.400 ;
        RECT 602.800 51.700 626.000 52.300 ;
        RECT 602.800 51.600 603.600 51.700 ;
        RECT 625.200 51.600 626.000 51.700 ;
        RECT 641.200 52.300 642.000 52.400 ;
        RECT 650.800 52.300 651.600 52.400 ;
        RECT 660.400 52.300 661.200 52.400 ;
        RECT 678.000 52.300 678.800 52.400 ;
        RECT 641.200 51.700 649.900 52.300 ;
        RECT 641.200 51.600 642.000 51.700 ;
        RECT 18.800 50.300 19.600 50.400 ;
        RECT 25.200 50.300 26.000 50.400 ;
        RECT 49.200 50.300 50.000 50.400 ;
        RECT 18.800 49.700 50.000 50.300 ;
        RECT 18.800 49.600 19.600 49.700 ;
        RECT 25.200 49.600 26.000 49.700 ;
        RECT 49.200 49.600 50.000 49.700 ;
        RECT 50.800 50.300 51.600 50.400 ;
        RECT 52.400 50.300 53.200 50.400 ;
        RECT 50.800 49.700 53.200 50.300 ;
        RECT 50.800 49.600 51.600 49.700 ;
        RECT 52.400 49.600 53.200 49.700 ;
        RECT 87.600 50.300 88.400 50.400 ;
        RECT 90.800 50.300 91.600 50.400 ;
        RECT 87.600 49.700 91.600 50.300 ;
        RECT 87.600 49.600 88.400 49.700 ;
        RECT 90.800 49.600 91.600 49.700 ;
        RECT 94.000 50.300 94.800 50.400 ;
        RECT 137.200 50.300 138.000 50.400 ;
        RECT 142.000 50.300 142.800 50.400 ;
        RECT 145.200 50.300 146.000 50.400 ;
        RECT 94.000 49.700 146.000 50.300 ;
        RECT 94.000 49.600 94.800 49.700 ;
        RECT 137.200 49.600 138.000 49.700 ;
        RECT 142.000 49.600 142.800 49.700 ;
        RECT 145.200 49.600 146.000 49.700 ;
        RECT 156.400 50.300 157.200 50.400 ;
        RECT 169.200 50.300 170.000 50.400 ;
        RECT 156.400 49.700 170.000 50.300 ;
        RECT 156.400 49.600 157.200 49.700 ;
        RECT 169.200 49.600 170.000 49.700 ;
        RECT 206.000 50.300 206.800 50.400 ;
        RECT 218.800 50.300 219.600 50.400 ;
        RECT 206.000 49.700 219.600 50.300 ;
        RECT 206.000 49.600 206.800 49.700 ;
        RECT 218.800 49.600 219.600 49.700 ;
        RECT 287.600 50.300 288.400 50.400 ;
        RECT 295.600 50.300 296.400 50.400 ;
        RECT 302.000 50.300 302.800 50.400 ;
        RECT 287.600 49.700 302.800 50.300 ;
        RECT 287.600 49.600 288.400 49.700 ;
        RECT 295.600 49.600 296.400 49.700 ;
        RECT 302.000 49.600 302.800 49.700 ;
        RECT 498.800 50.300 499.600 50.400 ;
        RECT 508.400 50.300 509.200 50.400 ;
        RECT 498.800 49.700 509.200 50.300 ;
        RECT 498.800 49.600 499.600 49.700 ;
        RECT 508.400 49.600 509.200 49.700 ;
        RECT 534.000 50.300 534.800 50.400 ;
        RECT 540.400 50.300 541.200 50.400 ;
        RECT 534.000 49.700 541.200 50.300 ;
        RECT 534.000 49.600 534.800 49.700 ;
        RECT 540.400 49.600 541.200 49.700 ;
        RECT 554.800 50.300 555.600 50.400 ;
        RECT 562.800 50.300 563.600 50.400 ;
        RECT 554.800 49.700 563.600 50.300 ;
        RECT 554.800 49.600 555.600 49.700 ;
        RECT 562.800 49.600 563.600 49.700 ;
        RECT 599.600 50.300 600.400 50.400 ;
        RECT 620.400 50.300 621.200 50.400 ;
        RECT 644.400 50.300 645.200 50.400 ;
        RECT 599.600 49.700 645.200 50.300 ;
        RECT 649.300 50.300 649.900 51.700 ;
        RECT 650.800 51.700 678.800 52.300 ;
        RECT 650.800 51.600 651.600 51.700 ;
        RECT 660.400 51.600 661.200 51.700 ;
        RECT 678.000 51.600 678.800 51.700 ;
        RECT 668.400 50.300 669.200 50.400 ;
        RECT 649.300 49.700 669.200 50.300 ;
        RECT 599.600 49.600 600.400 49.700 ;
        RECT 620.400 49.600 621.200 49.700 ;
        RECT 644.400 49.600 645.200 49.700 ;
        RECT 668.400 49.600 669.200 49.700 ;
        RECT 671.600 50.300 672.400 50.400 ;
        RECT 676.400 50.300 677.200 50.400 ;
        RECT 681.200 50.300 682.000 50.400 ;
        RECT 671.600 49.700 682.000 50.300 ;
        RECT 671.600 49.600 672.400 49.700 ;
        RECT 676.400 49.600 677.200 49.700 ;
        RECT 681.200 49.600 682.000 49.700 ;
        RECT 129.200 48.300 130.000 48.400 ;
        RECT 132.400 48.300 133.200 48.400 ;
        RECT 129.200 47.700 133.200 48.300 ;
        RECT 129.200 47.600 130.000 47.700 ;
        RECT 132.400 47.600 133.200 47.700 ;
        RECT 135.600 48.300 136.400 48.400 ;
        RECT 140.400 48.300 141.200 48.400 ;
        RECT 143.600 48.300 144.400 48.400 ;
        RECT 159.600 48.300 160.400 48.400 ;
        RECT 135.600 47.700 160.400 48.300 ;
        RECT 135.600 47.600 136.400 47.700 ;
        RECT 140.400 47.600 141.200 47.700 ;
        RECT 143.600 47.600 144.400 47.700 ;
        RECT 159.600 47.600 160.400 47.700 ;
        RECT 167.600 48.300 168.400 48.400 ;
        RECT 170.800 48.300 171.600 48.400 ;
        RECT 167.600 47.700 171.600 48.300 ;
        RECT 167.600 47.600 168.400 47.700 ;
        RECT 170.800 47.600 171.600 47.700 ;
        RECT 172.400 48.300 173.200 48.400 ;
        RECT 175.600 48.300 176.400 48.400 ;
        RECT 172.400 47.700 176.400 48.300 ;
        RECT 172.400 47.600 173.200 47.700 ;
        RECT 175.600 47.600 176.400 47.700 ;
        RECT 497.200 48.300 498.000 48.400 ;
        RECT 506.800 48.300 507.600 48.400 ;
        RECT 511.600 48.300 512.400 48.400 ;
        RECT 497.200 47.700 512.400 48.300 ;
        RECT 497.200 47.600 498.000 47.700 ;
        RECT 506.800 47.600 507.600 47.700 ;
        RECT 511.600 47.600 512.400 47.700 ;
        RECT 569.200 48.300 570.000 48.400 ;
        RECT 583.600 48.300 584.400 48.400 ;
        RECT 569.200 47.700 584.400 48.300 ;
        RECT 569.200 47.600 570.000 47.700 ;
        RECT 583.600 47.600 584.400 47.700 ;
        RECT 588.400 48.300 589.200 48.400 ;
        RECT 612.400 48.300 613.200 48.400 ;
        RECT 646.000 48.300 646.800 48.400 ;
        RECT 588.400 47.700 593.900 48.300 ;
        RECT 588.400 47.600 589.200 47.700 ;
        RECT 79.600 46.300 80.400 46.400 ;
        RECT 212.400 46.300 213.200 46.400 ;
        RECT 79.600 45.700 213.200 46.300 ;
        RECT 79.600 45.600 80.400 45.700 ;
        RECT 212.400 45.600 213.200 45.700 ;
        RECT 514.800 46.300 515.600 46.400 ;
        RECT 546.800 46.300 547.600 46.400 ;
        RECT 514.800 45.700 547.600 46.300 ;
        RECT 514.800 45.600 515.600 45.700 ;
        RECT 546.800 45.600 547.600 45.700 ;
        RECT 548.400 46.300 549.200 46.400 ;
        RECT 591.600 46.300 592.400 46.400 ;
        RECT 548.400 45.700 592.400 46.300 ;
        RECT 593.300 46.300 593.900 47.700 ;
        RECT 612.400 47.700 646.800 48.300 ;
        RECT 612.400 47.600 613.200 47.700 ;
        RECT 646.000 47.600 646.800 47.700 ;
        RECT 647.600 48.300 648.400 48.400 ;
        RECT 650.800 48.300 651.600 48.400 ;
        RECT 647.600 47.700 651.600 48.300 ;
        RECT 647.600 47.600 648.400 47.700 ;
        RECT 650.800 47.600 651.600 47.700 ;
        RECT 671.600 48.300 672.400 48.400 ;
        RECT 686.000 48.300 686.800 48.400 ;
        RECT 671.600 47.700 686.800 48.300 ;
        RECT 671.600 47.600 672.400 47.700 ;
        RECT 686.000 47.600 686.800 47.700 ;
        RECT 657.200 46.300 658.000 46.400 ;
        RECT 663.600 46.300 664.400 46.400 ;
        RECT 593.300 45.700 664.400 46.300 ;
        RECT 548.400 45.600 549.200 45.700 ;
        RECT 591.600 45.600 592.400 45.700 ;
        RECT 657.200 45.600 658.000 45.700 ;
        RECT 663.600 45.600 664.400 45.700 ;
        RECT 681.200 46.300 682.000 46.400 ;
        RECT 684.400 46.300 685.200 46.400 ;
        RECT 681.200 45.700 685.200 46.300 ;
        RECT 681.200 45.600 682.000 45.700 ;
        RECT 684.400 45.600 685.200 45.700 ;
        RECT 12.400 44.300 13.200 44.400 ;
        RECT 17.200 44.300 18.000 44.400 ;
        RECT 12.400 43.700 18.000 44.300 ;
        RECT 12.400 43.600 13.200 43.700 ;
        RECT 17.200 43.600 18.000 43.700 ;
        RECT 90.800 44.300 91.600 44.400 ;
        RECT 94.000 44.300 94.800 44.400 ;
        RECT 90.800 43.700 94.800 44.300 ;
        RECT 90.800 43.600 91.600 43.700 ;
        RECT 94.000 43.600 94.800 43.700 ;
        RECT 615.600 44.300 616.400 44.400 ;
        RECT 633.200 44.300 634.000 44.400 ;
        RECT 615.600 43.700 634.000 44.300 ;
        RECT 615.600 43.600 616.400 43.700 ;
        RECT 633.200 43.600 634.000 43.700 ;
        RECT 636.400 44.300 637.200 44.400 ;
        RECT 658.800 44.300 659.600 44.400 ;
        RECT 636.400 43.700 659.600 44.300 ;
        RECT 636.400 43.600 637.200 43.700 ;
        RECT 658.800 43.600 659.600 43.700 ;
        RECT 673.200 44.300 674.000 44.400 ;
        RECT 679.600 44.300 680.400 44.400 ;
        RECT 673.200 43.700 680.400 44.300 ;
        RECT 673.200 43.600 674.000 43.700 ;
        RECT 679.600 43.600 680.400 43.700 ;
        RECT 90.800 42.300 91.600 42.400 ;
        RECT 97.200 42.300 98.000 42.400 ;
        RECT 90.800 41.700 98.000 42.300 ;
        RECT 90.800 41.600 91.600 41.700 ;
        RECT 97.200 41.600 98.000 41.700 ;
        RECT 118.000 42.300 118.800 42.400 ;
        RECT 158.000 42.300 158.800 42.400 ;
        RECT 175.600 42.300 176.400 42.400 ;
        RECT 118.000 41.700 176.400 42.300 ;
        RECT 118.000 41.600 118.800 41.700 ;
        RECT 158.000 41.600 158.800 41.700 ;
        RECT 175.600 41.600 176.400 41.700 ;
        RECT 454.000 42.300 454.800 42.400 ;
        RECT 468.400 42.300 469.200 42.400 ;
        RECT 479.600 42.300 480.400 42.400 ;
        RECT 454.000 41.700 480.400 42.300 ;
        RECT 454.000 41.600 454.800 41.700 ;
        RECT 468.400 41.600 469.200 41.700 ;
        RECT 479.600 41.600 480.400 41.700 ;
        RECT 628.400 42.300 629.200 42.400 ;
        RECT 638.000 42.300 638.800 42.400 ;
        RECT 628.400 41.700 638.800 42.300 ;
        RECT 628.400 41.600 629.200 41.700 ;
        RECT 638.000 41.600 638.800 41.700 ;
        RECT 252.400 40.300 253.200 40.400 ;
        RECT 278.000 40.300 278.800 40.400 ;
        RECT 252.400 39.700 278.800 40.300 ;
        RECT 252.400 39.600 253.200 39.700 ;
        RECT 278.000 39.600 278.800 39.700 ;
        RECT 370.800 40.300 371.600 40.400 ;
        RECT 394.800 40.300 395.600 40.400 ;
        RECT 370.800 39.700 395.600 40.300 ;
        RECT 370.800 39.600 371.600 39.700 ;
        RECT 394.800 39.600 395.600 39.700 ;
        RECT 442.800 40.300 443.600 40.400 ;
        RECT 478.000 40.300 478.800 40.400 ;
        RECT 442.800 39.700 478.800 40.300 ;
        RECT 442.800 39.600 443.600 39.700 ;
        RECT 478.000 39.600 478.800 39.700 ;
        RECT 513.200 40.300 514.000 40.400 ;
        RECT 521.200 40.300 522.000 40.400 ;
        RECT 513.200 39.700 522.000 40.300 ;
        RECT 513.200 39.600 514.000 39.700 ;
        RECT 521.200 39.600 522.000 39.700 ;
        RECT 100.400 38.300 101.200 38.400 ;
        RECT 135.600 38.300 136.400 38.400 ;
        RECT 146.800 38.300 147.600 38.400 ;
        RECT 100.400 37.700 147.600 38.300 ;
        RECT 100.400 37.600 101.200 37.700 ;
        RECT 135.600 37.600 136.400 37.700 ;
        RECT 146.800 37.600 147.600 37.700 ;
        RECT 169.200 38.300 170.000 38.400 ;
        RECT 172.400 38.300 173.200 38.400 ;
        RECT 169.200 37.700 173.200 38.300 ;
        RECT 169.200 37.600 170.000 37.700 ;
        RECT 172.400 37.600 173.200 37.700 ;
        RECT 233.200 38.300 234.000 38.400 ;
        RECT 249.200 38.300 250.000 38.400 ;
        RECT 279.600 38.300 280.400 38.400 ;
        RECT 290.800 38.300 291.600 38.400 ;
        RECT 233.200 37.700 291.600 38.300 ;
        RECT 233.200 37.600 234.000 37.700 ;
        RECT 249.200 37.600 250.000 37.700 ;
        RECT 279.600 37.600 280.400 37.700 ;
        RECT 290.800 37.600 291.600 37.700 ;
        RECT 426.800 38.300 427.600 38.400 ;
        RECT 433.200 38.300 434.000 38.400 ;
        RECT 426.800 37.700 434.000 38.300 ;
        RECT 426.800 37.600 427.600 37.700 ;
        RECT 433.200 37.600 434.000 37.700 ;
        RECT 457.200 38.300 458.000 38.400 ;
        RECT 463.600 38.300 464.400 38.400 ;
        RECT 473.200 38.300 474.000 38.400 ;
        RECT 457.200 37.700 474.000 38.300 ;
        RECT 457.200 37.600 458.000 37.700 ;
        RECT 463.600 37.600 464.400 37.700 ;
        RECT 473.200 37.600 474.000 37.700 ;
        RECT 514.800 38.300 515.600 38.400 ;
        RECT 530.800 38.300 531.600 38.400 ;
        RECT 514.800 37.700 531.600 38.300 ;
        RECT 514.800 37.600 515.600 37.700 ;
        RECT 530.800 37.600 531.600 37.700 ;
        RECT 559.600 38.300 560.400 38.400 ;
        RECT 609.200 38.300 610.000 38.400 ;
        RECT 559.600 37.700 610.000 38.300 ;
        RECT 559.600 37.600 560.400 37.700 ;
        RECT 609.200 37.600 610.000 37.700 ;
        RECT 625.200 38.300 626.000 38.400 ;
        RECT 636.400 38.300 637.200 38.400 ;
        RECT 625.200 37.700 637.200 38.300 ;
        RECT 625.200 37.600 626.000 37.700 ;
        RECT 636.400 37.600 637.200 37.700 ;
        RECT 638.000 38.300 638.800 38.400 ;
        RECT 666.800 38.300 667.600 38.400 ;
        RECT 638.000 37.700 667.600 38.300 ;
        RECT 638.000 37.600 638.800 37.700 ;
        RECT 666.800 37.600 667.600 37.700 ;
        RECT 103.600 36.300 104.400 36.400 ;
        RECT 106.800 36.300 107.600 36.400 ;
        RECT 103.600 35.700 107.600 36.300 ;
        RECT 103.600 35.600 104.400 35.700 ;
        RECT 106.800 35.600 107.600 35.700 ;
        RECT 407.600 36.300 408.400 36.400 ;
        RECT 422.000 36.300 422.800 36.400 ;
        RECT 407.600 35.700 422.800 36.300 ;
        RECT 407.600 35.600 408.400 35.700 ;
        RECT 422.000 35.600 422.800 35.700 ;
        RECT 550.000 36.300 550.800 36.400 ;
        RECT 638.000 36.300 638.800 36.400 ;
        RECT 550.000 35.700 638.800 36.300 ;
        RECT 550.000 35.600 550.800 35.700 ;
        RECT 638.000 35.600 638.800 35.700 ;
        RECT 663.600 36.300 664.400 36.400 ;
        RECT 666.800 36.300 667.600 36.400 ;
        RECT 663.600 35.700 667.600 36.300 ;
        RECT 663.600 35.600 664.400 35.700 ;
        RECT 666.800 35.600 667.600 35.700 ;
        RECT 41.200 34.300 42.000 34.400 ;
        RECT 49.200 34.300 50.000 34.400 ;
        RECT 57.200 34.300 58.000 34.400 ;
        RECT 41.200 33.700 58.000 34.300 ;
        RECT 41.200 33.600 42.000 33.700 ;
        RECT 49.200 33.600 50.000 33.700 ;
        RECT 57.200 33.600 58.000 33.700 ;
        RECT 103.600 34.300 104.400 34.400 ;
        RECT 119.600 34.300 120.400 34.400 ;
        RECT 103.600 33.700 120.400 34.300 ;
        RECT 103.600 33.600 104.400 33.700 ;
        RECT 119.600 33.600 120.400 33.700 ;
        RECT 302.000 34.300 302.800 34.400 ;
        RECT 348.400 34.300 349.200 34.400 ;
        RECT 302.000 33.700 349.200 34.300 ;
        RECT 302.000 33.600 302.800 33.700 ;
        RECT 348.400 33.600 349.200 33.700 ;
        RECT 385.200 34.300 386.000 34.400 ;
        RECT 414.000 34.300 414.800 34.400 ;
        RECT 385.200 33.700 414.800 34.300 ;
        RECT 385.200 33.600 386.000 33.700 ;
        RECT 414.000 33.600 414.800 33.700 ;
        RECT 478.000 34.300 478.800 34.400 ;
        RECT 484.400 34.300 485.200 34.400 ;
        RECT 505.200 34.300 506.000 34.400 ;
        RECT 478.000 33.700 506.000 34.300 ;
        RECT 478.000 33.600 478.800 33.700 ;
        RECT 484.400 33.600 485.200 33.700 ;
        RECT 505.200 33.600 506.000 33.700 ;
        RECT 527.600 34.300 528.400 34.400 ;
        RECT 538.800 34.300 539.600 34.400 ;
        RECT 543.600 34.300 544.400 34.400 ;
        RECT 527.600 33.700 544.400 34.300 ;
        RECT 527.600 33.600 528.400 33.700 ;
        RECT 538.800 33.600 539.600 33.700 ;
        RECT 543.600 33.600 544.400 33.700 ;
        RECT 556.400 34.300 557.200 34.400 ;
        RECT 567.600 34.300 568.400 34.400 ;
        RECT 572.400 34.300 573.200 34.400 ;
        RECT 556.400 33.700 573.200 34.300 ;
        RECT 556.400 33.600 557.200 33.700 ;
        RECT 567.600 33.600 568.400 33.700 ;
        RECT 572.400 33.600 573.200 33.700 ;
        RECT 593.200 34.300 594.000 34.400 ;
        RECT 609.200 34.300 610.000 34.400 ;
        RECT 593.200 33.700 610.000 34.300 ;
        RECT 593.200 33.600 594.000 33.700 ;
        RECT 609.200 33.600 610.000 33.700 ;
        RECT 610.800 34.300 611.600 34.400 ;
        RECT 626.800 34.300 627.600 34.400 ;
        RECT 610.800 33.700 627.600 34.300 ;
        RECT 610.800 33.600 611.600 33.700 ;
        RECT 626.800 33.600 627.600 33.700 ;
        RECT 634.800 34.300 635.600 34.400 ;
        RECT 647.600 34.300 648.400 34.400 ;
        RECT 654.000 34.300 654.800 34.400 ;
        RECT 634.800 33.700 654.800 34.300 ;
        RECT 634.800 33.600 635.600 33.700 ;
        RECT 647.600 33.600 648.400 33.700 ;
        RECT 654.000 33.600 654.800 33.700 ;
        RECT 663.600 34.300 664.400 34.400 ;
        RECT 684.400 34.300 685.200 34.400 ;
        RECT 663.600 33.700 685.200 34.300 ;
        RECT 663.600 33.600 664.400 33.700 ;
        RECT 684.400 33.600 685.200 33.700 ;
        RECT 33.200 32.300 34.000 32.400 ;
        RECT 46.000 32.300 46.800 32.400 ;
        RECT 33.200 31.700 46.800 32.300 ;
        RECT 33.200 31.600 34.000 31.700 ;
        RECT 46.000 31.600 46.800 31.700 ;
        RECT 58.800 32.300 59.600 32.400 ;
        RECT 63.600 32.300 64.400 32.400 ;
        RECT 58.800 31.700 64.400 32.300 ;
        RECT 58.800 31.600 59.600 31.700 ;
        RECT 63.600 31.600 64.400 31.700 ;
        RECT 110.000 32.300 110.800 32.400 ;
        RECT 122.800 32.300 123.600 32.400 ;
        RECT 110.000 31.700 123.600 32.300 ;
        RECT 110.000 31.600 110.800 31.700 ;
        RECT 122.800 31.600 123.600 31.700 ;
        RECT 142.000 32.300 142.800 32.400 ;
        RECT 156.400 32.300 157.200 32.400 ;
        RECT 142.000 31.700 157.200 32.300 ;
        RECT 142.000 31.600 142.800 31.700 ;
        RECT 156.400 31.600 157.200 31.700 ;
        RECT 308.400 32.300 309.200 32.400 ;
        RECT 311.600 32.300 312.400 32.400 ;
        RECT 308.400 31.700 312.400 32.300 ;
        RECT 308.400 31.600 309.200 31.700 ;
        RECT 311.600 31.600 312.400 31.700 ;
        RECT 410.800 32.300 411.600 32.400 ;
        RECT 434.800 32.300 435.600 32.400 ;
        RECT 410.800 31.700 435.600 32.300 ;
        RECT 410.800 31.600 411.600 31.700 ;
        RECT 434.800 31.600 435.600 31.700 ;
        RECT 447.600 32.300 448.400 32.400 ;
        RECT 462.000 32.300 462.800 32.400 ;
        RECT 466.800 32.300 467.600 32.400 ;
        RECT 447.600 31.700 467.600 32.300 ;
        RECT 447.600 31.600 448.400 31.700 ;
        RECT 462.000 31.600 462.800 31.700 ;
        RECT 466.800 31.600 467.600 31.700 ;
        RECT 482.800 32.300 483.600 32.400 ;
        RECT 486.000 32.300 486.800 32.400 ;
        RECT 482.800 31.700 486.800 32.300 ;
        RECT 482.800 31.600 483.600 31.700 ;
        RECT 486.000 31.600 486.800 31.700 ;
        RECT 524.400 32.300 525.200 32.400 ;
        RECT 551.600 32.300 552.400 32.400 ;
        RECT 524.400 31.700 552.400 32.300 ;
        RECT 524.400 31.600 525.200 31.700 ;
        RECT 551.600 31.600 552.400 31.700 ;
        RECT 553.200 32.300 554.000 32.400 ;
        RECT 618.800 32.300 619.600 32.400 ;
        RECT 553.200 31.700 619.600 32.300 ;
        RECT 553.200 31.600 554.000 31.700 ;
        RECT 618.800 31.600 619.600 31.700 ;
        RECT 622.000 32.300 622.800 32.400 ;
        RECT 631.600 32.300 632.400 32.400 ;
        RECT 622.000 31.700 632.400 32.300 ;
        RECT 622.000 31.600 622.800 31.700 ;
        RECT 631.600 31.600 632.400 31.700 ;
        RECT 650.800 32.300 651.600 32.400 ;
        RECT 660.400 32.300 661.200 32.400 ;
        RECT 650.800 31.700 661.200 32.300 ;
        RECT 650.800 31.600 651.600 31.700 ;
        RECT 660.400 31.600 661.200 31.700 ;
        RECT 662.000 32.300 662.800 32.400 ;
        RECT 671.600 32.300 672.400 32.400 ;
        RECT 662.000 31.700 672.400 32.300 ;
        RECT 662.000 31.600 662.800 31.700 ;
        RECT 671.600 31.600 672.400 31.700 ;
        RECT 2.800 30.300 3.600 30.400 ;
        RECT 41.200 30.300 42.000 30.400 ;
        RECT 60.400 30.300 61.200 30.400 ;
        RECT 2.800 29.700 61.200 30.300 ;
        RECT 2.800 29.600 3.600 29.700 ;
        RECT 41.200 29.600 42.000 29.700 ;
        RECT 60.400 29.600 61.200 29.700 ;
        RECT 98.800 30.300 99.600 30.400 ;
        RECT 110.000 30.300 110.800 30.400 ;
        RECT 98.800 29.700 110.800 30.300 ;
        RECT 98.800 29.600 99.600 29.700 ;
        RECT 110.000 29.600 110.800 29.700 ;
        RECT 134.000 30.300 134.800 30.400 ;
        RECT 137.200 30.300 138.000 30.400 ;
        RECT 134.000 29.700 138.000 30.300 ;
        RECT 134.000 29.600 134.800 29.700 ;
        RECT 137.200 29.600 138.000 29.700 ;
        RECT 143.600 30.300 144.400 30.400 ;
        RECT 148.400 30.300 149.200 30.400 ;
        RECT 143.600 29.700 149.200 30.300 ;
        RECT 143.600 29.600 144.400 29.700 ;
        RECT 148.400 29.600 149.200 29.700 ;
        RECT 150.000 30.300 150.800 30.400 ;
        RECT 159.600 30.300 160.400 30.400 ;
        RECT 150.000 29.700 160.400 30.300 ;
        RECT 150.000 29.600 150.800 29.700 ;
        RECT 159.600 29.600 160.400 29.700 ;
        RECT 177.200 30.300 178.000 30.400 ;
        RECT 186.800 30.300 187.600 30.400 ;
        RECT 177.200 29.700 187.600 30.300 ;
        RECT 177.200 29.600 178.000 29.700 ;
        RECT 186.800 29.600 187.600 29.700 ;
        RECT 246.000 30.300 246.800 30.400 ;
        RECT 276.400 30.300 277.200 30.400 ;
        RECT 246.000 29.700 277.200 30.300 ;
        RECT 246.000 29.600 246.800 29.700 ;
        RECT 276.400 29.600 277.200 29.700 ;
        RECT 289.200 30.300 290.000 30.400 ;
        RECT 302.000 30.300 302.800 30.400 ;
        RECT 289.200 29.700 302.800 30.300 ;
        RECT 289.200 29.600 290.000 29.700 ;
        RECT 302.000 29.600 302.800 29.700 ;
        RECT 305.200 30.300 306.000 30.400 ;
        RECT 308.400 30.300 309.200 30.400 ;
        RECT 305.200 29.700 309.200 30.300 ;
        RECT 305.200 29.600 306.000 29.700 ;
        RECT 308.400 29.600 309.200 29.700 ;
        RECT 359.600 30.300 360.400 30.400 ;
        RECT 370.800 30.300 371.600 30.400 ;
        RECT 359.600 29.700 371.600 30.300 ;
        RECT 359.600 29.600 360.400 29.700 ;
        RECT 370.800 29.600 371.600 29.700 ;
        RECT 410.800 30.300 411.600 30.400 ;
        RECT 414.000 30.300 414.800 30.400 ;
        RECT 410.800 29.700 414.800 30.300 ;
        RECT 410.800 29.600 411.600 29.700 ;
        RECT 414.000 29.600 414.800 29.700 ;
        RECT 428.400 30.300 429.200 30.400 ;
        RECT 434.800 30.300 435.600 30.400 ;
        RECT 428.400 29.700 435.600 30.300 ;
        RECT 428.400 29.600 429.200 29.700 ;
        RECT 434.800 29.600 435.600 29.700 ;
        RECT 444.400 30.300 445.200 30.400 ;
        RECT 476.400 30.300 477.200 30.400 ;
        RECT 482.800 30.300 483.600 30.400 ;
        RECT 503.600 30.300 504.400 30.400 ;
        RECT 444.400 29.700 504.400 30.300 ;
        RECT 444.400 29.600 445.200 29.700 ;
        RECT 476.400 29.600 477.200 29.700 ;
        RECT 482.800 29.600 483.600 29.700 ;
        RECT 503.600 29.600 504.400 29.700 ;
        RECT 516.400 30.300 517.200 30.400 ;
        RECT 530.800 30.300 531.600 30.400 ;
        RECT 516.400 29.700 531.600 30.300 ;
        RECT 516.400 29.600 517.200 29.700 ;
        RECT 530.800 29.600 531.600 29.700 ;
        RECT 546.800 30.300 547.600 30.400 ;
        RECT 556.400 30.300 557.200 30.400 ;
        RECT 546.800 29.700 557.200 30.300 ;
        RECT 546.800 29.600 547.600 29.700 ;
        RECT 556.400 29.600 557.200 29.700 ;
        RECT 566.000 30.300 566.800 30.400 ;
        RECT 583.600 30.300 584.400 30.400 ;
        RECT 566.000 29.700 584.400 30.300 ;
        RECT 566.000 29.600 566.800 29.700 ;
        RECT 583.600 29.600 584.400 29.700 ;
        RECT 598.000 30.300 598.800 30.400 ;
        RECT 622.100 30.300 622.700 31.600 ;
        RECT 598.000 29.700 622.700 30.300 ;
        RECT 630.000 30.300 630.800 30.400 ;
        RECT 649.200 30.300 650.000 30.400 ;
        RECT 662.000 30.300 662.800 30.400 ;
        RECT 674.800 30.300 675.600 30.400 ;
        RECT 630.000 29.700 675.600 30.300 ;
        RECT 598.000 29.600 598.800 29.700 ;
        RECT 630.000 29.600 630.800 29.700 ;
        RECT 649.200 29.600 650.000 29.700 ;
        RECT 662.000 29.600 662.800 29.700 ;
        RECT 674.800 29.600 675.600 29.700 ;
        RECT 14.000 28.300 14.800 28.400 ;
        RECT 42.800 28.300 43.600 28.400 ;
        RECT 14.000 27.700 43.600 28.300 ;
        RECT 14.000 27.600 14.800 27.700 ;
        RECT 42.800 27.600 43.600 27.700 ;
        RECT 46.000 28.300 46.800 28.400 ;
        RECT 58.800 28.300 59.600 28.400 ;
        RECT 46.000 27.700 59.600 28.300 ;
        RECT 46.000 27.600 46.800 27.700 ;
        RECT 58.800 27.600 59.600 27.700 ;
        RECT 92.400 28.300 93.200 28.400 ;
        RECT 98.800 28.300 99.600 28.400 ;
        RECT 105.200 28.300 106.000 28.400 ;
        RECT 137.200 28.300 138.000 28.400 ;
        RECT 92.400 27.700 138.000 28.300 ;
        RECT 92.400 27.600 93.200 27.700 ;
        RECT 98.800 27.600 99.600 27.700 ;
        RECT 105.200 27.600 106.000 27.700 ;
        RECT 137.200 27.600 138.000 27.700 ;
        RECT 142.000 28.300 142.800 28.400 ;
        RECT 153.200 28.300 154.000 28.400 ;
        RECT 177.300 28.300 177.900 29.600 ;
        RECT 142.000 27.700 177.900 28.300 ;
        RECT 180.400 28.300 181.200 28.400 ;
        RECT 185.200 28.300 186.000 28.400 ;
        RECT 196.400 28.300 197.200 28.400 ;
        RECT 180.400 27.700 197.200 28.300 ;
        RECT 142.000 27.600 142.800 27.700 ;
        RECT 153.200 27.600 154.000 27.700 ;
        RECT 180.400 27.600 181.200 27.700 ;
        RECT 185.200 27.600 186.000 27.700 ;
        RECT 196.400 27.600 197.200 27.700 ;
        RECT 198.000 28.300 198.800 28.400 ;
        RECT 218.800 28.300 219.600 28.400 ;
        RECT 198.000 27.700 219.600 28.300 ;
        RECT 198.000 27.600 198.800 27.700 ;
        RECT 218.800 27.600 219.600 27.700 ;
        RECT 273.200 28.300 274.000 28.400 ;
        RECT 276.400 28.300 277.200 28.400 ;
        RECT 284.400 28.300 285.200 28.400 ;
        RECT 303.600 28.300 304.400 28.400 ;
        RECT 313.200 28.300 314.000 28.400 ;
        RECT 273.200 27.700 314.000 28.300 ;
        RECT 273.200 27.600 274.000 27.700 ;
        RECT 276.400 27.600 277.200 27.700 ;
        RECT 284.400 27.600 285.200 27.700 ;
        RECT 303.600 27.600 304.400 27.700 ;
        RECT 313.200 27.600 314.000 27.700 ;
        RECT 366.000 28.300 366.800 28.400 ;
        RECT 401.200 28.300 402.000 28.400 ;
        RECT 415.600 28.300 416.400 28.400 ;
        RECT 426.800 28.300 427.600 28.400 ;
        RECT 366.000 27.700 427.600 28.300 ;
        RECT 366.000 27.600 366.800 27.700 ;
        RECT 401.200 27.600 402.000 27.700 ;
        RECT 415.600 27.600 416.400 27.700 ;
        RECT 426.800 27.600 427.600 27.700 ;
        RECT 444.400 28.300 445.200 28.400 ;
        RECT 470.000 28.300 470.800 28.400 ;
        RECT 444.400 27.700 470.800 28.300 ;
        RECT 444.400 27.600 445.200 27.700 ;
        RECT 470.000 27.600 470.800 27.700 ;
        RECT 503.600 28.300 504.400 28.400 ;
        RECT 537.200 28.300 538.000 28.400 ;
        RECT 503.600 27.700 538.000 28.300 ;
        RECT 503.600 27.600 504.400 27.700 ;
        RECT 537.200 27.600 538.000 27.700 ;
        RECT 538.800 28.300 539.600 28.400 ;
        RECT 540.400 28.300 541.200 28.400 ;
        RECT 538.800 27.700 541.200 28.300 ;
        RECT 538.800 27.600 539.600 27.700 ;
        RECT 540.400 27.600 541.200 27.700 ;
        RECT 550.000 28.300 550.800 28.400 ;
        RECT 559.600 28.300 560.400 28.400 ;
        RECT 550.000 27.700 560.400 28.300 ;
        RECT 550.000 27.600 550.800 27.700 ;
        RECT 559.600 27.600 560.400 27.700 ;
        RECT 591.600 28.300 592.400 28.400 ;
        RECT 604.400 28.300 605.200 28.400 ;
        RECT 591.600 27.700 605.200 28.300 ;
        RECT 591.600 27.600 592.400 27.700 ;
        RECT 604.400 27.600 605.200 27.700 ;
        RECT 617.200 28.300 618.000 28.400 ;
        RECT 618.800 28.300 619.600 28.400 ;
        RECT 630.000 28.300 630.800 28.400 ;
        RECT 617.200 27.700 630.800 28.300 ;
        RECT 617.200 27.600 618.000 27.700 ;
        RECT 618.800 27.600 619.600 27.700 ;
        RECT 630.000 27.600 630.800 27.700 ;
        RECT 647.600 28.300 648.400 28.400 ;
        RECT 658.800 28.300 659.600 28.400 ;
        RECT 647.600 27.700 659.600 28.300 ;
        RECT 647.600 27.600 648.400 27.700 ;
        RECT 658.800 27.600 659.600 27.700 ;
        RECT 660.400 28.300 661.200 28.400 ;
        RECT 673.200 28.300 674.000 28.400 ;
        RECT 660.400 27.700 674.000 28.300 ;
        RECT 660.400 27.600 661.200 27.700 ;
        RECT 673.200 27.600 674.000 27.700 ;
        RECT 674.800 28.300 675.600 28.400 ;
        RECT 676.400 28.300 677.200 28.400 ;
        RECT 674.800 27.700 677.200 28.300 ;
        RECT 674.800 27.600 675.600 27.700 ;
        RECT 676.400 27.600 677.200 27.700 ;
        RECT 38.000 26.300 38.800 26.400 ;
        RECT 97.200 26.300 98.000 26.400 ;
        RECT 38.000 25.700 98.000 26.300 ;
        RECT 38.000 25.600 38.800 25.700 ;
        RECT 97.200 25.600 98.000 25.700 ;
        RECT 111.600 26.300 112.400 26.400 ;
        RECT 126.000 26.300 126.800 26.400 ;
        RECT 142.000 26.300 142.800 26.400 ;
        RECT 111.600 25.700 142.800 26.300 ;
        RECT 111.600 25.600 112.400 25.700 ;
        RECT 126.000 25.600 126.800 25.700 ;
        RECT 142.000 25.600 142.800 25.700 ;
        RECT 174.000 26.300 174.800 26.400 ;
        RECT 182.000 26.300 182.800 26.400 ;
        RECT 174.000 25.700 182.800 26.300 ;
        RECT 174.000 25.600 174.800 25.700 ;
        RECT 182.000 25.600 182.800 25.700 ;
        RECT 257.200 26.300 258.000 26.400 ;
        RECT 292.400 26.300 293.200 26.400 ;
        RECT 257.200 25.700 293.200 26.300 ;
        RECT 257.200 25.600 258.000 25.700 ;
        RECT 292.400 25.600 293.200 25.700 ;
        RECT 308.400 26.300 309.200 26.400 ;
        RECT 334.000 26.300 334.800 26.400 ;
        RECT 308.400 25.700 334.800 26.300 ;
        RECT 308.400 25.600 309.200 25.700 ;
        RECT 334.000 25.600 334.800 25.700 ;
        RECT 466.800 26.300 467.600 26.400 ;
        RECT 489.200 26.300 490.000 26.400 ;
        RECT 498.800 26.300 499.600 26.400 ;
        RECT 534.000 26.300 534.800 26.400 ;
        RECT 466.800 25.700 534.800 26.300 ;
        RECT 466.800 25.600 467.600 25.700 ;
        RECT 489.200 25.600 490.000 25.700 ;
        RECT 498.800 25.600 499.600 25.700 ;
        RECT 534.000 25.600 534.800 25.700 ;
        RECT 535.600 26.300 536.400 26.400 ;
        RECT 540.400 26.300 541.200 26.400 ;
        RECT 535.600 25.700 541.200 26.300 ;
        RECT 535.600 25.600 536.400 25.700 ;
        RECT 540.400 25.600 541.200 25.700 ;
        RECT 636.400 26.300 637.200 26.400 ;
        RECT 660.400 26.300 661.200 26.400 ;
        RECT 636.400 25.700 661.200 26.300 ;
        RECT 636.400 25.600 637.200 25.700 ;
        RECT 660.400 25.600 661.200 25.700 ;
        RECT 673.200 26.300 674.000 26.400 ;
        RECT 687.600 26.300 688.400 26.400 ;
        RECT 673.200 25.700 688.400 26.300 ;
        RECT 673.200 25.600 674.000 25.700 ;
        RECT 687.600 25.600 688.400 25.700 ;
        RECT 260.400 24.300 261.200 24.400 ;
        RECT 265.200 24.300 266.000 24.400 ;
        RECT 260.400 23.700 266.000 24.300 ;
        RECT 260.400 23.600 261.200 23.700 ;
        RECT 265.200 23.600 266.000 23.700 ;
        RECT 314.800 24.300 315.600 24.400 ;
        RECT 321.200 24.300 322.000 24.400 ;
        RECT 314.800 23.700 322.000 24.300 ;
        RECT 314.800 23.600 315.600 23.700 ;
        RECT 321.200 23.600 322.000 23.700 ;
        RECT 375.600 24.300 376.400 24.400 ;
        RECT 404.400 24.300 405.200 24.400 ;
        RECT 375.600 23.700 405.200 24.300 ;
        RECT 375.600 23.600 376.400 23.700 ;
        RECT 404.400 23.600 405.200 23.700 ;
        RECT 673.200 24.300 674.000 24.400 ;
        RECT 681.200 24.300 682.000 24.400 ;
        RECT 673.200 23.700 682.000 24.300 ;
        RECT 673.200 23.600 674.000 23.700 ;
        RECT 681.200 23.600 682.000 23.700 ;
        RECT 337.200 22.300 338.000 22.400 ;
        RECT 362.800 22.300 363.600 22.400 ;
        RECT 337.200 21.700 363.600 22.300 ;
        RECT 337.200 21.600 338.000 21.700 ;
        RECT 362.800 21.600 363.600 21.700 ;
        RECT 614.000 22.300 614.800 22.400 ;
        RECT 649.200 22.300 650.000 22.400 ;
        RECT 614.000 21.700 650.000 22.300 ;
        RECT 614.000 21.600 614.800 21.700 ;
        RECT 649.200 21.600 650.000 21.700 ;
        RECT 63.600 20.300 64.400 20.400 ;
        RECT 68.400 20.300 69.200 20.400 ;
        RECT 63.600 19.700 69.200 20.300 ;
        RECT 63.600 19.600 64.400 19.700 ;
        RECT 68.400 19.600 69.200 19.700 ;
        RECT 94.000 20.300 94.800 20.400 ;
        RECT 103.600 20.300 104.400 20.400 ;
        RECT 94.000 19.700 104.400 20.300 ;
        RECT 94.000 19.600 94.800 19.700 ;
        RECT 103.600 19.600 104.400 19.700 ;
        RECT 145.200 20.300 146.000 20.400 ;
        RECT 164.400 20.300 165.200 20.400 ;
        RECT 178.800 20.300 179.600 20.400 ;
        RECT 145.200 19.700 179.600 20.300 ;
        RECT 145.200 19.600 146.000 19.700 ;
        RECT 164.400 19.600 165.200 19.700 ;
        RECT 178.800 19.600 179.600 19.700 ;
        RECT 353.200 20.300 354.000 20.400 ;
        RECT 359.600 20.300 360.400 20.400 ;
        RECT 377.200 20.300 378.000 20.400 ;
        RECT 388.400 20.300 389.200 20.400 ;
        RECT 396.400 20.300 397.200 20.400 ;
        RECT 353.200 19.700 397.200 20.300 ;
        RECT 353.200 19.600 354.000 19.700 ;
        RECT 359.600 19.600 360.400 19.700 ;
        RECT 377.200 19.600 378.000 19.700 ;
        RECT 388.400 19.600 389.200 19.700 ;
        RECT 396.400 19.600 397.200 19.700 ;
        RECT 441.200 20.300 442.000 20.400 ;
        RECT 447.600 20.300 448.400 20.400 ;
        RECT 474.800 20.300 475.600 20.400 ;
        RECT 484.400 20.300 485.200 20.400 ;
        RECT 513.200 20.300 514.000 20.400 ;
        RECT 521.200 20.300 522.000 20.400 ;
        RECT 441.200 19.700 522.000 20.300 ;
        RECT 441.200 19.600 442.000 19.700 ;
        RECT 447.600 19.600 448.400 19.700 ;
        RECT 474.800 19.600 475.600 19.700 ;
        RECT 484.400 19.600 485.200 19.700 ;
        RECT 513.200 19.600 514.000 19.700 ;
        RECT 521.200 19.600 522.000 19.700 ;
        RECT 625.200 20.300 626.000 20.400 ;
        RECT 642.800 20.300 643.600 20.400 ;
        RECT 625.200 19.700 643.600 20.300 ;
        RECT 625.200 19.600 626.000 19.700 ;
        RECT 642.800 19.600 643.600 19.700 ;
        RECT 166.000 18.300 166.800 18.400 ;
        RECT 183.600 18.300 184.400 18.400 ;
        RECT 217.200 18.300 218.000 18.400 ;
        RECT 166.000 17.700 218.000 18.300 ;
        RECT 166.000 17.600 166.800 17.700 ;
        RECT 183.600 17.600 184.400 17.700 ;
        RECT 217.200 17.600 218.000 17.700 ;
        RECT 266.800 18.300 267.600 18.400 ;
        RECT 271.600 18.300 272.400 18.400 ;
        RECT 266.800 17.700 272.400 18.300 ;
        RECT 266.800 17.600 267.600 17.700 ;
        RECT 271.600 17.600 272.400 17.700 ;
        RECT 290.800 18.300 291.600 18.400 ;
        RECT 300.400 18.300 301.200 18.400 ;
        RECT 318.000 18.300 318.800 18.400 ;
        RECT 330.800 18.300 331.600 18.400 ;
        RECT 290.800 17.700 331.600 18.300 ;
        RECT 290.800 17.600 291.600 17.700 ;
        RECT 300.400 17.600 301.200 17.700 ;
        RECT 318.000 17.600 318.800 17.700 ;
        RECT 330.800 17.600 331.600 17.700 ;
        RECT 546.800 18.300 547.600 18.400 ;
        RECT 575.600 18.300 576.400 18.400 ;
        RECT 546.800 17.700 576.400 18.300 ;
        RECT 546.800 17.600 547.600 17.700 ;
        RECT 575.600 17.600 576.400 17.700 ;
        RECT 588.400 18.300 589.200 18.400 ;
        RECT 596.400 18.300 597.200 18.400 ;
        RECT 614.000 18.300 614.800 18.400 ;
        RECT 588.400 17.700 614.800 18.300 ;
        RECT 588.400 17.600 589.200 17.700 ;
        RECT 596.400 17.600 597.200 17.700 ;
        RECT 614.000 17.600 614.800 17.700 ;
        RECT 628.400 18.300 629.200 18.400 ;
        RECT 641.200 18.300 642.000 18.400 ;
        RECT 628.400 17.700 642.000 18.300 ;
        RECT 628.400 17.600 629.200 17.700 ;
        RECT 641.200 17.600 642.000 17.700 ;
        RECT 654.000 18.300 654.800 18.400 ;
        RECT 662.000 18.300 662.800 18.400 ;
        RECT 654.000 17.700 662.800 18.300 ;
        RECT 654.000 17.600 654.800 17.700 ;
        RECT 662.000 17.600 662.800 17.700 ;
        RECT 17.200 16.300 18.000 16.400 ;
        RECT 20.400 16.300 21.200 16.400 ;
        RECT 65.200 16.300 66.000 16.400 ;
        RECT 17.200 15.700 66.000 16.300 ;
        RECT 17.200 15.600 18.000 15.700 ;
        RECT 20.400 15.600 21.200 15.700 ;
        RECT 65.200 15.600 66.000 15.700 ;
        RECT 90.800 16.300 91.600 16.400 ;
        RECT 100.400 16.300 101.200 16.400 ;
        RECT 124.400 16.300 125.200 16.400 ;
        RECT 90.800 15.700 125.200 16.300 ;
        RECT 90.800 15.600 91.600 15.700 ;
        RECT 100.400 15.600 101.200 15.700 ;
        RECT 124.400 15.600 125.200 15.700 ;
        RECT 146.800 16.300 147.600 16.400 ;
        RECT 159.600 16.300 160.400 16.400 ;
        RECT 167.600 16.300 168.400 16.400 ;
        RECT 174.000 16.300 174.800 16.400 ;
        RECT 146.800 15.700 174.800 16.300 ;
        RECT 146.800 15.600 147.600 15.700 ;
        RECT 159.600 15.600 160.400 15.700 ;
        RECT 167.600 15.600 168.400 15.700 ;
        RECT 174.000 15.600 174.800 15.700 ;
        RECT 196.400 16.300 197.200 16.400 ;
        RECT 207.600 16.300 208.400 16.400 ;
        RECT 196.400 15.700 208.400 16.300 ;
        RECT 196.400 15.600 197.200 15.700 ;
        RECT 207.600 15.600 208.400 15.700 ;
        RECT 214.000 16.300 214.800 16.400 ;
        RECT 244.400 16.300 245.200 16.400 ;
        RECT 214.000 15.700 245.200 16.300 ;
        RECT 214.000 15.600 214.800 15.700 ;
        RECT 244.400 15.600 245.200 15.700 ;
        RECT 250.800 16.300 251.600 16.400 ;
        RECT 276.400 16.300 277.200 16.400 ;
        RECT 250.800 15.700 277.200 16.300 ;
        RECT 250.800 15.600 251.600 15.700 ;
        RECT 276.400 15.600 277.200 15.700 ;
        RECT 282.800 16.300 283.600 16.400 ;
        RECT 303.600 16.300 304.400 16.400 ;
        RECT 282.800 15.700 304.400 16.300 ;
        RECT 282.800 15.600 283.600 15.700 ;
        RECT 303.600 15.600 304.400 15.700 ;
        RECT 393.200 16.300 394.000 16.400 ;
        RECT 417.200 16.300 418.000 16.400 ;
        RECT 393.200 15.700 418.000 16.300 ;
        RECT 393.200 15.600 394.000 15.700 ;
        RECT 417.200 15.600 418.000 15.700 ;
        RECT 559.600 16.300 560.400 16.400 ;
        RECT 582.000 16.300 582.800 16.400 ;
        RECT 559.600 15.700 582.800 16.300 ;
        RECT 559.600 15.600 560.400 15.700 ;
        RECT 582.000 15.600 582.800 15.700 ;
        RECT 607.600 16.300 608.400 16.400 ;
        RECT 628.400 16.300 629.200 16.400 ;
        RECT 607.600 15.700 629.200 16.300 ;
        RECT 607.600 15.600 608.400 15.700 ;
        RECT 628.400 15.600 629.200 15.700 ;
        RECT 630.000 16.300 630.800 16.400 ;
        RECT 639.600 16.300 640.400 16.400 ;
        RECT 630.000 15.700 640.400 16.300 ;
        RECT 630.000 15.600 630.800 15.700 ;
        RECT 639.600 15.600 640.400 15.700 ;
        RECT 2.800 14.300 3.600 14.400 ;
        RECT 17.200 14.300 18.000 14.400 ;
        RECT 2.800 13.700 18.000 14.300 ;
        RECT 2.800 13.600 3.600 13.700 ;
        RECT 17.200 13.600 18.000 13.700 ;
        RECT 44.400 14.300 45.200 14.400 ;
        RECT 50.800 14.300 51.600 14.400 ;
        RECT 84.400 14.300 85.200 14.400 ;
        RECT 89.200 14.300 90.000 14.400 ;
        RECT 44.400 13.700 90.000 14.300 ;
        RECT 44.400 13.600 45.200 13.700 ;
        RECT 50.800 13.600 51.600 13.700 ;
        RECT 84.400 13.600 85.200 13.700 ;
        RECT 89.200 13.600 90.000 13.700 ;
        RECT 156.400 14.300 157.200 14.400 ;
        RECT 186.800 14.300 187.600 14.400 ;
        RECT 156.400 13.700 187.600 14.300 ;
        RECT 156.400 13.600 157.200 13.700 ;
        RECT 186.800 13.600 187.600 13.700 ;
        RECT 236.400 14.300 237.200 14.400 ;
        RECT 239.600 14.300 240.400 14.400 ;
        RECT 236.400 13.700 240.400 14.300 ;
        RECT 236.400 13.600 237.200 13.700 ;
        RECT 239.600 13.600 240.400 13.700 ;
        RECT 273.200 14.300 274.000 14.400 ;
        RECT 282.800 14.300 283.600 14.400 ;
        RECT 273.200 13.700 283.600 14.300 ;
        RECT 273.200 13.600 274.000 13.700 ;
        RECT 282.800 13.600 283.600 13.700 ;
        RECT 356.400 14.300 357.200 14.400 ;
        RECT 369.200 14.300 370.000 14.400 ;
        RECT 356.400 13.700 370.000 14.300 ;
        RECT 356.400 13.600 357.200 13.700 ;
        RECT 369.200 13.600 370.000 13.700 ;
        RECT 412.400 14.300 413.200 14.400 ;
        RECT 418.800 14.300 419.600 14.400 ;
        RECT 430.000 14.300 430.800 14.400 ;
        RECT 412.400 13.700 430.800 14.300 ;
        RECT 412.400 13.600 413.200 13.700 ;
        RECT 418.800 13.600 419.600 13.700 ;
        RECT 430.000 13.600 430.800 13.700 ;
        RECT 438.000 14.300 438.800 14.400 ;
        RECT 458.800 14.300 459.600 14.400 ;
        RECT 438.000 13.700 459.600 14.300 ;
        RECT 438.000 13.600 438.800 13.700 ;
        RECT 458.800 13.600 459.600 13.700 ;
        RECT 518.000 14.300 518.800 14.400 ;
        RECT 538.800 14.300 539.600 14.400 ;
        RECT 518.000 13.700 539.600 14.300 ;
        RECT 518.000 13.600 518.800 13.700 ;
        RECT 538.800 13.600 539.600 13.700 ;
        RECT 628.400 14.300 629.200 14.400 ;
        RECT 631.600 14.300 632.400 14.400 ;
        RECT 628.400 13.700 632.400 14.300 ;
        RECT 628.400 13.600 629.200 13.700 ;
        RECT 631.600 13.600 632.400 13.700 ;
        RECT 658.800 14.300 659.600 14.400 ;
        RECT 670.000 14.300 670.800 14.400 ;
        RECT 658.800 13.700 670.800 14.300 ;
        RECT 658.800 13.600 659.600 13.700 ;
        RECT 670.000 13.600 670.800 13.700 ;
        RECT 28.400 12.300 29.200 12.400 ;
        RECT 57.200 12.300 58.000 12.400 ;
        RECT 28.400 11.700 58.000 12.300 ;
        RECT 28.400 11.600 29.200 11.700 ;
        RECT 57.200 11.600 58.000 11.700 ;
        RECT 78.000 12.300 78.800 12.400 ;
        RECT 92.400 12.300 93.200 12.400 ;
        RECT 78.000 11.700 93.200 12.300 ;
        RECT 78.000 11.600 78.800 11.700 ;
        RECT 92.400 11.600 93.200 11.700 ;
        RECT 225.200 12.300 226.000 12.400 ;
        RECT 234.800 12.300 235.600 12.400 ;
        RECT 225.200 11.700 235.600 12.300 ;
        RECT 225.200 11.600 226.000 11.700 ;
        RECT 234.800 11.600 235.600 11.700 ;
        RECT 238.000 12.300 238.800 12.400 ;
        RECT 247.600 12.300 248.400 12.400 ;
        RECT 238.000 11.700 248.400 12.300 ;
        RECT 238.000 11.600 238.800 11.700 ;
        RECT 247.600 11.600 248.400 11.700 ;
        RECT 313.200 12.300 314.000 12.400 ;
        RECT 324.400 12.300 325.200 12.400 ;
        RECT 313.200 11.700 325.200 12.300 ;
        RECT 313.200 11.600 314.000 11.700 ;
        RECT 324.400 11.600 325.200 11.700 ;
        RECT 366.000 12.300 366.800 12.400 ;
        RECT 378.800 12.300 379.600 12.400 ;
        RECT 383.600 12.300 384.400 12.400 ;
        RECT 366.000 11.700 384.400 12.300 ;
        RECT 366.000 11.600 366.800 11.700 ;
        RECT 378.800 11.600 379.600 11.700 ;
        RECT 383.600 11.600 384.400 11.700 ;
        RECT 404.400 12.300 405.200 12.400 ;
        RECT 428.400 12.300 429.200 12.400 ;
        RECT 404.400 11.700 429.200 12.300 ;
        RECT 404.400 11.600 405.200 11.700 ;
        RECT 428.400 11.600 429.200 11.700 ;
        RECT 449.200 12.300 450.000 12.400 ;
        RECT 476.400 12.300 477.200 12.400 ;
        RECT 449.200 11.700 477.200 12.300 ;
        RECT 449.200 11.600 450.000 11.700 ;
        RECT 476.400 11.600 477.200 11.700 ;
        RECT 498.800 12.300 499.600 12.400 ;
        RECT 505.200 12.300 506.000 12.400 ;
        RECT 508.400 12.300 509.200 12.400 ;
        RECT 498.800 11.700 509.200 12.300 ;
        RECT 498.800 11.600 499.600 11.700 ;
        RECT 505.200 11.600 506.000 11.700 ;
        RECT 508.400 11.600 509.200 11.700 ;
        RECT 529.200 12.300 530.000 12.400 ;
        RECT 546.800 12.300 547.600 12.400 ;
        RECT 529.200 11.700 547.600 12.300 ;
        RECT 529.200 11.600 530.000 11.700 ;
        RECT 546.800 11.600 547.600 11.700 ;
        RECT 602.800 12.300 603.600 12.400 ;
        RECT 639.600 12.300 640.400 12.400 ;
        RECT 602.800 11.700 640.400 12.300 ;
        RECT 602.800 11.600 603.600 11.700 ;
        RECT 639.600 11.600 640.400 11.700 ;
        RECT 655.600 12.300 656.400 12.400 ;
        RECT 673.200 12.300 674.000 12.400 ;
        RECT 655.600 11.700 674.000 12.300 ;
        RECT 655.600 11.600 656.400 11.700 ;
        RECT 673.200 11.600 674.000 11.700 ;
        RECT 682.800 12.300 683.600 12.400 ;
        RECT 684.400 12.300 685.200 12.400 ;
        RECT 682.800 11.700 685.200 12.300 ;
        RECT 682.800 11.600 683.600 11.700 ;
        RECT 684.400 11.600 685.200 11.700 ;
        RECT 111.600 10.300 112.400 10.400 ;
        RECT 202.800 10.300 203.600 10.400 ;
        RECT 111.600 9.700 203.600 10.300 ;
        RECT 111.600 9.600 112.400 9.700 ;
        RECT 202.800 9.600 203.600 9.700 ;
        RECT 244.400 10.300 245.200 10.400 ;
        RECT 250.800 10.300 251.600 10.400 ;
        RECT 244.400 9.700 251.600 10.300 ;
        RECT 244.400 9.600 245.200 9.700 ;
        RECT 250.800 9.600 251.600 9.700 ;
        RECT 254.000 10.300 254.800 10.400 ;
        RECT 260.400 10.300 261.200 10.400 ;
        RECT 254.000 9.700 261.200 10.300 ;
        RECT 254.000 9.600 254.800 9.700 ;
        RECT 260.400 9.600 261.200 9.700 ;
        RECT 281.200 10.300 282.000 10.400 ;
        RECT 286.000 10.300 286.800 10.400 ;
        RECT 281.200 9.700 286.800 10.300 ;
        RECT 281.200 9.600 282.000 9.700 ;
        RECT 286.000 9.600 286.800 9.700 ;
        RECT 601.200 10.300 602.000 10.400 ;
        RECT 609.200 10.300 610.000 10.400 ;
        RECT 601.200 9.700 610.000 10.300 ;
        RECT 601.200 9.600 602.000 9.700 ;
        RECT 609.200 9.600 610.000 9.700 ;
        RECT 630.000 10.300 630.800 10.400 ;
        RECT 654.000 10.300 654.800 10.400 ;
        RECT 630.000 9.700 654.800 10.300 ;
        RECT 630.000 9.600 630.800 9.700 ;
        RECT 654.000 9.600 654.800 9.700 ;
        RECT 679.600 10.300 680.400 10.400 ;
        RECT 681.200 10.300 682.000 10.400 ;
        RECT 679.600 9.700 682.000 10.300 ;
        RECT 679.600 9.600 680.400 9.700 ;
        RECT 681.200 9.600 682.000 9.700 ;
        RECT 623.600 8.300 624.400 8.400 ;
        RECT 636.400 8.300 637.200 8.400 ;
        RECT 623.600 7.700 637.200 8.300 ;
        RECT 623.600 7.600 624.400 7.700 ;
        RECT 636.400 7.600 637.200 7.700 ;
      LAYER metal4 ;
        RECT 42.600 435.400 43.800 456.600 ;
        RECT 29.800 399.400 31.000 416.600 ;
        RECT 33.000 385.400 34.200 432.600 ;
        RECT 36.200 377.400 37.400 430.600 ;
        RECT 17.000 265.400 18.200 330.600 ;
        RECT 45.800 315.400 47.000 490.600 ;
        RECT 65.000 419.400 66.200 450.600 ;
        RECT 58.600 389.400 59.800 418.600 ;
        RECT 61.800 305.400 63.000 410.600 ;
        RECT 65.000 387.400 66.200 408.600 ;
        RECT 68.200 335.400 69.400 398.600 ;
        RECT 71.400 375.400 72.600 396.600 ;
        RECT 77.800 353.400 79.000 422.600 ;
        RECT 87.400 283.400 88.600 424.600 ;
        RECT 90.600 351.400 91.800 420.600 ;
        RECT 93.800 371.400 95.000 468.600 ;
        RECT 161.000 427.400 162.200 464.600 ;
        RECT 164.200 423.400 165.400 454.600 ;
        RECT 103.400 391.400 104.600 420.600 ;
        RECT 170.600 415.400 171.800 454.600 ;
        RECT 276.200 443.400 277.400 472.600 ;
        RECT 125.800 353.400 127.000 406.600 ;
        RECT 138.600 345.400 139.800 388.600 ;
        RECT 141.800 385.400 143.000 394.600 ;
        RECT 177.000 391.400 178.200 412.600 ;
        RECT 151.400 357.400 152.600 386.600 ;
        RECT 93.800 321.400 95.000 338.600 ;
        RECT 154.600 333.400 155.800 338.600 ;
        RECT 167.400 329.400 168.600 350.600 ;
        RECT 106.600 215.400 107.800 256.600 ;
        RECT 122.600 237.400 123.800 260.600 ;
        RECT 157.800 255.400 159.000 278.600 ;
        RECT 186.600 265.400 187.800 306.600 ;
        RECT 189.800 297.400 191.000 318.600 ;
        RECT 138.600 211.400 139.800 222.600 ;
        RECT 157.800 217.400 159.000 226.600 ;
        RECT 13.800 149.400 15.000 184.600 ;
        RECT 17.000 147.400 18.200 188.600 ;
        RECT 20.200 55.400 21.400 70.600 ;
        RECT 29.800 53.400 31.000 174.600 ;
        RECT 36.200 111.400 37.400 158.600 ;
        RECT 42.600 99.400 43.800 166.600 ;
        RECT 52.200 49.400 53.400 170.600 ;
        RECT 90.600 163.400 91.800 190.600 ;
        RECT 100.200 131.400 101.400 146.600 ;
        RECT 122.600 127.400 123.800 134.600 ;
        RECT 100.200 95.400 101.400 106.600 ;
        RECT 103.400 105.400 104.600 124.600 ;
        RECT 90.600 49.400 91.800 72.600 ;
        RECT 125.800 71.400 127.000 112.600 ;
        RECT 135.400 83.400 136.600 94.600 ;
        RECT 141.800 49.400 143.000 78.600 ;
        RECT 148.200 51.400 149.400 164.600 ;
        RECT 157.800 41.400 159.000 172.600 ;
        RECT 173.800 143.400 175.000 184.600 ;
        RECT 202.600 173.400 203.800 390.600 ;
        RECT 212.200 331.400 213.400 380.600 ;
        RECT 241.000 337.400 242.200 386.600 ;
        RECT 269.800 345.400 271.000 420.600 ;
        RECT 273.000 353.400 274.200 428.600 ;
        RECT 285.800 371.400 287.000 404.600 ;
        RECT 292.200 375.400 293.400 418.600 ;
        RECT 295.400 381.400 296.600 460.600 ;
        RECT 305.000 427.400 306.200 456.600 ;
        RECT 333.800 419.400 335.000 430.600 ;
        RECT 343.400 421.400 344.600 466.600 ;
        RECT 346.600 423.400 347.800 438.600 ;
        RECT 301.800 351.400 303.000 388.600 ;
        RECT 314.600 355.400 315.800 406.600 ;
        RECT 215.400 283.400 216.600 304.600 ;
        RECT 279.400 293.400 280.600 312.600 ;
        RECT 311.400 311.400 312.600 354.600 ;
        RECT 317.800 351.400 319.000 382.600 ;
        RECT 321.000 339.400 322.200 378.600 ;
        RECT 324.200 365.400 325.400 416.600 ;
        RECT 327.400 353.400 328.600 412.600 ;
        RECT 340.200 371.400 341.400 404.600 ;
        RECT 359.400 387.400 360.600 412.600 ;
        RECT 365.800 403.400 367.000 438.600 ;
        RECT 369.000 435.400 370.200 452.600 ;
        RECT 381.800 435.400 383.000 466.600 ;
        RECT 372.200 407.400 373.400 434.600 ;
        RECT 385.000 407.400 386.200 428.600 ;
        RECT 330.600 333.400 331.800 354.600 ;
        RECT 333.800 343.400 335.000 358.600 ;
        RECT 346.600 355.400 347.800 386.600 ;
        RECT 362.600 371.400 363.800 394.600 ;
        RECT 237.800 231.400 239.000 278.600 ;
        RECT 260.200 215.400 261.400 244.600 ;
        RECT 273.000 211.400 274.200 268.600 ;
        RECT 285.800 241.400 287.000 268.600 ;
        RECT 177.000 85.400 178.200 142.600 ;
        RECT 279.400 141.400 280.600 174.600 ;
        RECT 285.800 139.400 287.000 226.600 ;
        RECT 289.000 215.400 290.200 250.600 ;
        RECT 292.200 245.400 293.400 272.600 ;
        RECT 295.400 241.400 296.600 260.600 ;
        RECT 314.600 251.400 315.800 276.600 ;
        RECT 321.000 213.400 322.200 248.600 ;
        RECT 324.200 225.400 325.400 248.600 ;
        RECT 327.400 211.400 328.600 246.600 ;
        RECT 330.600 235.400 331.800 254.600 ;
        RECT 337.000 243.400 338.200 318.600 ;
        RECT 340.200 241.400 341.400 272.600 ;
        RECT 189.800 65.400 191.000 112.600 ;
        RECT 193.000 109.400 194.200 132.600 ;
        RECT 237.800 77.400 239.000 114.600 ;
        RECT 193.000 55.400 194.200 72.600 ;
        RECT 247.400 55.400 248.600 94.600 ;
        RECT 260.200 9.400 261.400 80.600 ;
        RECT 273.000 69.400 274.200 132.600 ;
        RECT 276.200 63.400 277.400 128.600 ;
        RECT 295.400 95.400 296.600 136.600 ;
        RECT 305.000 109.400 306.200 148.600 ;
        RECT 308.200 113.400 309.400 186.600 ;
        RECT 343.400 169.400 344.600 224.600 ;
        RECT 346.600 173.400 347.800 344.600 ;
        RECT 349.800 321.400 351.000 358.600 ;
        RECT 365.800 357.400 367.000 380.600 ;
        RECT 349.800 257.400 351.000 280.600 ;
        RECT 353.000 265.400 354.200 306.600 ;
        RECT 356.200 153.400 357.400 350.600 ;
        RECT 359.400 271.400 360.600 308.600 ;
        RECT 365.800 275.400 367.000 346.600 ;
        RECT 375.400 317.400 376.600 362.600 ;
        RECT 369.000 235.400 370.200 260.600 ;
        RECT 372.200 221.400 373.400 286.600 ;
        RECT 375.400 265.400 376.600 270.600 ;
        RECT 375.400 197.400 376.600 224.600 ;
        RECT 375.400 141.400 376.600 194.600 ;
        RECT 378.600 137.400 379.800 292.600 ;
        RECT 381.800 197.400 383.000 276.600 ;
        RECT 385.000 269.400 386.200 370.600 ;
        RECT 385.000 115.400 386.200 228.600 ;
        RECT 388.200 213.400 389.400 452.600 ;
        RECT 397.800 425.400 399.000 472.600 ;
        RECT 391.400 335.400 392.600 416.600 ;
        RECT 397.800 381.400 399.000 414.600 ;
        RECT 477.800 395.400 479.000 450.600 ;
        RECT 391.400 211.400 392.600 252.600 ;
        RECT 404.200 219.400 405.400 292.600 ;
        RECT 410.600 273.400 411.800 368.600 ;
        RECT 429.800 347.400 431.000 388.600 ;
        RECT 426.600 249.400 427.800 330.600 ;
        RECT 436.200 255.400 437.400 296.600 ;
        RECT 401.000 123.400 402.200 186.600 ;
        RECT 321.000 81.400 322.200 112.600 ;
        RECT 404.200 89.400 405.400 190.600 ;
        RECT 410.600 183.400 411.800 220.600 ;
        RECT 426.600 197.400 427.800 208.600 ;
        RECT 433.000 131.400 434.200 212.600 ;
        RECT 436.200 187.400 437.400 208.600 ;
        RECT 445.800 187.400 447.000 258.600 ;
        RECT 455.400 257.400 456.600 296.600 ;
        RECT 471.400 289.400 472.600 330.600 ;
        RECT 477.800 327.400 479.000 348.600 ;
        RECT 481.000 335.400 482.200 396.600 ;
        RECT 506.600 389.400 507.800 428.600 ;
        RECT 532.200 403.400 533.400 432.600 ;
        RECT 519.400 385.400 520.600 394.600 ;
        RECT 535.400 385.400 536.600 428.600 ;
        RECT 442.600 53.400 443.800 116.600 ;
        RECT 449.000 69.400 450.200 118.600 ;
        RECT 458.600 95.400 459.800 160.600 ;
        RECT 484.200 155.400 485.400 176.600 ;
        RECT 490.600 175.400 491.800 380.600 ;
        RECT 493.800 329.400 495.000 384.600 ;
        RECT 506.600 279.400 507.800 328.600 ;
        RECT 522.600 291.400 523.800 354.600 ;
        RECT 538.600 339.400 539.800 360.600 ;
        RECT 541.800 329.400 543.000 426.600 ;
        RECT 548.200 407.400 549.400 484.600 ;
        RECT 545.000 291.400 546.200 342.600 ;
        RECT 548.200 251.400 549.400 262.600 ;
        RECT 551.400 257.400 552.600 408.600 ;
        RECT 557.800 351.400 559.000 432.600 ;
        RECT 561.000 413.400 562.200 428.600 ;
        RECT 596.200 415.400 597.400 450.600 ;
        RECT 567.400 407.400 568.600 414.600 ;
        RECT 557.800 335.400 559.000 344.600 ;
        RECT 561.000 313.400 562.200 384.600 ;
        RECT 567.400 377.400 568.600 382.600 ;
        RECT 564.200 323.400 565.400 360.600 ;
        RECT 586.600 349.400 587.800 384.600 ;
        RECT 589.800 375.400 591.000 396.600 ;
        RECT 557.800 297.400 559.000 310.600 ;
        RECT 599.400 283.400 600.600 310.600 ;
        RECT 503.400 95.400 504.600 164.600 ;
        RECT 506.600 131.400 507.800 162.600 ;
        RECT 519.400 111.400 520.600 168.600 ;
        RECT 525.800 115.400 527.000 170.600 ;
        RECT 529.000 51.400 530.200 164.600 ;
        RECT 532.200 107.400 533.400 180.600 ;
        RECT 567.400 165.400 568.600 184.600 ;
        RECT 545.000 149.400 546.200 154.600 ;
        RECT 580.200 151.400 581.400 164.600 ;
        RECT 567.400 135.400 568.600 150.600 ;
        RECT 583.400 149.400 584.600 170.600 ;
        RECT 593.000 145.400 594.200 160.600 ;
        RECT 535.400 63.400 536.600 96.600 ;
        RECT 541.800 69.400 543.000 134.600 ;
        RECT 593.000 127.400 594.200 132.600 ;
        RECT 596.200 131.400 597.400 146.600 ;
        RECT 557.800 51.400 559.000 66.600 ;
        RECT 567.400 59.400 568.600 82.600 ;
        RECT 580.200 53.400 581.400 116.600 ;
        RECT 583.400 103.400 584.600 114.600 ;
        RECT 583.400 47.400 584.600 96.600 ;
        RECT 599.400 61.400 600.600 212.600 ;
        RECT 538.600 13.400 539.800 28.600 ;
        RECT 602.600 11.400 603.800 292.600 ;
        RECT 605.800 163.400 607.000 356.600 ;
        RECT 615.400 307.400 616.600 424.600 ;
        RECT 618.600 197.400 619.800 378.600 ;
        RECT 628.200 373.400 629.400 450.600 ;
        RECT 631.400 429.400 632.600 448.600 ;
        RECT 631.400 345.400 632.600 374.600 ;
        RECT 634.600 267.400 635.800 386.600 ;
        RECT 637.800 375.400 639.000 402.600 ;
        RECT 637.800 335.400 639.000 354.600 ;
        RECT 641.000 305.400 642.200 390.600 ;
        RECT 641.000 251.400 642.200 272.600 ;
        RECT 609.000 99.400 610.200 164.600 ;
        RECT 612.200 131.400 613.400 186.600 ;
        RECT 612.200 59.400 613.400 96.600 ;
        RECT 621.800 77.400 623.000 150.600 ;
        RECT 628.200 17.400 629.400 114.600 ;
        RECT 634.600 113.400 635.800 198.600 ;
        RECT 644.200 191.400 645.400 470.600 ;
        RECT 650.600 441.400 651.800 468.600 ;
        RECT 647.400 187.400 648.600 368.600 ;
        RECT 634.600 91.400 635.800 110.600 ;
        RECT 641.000 51.400 642.200 100.600 ;
        RECT 650.600 93.400 651.800 400.600 ;
        RECT 653.800 343.400 655.000 472.600 ;
        RECT 657.000 373.400 658.200 458.600 ;
        RECT 653.800 253.400 655.000 306.600 ;
        RECT 657.000 249.400 658.200 368.600 ;
        RECT 660.200 269.400 661.400 352.600 ;
        RECT 663.400 347.400 664.600 450.600 ;
        RECT 669.800 415.400 671.000 470.600 ;
        RECT 653.800 195.400 655.000 240.600 ;
        RECT 657.000 145.400 658.200 194.600 ;
        RECT 653.800 69.400 655.000 116.600 ;
        RECT 657.000 45.400 658.200 96.600 ;
        RECT 660.200 25.400 661.400 236.600 ;
        RECT 663.400 195.400 664.600 336.600 ;
        RECT 666.600 305.400 667.800 348.600 ;
        RECT 669.800 293.400 671.000 358.600 ;
        RECT 666.600 249.400 667.800 260.600 ;
        RECT 663.400 177.400 664.600 186.600 ;
        RECT 663.400 33.400 664.600 152.600 ;
        RECT 666.600 129.400 667.800 178.600 ;
        RECT 669.800 163.400 671.000 290.600 ;
        RECT 673.000 65.400 674.200 464.600 ;
        RECT 676.200 289.400 677.400 416.600 ;
        RECT 679.400 243.400 680.600 374.600 ;
        RECT 682.600 235.400 683.800 414.600 ;
        RECT 673.000 23.400 674.200 44.600 ;
        RECT 676.200 27.400 677.400 194.600 ;
        RECT 679.400 175.400 680.600 206.600 ;
        RECT 679.400 73.400 680.600 168.600 ;
        RECT 682.600 153.400 683.800 200.600 ;
        RECT 679.400 9.400 680.600 58.600 ;
        RECT 682.600 11.400 683.800 100.600 ;
        RECT 685.800 47.400 687.000 230.600 ;
  END
END noc_top
END LIBRARY


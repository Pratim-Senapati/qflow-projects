VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 1.900 4.000 ;
  SIZE 90.200 BY 68.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 4.400 52.400 5.200 59.800 ;
        RECT 1.200 41.600 2.000 50.400 ;
        RECT 4.400 50.200 5.000 52.400 ;
        RECT 7.600 52.300 8.400 53.200 ;
        RECT 12.400 52.300 13.200 52.400 ;
        RECT 7.600 51.700 13.200 52.300 ;
        RECT 7.600 51.600 8.400 51.700 ;
        RECT 12.400 51.600 13.200 51.700 ;
        RECT 43.400 50.800 44.200 51.000 ;
        RECT 17.200 50.200 44.200 50.800 ;
        RECT 4.400 44.300 5.200 50.200 ;
        RECT 17.200 49.600 18.000 50.200 ;
        RECT 20.400 50.000 21.400 50.200 ;
        RECT 6.000 44.300 6.800 49.000 ;
        RECT 12.400 46.300 13.200 46.400 ;
        RECT 12.400 46.200 14.700 46.300 ;
        RECT 12.400 45.700 14.800 46.200 ;
        RECT 12.400 45.600 13.200 45.700 ;
        RECT 4.400 43.700 6.800 44.300 ;
        RECT 4.400 42.200 5.200 43.700 ;
        RECT 6.000 41.600 6.800 43.700 ;
        RECT 14.000 41.600 14.800 45.700 ;
        RECT 17.200 41.600 18.000 46.200 ;
        RECT 20.400 41.600 21.200 46.200 ;
        RECT 26.800 41.600 27.600 46.200 ;
        RECT 30.000 41.600 30.800 46.200 ;
        RECT 38.000 41.600 38.800 46.200 ;
        RECT 41.200 41.600 42.000 46.200 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 47.600 41.600 48.400 46.200 ;
        RECT 50.800 41.600 51.800 48.800 ;
        RECT 57.000 42.200 58.000 48.800 ;
        RECT 57.000 41.600 57.800 42.200 ;
        RECT 66.800 41.600 67.600 49.000 ;
        RECT 71.600 41.600 72.400 49.000 ;
        RECT 76.400 41.600 77.200 49.000 ;
        RECT 81.200 41.600 82.000 46.200 ;
        RECT 0.400 40.400 86.000 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 4.400 35.800 5.200 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 14.000 35.800 14.800 40.400 ;
        RECT 17.200 35.800 18.000 40.400 ;
        RECT 25.200 35.800 26.000 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 42.800 33.200 43.800 40.400 ;
        RECT 49.000 39.800 49.800 40.400 ;
        RECT 49.000 33.200 50.000 39.800 ;
        RECT 52.400 35.800 53.200 40.400 ;
        RECT 4.400 31.800 5.200 32.400 ;
        RECT 7.800 31.800 8.600 32.000 ;
        RECT 58.800 31.800 59.600 40.400 ;
        RECT 68.400 33.000 69.200 40.400 ;
        RECT 71.600 35.800 72.400 40.400 ;
        RECT 74.800 36.200 75.600 40.400 ;
        RECT 79.600 33.000 80.400 40.400 ;
        RECT 4.400 31.200 31.400 31.800 ;
        RECT 30.600 31.000 31.400 31.200 ;
        RECT 30.600 10.800 31.400 11.000 ;
        RECT 80.200 10.800 81.000 11.000 ;
        RECT 4.400 10.200 31.400 10.800 ;
        RECT 54.000 10.200 81.000 10.800 ;
        RECT 4.400 9.600 5.200 10.200 ;
        RECT 7.800 10.000 8.600 10.200 ;
        RECT 54.000 9.600 54.800 10.200 ;
        RECT 57.200 10.000 58.200 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 14.000 1.600 14.800 6.200 ;
        RECT 17.200 1.600 18.000 6.200 ;
        RECT 25.200 1.600 26.000 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 42.800 1.600 43.600 9.000 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 54.000 1.600 54.800 6.200 ;
        RECT 57.200 1.600 58.000 6.200 ;
        RECT 63.600 1.600 64.400 6.200 ;
        RECT 66.800 1.600 67.600 6.200 ;
        RECT 74.800 1.600 75.600 6.200 ;
        RECT 78.000 1.600 78.800 6.200 ;
        RECT 81.200 1.600 82.000 6.200 ;
        RECT 84.400 1.600 85.200 6.200 ;
        RECT 0.400 0.400 86.000 1.600 ;
      LAYER via1 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 20.400 45.400 21.200 46.200 ;
        RECT 27.000 40.600 27.800 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 29.800 40.600 30.600 41.400 ;
        RECT 4.400 37.600 5.200 38.400 ;
        RECT 4.400 31.600 5.200 32.400 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 57.200 5.400 58.000 6.200 ;
        RECT 27.000 0.600 27.800 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 29.800 0.600 30.600 1.400 ;
      LAYER metal2 ;
        RECT 1.200 51.600 2.000 52.400 ;
        RECT 12.400 51.600 13.200 52.400 ;
        RECT 1.300 50.400 1.900 51.600 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 12.500 46.400 13.100 51.600 ;
        RECT 20.400 50.000 21.200 50.800 ;
        RECT 12.400 45.600 13.200 46.400 ;
        RECT 20.500 46.200 21.100 50.000 ;
        RECT 20.400 45.400 21.200 46.200 ;
        RECT 26.400 40.600 31.200 41.400 ;
        RECT 4.400 37.600 5.200 38.400 ;
        RECT 4.500 32.400 5.100 37.600 ;
        RECT 4.400 31.600 5.200 32.400 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 57.200 10.000 58.000 10.800 ;
        RECT 4.500 4.400 5.100 9.600 ;
        RECT 57.300 6.200 57.900 10.000 ;
        RECT 57.200 5.400 58.000 6.200 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 26.400 0.600 31.200 1.400 ;
      LAYER via2 ;
        RECT 27.000 40.600 27.800 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 29.800 40.600 30.600 41.400 ;
        RECT 27.000 0.600 27.800 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 29.800 0.600 30.600 1.400 ;
      LAYER metal3 ;
        RECT 1.200 52.300 2.000 52.400 ;
        RECT -1.900 51.700 2.000 52.300 ;
        RECT 1.200 51.600 2.000 51.700 ;
        RECT 26.400 40.400 31.200 41.600 ;
        RECT 26.400 0.400 31.200 1.600 ;
      LAYER via3 ;
        RECT 26.800 40.600 27.600 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 30.000 40.600 30.800 41.400 ;
        RECT 26.800 0.600 27.600 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 30.000 0.600 30.800 1.400 ;
      LAYER metal4 ;
        RECT 26.400 -4.000 31.200 64.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 60.400 86.000 61.600 ;
        RECT 1.200 55.800 2.000 60.400 ;
        RECT 6.000 55.800 6.800 60.400 ;
        RECT 17.200 55.800 18.000 60.400 ;
        RECT 26.800 57.800 27.600 60.400 ;
        RECT 30.000 57.800 30.800 60.400 ;
        RECT 41.200 55.800 42.000 60.400 ;
        RECT 47.600 57.800 48.400 60.400 ;
        RECT 50.800 56.400 51.800 60.400 ;
        RECT 57.000 59.800 57.800 60.400 ;
        RECT 57.000 56.400 58.000 59.800 ;
        RECT 66.800 58.300 67.600 60.400 ;
        RECT 68.400 58.300 69.200 59.800 ;
        RECT 66.800 57.700 69.200 58.300 ;
        RECT 66.800 55.800 67.600 57.700 ;
        RECT 65.200 51.600 66.000 53.200 ;
        RECT 68.400 52.400 69.200 57.700 ;
        RECT 71.600 55.800 72.400 60.400 ;
        RECT 76.400 55.800 77.200 60.400 ;
        RECT 81.200 57.800 82.000 60.400 ;
        RECT 68.600 50.200 69.200 52.400 ;
        RECT 68.400 42.200 69.200 50.200 ;
        RECT 4.400 21.600 5.200 26.200 ;
        RECT 14.000 21.600 14.800 24.200 ;
        RECT 17.200 21.600 18.000 24.200 ;
        RECT 28.400 21.600 29.200 26.200 ;
        RECT 34.800 21.600 35.600 24.200 ;
        RECT 42.800 21.600 43.800 25.600 ;
        RECT 49.000 22.200 50.000 25.600 ;
        RECT 49.000 21.600 49.800 22.200 ;
        RECT 52.400 21.600 53.200 24.200 ;
        RECT 55.600 21.600 56.400 24.200 ;
        RECT 58.800 21.600 59.600 24.200 ;
        RECT 65.200 21.600 66.000 24.200 ;
        RECT 69.400 21.600 70.200 26.200 ;
        RECT 71.600 21.600 72.400 28.200 ;
        RECT 79.600 21.600 80.400 26.200 ;
        RECT 0.400 20.400 86.000 21.600 ;
        RECT 4.400 15.800 5.200 20.400 ;
        RECT 14.000 17.800 14.800 20.400 ;
        RECT 17.200 17.800 18.000 20.400 ;
        RECT 28.400 15.800 29.200 20.400 ;
        RECT 34.800 17.800 35.600 20.400 ;
        RECT 42.800 15.800 43.600 20.400 ;
        RECT 54.000 15.800 54.800 20.400 ;
        RECT 63.600 17.800 64.400 20.400 ;
        RECT 66.800 17.800 67.600 20.400 ;
        RECT 78.000 15.800 78.800 20.400 ;
        RECT 84.400 17.800 85.200 20.400 ;
      LAYER via1 ;
        RECT 55.800 60.600 56.600 61.400 ;
        RECT 57.200 60.600 58.000 61.400 ;
        RECT 58.600 60.600 59.400 61.400 ;
        RECT 55.800 20.600 56.600 21.400 ;
        RECT 57.200 20.600 58.000 21.400 ;
        RECT 58.600 20.600 59.400 21.400 ;
      LAYER metal2 ;
        RECT 60.500 63.700 62.700 64.300 ;
        RECT 55.200 60.600 60.000 61.400 ;
        RECT 62.100 56.400 62.700 63.700 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 65.200 56.300 66.000 56.400 ;
        RECT 66.800 56.300 67.600 56.600 ;
        RECT 65.200 55.800 67.600 56.300 ;
        RECT 65.200 55.700 67.500 55.800 ;
        RECT 65.200 55.600 66.000 55.700 ;
        RECT 65.300 52.400 65.900 55.600 ;
        RECT 65.200 51.600 66.000 52.400 ;
        RECT 55.200 20.600 60.000 21.400 ;
      LAYER via2 ;
        RECT 55.800 60.600 56.600 61.400 ;
        RECT 57.200 60.600 58.000 61.400 ;
        RECT 58.600 60.600 59.400 61.400 ;
        RECT 55.800 20.600 56.600 21.400 ;
        RECT 57.200 20.600 58.000 21.400 ;
        RECT 58.600 20.600 59.400 21.400 ;
      LAYER metal3 ;
        RECT 55.200 60.400 60.000 61.600 ;
        RECT 62.000 56.300 62.800 56.400 ;
        RECT 65.200 56.300 66.000 56.400 ;
        RECT 62.000 55.700 66.000 56.300 ;
        RECT 62.000 55.600 62.800 55.700 ;
        RECT 65.200 55.600 66.000 55.700 ;
        RECT 55.200 20.400 60.000 21.600 ;
      LAYER via3 ;
        RECT 55.600 60.600 56.400 61.400 ;
        RECT 57.200 60.600 58.000 61.400 ;
        RECT 58.800 60.600 59.600 61.400 ;
        RECT 55.600 20.600 56.400 21.400 ;
        RECT 57.200 20.600 58.000 21.400 ;
        RECT 58.800 20.600 59.600 21.400 ;
      LAYER metal4 ;
        RECT 55.200 -4.000 60.000 64.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 30.000 55.600 31.600 56.400 ;
        RECT 17.200 25.600 18.800 26.400 ;
        RECT 17.200 15.600 18.800 16.400 ;
        RECT 66.800 15.600 68.400 16.400 ;
      LAYER metal2 ;
        RECT 30.100 63.700 32.300 64.300 ;
        RECT 30.100 56.400 30.700 63.700 ;
        RECT 30.000 55.600 30.800 56.400 ;
        RECT 30.100 50.400 30.700 55.600 ;
        RECT 17.200 49.600 18.000 50.400 ;
        RECT 30.000 49.600 30.800 50.400 ;
        RECT 17.300 26.400 17.900 49.600 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 17.300 16.400 17.900 25.600 ;
        RECT 17.200 15.600 18.000 16.400 ;
        RECT 66.800 15.600 67.600 16.400 ;
      LAYER metal3 ;
        RECT 17.200 50.300 18.000 50.400 ;
        RECT 30.000 50.300 30.800 50.400 ;
        RECT 17.200 49.700 30.800 50.300 ;
        RECT 17.200 49.600 18.000 49.700 ;
        RECT 30.000 49.600 30.800 49.700 ;
        RECT 17.200 16.300 18.000 16.400 ;
        RECT 66.800 16.300 67.600 16.400 ;
        RECT 17.200 15.700 67.600 16.300 ;
        RECT 17.200 15.600 18.000 15.700 ;
        RECT 66.800 15.600 67.600 15.700 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 1.200 53.600 2.000 55.200 ;
      LAYER metal2 ;
        RECT 1.200 53.600 2.000 54.400 ;
      LAYER metal3 ;
        RECT 1.200 53.600 2.000 54.400 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -1.900 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
      LAYER metal4 ;
        RECT 1.000 49.400 2.200 54.600 ;
    END
  END rst
  PIN count[0]
    PORT
      LAYER metal1 ;
        RECT 78.000 52.400 78.800 59.800 ;
        RECT 78.200 50.200 78.800 52.400 ;
        RECT 78.000 42.200 78.800 50.200 ;
      LAYER via1 ;
        RECT 78.000 57.600 78.800 58.400 ;
      LAYER metal2 ;
        RECT 76.500 63.700 78.700 64.300 ;
        RECT 78.100 58.400 78.700 63.700 ;
        RECT 78.000 57.600 78.800 58.400 ;
    END
  END count[0]
  PIN count[1]
    PORT
      LAYER metal1 ;
        RECT 73.200 52.400 74.000 59.800 ;
        RECT 73.400 50.200 74.000 52.400 ;
        RECT 73.200 42.200 74.000 50.200 ;
      LAYER via1 ;
        RECT 73.200 57.600 74.000 58.400 ;
      LAYER metal2 ;
        RECT 71.700 63.700 73.900 64.300 ;
        RECT 73.300 58.400 73.900 63.700 ;
        RECT 73.200 57.600 74.000 58.400 ;
    END
  END count[1]
  PIN count[2]
    PORT
      LAYER metal1 ;
        RECT 81.200 31.800 82.000 39.800 ;
        RECT 81.400 29.600 82.000 31.800 ;
        RECT 81.200 28.300 82.000 29.600 ;
        RECT 84.400 28.300 85.200 28.400 ;
        RECT 81.200 27.700 85.200 28.300 ;
        RECT 81.200 22.200 82.000 27.700 ;
        RECT 84.400 27.600 85.200 27.700 ;
      LAYER metal2 ;
        RECT 84.400 29.600 85.200 30.400 ;
        RECT 84.500 28.400 85.100 29.600 ;
        RECT 84.400 27.600 85.200 28.400 ;
      LAYER metal3 ;
        RECT 84.400 30.300 85.200 30.400 ;
        RECT 84.400 29.700 88.300 30.300 ;
        RECT 84.400 29.600 85.200 29.700 ;
    END
  END count[2]
  PIN count[3]
    PORT
      LAYER metal1 ;
        RECT 41.200 12.400 42.000 19.800 ;
        RECT 41.200 10.200 41.800 12.400 ;
        RECT 41.200 2.200 42.000 10.200 ;
      LAYER via1 ;
        RECT 41.200 3.600 42.000 4.400 ;
      LAYER metal2 ;
        RECT 41.200 3.600 42.000 4.400 ;
        RECT 41.300 -1.700 41.900 3.600 ;
        RECT 41.300 -2.300 43.500 -1.700 ;
    END
  END count[3]
  OBS
      LAYER metal1 ;
        RECT 2.800 42.200 3.600 59.800 ;
        RECT 7.600 55.200 8.400 59.800 ;
        RECT 6.200 54.600 8.400 55.200 ;
        RECT 6.200 51.600 6.800 54.600 ;
        RECT 5.600 50.800 6.800 51.600 ;
        RECT 6.200 50.200 6.800 50.800 ;
        RECT 14.000 53.800 14.800 59.800 ;
        RECT 20.400 56.600 21.200 59.800 ;
        RECT 22.000 57.000 22.800 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 25.200 57.000 26.000 59.800 ;
        RECT 28.400 57.000 29.200 59.800 ;
        RECT 31.600 57.000 32.400 59.800 ;
        RECT 33.200 57.000 34.000 59.800 ;
        RECT 34.800 57.000 35.600 59.800 ;
        RECT 36.400 57.000 37.200 59.800 ;
        RECT 18.600 55.800 21.200 56.600 ;
        RECT 38.000 56.600 38.800 59.800 ;
        RECT 24.600 55.800 29.200 56.400 ;
        RECT 18.600 55.200 19.400 55.800 ;
        RECT 16.400 54.400 19.400 55.200 ;
        RECT 14.000 53.000 22.800 53.800 ;
        RECT 24.600 53.400 25.400 55.800 ;
        RECT 28.400 55.600 29.200 55.800 ;
        RECT 34.600 55.600 35.600 56.400 ;
        RECT 38.000 55.800 40.400 56.600 ;
        RECT 26.800 53.600 27.600 55.200 ;
        RECT 28.400 54.800 29.200 55.000 ;
        RECT 28.400 54.200 32.800 54.800 ;
        RECT 32.000 54.000 32.800 54.200 ;
        RECT 6.200 49.600 8.400 50.200 ;
        RECT 7.600 42.200 8.400 49.600 ;
        RECT 14.000 47.400 14.800 53.000 ;
        RECT 23.400 52.600 25.400 53.400 ;
        RECT 29.200 52.600 32.400 53.400 ;
        RECT 34.800 52.800 35.600 55.600 ;
        RECT 39.600 55.200 40.400 55.800 ;
        RECT 39.600 54.600 41.400 55.200 ;
        RECT 40.600 53.400 41.400 54.600 ;
        RECT 44.400 54.600 45.200 59.800 ;
        RECT 46.000 56.000 46.800 59.800 ;
        RECT 46.000 55.200 47.000 56.000 ;
        RECT 49.200 55.800 50.000 59.800 ;
        RECT 53.600 56.200 55.200 59.800 ;
        RECT 49.200 55.200 51.600 55.800 ;
        RECT 44.400 54.000 45.600 54.600 ;
        RECT 40.600 52.600 44.400 53.400 ;
        RECT 15.400 52.000 16.200 52.200 ;
        RECT 17.200 52.000 18.000 52.400 ;
        RECT 20.400 52.000 21.200 52.400 ;
        RECT 38.000 52.000 38.800 52.600 ;
        RECT 45.000 52.000 45.600 54.000 ;
        RECT 15.400 51.400 38.800 52.000 ;
        RECT 44.800 51.400 45.600 52.000 ;
        RECT 46.200 54.300 47.000 55.200 ;
        RECT 50.800 55.000 51.600 55.200 ;
        RECT 52.200 54.800 53.000 55.600 ;
        RECT 52.200 54.400 52.800 54.800 ;
        RECT 49.200 54.300 50.800 54.400 ;
        RECT 46.200 53.700 50.800 54.300 ;
        RECT 44.800 49.600 45.400 51.400 ;
        RECT 46.200 50.800 47.000 53.700 ;
        RECT 49.200 53.600 50.800 53.700 ;
        RECT 52.000 53.600 52.800 54.400 ;
        RECT 53.600 54.200 54.200 56.200 ;
        RECT 58.800 55.800 59.600 59.800 ;
        RECT 54.800 54.800 56.400 55.600 ;
        RECT 57.000 55.200 59.600 55.800 ;
        RECT 65.200 55.200 66.000 59.800 ;
        RECT 70.000 55.200 70.800 59.800 ;
        RECT 74.800 55.200 75.600 59.800 ;
        RECT 57.000 55.000 57.800 55.200 ;
        RECT 65.200 54.600 67.400 55.200 ;
        RECT 70.000 54.600 72.200 55.200 ;
        RECT 74.800 54.600 77.000 55.200 ;
        RECT 58.000 54.200 59.600 54.400 ;
        RECT 53.600 53.600 54.600 54.200 ;
        RECT 57.400 54.000 59.600 54.200 ;
        RECT 23.600 49.400 24.400 49.600 ;
        RECT 19.000 49.000 24.400 49.400 ;
        RECT 18.200 48.800 24.400 49.000 ;
        RECT 25.400 49.000 34.000 49.600 ;
        RECT 15.600 48.000 17.200 48.800 ;
        RECT 18.200 48.200 19.600 48.800 ;
        RECT 25.400 48.200 26.000 49.000 ;
        RECT 33.200 48.800 34.000 49.000 ;
        RECT 36.400 49.000 45.400 49.600 ;
        RECT 36.400 48.800 37.200 49.000 ;
        RECT 16.600 47.600 17.200 48.000 ;
        RECT 20.200 47.600 26.000 48.200 ;
        RECT 26.600 47.600 29.200 48.400 ;
        RECT 14.000 46.800 16.000 47.400 ;
        RECT 16.600 46.800 20.800 47.600 ;
        RECT 15.400 46.200 16.000 46.800 ;
        RECT 15.400 45.600 16.400 46.200 ;
        RECT 15.600 42.200 16.400 45.600 ;
        RECT 18.800 42.200 19.600 46.800 ;
        RECT 22.000 42.200 22.800 45.000 ;
        RECT 23.600 42.200 24.400 45.000 ;
        RECT 25.200 42.200 26.000 47.000 ;
        RECT 28.400 42.200 29.200 47.000 ;
        RECT 31.600 42.200 32.400 48.400 ;
        RECT 39.600 47.600 42.200 48.400 ;
        RECT 34.800 46.800 39.000 47.600 ;
        RECT 33.200 42.200 34.000 45.000 ;
        RECT 34.800 42.200 35.600 45.000 ;
        RECT 36.400 42.200 37.200 45.000 ;
        RECT 39.600 42.200 40.400 47.600 ;
        RECT 44.800 47.400 45.400 49.000 ;
        RECT 42.800 46.800 45.400 47.400 ;
        RECT 46.000 50.000 47.000 50.800 ;
        RECT 54.000 52.400 54.600 53.600 ;
        RECT 55.200 53.600 59.600 54.000 ;
        RECT 55.200 53.400 58.000 53.600 ;
        RECT 55.200 53.200 56.000 53.400 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 56.600 52.200 57.400 52.400 ;
        RECT 55.800 51.600 57.400 52.200 ;
        RECT 66.800 51.600 67.400 54.600 ;
        RECT 70.000 51.600 70.800 53.200 ;
        RECT 71.600 51.600 72.200 54.600 ;
        RECT 74.800 51.600 75.600 53.200 ;
        RECT 76.400 51.600 77.000 54.600 ;
        RECT 54.000 50.200 54.600 51.600 ;
        RECT 55.800 51.400 56.600 51.600 ;
        RECT 66.800 50.800 68.000 51.600 ;
        RECT 71.600 50.800 72.800 51.600 ;
        RECT 76.400 50.800 77.600 51.600 ;
        RECT 66.800 50.200 67.400 50.800 ;
        RECT 71.600 50.200 72.200 50.800 ;
        RECT 76.400 50.200 77.000 50.800 ;
        RECT 42.800 42.200 43.600 46.800 ;
        RECT 46.000 42.200 46.800 50.000 ;
        RECT 49.200 49.600 51.600 50.200 ;
        RECT 49.200 42.200 50.000 49.600 ;
        RECT 50.800 49.400 51.600 49.600 ;
        RECT 53.600 42.200 55.200 50.200 ;
        RECT 57.000 49.600 59.600 50.200 ;
        RECT 57.000 49.400 57.800 49.600 ;
        RECT 58.800 42.200 59.600 49.600 ;
        RECT 65.200 49.600 67.400 50.200 ;
        RECT 70.000 49.600 72.200 50.200 ;
        RECT 74.800 49.600 77.000 50.200 ;
        RECT 65.200 42.200 66.000 49.600 ;
        RECT 70.000 42.200 70.800 49.600 ;
        RECT 74.800 42.200 75.600 49.600 ;
        RECT 79.600 42.200 80.400 59.800 ;
        RECT 81.200 55.600 82.000 57.200 ;
        RECT 2.800 36.400 3.600 39.800 ;
        RECT 2.600 35.800 3.600 36.400 ;
        RECT 2.600 35.200 3.200 35.800 ;
        RECT 6.000 35.200 6.800 39.800 ;
        RECT 9.200 37.000 10.000 39.800 ;
        RECT 10.800 37.000 11.600 39.800 ;
        RECT 1.200 34.600 3.200 35.200 ;
        RECT 1.200 29.000 2.000 34.600 ;
        RECT 3.800 34.400 8.000 35.200 ;
        RECT 12.400 35.000 13.200 39.800 ;
        RECT 15.600 35.000 16.400 39.800 ;
        RECT 3.800 34.000 4.400 34.400 ;
        RECT 2.800 33.200 4.400 34.000 ;
        RECT 7.400 33.800 13.200 34.400 ;
        RECT 5.400 33.200 6.800 33.800 ;
        RECT 5.400 33.000 11.600 33.200 ;
        RECT 6.200 32.600 11.600 33.000 ;
        RECT 10.800 32.400 11.600 32.600 ;
        RECT 12.600 33.000 13.200 33.800 ;
        RECT 13.800 33.600 16.400 34.400 ;
        RECT 18.800 33.600 19.600 39.800 ;
        RECT 20.400 37.000 21.200 39.800 ;
        RECT 22.000 37.000 22.800 39.800 ;
        RECT 23.600 37.000 24.400 39.800 ;
        RECT 22.000 34.400 26.200 35.200 ;
        RECT 26.800 34.400 27.600 39.800 ;
        RECT 30.000 35.200 30.800 39.800 ;
        RECT 30.000 34.600 32.600 35.200 ;
        RECT 26.800 33.600 29.400 34.400 ;
        RECT 20.400 33.000 21.200 33.200 ;
        RECT 12.600 32.400 21.200 33.000 ;
        RECT 23.600 33.000 24.400 33.200 ;
        RECT 32.000 33.000 32.600 34.600 ;
        RECT 23.600 32.400 32.600 33.000 ;
        RECT 32.000 30.600 32.600 32.400 ;
        RECT 33.200 32.000 34.000 39.800 ;
        RECT 41.200 32.400 42.000 39.800 ;
        RECT 42.800 32.400 43.600 32.600 ;
        RECT 45.600 32.400 47.200 39.800 ;
        RECT 33.200 31.200 34.200 32.000 ;
        RECT 41.200 31.800 43.600 32.400 ;
        RECT 45.200 31.800 47.200 32.400 ;
        RECT 49.400 32.400 50.200 32.600 ;
        RECT 50.800 32.400 51.600 39.800 ;
        RECT 49.400 31.800 51.600 32.400 ;
        RECT 2.600 30.000 26.000 30.600 ;
        RECT 32.000 30.000 32.800 30.600 ;
        RECT 2.600 29.800 3.400 30.000 ;
        RECT 4.400 29.600 5.200 30.000 ;
        RECT 7.600 29.600 8.400 30.000 ;
        RECT 25.200 29.400 26.000 30.000 ;
        RECT 1.200 28.200 10.000 29.000 ;
        RECT 10.600 28.600 12.600 29.400 ;
        RECT 16.400 28.600 19.600 29.400 ;
        RECT 1.200 22.200 2.000 28.200 ;
        RECT 3.600 26.800 6.600 27.600 ;
        RECT 5.800 26.200 6.600 26.800 ;
        RECT 11.800 26.200 12.600 28.600 ;
        RECT 14.000 26.800 14.800 28.400 ;
        RECT 19.200 27.800 20.000 28.000 ;
        RECT 15.600 27.200 20.000 27.800 ;
        RECT 15.600 27.000 16.400 27.200 ;
        RECT 22.000 26.400 22.800 29.200 ;
        RECT 27.800 28.600 31.600 29.400 ;
        RECT 27.800 27.400 28.600 28.600 ;
        RECT 32.200 28.000 32.800 30.000 ;
        RECT 15.600 26.200 16.400 26.400 ;
        RECT 5.800 25.400 8.400 26.200 ;
        RECT 11.800 25.600 16.400 26.200 ;
        RECT 21.800 25.600 22.800 26.400 ;
        RECT 26.800 26.800 28.600 27.400 ;
        RECT 31.600 27.400 32.800 28.000 ;
        RECT 26.800 26.200 27.600 26.800 ;
        RECT 7.600 22.200 8.400 25.400 ;
        RECT 25.200 25.400 27.600 26.200 ;
        RECT 9.200 22.200 10.000 25.000 ;
        RECT 10.800 22.200 11.600 25.000 ;
        RECT 12.400 22.200 13.200 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 18.800 22.200 19.600 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 22.000 22.200 22.800 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.400 ;
        RECT 31.600 22.200 32.400 27.400 ;
        RECT 33.400 26.800 34.200 31.200 ;
        RECT 45.200 30.400 45.800 31.800 ;
        RECT 49.400 31.200 50.000 31.800 ;
        RECT 46.600 30.600 50.000 31.200 ;
        RECT 46.600 30.400 47.400 30.600 ;
        RECT 44.400 29.800 45.800 30.400 ;
        RECT 54.000 30.300 54.800 39.800 ;
        RECT 56.200 32.600 57.000 39.800 ;
        RECT 56.200 31.800 58.000 32.600 ;
        RECT 65.200 31.800 66.000 39.800 ;
        RECT 66.800 32.400 67.600 39.800 ;
        RECT 70.000 32.400 70.800 39.800 ;
        RECT 73.200 35.800 74.000 39.800 ;
        RECT 73.400 35.600 74.000 35.800 ;
        RECT 76.400 35.800 77.200 39.800 ;
        RECT 76.400 35.600 77.000 35.800 ;
        RECT 73.400 35.000 77.000 35.600 ;
        RECT 74.800 32.800 75.600 34.400 ;
        RECT 76.400 32.400 77.000 35.000 ;
        RECT 78.000 32.400 78.800 39.800 ;
        RECT 66.800 31.800 70.800 32.400 ;
        RECT 55.600 30.300 56.400 31.200 ;
        RECT 48.800 29.800 49.600 30.000 ;
        RECT 44.400 29.600 46.200 29.800 ;
        RECT 45.200 29.200 46.200 29.600 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 41.200 28.300 42.800 28.400 ;
        RECT 39.600 27.700 42.800 28.300 ;
        RECT 39.600 27.600 40.400 27.700 ;
        RECT 41.200 27.600 42.800 27.700 ;
        RECT 44.000 27.600 44.800 28.400 ;
        RECT 44.200 27.200 44.800 27.600 ;
        RECT 42.800 26.800 43.600 27.000 ;
        RECT 33.200 26.000 34.200 26.800 ;
        RECT 41.200 26.200 43.600 26.800 ;
        RECT 44.200 26.400 45.000 27.200 ;
        RECT 33.200 22.200 34.000 26.000 ;
        RECT 41.200 22.200 42.000 26.200 ;
        RECT 45.600 25.800 46.200 29.200 ;
        RECT 47.000 29.200 49.600 29.800 ;
        RECT 54.000 29.700 56.400 30.300 ;
        RECT 47.000 28.600 47.600 29.200 ;
        RECT 46.800 27.800 47.600 28.600 ;
        RECT 50.000 28.300 51.600 28.400 ;
        RECT 50.000 28.200 53.100 28.300 ;
        RECT 48.200 27.700 53.100 28.200 ;
        RECT 48.200 27.600 51.600 27.700 ;
        RECT 48.200 27.200 48.800 27.600 ;
        RECT 46.800 26.600 48.800 27.200 ;
        RECT 49.400 26.800 50.200 27.000 ;
        RECT 46.800 26.400 48.400 26.600 ;
        RECT 49.400 26.200 51.600 26.800 ;
        RECT 52.500 26.400 53.100 27.700 ;
        RECT 45.600 24.400 47.200 25.800 ;
        RECT 44.400 23.600 47.200 24.400 ;
        RECT 45.600 22.200 47.200 23.600 ;
        RECT 50.800 22.200 51.600 26.200 ;
        RECT 52.400 24.800 53.200 26.400 ;
        RECT 54.000 22.200 54.800 29.700 ;
        RECT 55.600 29.600 56.400 29.700 ;
        RECT 57.200 28.400 57.800 31.800 ;
        RECT 65.400 30.400 66.000 31.800 ;
        RECT 69.200 30.400 70.000 30.800 ;
        RECT 65.200 29.800 67.600 30.400 ;
        RECT 69.200 30.300 70.800 30.400 ;
        RECT 71.600 30.300 72.400 32.400 ;
        RECT 76.400 31.600 77.200 32.400 ;
        RECT 78.000 31.800 80.200 32.400 ;
        RECT 69.200 29.800 72.400 30.300 ;
        RECT 65.200 29.600 66.000 29.800 ;
        RECT 55.600 28.300 56.400 28.400 ;
        RECT 57.200 28.300 58.000 28.400 ;
        RECT 67.000 28.300 67.600 29.800 ;
        RECT 70.000 29.700 72.400 29.800 ;
        RECT 70.000 29.600 70.800 29.700 ;
        RECT 73.200 29.600 74.800 30.400 ;
        RECT 55.600 27.700 58.000 28.300 ;
        RECT 55.600 27.600 56.400 27.700 ;
        RECT 57.200 27.600 58.000 27.700 ;
        RECT 62.100 27.700 67.600 28.300 ;
        RECT 57.200 24.200 57.800 27.600 ;
        RECT 58.800 26.300 59.600 26.400 ;
        RECT 62.100 26.300 62.700 27.700 ;
        RECT 58.800 25.700 62.700 26.300 ;
        RECT 58.800 24.800 59.600 25.700 ;
        RECT 65.200 25.600 66.000 26.400 ;
        RECT 67.000 26.200 67.600 27.700 ;
        RECT 68.400 28.300 69.200 29.200 ;
        RECT 76.400 28.400 77.000 31.600 ;
        RECT 79.600 31.200 80.200 31.800 ;
        RECT 79.600 30.400 80.800 31.200 ;
        RECT 78.000 28.800 78.800 30.400 ;
        RECT 70.000 28.300 70.800 28.400 ;
        RECT 68.400 27.700 70.800 28.300 ;
        RECT 75.400 28.200 77.000 28.400 ;
        RECT 68.400 27.600 69.200 27.700 ;
        RECT 70.000 27.600 70.800 27.700 ;
        RECT 75.200 27.800 77.000 28.200 ;
        RECT 75.200 26.400 76.000 27.800 ;
        RECT 79.600 27.400 80.200 30.400 ;
        RECT 65.400 24.800 66.200 25.600 ;
        RECT 57.200 22.200 58.000 24.200 ;
        RECT 66.800 22.200 67.600 26.200 ;
        RECT 74.800 25.600 76.000 26.400 ;
        RECT 75.200 22.200 76.000 25.600 ;
        RECT 78.000 26.800 80.200 27.400 ;
        RECT 78.000 22.200 78.800 26.800 ;
        RECT 1.200 13.800 2.000 19.800 ;
        RECT 7.600 16.600 8.400 19.800 ;
        RECT 9.200 17.000 10.000 19.800 ;
        RECT 10.800 17.000 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 5.800 15.800 8.400 16.600 ;
        RECT 25.200 16.600 26.000 19.800 ;
        RECT 11.800 15.800 16.400 16.400 ;
        RECT 5.800 15.200 6.600 15.800 ;
        RECT 3.600 14.400 6.600 15.200 ;
        RECT 1.200 13.000 10.000 13.800 ;
        RECT 11.800 13.400 12.600 15.800 ;
        RECT 15.600 15.600 16.400 15.800 ;
        RECT 21.800 15.600 22.800 16.400 ;
        RECT 25.200 15.800 27.600 16.600 ;
        RECT 14.000 13.600 14.800 15.200 ;
        RECT 15.600 14.800 16.400 15.000 ;
        RECT 15.600 14.200 20.000 14.800 ;
        RECT 19.200 14.000 20.000 14.200 ;
        RECT 1.200 7.400 2.000 13.000 ;
        RECT 10.600 12.600 12.600 13.400 ;
        RECT 16.400 12.600 19.600 13.400 ;
        RECT 22.000 12.800 22.800 15.600 ;
        RECT 26.800 15.200 27.600 15.800 ;
        RECT 26.800 14.600 28.600 15.200 ;
        RECT 27.800 13.400 28.600 14.600 ;
        RECT 31.600 14.600 32.400 19.800 ;
        RECT 33.200 16.300 34.000 19.800 ;
        RECT 39.600 16.300 40.400 16.400 ;
        RECT 33.200 15.700 40.400 16.300 ;
        RECT 33.200 15.200 34.200 15.700 ;
        RECT 39.600 15.600 40.400 15.700 ;
        RECT 44.400 15.200 45.200 19.800 ;
        RECT 31.600 14.000 32.800 14.600 ;
        RECT 27.800 12.600 31.600 13.400 ;
        RECT 2.600 12.000 3.400 12.200 ;
        RECT 4.400 12.000 5.200 12.400 ;
        RECT 7.600 12.000 8.400 12.400 ;
        RECT 25.200 12.000 26.000 12.600 ;
        RECT 32.200 12.000 32.800 14.000 ;
        RECT 2.600 11.400 26.000 12.000 ;
        RECT 32.000 11.400 32.800 12.000 ;
        RECT 32.000 9.600 32.600 11.400 ;
        RECT 33.400 10.800 34.200 15.200 ;
        RECT 43.000 14.600 45.200 15.200 ;
        RECT 43.000 11.600 43.600 14.600 ;
        RECT 50.800 13.800 51.600 19.800 ;
        RECT 57.200 16.600 58.000 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 60.400 17.000 61.200 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 65.200 17.000 66.000 19.800 ;
        RECT 68.400 17.000 69.200 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 71.600 17.000 72.400 19.800 ;
        RECT 73.200 17.000 74.000 19.800 ;
        RECT 55.400 15.800 58.000 16.600 ;
        RECT 74.800 16.600 75.600 19.800 ;
        RECT 61.400 15.800 66.000 16.400 ;
        RECT 55.400 15.200 56.200 15.800 ;
        RECT 53.200 14.400 56.200 15.200 ;
        RECT 44.400 11.600 45.200 13.200 ;
        RECT 50.800 13.000 59.600 13.800 ;
        RECT 61.400 13.400 62.200 15.800 ;
        RECT 65.200 15.600 66.000 15.800 ;
        RECT 71.400 15.600 72.400 16.400 ;
        RECT 74.800 15.800 77.200 16.600 ;
        RECT 63.600 13.600 64.400 15.200 ;
        RECT 65.200 14.800 66.000 15.000 ;
        RECT 65.200 14.200 69.600 14.800 ;
        RECT 68.800 14.000 69.600 14.200 ;
        RECT 42.400 10.800 43.600 11.600 ;
        RECT 10.800 9.400 11.600 9.600 ;
        RECT 6.200 9.000 11.600 9.400 ;
        RECT 5.400 8.800 11.600 9.000 ;
        RECT 12.600 9.000 21.200 9.600 ;
        RECT 2.800 8.000 4.400 8.800 ;
        RECT 5.400 8.200 6.800 8.800 ;
        RECT 12.600 8.200 13.200 9.000 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 23.600 9.000 32.600 9.600 ;
        RECT 23.600 8.800 24.400 9.000 ;
        RECT 3.800 7.600 4.400 8.000 ;
        RECT 7.400 7.600 13.200 8.200 ;
        RECT 13.800 7.600 16.400 8.400 ;
        RECT 1.200 6.800 3.200 7.400 ;
        RECT 3.800 6.800 8.000 7.600 ;
        RECT 2.600 6.200 3.200 6.800 ;
        RECT 2.600 5.600 3.600 6.200 ;
        RECT 2.800 2.200 3.600 5.600 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 5.000 ;
        RECT 10.800 2.200 11.600 5.000 ;
        RECT 12.400 2.200 13.200 7.000 ;
        RECT 15.600 2.200 16.400 7.000 ;
        RECT 18.800 2.200 19.600 8.400 ;
        RECT 26.800 7.600 29.400 8.400 ;
        RECT 22.000 6.800 26.200 7.600 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 5.000 ;
        RECT 23.600 2.200 24.400 5.000 ;
        RECT 26.800 2.200 27.600 7.600 ;
        RECT 32.000 7.400 32.600 9.000 ;
        RECT 30.000 6.800 32.600 7.400 ;
        RECT 33.200 10.000 34.200 10.800 ;
        RECT 43.000 10.200 43.600 10.800 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.200 2.200 34.000 10.000 ;
        RECT 43.000 9.600 45.200 10.200 ;
        RECT 44.400 2.200 45.200 9.600 ;
        RECT 50.800 7.400 51.600 13.000 ;
        RECT 60.200 12.600 62.200 13.400 ;
        RECT 66.000 12.600 69.200 13.400 ;
        RECT 71.600 12.800 72.400 15.600 ;
        RECT 76.400 15.200 77.200 15.800 ;
        RECT 76.400 14.600 78.200 15.200 ;
        RECT 77.400 13.400 78.200 14.600 ;
        RECT 81.200 14.600 82.000 19.800 ;
        RECT 82.800 16.000 83.600 19.800 ;
        RECT 82.800 15.200 83.800 16.000 ;
        RECT 81.200 14.000 82.400 14.600 ;
        RECT 77.400 12.600 81.200 13.400 ;
        RECT 52.200 12.000 53.000 12.200 ;
        RECT 54.000 12.000 54.800 12.400 ;
        RECT 57.200 12.000 58.000 12.400 ;
        RECT 74.800 12.000 75.600 12.600 ;
        RECT 81.800 12.000 82.400 14.000 ;
        RECT 52.200 11.400 75.600 12.000 ;
        RECT 81.600 11.400 82.400 12.000 ;
        RECT 81.600 9.600 82.200 11.400 ;
        RECT 83.000 10.800 83.800 15.200 ;
        RECT 60.400 9.400 61.200 9.600 ;
        RECT 55.800 9.000 61.200 9.400 ;
        RECT 55.000 8.800 61.200 9.000 ;
        RECT 62.200 9.000 70.800 9.600 ;
        RECT 52.400 8.000 54.000 8.800 ;
        RECT 55.000 8.200 56.400 8.800 ;
        RECT 62.200 8.200 62.800 9.000 ;
        RECT 70.000 8.800 70.800 9.000 ;
        RECT 73.200 9.000 82.200 9.600 ;
        RECT 73.200 8.800 74.000 9.000 ;
        RECT 53.400 7.600 54.000 8.000 ;
        RECT 57.000 7.600 62.800 8.200 ;
        RECT 63.400 7.600 66.000 8.400 ;
        RECT 50.800 6.800 52.800 7.400 ;
        RECT 53.400 6.800 57.600 7.600 ;
        RECT 52.200 6.200 52.800 6.800 ;
        RECT 52.200 5.600 53.200 6.200 ;
        RECT 52.400 2.200 53.200 5.600 ;
        RECT 55.600 2.200 56.400 6.800 ;
        RECT 58.800 2.200 59.600 5.000 ;
        RECT 60.400 2.200 61.200 5.000 ;
        RECT 62.000 2.200 62.800 7.000 ;
        RECT 65.200 2.200 66.000 7.000 ;
        RECT 68.400 2.200 69.200 8.400 ;
        RECT 76.400 7.600 79.000 8.400 ;
        RECT 71.600 6.800 75.800 7.600 ;
        RECT 70.000 2.200 70.800 5.000 ;
        RECT 71.600 2.200 72.400 5.000 ;
        RECT 73.200 2.200 74.000 5.000 ;
        RECT 76.400 2.200 77.200 7.600 ;
        RECT 81.600 7.400 82.200 9.000 ;
        RECT 79.600 6.800 82.200 7.400 ;
        RECT 82.800 10.000 83.800 10.800 ;
        RECT 79.600 2.200 80.400 6.800 ;
        RECT 82.800 2.200 83.600 10.000 ;
      LAYER via1 ;
        RECT 22.000 53.000 22.800 53.800 ;
        RECT 2.800 43.600 3.600 44.400 ;
        RECT 31.600 52.600 32.400 53.400 ;
        RECT 54.000 57.600 54.800 58.400 ;
        RECT 17.200 51.600 18.000 52.400 ;
        RECT 55.600 54.800 56.400 55.600 ;
        RECT 23.600 48.800 24.400 49.600 ;
        RECT 28.400 47.600 29.200 48.400 ;
        RECT 25.200 46.200 26.000 47.000 ;
        RECT 22.000 44.200 22.800 45.000 ;
        RECT 23.600 44.200 24.400 45.000 ;
        RECT 28.400 46.200 29.200 47.000 ;
        RECT 31.600 46.200 32.400 47.000 ;
        RECT 33.200 44.200 34.000 45.000 ;
        RECT 34.800 44.200 35.600 45.000 ;
        RECT 36.400 44.200 37.200 45.000 ;
        RECT 58.800 53.600 59.600 54.400 ;
        RECT 79.600 43.600 80.400 44.400 ;
        RECT 18.800 35.000 19.600 35.800 ;
        RECT 15.600 33.600 16.400 34.400 ;
        RECT 20.400 32.400 21.200 33.200 ;
        RECT 33.200 33.600 34.000 34.400 ;
        RECT 42.800 31.800 43.600 32.600 ;
        RECT 9.200 28.200 10.000 29.000 ;
        RECT 18.800 28.600 19.600 29.400 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 9.200 24.200 10.000 25.000 ;
        RECT 10.800 24.200 11.600 25.000 ;
        RECT 12.400 24.200 13.200 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 18.800 24.200 19.600 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 22.000 24.200 22.800 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 74.800 33.600 75.600 34.400 ;
        RECT 42.800 26.200 43.600 27.000 ;
        RECT 47.600 26.400 48.400 27.200 ;
        RECT 71.600 31.600 72.400 32.400 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 9.200 13.000 10.000 13.800 ;
        RECT 18.800 12.600 19.600 13.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 58.800 13.000 59.600 13.800 ;
        RECT 10.800 8.800 11.600 9.600 ;
        RECT 15.600 7.600 16.400 8.400 ;
        RECT 12.400 6.200 13.200 7.000 ;
        RECT 9.200 4.200 10.000 5.000 ;
        RECT 10.800 4.200 11.600 5.000 ;
        RECT 15.600 6.200 16.400 7.000 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 22.000 4.200 22.800 5.000 ;
        RECT 23.600 4.200 24.400 5.000 ;
        RECT 68.400 12.600 69.200 13.400 ;
        RECT 82.800 17.600 83.600 18.400 ;
        RECT 54.000 11.600 54.800 12.400 ;
        RECT 60.400 8.800 61.200 9.600 ;
        RECT 65.200 7.600 66.000 8.400 ;
        RECT 62.000 6.200 62.800 7.000 ;
        RECT 58.800 4.200 59.600 5.000 ;
        RECT 60.400 4.200 61.200 5.000 ;
        RECT 65.200 6.200 66.000 7.000 ;
        RECT 68.400 6.200 69.200 7.000 ;
        RECT 70.000 4.200 70.800 5.000 ;
        RECT 71.600 4.200 72.400 5.000 ;
        RECT 73.200 4.200 74.000 5.000 ;
      LAYER metal2 ;
        RECT 2.800 51.600 3.600 52.400 ;
        RECT 17.200 51.600 18.000 52.400 ;
        RECT 2.900 44.400 3.500 51.600 ;
        RECT 2.800 43.600 3.600 44.400 ;
        RECT 22.000 44.200 22.800 57.800 ;
        RECT 23.600 44.200 24.400 57.800 ;
        RECT 25.200 46.200 26.000 57.800 ;
        RECT 26.800 57.600 27.600 58.400 ;
        RECT 26.900 54.400 27.500 57.600 ;
        RECT 26.800 53.600 27.600 54.400 ;
        RECT 28.400 46.200 29.200 57.800 ;
        RECT 31.600 46.200 32.400 57.800 ;
        RECT 33.200 44.200 34.000 57.800 ;
        RECT 34.800 44.200 35.600 57.800 ;
        RECT 36.400 44.200 37.200 57.800 ;
        RECT 54.000 57.600 54.800 58.400 ;
        RECT 50.800 55.000 51.600 55.800 ;
        RECT 57.000 55.600 57.800 55.800 ;
        RECT 81.200 55.600 82.000 56.400 ;
        RECT 52.200 55.000 57.800 55.600 ;
        RECT 49.200 53.600 50.000 54.400 ;
        RECT 50.800 54.200 51.400 55.000 ;
        RECT 52.200 54.800 53.000 55.000 ;
        RECT 55.600 54.800 56.400 55.000 ;
        RECT 50.800 53.600 56.400 54.200 ;
        RECT 50.800 50.200 51.400 53.600 ;
        RECT 55.800 52.200 56.400 53.600 ;
        RECT 55.800 51.400 56.600 52.200 ;
        RECT 57.200 50.200 57.800 55.000 ;
        RECT 58.800 53.600 59.600 54.400 ;
        RECT 70.000 53.600 70.800 54.400 ;
        RECT 58.900 52.400 59.500 53.600 ;
        RECT 70.100 52.400 70.700 53.600 ;
        RECT 81.300 52.400 81.900 55.600 ;
        RECT 58.800 51.600 59.600 52.400 ;
        RECT 70.000 51.600 70.800 52.400 ;
        RECT 71.600 51.600 72.400 52.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 81.200 52.300 82.000 52.400 ;
        RECT 81.200 51.700 83.500 52.300 ;
        RECT 81.200 51.600 82.000 51.700 ;
        RECT 50.800 49.400 51.600 50.200 ;
        RECT 57.000 49.400 57.800 50.200 ;
        RECT 2.900 30.300 3.500 43.600 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 2.900 29.700 5.200 30.300 ;
        RECT 4.400 29.600 5.200 29.700 ;
        RECT 4.500 12.400 5.100 29.600 ;
        RECT 9.200 24.200 10.000 37.800 ;
        RECT 10.800 24.200 11.600 37.800 ;
        RECT 12.400 24.200 13.200 35.800 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 15.600 24.200 16.400 35.800 ;
        RECT 18.800 24.200 19.600 35.800 ;
        RECT 20.400 24.200 21.200 37.800 ;
        RECT 22.000 24.200 22.800 37.800 ;
        RECT 23.600 24.200 24.400 37.800 ;
        RECT 33.200 33.600 34.000 34.400 ;
        RECT 65.200 33.600 66.000 34.400 ;
        RECT 42.800 31.800 43.600 32.600 ;
        RECT 49.400 31.800 50.200 32.600 ;
        RECT 42.800 28.400 43.400 31.800 ;
        RECT 46.800 28.400 47.600 28.600 ;
        RECT 39.600 27.600 40.400 28.400 ;
        RECT 42.800 27.800 47.600 28.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 9.200 4.200 10.000 17.800 ;
        RECT 10.800 4.200 11.600 17.800 ;
        RECT 12.400 6.200 13.200 17.800 ;
        RECT 14.000 17.600 14.800 18.400 ;
        RECT 14.100 14.400 14.700 17.600 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 15.600 6.200 16.400 17.800 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 4.200 22.800 17.800 ;
        RECT 23.600 4.200 24.400 17.800 ;
        RECT 39.700 16.400 40.300 27.600 ;
        RECT 42.800 27.000 43.400 27.800 ;
        RECT 44.200 27.000 45.000 27.200 ;
        RECT 47.600 27.000 48.400 27.200 ;
        RECT 49.600 27.000 50.200 31.800 ;
        RECT 55.600 27.600 56.400 28.400 ;
        RECT 42.800 26.200 43.600 27.000 ;
        RECT 44.200 26.400 48.400 27.000 ;
        RECT 47.600 25.600 48.400 26.400 ;
        RECT 49.400 26.200 50.200 27.000 ;
        RECT 65.300 26.400 65.900 33.600 ;
        RECT 70.100 30.400 70.700 51.600 ;
        RECT 71.700 32.400 72.300 51.600 ;
        RECT 79.600 43.600 80.400 44.400 ;
        RECT 74.800 33.600 75.600 34.400 ;
        RECT 78.000 33.600 78.800 34.400 ;
        RECT 71.600 31.600 72.400 32.400 ;
        RECT 78.100 30.400 78.700 33.600 ;
        RECT 70.000 29.600 70.800 30.400 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 70.100 28.400 70.700 29.600 ;
        RECT 70.000 27.600 70.800 28.400 ;
        RECT 65.200 25.600 66.000 26.400 ;
        RECT 74.800 25.600 75.600 26.400 ;
        RECT 44.400 23.600 45.200 24.400 ;
        RECT 44.500 18.400 45.100 23.600 ;
        RECT 44.400 17.600 45.200 18.400 ;
        RECT 39.600 15.600 40.400 16.400 ;
        RECT 25.200 13.600 26.000 14.400 ;
        RECT 25.300 12.400 25.900 13.600 ;
        RECT 39.700 12.400 40.300 15.600 ;
        RECT 54.000 13.600 54.800 14.400 ;
        RECT 54.100 12.400 54.700 13.600 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 39.600 11.600 40.400 12.400 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 54.000 11.600 54.800 12.400 ;
        RECT 58.800 4.200 59.600 17.800 ;
        RECT 60.400 4.200 61.200 17.800 ;
        RECT 62.000 6.200 62.800 17.800 ;
        RECT 63.600 13.600 64.400 14.400 ;
        RECT 65.200 6.200 66.000 17.800 ;
        RECT 68.400 6.200 69.200 17.800 ;
        RECT 70.000 4.200 70.800 17.800 ;
        RECT 71.600 4.200 72.400 17.800 ;
        RECT 73.200 4.200 74.000 17.800 ;
        RECT 79.700 14.400 80.300 43.600 ;
        RECT 82.900 18.400 83.500 51.700 ;
        RECT 82.800 17.600 83.600 18.400 ;
        RECT 79.600 13.600 80.400 14.400 ;
      LAYER metal3 ;
        RECT 26.800 58.300 27.600 58.400 ;
        RECT 54.000 58.300 54.800 58.400 ;
        RECT 26.800 57.700 54.800 58.300 ;
        RECT 26.800 57.600 27.600 57.700 ;
        RECT 54.000 57.600 54.800 57.700 ;
        RECT 49.200 54.300 50.000 54.400 ;
        RECT 70.000 54.300 70.800 54.400 ;
        RECT 49.200 53.700 70.800 54.300 ;
        RECT 49.200 53.600 50.000 53.700 ;
        RECT 70.000 53.600 70.800 53.700 ;
        RECT 2.800 52.300 3.600 52.400 ;
        RECT 17.200 52.300 18.000 52.400 ;
        RECT 2.800 51.700 18.000 52.300 ;
        RECT 2.800 51.600 3.600 51.700 ;
        RECT 17.200 51.600 18.000 51.700 ;
        RECT 58.800 52.300 59.600 52.400 ;
        RECT 71.600 52.300 72.400 52.400 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 81.200 52.300 82.000 52.400 ;
        RECT 58.800 51.700 82.000 52.300 ;
        RECT 58.800 51.600 59.600 51.700 ;
        RECT 71.600 51.600 72.400 51.700 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 81.200 51.600 82.000 51.700 ;
        RECT 33.200 34.300 34.000 34.400 ;
        RECT 65.200 34.300 66.000 34.400 ;
        RECT 74.800 34.300 75.600 34.400 ;
        RECT 78.000 34.300 78.800 34.400 ;
        RECT 33.200 33.700 78.800 34.300 ;
        RECT 33.200 33.600 34.000 33.700 ;
        RECT 65.200 33.600 66.000 33.700 ;
        RECT 74.800 33.600 75.600 33.700 ;
        RECT 78.000 33.600 78.800 33.700 ;
        RECT 70.000 30.300 70.800 30.400 ;
        RECT 73.200 30.300 74.000 30.400 ;
        RECT 70.000 29.700 74.000 30.300 ;
        RECT 70.000 29.600 70.800 29.700 ;
        RECT 73.200 29.600 74.000 29.700 ;
        RECT 14.000 28.300 14.800 28.400 ;
        RECT 55.600 28.300 56.400 28.400 ;
        RECT 14.000 27.700 56.400 28.300 ;
        RECT 14.000 27.600 14.800 27.700 ;
        RECT 55.600 27.600 56.400 27.700 ;
        RECT 47.600 26.300 48.400 26.400 ;
        RECT 74.800 26.300 75.600 26.400 ;
        RECT 47.600 25.700 75.600 26.300 ;
        RECT 47.600 25.600 48.400 25.700 ;
        RECT 74.800 25.600 75.600 25.700 ;
        RECT 14.000 18.300 14.800 18.400 ;
        RECT 44.400 18.300 45.200 18.400 ;
        RECT 14.000 17.700 45.200 18.300 ;
        RECT 14.000 17.600 14.800 17.700 ;
        RECT 44.400 17.600 45.200 17.700 ;
        RECT 25.200 14.300 26.000 14.400 ;
        RECT 54.000 14.300 54.800 14.400 ;
        RECT 25.200 13.700 54.800 14.300 ;
        RECT 25.200 13.600 26.000 13.700 ;
        RECT 54.000 13.600 54.800 13.700 ;
        RECT 63.600 14.300 64.400 14.400 ;
        RECT 79.600 14.300 80.400 14.400 ;
        RECT 63.600 13.700 80.400 14.300 ;
        RECT 63.600 13.600 64.400 13.700 ;
        RECT 79.600 13.600 80.400 13.700 ;
        RECT 39.600 12.300 40.400 12.400 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 39.600 11.700 45.200 12.300 ;
        RECT 39.600 11.600 40.400 11.700 ;
        RECT 44.400 11.600 45.200 11.700 ;
  END
END counter
END LIBRARY


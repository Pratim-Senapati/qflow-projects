magic
tech scmos
timestamp 1739818576
<< metal1 >>
rect 3 1010 1497 1497
rect 3 520 1500 1010
rect 3 489 1497 520
rect 3 3 1500 489
rect 490 0 979 3
rect 1011 0 1500 3
<< metal2 >>
rect 3 1010 1497 1497
rect 3 648 1500 1010
rect 3 626 1497 648
rect 3 520 1500 626
rect 3 489 1497 520
rect 3 384 1500 489
rect 3 362 1497 384
rect 3 3 1500 362
rect 490 0 852 3
rect 874 0 979 3
rect 1011 0 1116 3
rect 1138 0 1500 3
<< metal3 >>
rect 3 3 1497 1497
<< metal4 >>
rect 3 3 1497 1497
<< properties >>
string LEFsite corner
string LEFclass ENDCAP TOPLEFT
string FIXED_BBOX 0 0 1500 1500
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>

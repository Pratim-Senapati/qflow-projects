magic
tech scmos
timestamp 0
<< properties >>
string LEFclass CORE
string FIXED_BBOX 0 0 8 100
string LEFsymmetry Y
string LEFview TRUE
<< end >>
